module rvclkhdr(
  output  io_l1clk,
  input   io_clk,
  input   io_en,
  input   io_scan_mode
);
  wire  clkhdr_Q; // @[lib.scala 334:26]
  wire  clkhdr_CK; // @[lib.scala 334:26]
  wire  clkhdr_EN; // @[lib.scala 334:26]
  wire  clkhdr_SE; // @[lib.scala 334:26]
  gated_latch clkhdr ( // @[lib.scala 334:26]
    .Q(clkhdr_Q),
    .CK(clkhdr_CK),
    .EN(clkhdr_EN),
    .SE(clkhdr_SE)
  );
  assign io_l1clk = clkhdr_Q; // @[lib.scala 335:14]
  assign clkhdr_CK = io_clk; // @[lib.scala 336:18]
  assign clkhdr_EN = io_en; // @[lib.scala 337:18]
  assign clkhdr_SE = io_scan_mode; // @[lib.scala 338:18]
endmodule
module ifu_mem_ctl(
  input         clock,
  input         reset,
  input         io_free_clk,
  input         io_active_clk,
  input         io_exu_flush_final,
  input         io_dec_mem_ctrl_dec_tlu_flush_err_wb,
  input         io_dec_mem_ctrl_dec_tlu_i0_commit_cmt,
  input         io_dec_mem_ctrl_dec_tlu_force_halt,
  input         io_dec_mem_ctrl_dec_tlu_fence_i_wb,
  input  [70:0] io_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_wrdata,
  input  [16:0] io_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_dicawics,
  input         io_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_rd_valid,
  input         io_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_wr_valid,
  input         io_dec_mem_ctrl_dec_tlu_core_ecc_disable,
  output        io_dec_mem_ctrl_ifu_pmu_ic_miss,
  output        io_dec_mem_ctrl_ifu_pmu_ic_hit,
  output        io_dec_mem_ctrl_ifu_pmu_bus_error,
  output        io_dec_mem_ctrl_ifu_pmu_bus_busy,
  output        io_dec_mem_ctrl_ifu_ic_error_start,
  output        io_dec_mem_ctrl_ifu_iccm_rd_ecc_single_err,
  output [70:0] io_dec_mem_ctrl_ifu_ic_debug_rd_data,
  output        io_dec_mem_ctrl_ifu_ic_debug_rd_data_valid,
  output        io_dec_mem_ctrl_ifu_miss_state_idle,
  input  [30:0] io_ifc_fetch_addr_bf,
  input         io_ifc_fetch_uncacheable_bf,
  input         io_ifc_fetch_req_bf,
  input         io_ifc_fetch_req_bf_raw,
  input         io_ifc_iccm_access_bf,
  input         io_ifc_region_acc_fault_bf,
  input         io_ifc_dma_access_ok,
  input         io_ifu_bp_hit_taken_f,
  input         io_ifu_bp_inst_mask_f,
  output        io_ifu_axi_ar_valid,
  output [31:0] io_ifu_axi_ar_bits_addr,
  input         io_ifu_bus_clk_en,
  input         io_dma_mem_ctl_dma_iccm_req,
  input  [31:0] io_dma_mem_ctl_dma_mem_addr,
  input  [2:0]  io_dma_mem_ctl_dma_mem_sz,
  input         io_dma_mem_ctl_dma_mem_write,
  input  [63:0] io_dma_mem_ctl_dma_mem_wdata,
  input  [2:0]  io_dma_mem_ctl_dma_mem_tag,
  output [14:0] io_iccm_rw_addr,
  output        io_iccm_buf_correct_ecc,
  output        io_iccm_correction_state,
  output        io_iccm_wren,
  output        io_iccm_rden,
  output [2:0]  io_iccm_wr_size,
  output [77:0] io_iccm_wr_data,
  input  [63:0] io_iccm_rd_data,
  input  [77:0] io_iccm_rd_data_ecc,
  output [30:0] io_ic_rw_addr,
  output [1:0]  io_ic_tag_valid,
  output        io_ic_rd_en,
  output [70:0] io_ic_debug_wr_data,
  output [9:0]  io_ic_debug_addr,
  input  [63:0] io_ic_rd_data,
  input  [70:0] io_ic_debug_rd_data,
  input  [25:0] io_ic_tag_debug_rd_data,
  input  [1:0]  io_ic_eccerr,
  input  [1:0]  io_ic_rd_hit,
  input         io_ic_tag_perr,
  output        io_ic_debug_rd_en,
  output        io_ic_debug_wr_en,
  output        io_ic_debug_tag_array,
  output [1:0]  io_ic_debug_way,
  output [63:0] io_ic_premux_data,
  output        io_ic_sel_premux_data,
  input  [1:0]  io_ifu_fetch_val,
  output        io_ifu_ic_mb_empty,
  output        io_ic_dma_active,
  output        io_iccm_dma_ecc_error,
  output        io_iccm_dma_rvalid,
  output [63:0] io_iccm_dma_rdata,
  output [2:0]  io_iccm_dma_rtag,
  output        io_iccm_ready,
  input         io_dec_tlu_flush_lower_wb,
  output        io_iccm_rd_ecc_double_err,
  output        io_iccm_dma_sb_error,
  output        io_ic_hit_f,
  output        io_ic_access_fault_f,
  output [1:0]  io_ic_access_fault_type_f,
  output        io_ifu_async_error_start,
  output [1:0]  io_ic_fetch_val_f,
  output [31:0] io_ic_data_f,
  input         io_scan_mode
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [95:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [63:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [63:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
`endif // RANDOMIZE_REG_INIT
  wire  rvclkhdr_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_1_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_1_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_1_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_1_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_2_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_2_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_2_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_2_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_3_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_3_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_3_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_3_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_4_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_4_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_4_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_4_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_5_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_5_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_5_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_5_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_6_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_6_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_6_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_6_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_7_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_7_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_7_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_7_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_8_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_8_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_8_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_8_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_9_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_9_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_9_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_9_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_10_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_10_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_10_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_10_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_11_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_11_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_11_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_11_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_12_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_12_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_12_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_12_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_13_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_13_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_13_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_13_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_14_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_14_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_14_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_14_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_15_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_15_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_15_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_15_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_16_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_16_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_16_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_16_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_17_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_17_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_17_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_17_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_18_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_18_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_18_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_18_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_19_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_19_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_19_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_19_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_20_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_20_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_20_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_20_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_21_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_21_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_21_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_21_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_22_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_22_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_22_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_22_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_23_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_23_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_23_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_23_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_24_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_24_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_24_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_24_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_25_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_25_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_25_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_25_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_26_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_26_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_26_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_26_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_27_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_27_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_27_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_27_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_28_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_28_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_28_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_28_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_29_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_29_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_29_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_29_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_30_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_30_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_30_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_30_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_31_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_31_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_31_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_31_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_32_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_32_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_32_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_32_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_33_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_33_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_33_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_33_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_34_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_34_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_34_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_34_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_35_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_35_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_35_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_35_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_36_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_36_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_36_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_36_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_37_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_37_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_37_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_37_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_38_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_38_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_38_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_38_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_39_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_39_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_39_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_39_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_40_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_40_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_40_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_40_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_41_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_41_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_41_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_41_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_42_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_42_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_42_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_42_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_43_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_43_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_43_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_43_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_44_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_44_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_44_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_44_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_45_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_45_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_45_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_45_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_46_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_46_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_46_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_46_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_47_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_47_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_47_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_47_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_48_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_48_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_48_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_48_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_49_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_49_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_49_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_49_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_50_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_50_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_50_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_50_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_51_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_51_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_51_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_51_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_52_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_52_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_52_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_52_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_53_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_53_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_53_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_53_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_54_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_54_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_54_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_54_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_55_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_55_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_55_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_55_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_56_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_56_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_56_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_56_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_57_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_57_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_57_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_57_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_58_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_58_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_58_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_58_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_59_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_59_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_59_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_59_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_60_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_60_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_60_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_60_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_61_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_61_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_61_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_61_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_62_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_62_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_62_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_62_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_63_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_63_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_63_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_63_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_64_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_64_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_64_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_64_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_65_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_65_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_65_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_65_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_66_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_66_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_66_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_66_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_67_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_67_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_67_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_67_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_68_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_68_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_68_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_68_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_69_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_69_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_69_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_69_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_70_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_70_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_70_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_70_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_71_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_71_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_71_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_71_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_72_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_72_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_72_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_72_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_73_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_73_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_73_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_73_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_74_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_74_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_74_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_74_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_75_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_75_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_75_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_75_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_76_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_76_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_76_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_76_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_77_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_77_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_77_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_77_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_78_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_78_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_78_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_78_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_79_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_79_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_79_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_79_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_80_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_80_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_80_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_80_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_81_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_81_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_81_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_81_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_82_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_82_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_82_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_82_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_83_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_83_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_83_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_83_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_84_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_84_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_84_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_84_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_85_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_85_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_85_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_85_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_86_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_86_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_86_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_86_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_87_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_87_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_87_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_87_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_88_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_88_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_88_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_88_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_89_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_89_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_89_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_89_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_90_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_90_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_90_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_90_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_91_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_91_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_91_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_91_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_92_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_92_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_92_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_92_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_93_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_93_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_93_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_93_io_scan_mode; // @[lib.scala 343:22]
  reg  flush_final_f; // @[ifu_mem_ctl.scala 90:53]
  reg  ifc_fetch_req_f_raw; // @[ifu_mem_ctl.scala 227:61]
  wire  _T_319 = ~io_exu_flush_final; // @[ifu_mem_ctl.scala 228:44]
  wire  ifc_fetch_req_f = ifc_fetch_req_f_raw & _T_319; // @[ifu_mem_ctl.scala 228:42]
  wire  _T = io_ifc_fetch_req_bf_raw | ifc_fetch_req_f; // @[ifu_mem_ctl.scala 91:53]
  reg [2:0] miss_state; // @[Reg.scala 27:20]
  wire  miss_pending = miss_state != 3'h0; // @[ifu_mem_ctl.scala 159:30]
  wire  _T_1 = _T | miss_pending; // @[ifu_mem_ctl.scala 91:71]
  wire  debug_c1_clken = io_ic_debug_rd_en | io_ic_debug_wr_en; // @[ifu_mem_ctl.scala 92:42]
  wire [3:0] ic_fetch_val_int_f = {2'h0,io_ic_fetch_val_f}; // @[Cat.scala 29:58]
  reg [30:0] ifu_fetch_addr_int_f; // @[ifu_mem_ctl.scala 214:63]
  wire [4:0] _GEN_435 = {{1'd0}, ic_fetch_val_int_f}; // @[ifu_mem_ctl.scala 602:53]
  wire [4:0] ic_fetch_val_shift_right = _GEN_435 << ifu_fetch_addr_int_f[0]; // @[ifu_mem_ctl.scala 602:53]
  wire  _T_3129 = |ic_fetch_val_shift_right[3:2]; // @[ifu_mem_ctl.scala 605:91]
  wire  _T_3131 = _T_3129 & _T_319; // @[ifu_mem_ctl.scala 605:95]
  reg  ifc_iccm_access_f; // @[ifu_mem_ctl.scala 229:60]
  wire  fetch_req_iccm_f = ifc_fetch_req_f & ifc_iccm_access_f; // @[ifu_mem_ctl.scala 181:46]
  wire  _T_3132 = _T_3131 & fetch_req_iccm_f; // @[ifu_mem_ctl.scala 605:117]
  reg  iccm_dma_rvalid_in; // @[ifu_mem_ctl.scala 591:59]
  wire  _T_3133 = _T_3132 | iccm_dma_rvalid_in; // @[ifu_mem_ctl.scala 605:134]
  wire  _T_3134 = ~io_dec_mem_ctrl_dec_tlu_core_ecc_disable; // @[ifu_mem_ctl.scala 605:158]
  wire  _T_3135 = _T_3133 & _T_3134; // @[ifu_mem_ctl.scala 605:156]
  wire  _T_3121 = |ic_fetch_val_shift_right[1:0]; // @[ifu_mem_ctl.scala 605:91]
  wire  _T_3123 = _T_3121 & _T_319; // @[ifu_mem_ctl.scala 605:95]
  wire  _T_3124 = _T_3123 & fetch_req_iccm_f; // @[ifu_mem_ctl.scala 605:117]
  wire  _T_3125 = _T_3124 | iccm_dma_rvalid_in; // @[ifu_mem_ctl.scala 605:134]
  wire  _T_3127 = _T_3125 & _T_3134; // @[ifu_mem_ctl.scala 605:156]
  wire [1:0] iccm_ecc_word_enable = {_T_3135,_T_3127}; // @[Cat.scala 29:58]
  wire  _T_3620 = ^io_iccm_rd_data_ecc[70:39]; // @[lib.scala 193:30]
  wire  _T_3621 = ^io_iccm_rd_data_ecc[77:71]; // @[lib.scala 193:44]
  wire  _T_3622 = _T_3620 ^ _T_3621; // @[lib.scala 193:35]
  wire [5:0] _T_3630 = {io_iccm_rd_data_ecc[70],io_iccm_rd_data_ecc[69],io_iccm_rd_data_ecc[68],io_iccm_rd_data_ecc[67],io_iccm_rd_data_ecc[66],io_iccm_rd_data_ecc[65]}; // @[lib.scala 193:76]
  wire  _T_3631 = ^_T_3630; // @[lib.scala 193:83]
  wire  _T_3632 = io_iccm_rd_data_ecc[76] ^ _T_3631; // @[lib.scala 193:71]
  wire [6:0] _T_3639 = {io_iccm_rd_data_ecc[56],io_iccm_rd_data_ecc[55],io_iccm_rd_data_ecc[54],io_iccm_rd_data_ecc[53],io_iccm_rd_data_ecc[52],io_iccm_rd_data_ecc[51],io_iccm_rd_data_ecc[50]}; // @[lib.scala 193:103]
  wire [14:0] _T_3647 = {io_iccm_rd_data_ecc[64],io_iccm_rd_data_ecc[63],io_iccm_rd_data_ecc[62],io_iccm_rd_data_ecc[61],io_iccm_rd_data_ecc[60],io_iccm_rd_data_ecc[59],io_iccm_rd_data_ecc[58],io_iccm_rd_data_ecc[57],_T_3639}; // @[lib.scala 193:103]
  wire  _T_3648 = ^_T_3647; // @[lib.scala 193:110]
  wire  _T_3649 = io_iccm_rd_data_ecc[75] ^ _T_3648; // @[lib.scala 193:98]
  wire [6:0] _T_3656 = {io_iccm_rd_data_ecc[49],io_iccm_rd_data_ecc[48],io_iccm_rd_data_ecc[47],io_iccm_rd_data_ecc[46],io_iccm_rd_data_ecc[45],io_iccm_rd_data_ecc[44],io_iccm_rd_data_ecc[43]}; // @[lib.scala 193:130]
  wire [14:0] _T_3664 = {io_iccm_rd_data_ecc[64],io_iccm_rd_data_ecc[63],io_iccm_rd_data_ecc[62],io_iccm_rd_data_ecc[61],io_iccm_rd_data_ecc[60],io_iccm_rd_data_ecc[59],io_iccm_rd_data_ecc[58],io_iccm_rd_data_ecc[57],_T_3656}; // @[lib.scala 193:130]
  wire  _T_3665 = ^_T_3664; // @[lib.scala 193:137]
  wire  _T_3666 = io_iccm_rd_data_ecc[74] ^ _T_3665; // @[lib.scala 193:125]
  wire [8:0] _T_3675 = {io_iccm_rd_data_ecc[54],io_iccm_rd_data_ecc[53],io_iccm_rd_data_ecc[49],io_iccm_rd_data_ecc[48],io_iccm_rd_data_ecc[47],io_iccm_rd_data_ecc[46],io_iccm_rd_data_ecc[42],io_iccm_rd_data_ecc[41],io_iccm_rd_data_ecc[40]}; // @[lib.scala 193:157]
  wire [17:0] _T_3684 = {io_iccm_rd_data_ecc[70],io_iccm_rd_data_ecc[69],io_iccm_rd_data_ecc[68],io_iccm_rd_data_ecc[64],io_iccm_rd_data_ecc[63],io_iccm_rd_data_ecc[62],io_iccm_rd_data_ecc[61],io_iccm_rd_data_ecc[56],io_iccm_rd_data_ecc[55],_T_3675}; // @[lib.scala 193:157]
  wire  _T_3685 = ^_T_3684; // @[lib.scala 193:164]
  wire  _T_3686 = io_iccm_rd_data_ecc[73] ^ _T_3685; // @[lib.scala 193:152]
  wire [8:0] _T_3695 = {io_iccm_rd_data_ecc[52],io_iccm_rd_data_ecc[51],io_iccm_rd_data_ecc[49],io_iccm_rd_data_ecc[48],io_iccm_rd_data_ecc[45],io_iccm_rd_data_ecc[44],io_iccm_rd_data_ecc[42],io_iccm_rd_data_ecc[41],io_iccm_rd_data_ecc[39]}; // @[lib.scala 193:184]
  wire [17:0] _T_3704 = {io_iccm_rd_data_ecc[70],io_iccm_rd_data_ecc[67],io_iccm_rd_data_ecc[66],io_iccm_rd_data_ecc[64],io_iccm_rd_data_ecc[63],io_iccm_rd_data_ecc[60],io_iccm_rd_data_ecc[59],io_iccm_rd_data_ecc[56],io_iccm_rd_data_ecc[55],_T_3695}; // @[lib.scala 193:184]
  wire  _T_3705 = ^_T_3704; // @[lib.scala 193:191]
  wire  _T_3706 = io_iccm_rd_data_ecc[72] ^ _T_3705; // @[lib.scala 193:179]
  wire [8:0] _T_3715 = {io_iccm_rd_data_ecc[52],io_iccm_rd_data_ecc[50],io_iccm_rd_data_ecc[49],io_iccm_rd_data_ecc[47],io_iccm_rd_data_ecc[45],io_iccm_rd_data_ecc[43],io_iccm_rd_data_ecc[42],io_iccm_rd_data_ecc[40],io_iccm_rd_data_ecc[39]}; // @[lib.scala 193:211]
  wire [17:0] _T_3724 = {io_iccm_rd_data_ecc[69],io_iccm_rd_data_ecc[67],io_iccm_rd_data_ecc[65],io_iccm_rd_data_ecc[64],io_iccm_rd_data_ecc[62],io_iccm_rd_data_ecc[60],io_iccm_rd_data_ecc[58],io_iccm_rd_data_ecc[56],io_iccm_rd_data_ecc[54],_T_3715}; // @[lib.scala 193:211]
  wire  _T_3725 = ^_T_3724; // @[lib.scala 193:218]
  wire  _T_3726 = io_iccm_rd_data_ecc[71] ^ _T_3725; // @[lib.scala 193:206]
  wire [6:0] _T_3732 = {_T_3622,_T_3632,_T_3649,_T_3666,_T_3686,_T_3706,_T_3726}; // @[Cat.scala 29:58]
  wire  _T_3733 = _T_3732 != 7'h0; // @[lib.scala 194:44]
  wire  _T_3734 = iccm_ecc_word_enable[1] & _T_3733; // @[lib.scala 194:32]
  wire  _T_3736 = _T_3734 & _T_3732[6]; // @[lib.scala 194:53]
  wire  _T_3235 = ^io_iccm_rd_data_ecc[31:0]; // @[lib.scala 193:30]
  wire  _T_3236 = ^io_iccm_rd_data_ecc[38:32]; // @[lib.scala 193:44]
  wire  _T_3237 = _T_3235 ^ _T_3236; // @[lib.scala 193:35]
  wire [5:0] _T_3245 = {io_iccm_rd_data_ecc[31],io_iccm_rd_data_ecc[30],io_iccm_rd_data_ecc[29],io_iccm_rd_data_ecc[28],io_iccm_rd_data_ecc[27],io_iccm_rd_data_ecc[26]}; // @[lib.scala 193:76]
  wire  _T_3246 = ^_T_3245; // @[lib.scala 193:83]
  wire  _T_3247 = io_iccm_rd_data_ecc[37] ^ _T_3246; // @[lib.scala 193:71]
  wire [6:0] _T_3254 = {io_iccm_rd_data_ecc[17],io_iccm_rd_data_ecc[16],io_iccm_rd_data_ecc[15],io_iccm_rd_data_ecc[14],io_iccm_rd_data_ecc[13],io_iccm_rd_data_ecc[12],io_iccm_rd_data_ecc[11]}; // @[lib.scala 193:103]
  wire [14:0] _T_3262 = {io_iccm_rd_data_ecc[25],io_iccm_rd_data_ecc[24],io_iccm_rd_data_ecc[23],io_iccm_rd_data_ecc[22],io_iccm_rd_data_ecc[21],io_iccm_rd_data_ecc[20],io_iccm_rd_data_ecc[19],io_iccm_rd_data_ecc[18],_T_3254}; // @[lib.scala 193:103]
  wire  _T_3263 = ^_T_3262; // @[lib.scala 193:110]
  wire  _T_3264 = io_iccm_rd_data_ecc[36] ^ _T_3263; // @[lib.scala 193:98]
  wire [6:0] _T_3271 = {io_iccm_rd_data_ecc[10],io_iccm_rd_data_ecc[9],io_iccm_rd_data_ecc[8],io_iccm_rd_data_ecc[7],io_iccm_rd_data_ecc[6],io_iccm_rd_data_ecc[5],io_iccm_rd_data_ecc[4]}; // @[lib.scala 193:130]
  wire [14:0] _T_3279 = {io_iccm_rd_data_ecc[25],io_iccm_rd_data_ecc[24],io_iccm_rd_data_ecc[23],io_iccm_rd_data_ecc[22],io_iccm_rd_data_ecc[21],io_iccm_rd_data_ecc[20],io_iccm_rd_data_ecc[19],io_iccm_rd_data_ecc[18],_T_3271}; // @[lib.scala 193:130]
  wire  _T_3280 = ^_T_3279; // @[lib.scala 193:137]
  wire  _T_3281 = io_iccm_rd_data_ecc[35] ^ _T_3280; // @[lib.scala 193:125]
  wire [8:0] _T_3290 = {io_iccm_rd_data_ecc[15],io_iccm_rd_data_ecc[14],io_iccm_rd_data_ecc[10],io_iccm_rd_data_ecc[9],io_iccm_rd_data_ecc[8],io_iccm_rd_data_ecc[7],io_iccm_rd_data_ecc[3],io_iccm_rd_data_ecc[2],io_iccm_rd_data_ecc[1]}; // @[lib.scala 193:157]
  wire [17:0] _T_3299 = {io_iccm_rd_data_ecc[31],io_iccm_rd_data_ecc[30],io_iccm_rd_data_ecc[29],io_iccm_rd_data_ecc[25],io_iccm_rd_data_ecc[24],io_iccm_rd_data_ecc[23],io_iccm_rd_data_ecc[22],io_iccm_rd_data_ecc[17],io_iccm_rd_data_ecc[16],_T_3290}; // @[lib.scala 193:157]
  wire  _T_3300 = ^_T_3299; // @[lib.scala 193:164]
  wire  _T_3301 = io_iccm_rd_data_ecc[34] ^ _T_3300; // @[lib.scala 193:152]
  wire [8:0] _T_3310 = {io_iccm_rd_data_ecc[13],io_iccm_rd_data_ecc[12],io_iccm_rd_data_ecc[10],io_iccm_rd_data_ecc[9],io_iccm_rd_data_ecc[6],io_iccm_rd_data_ecc[5],io_iccm_rd_data_ecc[3],io_iccm_rd_data_ecc[2],io_iccm_rd_data_ecc[0]}; // @[lib.scala 193:184]
  wire [17:0] _T_3319 = {io_iccm_rd_data_ecc[31],io_iccm_rd_data_ecc[28],io_iccm_rd_data_ecc[27],io_iccm_rd_data_ecc[25],io_iccm_rd_data_ecc[24],io_iccm_rd_data_ecc[21],io_iccm_rd_data_ecc[20],io_iccm_rd_data_ecc[17],io_iccm_rd_data_ecc[16],_T_3310}; // @[lib.scala 193:184]
  wire  _T_3320 = ^_T_3319; // @[lib.scala 193:191]
  wire  _T_3321 = io_iccm_rd_data_ecc[33] ^ _T_3320; // @[lib.scala 193:179]
  wire [8:0] _T_3330 = {io_iccm_rd_data_ecc[13],io_iccm_rd_data_ecc[11],io_iccm_rd_data_ecc[10],io_iccm_rd_data_ecc[8],io_iccm_rd_data_ecc[6],io_iccm_rd_data_ecc[4],io_iccm_rd_data_ecc[3],io_iccm_rd_data_ecc[1],io_iccm_rd_data_ecc[0]}; // @[lib.scala 193:211]
  wire [17:0] _T_3339 = {io_iccm_rd_data_ecc[30],io_iccm_rd_data_ecc[28],io_iccm_rd_data_ecc[26],io_iccm_rd_data_ecc[25],io_iccm_rd_data_ecc[23],io_iccm_rd_data_ecc[21],io_iccm_rd_data_ecc[19],io_iccm_rd_data_ecc[17],io_iccm_rd_data_ecc[15],_T_3330}; // @[lib.scala 193:211]
  wire  _T_3340 = ^_T_3339; // @[lib.scala 193:218]
  wire  _T_3341 = io_iccm_rd_data_ecc[32] ^ _T_3340; // @[lib.scala 193:206]
  wire [6:0] _T_3347 = {_T_3237,_T_3247,_T_3264,_T_3281,_T_3301,_T_3321,_T_3341}; // @[Cat.scala 29:58]
  wire  _T_3348 = _T_3347 != 7'h0; // @[lib.scala 194:44]
  wire  _T_3349 = iccm_ecc_word_enable[0] & _T_3348; // @[lib.scala 194:32]
  wire  _T_3351 = _T_3349 & _T_3347[6]; // @[lib.scala 194:53]
  wire [1:0] iccm_single_ecc_error = {_T_3736,_T_3351}; // @[Cat.scala 29:58]
  wire  _T_3 = |iccm_single_ecc_error; // @[ifu_mem_ctl.scala 95:52]
  reg  dma_iccm_req_f; // @[ifu_mem_ctl.scala 568:51]
  wire  _T_6 = io_dec_mem_ctrl_ifu_iccm_rd_ecc_single_err | io_dec_mem_ctrl_ifu_ic_error_start; // @[ifu_mem_ctl.scala 96:74]
  reg [2:0] perr_state; // @[Reg.scala 27:20]
  wire  _T_7 = perr_state == 3'h4; // @[ifu_mem_ctl.scala 97:54]
  wire  iccm_correct_ecc = perr_state == 3'h3; // @[ifu_mem_ctl.scala 392:34]
  wire  _T_8 = iccm_correct_ecc | _T_7; // @[ifu_mem_ctl.scala 97:40]
  reg [1:0] err_stop_state; // @[Reg.scala 27:20]
  wire  _T_9 = err_stop_state == 2'h3; // @[ifu_mem_ctl.scala 97:90]
  wire  _T_10 = _T_8 | _T_9; // @[ifu_mem_ctl.scala 97:72]
  wire  _T_2526 = 2'h0 == err_stop_state; // @[Conditional.scala 37:30]
  wire  _T_2531 = 2'h1 == err_stop_state; // @[Conditional.scala 37:30]
  wire  _T_2551 = io_ifu_fetch_val == 2'h3; // @[ifu_mem_ctl.scala 441:48]
  wire  two_byte_instr = io_ic_data_f[1:0] != 2'h3; // @[ifu_mem_ctl.scala 306:42]
  wire  _T_2553 = io_ifu_fetch_val[0] & two_byte_instr; // @[ifu_mem_ctl.scala 441:79]
  wire  _T_2554 = _T_2551 | _T_2553; // @[ifu_mem_ctl.scala 441:56]
  wire  _T_2555 = io_exu_flush_final | io_dec_mem_ctrl_dec_tlu_i0_commit_cmt; // @[ifu_mem_ctl.scala 441:122]
  wire  _T_2556 = ~_T_2555; // @[ifu_mem_ctl.scala 441:101]
  wire  _T_2557 = _T_2554 & _T_2556; // @[ifu_mem_ctl.scala 441:99]
  wire  _T_2558 = 2'h2 == err_stop_state; // @[Conditional.scala 37:30]
  wire  _T_2572 = io_ifu_fetch_val[0] & _T_319; // @[ifu_mem_ctl.scala 448:45]
  wire  _T_2573 = ~io_dec_mem_ctrl_dec_tlu_i0_commit_cmt; // @[ifu_mem_ctl.scala 448:69]
  wire  _T_2574 = _T_2572 & _T_2573; // @[ifu_mem_ctl.scala 448:67]
  wire  _T_2575 = 2'h3 == err_stop_state; // @[Conditional.scala 37:30]
  wire  _GEN_37 = _T_2558 ? _T_2574 : _T_2575; // @[Conditional.scala 39:67]
  wire  _GEN_41 = _T_2531 ? _T_2557 : _GEN_37; // @[Conditional.scala 39:67]
  wire  err_stop_fetch = _T_2526 ? 1'h0 : _GEN_41; // @[Conditional.scala 40:58]
  wire  _T_11 = _T_10 | err_stop_fetch; // @[ifu_mem_ctl.scala 97:112]
  wire  _T_227 = |io_ic_rd_hit; // @[ifu_mem_ctl.scala 189:37]
  wire  _T_228 = ~_T_227; // @[ifu_mem_ctl.scala 189:23]
  reg  reset_all_tags; // @[ifu_mem_ctl.scala 637:53]
  wire  _T_229 = _T_228 | reset_all_tags; // @[ifu_mem_ctl.scala 189:41]
  wire  _T_207 = ~ifc_iccm_access_f; // @[ifu_mem_ctl.scala 180:48]
  wire  _T_208 = ifc_fetch_req_f & _T_207; // @[ifu_mem_ctl.scala 180:46]
  reg  ifc_region_acc_fault_final_f; // @[ifu_mem_ctl.scala 231:71]
  wire  _T_209 = ~ifc_region_acc_fault_final_f; // @[ifu_mem_ctl.scala 180:69]
  wire  fetch_req_icache_f = _T_208 & _T_209; // @[ifu_mem_ctl.scala 180:67]
  wire  _T_230 = _T_229 & fetch_req_icache_f; // @[ifu_mem_ctl.scala 189:59]
  wire  _T_231 = ~miss_pending; // @[ifu_mem_ctl.scala 189:82]
  wire  _T_232 = _T_230 & _T_231; // @[ifu_mem_ctl.scala 189:80]
  wire  ic_act_miss_f = _T_232 & _T_209; // @[ifu_mem_ctl.scala 189:114]
  reg  uncacheable_miss_ff; // @[ifu_mem_ctl.scala 216:62]
  wire  _T_2623 = ~io_dec_mem_ctrl_dec_tlu_force_halt; // @[ifu_mem_ctl.scala 528:72]
  wire  _T_17 = ~uncacheable_miss_ff; // @[ifu_mem_ctl.scala 100:5]
  wire  _T_24 = 3'h0 == miss_state; // @[Conditional.scala 37:30]
  wire  _T_26 = ic_act_miss_f & _T_319; // @[ifu_mem_ctl.scala 106:43]
  wire [2:0] _T_28 = _T_26 ? 3'h1 : 3'h2; // @[ifu_mem_ctl.scala 106:27]
  wire  _T_31 = 3'h1 == miss_state; // @[Conditional.scala 37:30]
  wire [4:0] byp_fetch_index = ifu_fetch_addr_int_f[4:0]; // @[ifu_mem_ctl.scala 343:45]
  wire  _T_2155 = byp_fetch_index[4:2] == 3'h0; // @[ifu_mem_ctl.scala 364:127]
  reg [7:0] ic_miss_buff_data_valid; // @[ifu_mem_ctl.scala 320:60]
  wire  _T_2186 = _T_2155 & ic_miss_buff_data_valid[0]; // @[Mux.scala 27:72]
  wire  _T_2159 = byp_fetch_index[4:2] == 3'h1; // @[ifu_mem_ctl.scala 364:127]
  wire  _T_2187 = _T_2159 & ic_miss_buff_data_valid[1]; // @[Mux.scala 27:72]
  wire  _T_2194 = _T_2186 | _T_2187; // @[Mux.scala 27:72]
  wire  _T_2163 = byp_fetch_index[4:2] == 3'h2; // @[ifu_mem_ctl.scala 364:127]
  wire  _T_2188 = _T_2163 & ic_miss_buff_data_valid[2]; // @[Mux.scala 27:72]
  wire  _T_2195 = _T_2194 | _T_2188; // @[Mux.scala 27:72]
  wire  _T_2167 = byp_fetch_index[4:2] == 3'h3; // @[ifu_mem_ctl.scala 364:127]
  wire  _T_2189 = _T_2167 & ic_miss_buff_data_valid[3]; // @[Mux.scala 27:72]
  wire  _T_2196 = _T_2195 | _T_2189; // @[Mux.scala 27:72]
  wire  _T_2171 = byp_fetch_index[4:2] == 3'h4; // @[ifu_mem_ctl.scala 364:127]
  wire  _T_2190 = _T_2171 & ic_miss_buff_data_valid[4]; // @[Mux.scala 27:72]
  wire  _T_2197 = _T_2196 | _T_2190; // @[Mux.scala 27:72]
  wire  _T_2175 = byp_fetch_index[4:2] == 3'h5; // @[ifu_mem_ctl.scala 364:127]
  wire  _T_2191 = _T_2175 & ic_miss_buff_data_valid[5]; // @[Mux.scala 27:72]
  wire  _T_2198 = _T_2197 | _T_2191; // @[Mux.scala 27:72]
  wire  _T_2179 = byp_fetch_index[4:2] == 3'h6; // @[ifu_mem_ctl.scala 364:127]
  wire  _T_2192 = _T_2179 & ic_miss_buff_data_valid[6]; // @[Mux.scala 27:72]
  wire  _T_2199 = _T_2198 | _T_2192; // @[Mux.scala 27:72]
  wire  _T_2183 = byp_fetch_index[4:2] == 3'h7; // @[ifu_mem_ctl.scala 364:127]
  wire  _T_2193 = _T_2183 & ic_miss_buff_data_valid[7]; // @[Mux.scala 27:72]
  wire  ic_miss_buff_data_valid_bypass_index = _T_2199 | _T_2193; // @[Mux.scala 27:72]
  wire  _T_2241 = ~byp_fetch_index[1]; // @[ifu_mem_ctl.scala 366:69]
  wire  _T_2242 = ic_miss_buff_data_valid_bypass_index & _T_2241; // @[ifu_mem_ctl.scala 366:67]
  wire  _T_2244 = ~byp_fetch_index[0]; // @[ifu_mem_ctl.scala 366:91]
  wire  _T_2245 = _T_2242 & _T_2244; // @[ifu_mem_ctl.scala 366:89]
  wire  _T_2250 = _T_2242 & byp_fetch_index[0]; // @[ifu_mem_ctl.scala 367:65]
  wire  _T_2251 = _T_2245 | _T_2250; // @[ifu_mem_ctl.scala 366:112]
  wire  _T_2253 = ic_miss_buff_data_valid_bypass_index & byp_fetch_index[1]; // @[ifu_mem_ctl.scala 368:43]
  wire  _T_2256 = _T_2253 & _T_2244; // @[ifu_mem_ctl.scala 368:65]
  wire  _T_2257 = _T_2251 | _T_2256; // @[ifu_mem_ctl.scala 367:88]
  wire  _T_2261 = _T_2253 & byp_fetch_index[0]; // @[ifu_mem_ctl.scala 369:65]
  wire [2:0] byp_fetch_index_inc = ifu_fetch_addr_int_f[4:2] + 3'h1; // @[ifu_mem_ctl.scala 346:75]
  wire  _T_2201 = byp_fetch_index_inc == 3'h0; // @[ifu_mem_ctl.scala 365:110]
  wire  _T_2225 = _T_2201 & ic_miss_buff_data_valid[0]; // @[Mux.scala 27:72]
  wire  _T_2204 = byp_fetch_index_inc == 3'h1; // @[ifu_mem_ctl.scala 365:110]
  wire  _T_2226 = _T_2204 & ic_miss_buff_data_valid[1]; // @[Mux.scala 27:72]
  wire  _T_2233 = _T_2225 | _T_2226; // @[Mux.scala 27:72]
  wire  _T_2207 = byp_fetch_index_inc == 3'h2; // @[ifu_mem_ctl.scala 365:110]
  wire  _T_2227 = _T_2207 & ic_miss_buff_data_valid[2]; // @[Mux.scala 27:72]
  wire  _T_2234 = _T_2233 | _T_2227; // @[Mux.scala 27:72]
  wire  _T_2210 = byp_fetch_index_inc == 3'h3; // @[ifu_mem_ctl.scala 365:110]
  wire  _T_2228 = _T_2210 & ic_miss_buff_data_valid[3]; // @[Mux.scala 27:72]
  wire  _T_2235 = _T_2234 | _T_2228; // @[Mux.scala 27:72]
  wire  _T_2213 = byp_fetch_index_inc == 3'h4; // @[ifu_mem_ctl.scala 365:110]
  wire  _T_2229 = _T_2213 & ic_miss_buff_data_valid[4]; // @[Mux.scala 27:72]
  wire  _T_2236 = _T_2235 | _T_2229; // @[Mux.scala 27:72]
  wire  _T_2216 = byp_fetch_index_inc == 3'h5; // @[ifu_mem_ctl.scala 365:110]
  wire  _T_2230 = _T_2216 & ic_miss_buff_data_valid[5]; // @[Mux.scala 27:72]
  wire  _T_2237 = _T_2236 | _T_2230; // @[Mux.scala 27:72]
  wire  _T_2219 = byp_fetch_index_inc == 3'h6; // @[ifu_mem_ctl.scala 365:110]
  wire  _T_2231 = _T_2219 & ic_miss_buff_data_valid[6]; // @[Mux.scala 27:72]
  wire  _T_2238 = _T_2237 | _T_2231; // @[Mux.scala 27:72]
  wire  _T_2222 = byp_fetch_index_inc == 3'h7; // @[ifu_mem_ctl.scala 365:110]
  wire  _T_2232 = _T_2222 & ic_miss_buff_data_valid[7]; // @[Mux.scala 27:72]
  wire  ic_miss_buff_data_valid_inc_bypass_index = _T_2238 | _T_2232; // @[Mux.scala 27:72]
  wire  _T_2262 = _T_2261 & ic_miss_buff_data_valid_inc_bypass_index; // @[ifu_mem_ctl.scala 369:87]
  wire  _T_2263 = _T_2257 | _T_2262; // @[ifu_mem_ctl.scala 368:88]
  wire  _T_2267 = ic_miss_buff_data_valid_bypass_index & _T_2183; // @[ifu_mem_ctl.scala 370:43]
  wire  miss_buff_hit_unq_f = _T_2263 | _T_2267; // @[ifu_mem_ctl.scala 369:131]
  wire  _T_2283 = miss_state == 3'h4; // @[ifu_mem_ctl.scala 375:55]
  wire  _T_2284 = miss_state == 3'h1; // @[ifu_mem_ctl.scala 375:87]
  wire  _T_2285 = _T_2283 | _T_2284; // @[ifu_mem_ctl.scala 375:74]
  wire  crit_byp_hit_f = miss_buff_hit_unq_f & _T_2285; // @[ifu_mem_ctl.scala 375:41]
  wire  _T_2268 = miss_state == 3'h6; // @[ifu_mem_ctl.scala 372:30]
  reg [30:0] imb_ff; // @[ifu_mem_ctl.scala 217:49]
  wire  miss_wrap_f = imb_ff[5] != ifu_fetch_addr_int_f[5]; // @[ifu_mem_ctl.scala 363:51]
  wire  _T_2269 = ~miss_wrap_f; // @[ifu_mem_ctl.scala 372:68]
  wire  _T_2270 = miss_buff_hit_unq_f & _T_2269; // @[ifu_mem_ctl.scala 372:66]
  wire  stream_hit_f = _T_2268 & _T_2270; // @[ifu_mem_ctl.scala 372:43]
  wire  _T_215 = crit_byp_hit_f | stream_hit_f; // @[ifu_mem_ctl.scala 184:35]
  wire  _T_216 = _T_215 & fetch_req_icache_f; // @[ifu_mem_ctl.scala 184:52]
  wire  ic_byp_hit_f = _T_216 & miss_pending; // @[ifu_mem_ctl.scala 184:73]
  wire  _T_40 = ic_byp_hit_f & uncacheable_miss_ff; // @[ifu_mem_ctl.scala 111:53]
  wire  _T_54 = ic_byp_hit_f & _T_319; // @[ifu_mem_ctl.scala 114:33]
  wire  ifu_bp_hit_taken_q_f = io_ifu_bp_hit_taken_f & io_ic_hit_f; // @[ifu_mem_ctl.scala 102:52]
  wire  _T_58 = ~ifu_bp_hit_taken_q_f; // @[ifu_mem_ctl.scala 114:91]
  wire  _T_59 = _T_54 & _T_58; // @[ifu_mem_ctl.scala 114:89]
  wire  _T_61 = _T_59 & _T_17; // @[ifu_mem_ctl.scala 114:113]
  wire  _T_81 = io_exu_flush_final | ifu_bp_hit_taken_q_f; // @[ifu_mem_ctl.scala 117:44]
  wire [2:0] _T_86 = _T_81 ? 3'h2 : 3'h0; // @[ifu_mem_ctl.scala 117:22]
  wire [2:0] _T_89 = _T_61 ? 3'h6 : _T_86; // @[ifu_mem_ctl.scala 114:18]
  wire [2:0] _T_92 = _T_40 ? 3'h3 : _T_89; // @[ifu_mem_ctl.scala 111:12]
  wire [2:0] _T_93 = io_dec_mem_ctrl_dec_tlu_force_halt ? 3'h0 : _T_92; // @[ifu_mem_ctl.scala 110:27]
  wire  _T_102 = 3'h4 == miss_state; // @[Conditional.scala 37:30]
  wire  _T_106 = 3'h6 == miss_state; // @[Conditional.scala 37:30]
  wire  _T_2280 = byp_fetch_index[4:1] == 4'hf; // @[ifu_mem_ctl.scala 374:60]
  wire  _T_2281 = _T_2280 & ifc_fetch_req_f; // @[ifu_mem_ctl.scala 374:94]
  wire  stream_eol_f = _T_2281 & stream_hit_f; // @[ifu_mem_ctl.scala 374:112]
  wire  _T_108 = _T_81 | stream_eol_f; // @[ifu_mem_ctl.scala 125:72]
  wire  _T_113 = _T_108 & _T_2623; // @[ifu_mem_ctl.scala 125:122]
  wire [2:0] _T_115 = _T_113 ? 3'h2 : 3'h0; // @[ifu_mem_ctl.scala 125:27]
  wire  _T_121 = 3'h3 == miss_state; // @[Conditional.scala 37:30]
  wire  _T_126 = io_exu_flush_final & _T_2623; // @[ifu_mem_ctl.scala 129:82]
  wire [2:0] _T_128 = _T_126 ? 3'h2 : 3'h0; // @[ifu_mem_ctl.scala 129:27]
  wire  _T_132 = 3'h2 == miss_state; // @[Conditional.scala 37:30]
  wire  _T_236 = io_ic_rd_hit == 2'h0; // @[ifu_mem_ctl.scala 190:28]
  wire  _T_237 = _T_236 | reset_all_tags; // @[ifu_mem_ctl.scala 190:42]
  wire  _T_238 = _T_237 & fetch_req_icache_f; // @[ifu_mem_ctl.scala 190:60]
  wire  _T_239 = miss_state == 3'h2; // @[ifu_mem_ctl.scala 190:94]
  wire  _T_240 = _T_238 & _T_239; // @[ifu_mem_ctl.scala 190:81]
  wire  _T_243 = imb_ff[30:5] != ifu_fetch_addr_int_f[30:5]; // @[ifu_mem_ctl.scala 191:39]
  wire  _T_244 = _T_240 & _T_243; // @[ifu_mem_ctl.scala 190:111]
  wire  _T_246 = _T_244 & _T_17; // @[ifu_mem_ctl.scala 191:91]
  reg  sel_mb_addr_ff; // @[ifu_mem_ctl.scala 245:51]
  wire  _T_247 = ~sel_mb_addr_ff; // @[ifu_mem_ctl.scala 191:116]
  wire  _T_248 = _T_246 & _T_247; // @[ifu_mem_ctl.scala 191:114]
  wire  ic_miss_under_miss_f = _T_248 & _T_209; // @[ifu_mem_ctl.scala 191:132]
  wire  _T_137 = ic_miss_under_miss_f & _T_2623; // @[ifu_mem_ctl.scala 133:84]
  wire  _T_256 = _T_230 & _T_239; // @[ifu_mem_ctl.scala 192:85]
  wire  _T_259 = imb_ff[30:5] == ifu_fetch_addr_int_f[30:5]; // @[ifu_mem_ctl.scala 193:39]
  wire  _T_260 = _T_259 | uncacheable_miss_ff; // @[ifu_mem_ctl.scala 193:91]
  wire  ic_ignore_2nd_miss_f = _T_256 & _T_260; // @[ifu_mem_ctl.scala 192:117]
  wire  _T_143 = ic_ignore_2nd_miss_f & _T_2623; // @[ifu_mem_ctl.scala 134:69]
  wire [2:0] _T_145 = _T_143 ? 3'h7 : 3'h0; // @[ifu_mem_ctl.scala 134:12]
  wire [2:0] _T_146 = _T_137 ? 3'h5 : _T_145; // @[ifu_mem_ctl.scala 133:27]
  wire  _T_151 = 3'h5 == miss_state; // @[Conditional.scala 37:30]
  wire [2:0] _T_155 = io_exu_flush_final ? 3'h2 : 3'h1; // @[ifu_mem_ctl.scala 138:75]
  wire [2:0] _T_156 = io_dec_mem_ctrl_dec_tlu_force_halt ? 3'h0 : _T_155; // @[ifu_mem_ctl.scala 138:27]
  wire  _T_160 = 3'h7 == miss_state; // @[Conditional.scala 37:30]
  wire [2:0] _T_164 = io_exu_flush_final ? 3'h2 : 3'h0; // @[ifu_mem_ctl.scala 143:75]
  wire [2:0] _T_165 = io_dec_mem_ctrl_dec_tlu_force_halt ? 3'h0 : _T_164; // @[ifu_mem_ctl.scala 143:27]
  wire [2:0] _GEN_0 = _T_160 ? _T_165 : 3'h0; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_2 = _T_151 ? _T_156 : _GEN_0; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_4 = _T_132 ? _T_146 : _GEN_2; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_6 = _T_121 ? _T_128 : _GEN_4; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_8 = _T_106 ? _T_115 : _GEN_6; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_10 = _T_102 ? 3'h0 : _GEN_8; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_12 = _T_31 ? _T_93 : _GEN_10; // @[Conditional.scala 39:67]
  wire [2:0] miss_nxtstate = _T_24 ? _T_28 : _GEN_12; // @[Conditional.scala 40:58]
  wire  _T_30 = ic_act_miss_f & _T_2623; // @[ifu_mem_ctl.scala 107:38]
  wire  _T_94 = io_dec_mem_ctrl_dec_tlu_force_halt | io_exu_flush_final; // @[ifu_mem_ctl.scala 118:59]
  wire  _T_95 = _T_94 | ic_byp_hit_f; // @[ifu_mem_ctl.scala 118:80]
  wire  _T_96 = _T_95 | ifu_bp_hit_taken_q_f; // @[ifu_mem_ctl.scala 118:95]
  wire  _T_103 = io_exu_flush_final | flush_final_f; // @[ifu_mem_ctl.scala 122:43]
  wire  _T_104 = _T_103 | ic_byp_hit_f; // @[ifu_mem_ctl.scala 122:59]
  wire  _T_105 = _T_104 | io_dec_mem_ctrl_dec_tlu_force_halt; // @[ifu_mem_ctl.scala 122:74]
  wire  _T_120 = _T_108 | io_dec_mem_ctrl_dec_tlu_force_halt; // @[ifu_mem_ctl.scala 126:118]
  wire  _T_131 = io_exu_flush_final | io_dec_mem_ctrl_dec_tlu_force_halt; // @[ifu_mem_ctl.scala 130:76]
  wire  _T_149 = ic_miss_under_miss_f | ic_ignore_2nd_miss_f; // @[ifu_mem_ctl.scala 135:78]
  wire  _T_150 = _T_149 | io_dec_mem_ctrl_dec_tlu_force_halt; // @[ifu_mem_ctl.scala 135:101]
  wire  _GEN_1 = _T_160 & _T_131; // @[Conditional.scala 39:67]
  wire  _GEN_3 = _T_151 ? _T_131 : _GEN_1; // @[Conditional.scala 39:67]
  wire  _GEN_5 = _T_132 ? _T_150 : _GEN_3; // @[Conditional.scala 39:67]
  wire  _GEN_7 = _T_121 ? _T_131 : _GEN_5; // @[Conditional.scala 39:67]
  wire  _GEN_9 = _T_106 ? _T_120 : _GEN_7; // @[Conditional.scala 39:67]
  wire  _GEN_11 = _T_102 ? _T_105 : _GEN_9; // @[Conditional.scala 39:67]
  wire  _GEN_13 = _T_31 ? _T_96 : _GEN_11; // @[Conditional.scala 39:67]
  wire  miss_state_en = _T_24 ? _T_30 : _GEN_13; // @[Conditional.scala 40:58]
  wire  _T_174 = ~flush_final_f; // @[ifu_mem_ctl.scala 160:95]
  wire  _T_175 = _T_2283 & _T_174; // @[ifu_mem_ctl.scala 160:93]
  wire  crit_wd_byp_ok_ff = _T_2284 | _T_175; // @[ifu_mem_ctl.scala 160:58]
  wire  _T_180 = _T_2283 & io_exu_flush_final; // @[ifu_mem_ctl.scala 161:106]
  wire  _T_181 = ~_T_180; // @[ifu_mem_ctl.scala 161:72]
  wire  _T_182 = miss_pending & _T_181; // @[ifu_mem_ctl.scala 161:70]
  wire  _T_184 = _T_2283 & crit_byp_hit_f; // @[ifu_mem_ctl.scala 162:57]
  wire  _T_185 = ~_T_184; // @[ifu_mem_ctl.scala 162:23]
  wire  _T_186 = _T_182 & _T_185; // @[ifu_mem_ctl.scala 161:128]
  wire  _T_187 = _T_186 | ic_act_miss_f; // @[ifu_mem_ctl.scala 162:77]
  wire  _T_188 = miss_nxtstate == 3'h4; // @[ifu_mem_ctl.scala 163:36]
  wire  _T_189 = miss_pending & _T_188; // @[ifu_mem_ctl.scala 163:19]
  wire  sel_hold_imb = _T_187 | _T_189; // @[ifu_mem_ctl.scala 162:93]
  reg [6:0] ifu_ic_rw_int_addr_ff; // @[ifu_mem_ctl.scala 669:14]
  wire  _T_4671 = ifu_ic_rw_int_addr_ff == 7'h0; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_0; // @[Reg.scala 27:20]
  wire  _T_4799 = _T_4671 & way_status_out_0; // @[Mux.scala 27:72]
  wire  _T_4672 = ifu_ic_rw_int_addr_ff == 7'h1; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_1; // @[Reg.scala 27:20]
  wire  _T_4800 = _T_4672 & way_status_out_1; // @[Mux.scala 27:72]
  wire  _T_4927 = _T_4799 | _T_4800; // @[Mux.scala 27:72]
  wire  _T_4673 = ifu_ic_rw_int_addr_ff == 7'h2; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_2; // @[Reg.scala 27:20]
  wire  _T_4801 = _T_4673 & way_status_out_2; // @[Mux.scala 27:72]
  wire  _T_4928 = _T_4927 | _T_4801; // @[Mux.scala 27:72]
  wire  _T_4674 = ifu_ic_rw_int_addr_ff == 7'h3; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_3; // @[Reg.scala 27:20]
  wire  _T_4802 = _T_4674 & way_status_out_3; // @[Mux.scala 27:72]
  wire  _T_4929 = _T_4928 | _T_4802; // @[Mux.scala 27:72]
  wire  _T_4675 = ifu_ic_rw_int_addr_ff == 7'h4; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_4; // @[Reg.scala 27:20]
  wire  _T_4803 = _T_4675 & way_status_out_4; // @[Mux.scala 27:72]
  wire  _T_4930 = _T_4929 | _T_4803; // @[Mux.scala 27:72]
  wire  _T_4676 = ifu_ic_rw_int_addr_ff == 7'h5; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_5; // @[Reg.scala 27:20]
  wire  _T_4804 = _T_4676 & way_status_out_5; // @[Mux.scala 27:72]
  wire  _T_4931 = _T_4930 | _T_4804; // @[Mux.scala 27:72]
  wire  _T_4677 = ifu_ic_rw_int_addr_ff == 7'h6; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_6; // @[Reg.scala 27:20]
  wire  _T_4805 = _T_4677 & way_status_out_6; // @[Mux.scala 27:72]
  wire  _T_4932 = _T_4931 | _T_4805; // @[Mux.scala 27:72]
  wire  _T_4678 = ifu_ic_rw_int_addr_ff == 7'h7; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_7; // @[Reg.scala 27:20]
  wire  _T_4806 = _T_4678 & way_status_out_7; // @[Mux.scala 27:72]
  wire  _T_4933 = _T_4932 | _T_4806; // @[Mux.scala 27:72]
  wire  _T_4679 = ifu_ic_rw_int_addr_ff == 7'h8; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_8; // @[Reg.scala 27:20]
  wire  _T_4807 = _T_4679 & way_status_out_8; // @[Mux.scala 27:72]
  wire  _T_4934 = _T_4933 | _T_4807; // @[Mux.scala 27:72]
  wire  _T_4680 = ifu_ic_rw_int_addr_ff == 7'h9; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_9; // @[Reg.scala 27:20]
  wire  _T_4808 = _T_4680 & way_status_out_9; // @[Mux.scala 27:72]
  wire  _T_4935 = _T_4934 | _T_4808; // @[Mux.scala 27:72]
  wire  _T_4681 = ifu_ic_rw_int_addr_ff == 7'ha; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_10; // @[Reg.scala 27:20]
  wire  _T_4809 = _T_4681 & way_status_out_10; // @[Mux.scala 27:72]
  wire  _T_4936 = _T_4935 | _T_4809; // @[Mux.scala 27:72]
  wire  _T_4682 = ifu_ic_rw_int_addr_ff == 7'hb; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_11; // @[Reg.scala 27:20]
  wire  _T_4810 = _T_4682 & way_status_out_11; // @[Mux.scala 27:72]
  wire  _T_4937 = _T_4936 | _T_4810; // @[Mux.scala 27:72]
  wire  _T_4683 = ifu_ic_rw_int_addr_ff == 7'hc; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_12; // @[Reg.scala 27:20]
  wire  _T_4811 = _T_4683 & way_status_out_12; // @[Mux.scala 27:72]
  wire  _T_4938 = _T_4937 | _T_4811; // @[Mux.scala 27:72]
  wire  _T_4684 = ifu_ic_rw_int_addr_ff == 7'hd; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_13; // @[Reg.scala 27:20]
  wire  _T_4812 = _T_4684 & way_status_out_13; // @[Mux.scala 27:72]
  wire  _T_4939 = _T_4938 | _T_4812; // @[Mux.scala 27:72]
  wire  _T_4685 = ifu_ic_rw_int_addr_ff == 7'he; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_14; // @[Reg.scala 27:20]
  wire  _T_4813 = _T_4685 & way_status_out_14; // @[Mux.scala 27:72]
  wire  _T_4940 = _T_4939 | _T_4813; // @[Mux.scala 27:72]
  wire  _T_4686 = ifu_ic_rw_int_addr_ff == 7'hf; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_15; // @[Reg.scala 27:20]
  wire  _T_4814 = _T_4686 & way_status_out_15; // @[Mux.scala 27:72]
  wire  _T_4941 = _T_4940 | _T_4814; // @[Mux.scala 27:72]
  wire  _T_4687 = ifu_ic_rw_int_addr_ff == 7'h10; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_16; // @[Reg.scala 27:20]
  wire  _T_4815 = _T_4687 & way_status_out_16; // @[Mux.scala 27:72]
  wire  _T_4942 = _T_4941 | _T_4815; // @[Mux.scala 27:72]
  wire  _T_4688 = ifu_ic_rw_int_addr_ff == 7'h11; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_17; // @[Reg.scala 27:20]
  wire  _T_4816 = _T_4688 & way_status_out_17; // @[Mux.scala 27:72]
  wire  _T_4943 = _T_4942 | _T_4816; // @[Mux.scala 27:72]
  wire  _T_4689 = ifu_ic_rw_int_addr_ff == 7'h12; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_18; // @[Reg.scala 27:20]
  wire  _T_4817 = _T_4689 & way_status_out_18; // @[Mux.scala 27:72]
  wire  _T_4944 = _T_4943 | _T_4817; // @[Mux.scala 27:72]
  wire  _T_4690 = ifu_ic_rw_int_addr_ff == 7'h13; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_19; // @[Reg.scala 27:20]
  wire  _T_4818 = _T_4690 & way_status_out_19; // @[Mux.scala 27:72]
  wire  _T_4945 = _T_4944 | _T_4818; // @[Mux.scala 27:72]
  wire  _T_4691 = ifu_ic_rw_int_addr_ff == 7'h14; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_20; // @[Reg.scala 27:20]
  wire  _T_4819 = _T_4691 & way_status_out_20; // @[Mux.scala 27:72]
  wire  _T_4946 = _T_4945 | _T_4819; // @[Mux.scala 27:72]
  wire  _T_4692 = ifu_ic_rw_int_addr_ff == 7'h15; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_21; // @[Reg.scala 27:20]
  wire  _T_4820 = _T_4692 & way_status_out_21; // @[Mux.scala 27:72]
  wire  _T_4947 = _T_4946 | _T_4820; // @[Mux.scala 27:72]
  wire  _T_4693 = ifu_ic_rw_int_addr_ff == 7'h16; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_22; // @[Reg.scala 27:20]
  wire  _T_4821 = _T_4693 & way_status_out_22; // @[Mux.scala 27:72]
  wire  _T_4948 = _T_4947 | _T_4821; // @[Mux.scala 27:72]
  wire  _T_4694 = ifu_ic_rw_int_addr_ff == 7'h17; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_23; // @[Reg.scala 27:20]
  wire  _T_4822 = _T_4694 & way_status_out_23; // @[Mux.scala 27:72]
  wire  _T_4949 = _T_4948 | _T_4822; // @[Mux.scala 27:72]
  wire  _T_4695 = ifu_ic_rw_int_addr_ff == 7'h18; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_24; // @[Reg.scala 27:20]
  wire  _T_4823 = _T_4695 & way_status_out_24; // @[Mux.scala 27:72]
  wire  _T_4950 = _T_4949 | _T_4823; // @[Mux.scala 27:72]
  wire  _T_4696 = ifu_ic_rw_int_addr_ff == 7'h19; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_25; // @[Reg.scala 27:20]
  wire  _T_4824 = _T_4696 & way_status_out_25; // @[Mux.scala 27:72]
  wire  _T_4951 = _T_4950 | _T_4824; // @[Mux.scala 27:72]
  wire  _T_4697 = ifu_ic_rw_int_addr_ff == 7'h1a; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_26; // @[Reg.scala 27:20]
  wire  _T_4825 = _T_4697 & way_status_out_26; // @[Mux.scala 27:72]
  wire  _T_4952 = _T_4951 | _T_4825; // @[Mux.scala 27:72]
  wire  _T_4698 = ifu_ic_rw_int_addr_ff == 7'h1b; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_27; // @[Reg.scala 27:20]
  wire  _T_4826 = _T_4698 & way_status_out_27; // @[Mux.scala 27:72]
  wire  _T_4953 = _T_4952 | _T_4826; // @[Mux.scala 27:72]
  wire  _T_4699 = ifu_ic_rw_int_addr_ff == 7'h1c; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_28; // @[Reg.scala 27:20]
  wire  _T_4827 = _T_4699 & way_status_out_28; // @[Mux.scala 27:72]
  wire  _T_4954 = _T_4953 | _T_4827; // @[Mux.scala 27:72]
  wire  _T_4700 = ifu_ic_rw_int_addr_ff == 7'h1d; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_29; // @[Reg.scala 27:20]
  wire  _T_4828 = _T_4700 & way_status_out_29; // @[Mux.scala 27:72]
  wire  _T_4955 = _T_4954 | _T_4828; // @[Mux.scala 27:72]
  wire  _T_4701 = ifu_ic_rw_int_addr_ff == 7'h1e; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_30; // @[Reg.scala 27:20]
  wire  _T_4829 = _T_4701 & way_status_out_30; // @[Mux.scala 27:72]
  wire  _T_4956 = _T_4955 | _T_4829; // @[Mux.scala 27:72]
  wire  _T_4702 = ifu_ic_rw_int_addr_ff == 7'h1f; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_31; // @[Reg.scala 27:20]
  wire  _T_4830 = _T_4702 & way_status_out_31; // @[Mux.scala 27:72]
  wire  _T_4957 = _T_4956 | _T_4830; // @[Mux.scala 27:72]
  wire  _T_4703 = ifu_ic_rw_int_addr_ff == 7'h20; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_32; // @[Reg.scala 27:20]
  wire  _T_4831 = _T_4703 & way_status_out_32; // @[Mux.scala 27:72]
  wire  _T_4958 = _T_4957 | _T_4831; // @[Mux.scala 27:72]
  wire  _T_4704 = ifu_ic_rw_int_addr_ff == 7'h21; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_33; // @[Reg.scala 27:20]
  wire  _T_4832 = _T_4704 & way_status_out_33; // @[Mux.scala 27:72]
  wire  _T_4959 = _T_4958 | _T_4832; // @[Mux.scala 27:72]
  wire  _T_4705 = ifu_ic_rw_int_addr_ff == 7'h22; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_34; // @[Reg.scala 27:20]
  wire  _T_4833 = _T_4705 & way_status_out_34; // @[Mux.scala 27:72]
  wire  _T_4960 = _T_4959 | _T_4833; // @[Mux.scala 27:72]
  wire  _T_4706 = ifu_ic_rw_int_addr_ff == 7'h23; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_35; // @[Reg.scala 27:20]
  wire  _T_4834 = _T_4706 & way_status_out_35; // @[Mux.scala 27:72]
  wire  _T_4961 = _T_4960 | _T_4834; // @[Mux.scala 27:72]
  wire  _T_4707 = ifu_ic_rw_int_addr_ff == 7'h24; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_36; // @[Reg.scala 27:20]
  wire  _T_4835 = _T_4707 & way_status_out_36; // @[Mux.scala 27:72]
  wire  _T_4962 = _T_4961 | _T_4835; // @[Mux.scala 27:72]
  wire  _T_4708 = ifu_ic_rw_int_addr_ff == 7'h25; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_37; // @[Reg.scala 27:20]
  wire  _T_4836 = _T_4708 & way_status_out_37; // @[Mux.scala 27:72]
  wire  _T_4963 = _T_4962 | _T_4836; // @[Mux.scala 27:72]
  wire  _T_4709 = ifu_ic_rw_int_addr_ff == 7'h26; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_38; // @[Reg.scala 27:20]
  wire  _T_4837 = _T_4709 & way_status_out_38; // @[Mux.scala 27:72]
  wire  _T_4964 = _T_4963 | _T_4837; // @[Mux.scala 27:72]
  wire  _T_4710 = ifu_ic_rw_int_addr_ff == 7'h27; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_39; // @[Reg.scala 27:20]
  wire  _T_4838 = _T_4710 & way_status_out_39; // @[Mux.scala 27:72]
  wire  _T_4965 = _T_4964 | _T_4838; // @[Mux.scala 27:72]
  wire  _T_4711 = ifu_ic_rw_int_addr_ff == 7'h28; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_40; // @[Reg.scala 27:20]
  wire  _T_4839 = _T_4711 & way_status_out_40; // @[Mux.scala 27:72]
  wire  _T_4966 = _T_4965 | _T_4839; // @[Mux.scala 27:72]
  wire  _T_4712 = ifu_ic_rw_int_addr_ff == 7'h29; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_41; // @[Reg.scala 27:20]
  wire  _T_4840 = _T_4712 & way_status_out_41; // @[Mux.scala 27:72]
  wire  _T_4967 = _T_4966 | _T_4840; // @[Mux.scala 27:72]
  wire  _T_4713 = ifu_ic_rw_int_addr_ff == 7'h2a; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_42; // @[Reg.scala 27:20]
  wire  _T_4841 = _T_4713 & way_status_out_42; // @[Mux.scala 27:72]
  wire  _T_4968 = _T_4967 | _T_4841; // @[Mux.scala 27:72]
  wire  _T_4714 = ifu_ic_rw_int_addr_ff == 7'h2b; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_43; // @[Reg.scala 27:20]
  wire  _T_4842 = _T_4714 & way_status_out_43; // @[Mux.scala 27:72]
  wire  _T_4969 = _T_4968 | _T_4842; // @[Mux.scala 27:72]
  wire  _T_4715 = ifu_ic_rw_int_addr_ff == 7'h2c; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_44; // @[Reg.scala 27:20]
  wire  _T_4843 = _T_4715 & way_status_out_44; // @[Mux.scala 27:72]
  wire  _T_4970 = _T_4969 | _T_4843; // @[Mux.scala 27:72]
  wire  _T_4716 = ifu_ic_rw_int_addr_ff == 7'h2d; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_45; // @[Reg.scala 27:20]
  wire  _T_4844 = _T_4716 & way_status_out_45; // @[Mux.scala 27:72]
  wire  _T_4971 = _T_4970 | _T_4844; // @[Mux.scala 27:72]
  wire  _T_4717 = ifu_ic_rw_int_addr_ff == 7'h2e; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_46; // @[Reg.scala 27:20]
  wire  _T_4845 = _T_4717 & way_status_out_46; // @[Mux.scala 27:72]
  wire  _T_4972 = _T_4971 | _T_4845; // @[Mux.scala 27:72]
  wire  _T_4718 = ifu_ic_rw_int_addr_ff == 7'h2f; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_47; // @[Reg.scala 27:20]
  wire  _T_4846 = _T_4718 & way_status_out_47; // @[Mux.scala 27:72]
  wire  _T_4973 = _T_4972 | _T_4846; // @[Mux.scala 27:72]
  wire  _T_4719 = ifu_ic_rw_int_addr_ff == 7'h30; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_48; // @[Reg.scala 27:20]
  wire  _T_4847 = _T_4719 & way_status_out_48; // @[Mux.scala 27:72]
  wire  _T_4974 = _T_4973 | _T_4847; // @[Mux.scala 27:72]
  wire  _T_4720 = ifu_ic_rw_int_addr_ff == 7'h31; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_49; // @[Reg.scala 27:20]
  wire  _T_4848 = _T_4720 & way_status_out_49; // @[Mux.scala 27:72]
  wire  _T_4975 = _T_4974 | _T_4848; // @[Mux.scala 27:72]
  wire  _T_4721 = ifu_ic_rw_int_addr_ff == 7'h32; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_50; // @[Reg.scala 27:20]
  wire  _T_4849 = _T_4721 & way_status_out_50; // @[Mux.scala 27:72]
  wire  _T_4976 = _T_4975 | _T_4849; // @[Mux.scala 27:72]
  wire  _T_4722 = ifu_ic_rw_int_addr_ff == 7'h33; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_51; // @[Reg.scala 27:20]
  wire  _T_4850 = _T_4722 & way_status_out_51; // @[Mux.scala 27:72]
  wire  _T_4977 = _T_4976 | _T_4850; // @[Mux.scala 27:72]
  wire  _T_4723 = ifu_ic_rw_int_addr_ff == 7'h34; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_52; // @[Reg.scala 27:20]
  wire  _T_4851 = _T_4723 & way_status_out_52; // @[Mux.scala 27:72]
  wire  _T_4978 = _T_4977 | _T_4851; // @[Mux.scala 27:72]
  wire  _T_4724 = ifu_ic_rw_int_addr_ff == 7'h35; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_53; // @[Reg.scala 27:20]
  wire  _T_4852 = _T_4724 & way_status_out_53; // @[Mux.scala 27:72]
  wire  _T_4979 = _T_4978 | _T_4852; // @[Mux.scala 27:72]
  wire  _T_4725 = ifu_ic_rw_int_addr_ff == 7'h36; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_54; // @[Reg.scala 27:20]
  wire  _T_4853 = _T_4725 & way_status_out_54; // @[Mux.scala 27:72]
  wire  _T_4980 = _T_4979 | _T_4853; // @[Mux.scala 27:72]
  wire  _T_4726 = ifu_ic_rw_int_addr_ff == 7'h37; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_55; // @[Reg.scala 27:20]
  wire  _T_4854 = _T_4726 & way_status_out_55; // @[Mux.scala 27:72]
  wire  _T_4981 = _T_4980 | _T_4854; // @[Mux.scala 27:72]
  wire  _T_4727 = ifu_ic_rw_int_addr_ff == 7'h38; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_56; // @[Reg.scala 27:20]
  wire  _T_4855 = _T_4727 & way_status_out_56; // @[Mux.scala 27:72]
  wire  _T_4982 = _T_4981 | _T_4855; // @[Mux.scala 27:72]
  wire  _T_4728 = ifu_ic_rw_int_addr_ff == 7'h39; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_57; // @[Reg.scala 27:20]
  wire  _T_4856 = _T_4728 & way_status_out_57; // @[Mux.scala 27:72]
  wire  _T_4983 = _T_4982 | _T_4856; // @[Mux.scala 27:72]
  wire  _T_4729 = ifu_ic_rw_int_addr_ff == 7'h3a; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_58; // @[Reg.scala 27:20]
  wire  _T_4857 = _T_4729 & way_status_out_58; // @[Mux.scala 27:72]
  wire  _T_4984 = _T_4983 | _T_4857; // @[Mux.scala 27:72]
  wire  _T_4730 = ifu_ic_rw_int_addr_ff == 7'h3b; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_59; // @[Reg.scala 27:20]
  wire  _T_4858 = _T_4730 & way_status_out_59; // @[Mux.scala 27:72]
  wire  _T_4985 = _T_4984 | _T_4858; // @[Mux.scala 27:72]
  wire  _T_4731 = ifu_ic_rw_int_addr_ff == 7'h3c; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_60; // @[Reg.scala 27:20]
  wire  _T_4859 = _T_4731 & way_status_out_60; // @[Mux.scala 27:72]
  wire  _T_4986 = _T_4985 | _T_4859; // @[Mux.scala 27:72]
  wire  _T_4732 = ifu_ic_rw_int_addr_ff == 7'h3d; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_61; // @[Reg.scala 27:20]
  wire  _T_4860 = _T_4732 & way_status_out_61; // @[Mux.scala 27:72]
  wire  _T_4987 = _T_4986 | _T_4860; // @[Mux.scala 27:72]
  wire  _T_4733 = ifu_ic_rw_int_addr_ff == 7'h3e; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_62; // @[Reg.scala 27:20]
  wire  _T_4861 = _T_4733 & way_status_out_62; // @[Mux.scala 27:72]
  wire  _T_4988 = _T_4987 | _T_4861; // @[Mux.scala 27:72]
  wire  _T_4734 = ifu_ic_rw_int_addr_ff == 7'h3f; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_63; // @[Reg.scala 27:20]
  wire  _T_4862 = _T_4734 & way_status_out_63; // @[Mux.scala 27:72]
  wire  _T_4989 = _T_4988 | _T_4862; // @[Mux.scala 27:72]
  wire  _T_4735 = ifu_ic_rw_int_addr_ff == 7'h40; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_64; // @[Reg.scala 27:20]
  wire  _T_4863 = _T_4735 & way_status_out_64; // @[Mux.scala 27:72]
  wire  _T_4990 = _T_4989 | _T_4863; // @[Mux.scala 27:72]
  wire  _T_4736 = ifu_ic_rw_int_addr_ff == 7'h41; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_65; // @[Reg.scala 27:20]
  wire  _T_4864 = _T_4736 & way_status_out_65; // @[Mux.scala 27:72]
  wire  _T_4991 = _T_4990 | _T_4864; // @[Mux.scala 27:72]
  wire  _T_4737 = ifu_ic_rw_int_addr_ff == 7'h42; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_66; // @[Reg.scala 27:20]
  wire  _T_4865 = _T_4737 & way_status_out_66; // @[Mux.scala 27:72]
  wire  _T_4992 = _T_4991 | _T_4865; // @[Mux.scala 27:72]
  wire  _T_4738 = ifu_ic_rw_int_addr_ff == 7'h43; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_67; // @[Reg.scala 27:20]
  wire  _T_4866 = _T_4738 & way_status_out_67; // @[Mux.scala 27:72]
  wire  _T_4993 = _T_4992 | _T_4866; // @[Mux.scala 27:72]
  wire  _T_4739 = ifu_ic_rw_int_addr_ff == 7'h44; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_68; // @[Reg.scala 27:20]
  wire  _T_4867 = _T_4739 & way_status_out_68; // @[Mux.scala 27:72]
  wire  _T_4994 = _T_4993 | _T_4867; // @[Mux.scala 27:72]
  wire  _T_4740 = ifu_ic_rw_int_addr_ff == 7'h45; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_69; // @[Reg.scala 27:20]
  wire  _T_4868 = _T_4740 & way_status_out_69; // @[Mux.scala 27:72]
  wire  _T_4995 = _T_4994 | _T_4868; // @[Mux.scala 27:72]
  wire  _T_4741 = ifu_ic_rw_int_addr_ff == 7'h46; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_70; // @[Reg.scala 27:20]
  wire  _T_4869 = _T_4741 & way_status_out_70; // @[Mux.scala 27:72]
  wire  _T_4996 = _T_4995 | _T_4869; // @[Mux.scala 27:72]
  wire  _T_4742 = ifu_ic_rw_int_addr_ff == 7'h47; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_71; // @[Reg.scala 27:20]
  wire  _T_4870 = _T_4742 & way_status_out_71; // @[Mux.scala 27:72]
  wire  _T_4997 = _T_4996 | _T_4870; // @[Mux.scala 27:72]
  wire  _T_4743 = ifu_ic_rw_int_addr_ff == 7'h48; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_72; // @[Reg.scala 27:20]
  wire  _T_4871 = _T_4743 & way_status_out_72; // @[Mux.scala 27:72]
  wire  _T_4998 = _T_4997 | _T_4871; // @[Mux.scala 27:72]
  wire  _T_4744 = ifu_ic_rw_int_addr_ff == 7'h49; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_73; // @[Reg.scala 27:20]
  wire  _T_4872 = _T_4744 & way_status_out_73; // @[Mux.scala 27:72]
  wire  _T_4999 = _T_4998 | _T_4872; // @[Mux.scala 27:72]
  wire  _T_4745 = ifu_ic_rw_int_addr_ff == 7'h4a; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_74; // @[Reg.scala 27:20]
  wire  _T_4873 = _T_4745 & way_status_out_74; // @[Mux.scala 27:72]
  wire  _T_5000 = _T_4999 | _T_4873; // @[Mux.scala 27:72]
  wire  _T_4746 = ifu_ic_rw_int_addr_ff == 7'h4b; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_75; // @[Reg.scala 27:20]
  wire  _T_4874 = _T_4746 & way_status_out_75; // @[Mux.scala 27:72]
  wire  _T_5001 = _T_5000 | _T_4874; // @[Mux.scala 27:72]
  wire  _T_4747 = ifu_ic_rw_int_addr_ff == 7'h4c; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_76; // @[Reg.scala 27:20]
  wire  _T_4875 = _T_4747 & way_status_out_76; // @[Mux.scala 27:72]
  wire  _T_5002 = _T_5001 | _T_4875; // @[Mux.scala 27:72]
  wire  _T_4748 = ifu_ic_rw_int_addr_ff == 7'h4d; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_77; // @[Reg.scala 27:20]
  wire  _T_4876 = _T_4748 & way_status_out_77; // @[Mux.scala 27:72]
  wire  _T_5003 = _T_5002 | _T_4876; // @[Mux.scala 27:72]
  wire  _T_4749 = ifu_ic_rw_int_addr_ff == 7'h4e; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_78; // @[Reg.scala 27:20]
  wire  _T_4877 = _T_4749 & way_status_out_78; // @[Mux.scala 27:72]
  wire  _T_5004 = _T_5003 | _T_4877; // @[Mux.scala 27:72]
  wire  _T_4750 = ifu_ic_rw_int_addr_ff == 7'h4f; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_79; // @[Reg.scala 27:20]
  wire  _T_4878 = _T_4750 & way_status_out_79; // @[Mux.scala 27:72]
  wire  _T_5005 = _T_5004 | _T_4878; // @[Mux.scala 27:72]
  wire  _T_4751 = ifu_ic_rw_int_addr_ff == 7'h50; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_80; // @[Reg.scala 27:20]
  wire  _T_4879 = _T_4751 & way_status_out_80; // @[Mux.scala 27:72]
  wire  _T_5006 = _T_5005 | _T_4879; // @[Mux.scala 27:72]
  wire  _T_4752 = ifu_ic_rw_int_addr_ff == 7'h51; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_81; // @[Reg.scala 27:20]
  wire  _T_4880 = _T_4752 & way_status_out_81; // @[Mux.scala 27:72]
  wire  _T_5007 = _T_5006 | _T_4880; // @[Mux.scala 27:72]
  wire  _T_4753 = ifu_ic_rw_int_addr_ff == 7'h52; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_82; // @[Reg.scala 27:20]
  wire  _T_4881 = _T_4753 & way_status_out_82; // @[Mux.scala 27:72]
  wire  _T_5008 = _T_5007 | _T_4881; // @[Mux.scala 27:72]
  wire  _T_4754 = ifu_ic_rw_int_addr_ff == 7'h53; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_83; // @[Reg.scala 27:20]
  wire  _T_4882 = _T_4754 & way_status_out_83; // @[Mux.scala 27:72]
  wire  _T_5009 = _T_5008 | _T_4882; // @[Mux.scala 27:72]
  wire  _T_4755 = ifu_ic_rw_int_addr_ff == 7'h54; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_84; // @[Reg.scala 27:20]
  wire  _T_4883 = _T_4755 & way_status_out_84; // @[Mux.scala 27:72]
  wire  _T_5010 = _T_5009 | _T_4883; // @[Mux.scala 27:72]
  wire  _T_4756 = ifu_ic_rw_int_addr_ff == 7'h55; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_85; // @[Reg.scala 27:20]
  wire  _T_4884 = _T_4756 & way_status_out_85; // @[Mux.scala 27:72]
  wire  _T_5011 = _T_5010 | _T_4884; // @[Mux.scala 27:72]
  wire  _T_4757 = ifu_ic_rw_int_addr_ff == 7'h56; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_86; // @[Reg.scala 27:20]
  wire  _T_4885 = _T_4757 & way_status_out_86; // @[Mux.scala 27:72]
  wire  _T_5012 = _T_5011 | _T_4885; // @[Mux.scala 27:72]
  wire  _T_4758 = ifu_ic_rw_int_addr_ff == 7'h57; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_87; // @[Reg.scala 27:20]
  wire  _T_4886 = _T_4758 & way_status_out_87; // @[Mux.scala 27:72]
  wire  _T_5013 = _T_5012 | _T_4886; // @[Mux.scala 27:72]
  wire  _T_4759 = ifu_ic_rw_int_addr_ff == 7'h58; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_88; // @[Reg.scala 27:20]
  wire  _T_4887 = _T_4759 & way_status_out_88; // @[Mux.scala 27:72]
  wire  _T_5014 = _T_5013 | _T_4887; // @[Mux.scala 27:72]
  wire  _T_4760 = ifu_ic_rw_int_addr_ff == 7'h59; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_89; // @[Reg.scala 27:20]
  wire  _T_4888 = _T_4760 & way_status_out_89; // @[Mux.scala 27:72]
  wire  _T_5015 = _T_5014 | _T_4888; // @[Mux.scala 27:72]
  wire  _T_4761 = ifu_ic_rw_int_addr_ff == 7'h5a; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_90; // @[Reg.scala 27:20]
  wire  _T_4889 = _T_4761 & way_status_out_90; // @[Mux.scala 27:72]
  wire  _T_5016 = _T_5015 | _T_4889; // @[Mux.scala 27:72]
  wire  _T_4762 = ifu_ic_rw_int_addr_ff == 7'h5b; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_91; // @[Reg.scala 27:20]
  wire  _T_4890 = _T_4762 & way_status_out_91; // @[Mux.scala 27:72]
  wire  _T_5017 = _T_5016 | _T_4890; // @[Mux.scala 27:72]
  wire  _T_4763 = ifu_ic_rw_int_addr_ff == 7'h5c; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_92; // @[Reg.scala 27:20]
  wire  _T_4891 = _T_4763 & way_status_out_92; // @[Mux.scala 27:72]
  wire  _T_5018 = _T_5017 | _T_4891; // @[Mux.scala 27:72]
  wire  _T_4764 = ifu_ic_rw_int_addr_ff == 7'h5d; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_93; // @[Reg.scala 27:20]
  wire  _T_4892 = _T_4764 & way_status_out_93; // @[Mux.scala 27:72]
  wire  _T_5019 = _T_5018 | _T_4892; // @[Mux.scala 27:72]
  wire  _T_4765 = ifu_ic_rw_int_addr_ff == 7'h5e; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_94; // @[Reg.scala 27:20]
  wire  _T_4893 = _T_4765 & way_status_out_94; // @[Mux.scala 27:72]
  wire  _T_5020 = _T_5019 | _T_4893; // @[Mux.scala 27:72]
  wire  _T_4766 = ifu_ic_rw_int_addr_ff == 7'h5f; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_95; // @[Reg.scala 27:20]
  wire  _T_4894 = _T_4766 & way_status_out_95; // @[Mux.scala 27:72]
  wire  _T_5021 = _T_5020 | _T_4894; // @[Mux.scala 27:72]
  wire  _T_4767 = ifu_ic_rw_int_addr_ff == 7'h60; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_96; // @[Reg.scala 27:20]
  wire  _T_4895 = _T_4767 & way_status_out_96; // @[Mux.scala 27:72]
  wire  _T_5022 = _T_5021 | _T_4895; // @[Mux.scala 27:72]
  wire  _T_4768 = ifu_ic_rw_int_addr_ff == 7'h61; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_97; // @[Reg.scala 27:20]
  wire  _T_4896 = _T_4768 & way_status_out_97; // @[Mux.scala 27:72]
  wire  _T_5023 = _T_5022 | _T_4896; // @[Mux.scala 27:72]
  wire  _T_4769 = ifu_ic_rw_int_addr_ff == 7'h62; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_98; // @[Reg.scala 27:20]
  wire  _T_4897 = _T_4769 & way_status_out_98; // @[Mux.scala 27:72]
  wire  _T_5024 = _T_5023 | _T_4897; // @[Mux.scala 27:72]
  wire  _T_4770 = ifu_ic_rw_int_addr_ff == 7'h63; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_99; // @[Reg.scala 27:20]
  wire  _T_4898 = _T_4770 & way_status_out_99; // @[Mux.scala 27:72]
  wire  _T_5025 = _T_5024 | _T_4898; // @[Mux.scala 27:72]
  wire  _T_4771 = ifu_ic_rw_int_addr_ff == 7'h64; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_100; // @[Reg.scala 27:20]
  wire  _T_4899 = _T_4771 & way_status_out_100; // @[Mux.scala 27:72]
  wire  _T_5026 = _T_5025 | _T_4899; // @[Mux.scala 27:72]
  wire  _T_4772 = ifu_ic_rw_int_addr_ff == 7'h65; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_101; // @[Reg.scala 27:20]
  wire  _T_4900 = _T_4772 & way_status_out_101; // @[Mux.scala 27:72]
  wire  _T_5027 = _T_5026 | _T_4900; // @[Mux.scala 27:72]
  wire  _T_4773 = ifu_ic_rw_int_addr_ff == 7'h66; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_102; // @[Reg.scala 27:20]
  wire  _T_4901 = _T_4773 & way_status_out_102; // @[Mux.scala 27:72]
  wire  _T_5028 = _T_5027 | _T_4901; // @[Mux.scala 27:72]
  wire  _T_4774 = ifu_ic_rw_int_addr_ff == 7'h67; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_103; // @[Reg.scala 27:20]
  wire  _T_4902 = _T_4774 & way_status_out_103; // @[Mux.scala 27:72]
  wire  _T_5029 = _T_5028 | _T_4902; // @[Mux.scala 27:72]
  wire  _T_4775 = ifu_ic_rw_int_addr_ff == 7'h68; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_104; // @[Reg.scala 27:20]
  wire  _T_4903 = _T_4775 & way_status_out_104; // @[Mux.scala 27:72]
  wire  _T_5030 = _T_5029 | _T_4903; // @[Mux.scala 27:72]
  wire  _T_4776 = ifu_ic_rw_int_addr_ff == 7'h69; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_105; // @[Reg.scala 27:20]
  wire  _T_4904 = _T_4776 & way_status_out_105; // @[Mux.scala 27:72]
  wire  _T_5031 = _T_5030 | _T_4904; // @[Mux.scala 27:72]
  wire  _T_4777 = ifu_ic_rw_int_addr_ff == 7'h6a; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_106; // @[Reg.scala 27:20]
  wire  _T_4905 = _T_4777 & way_status_out_106; // @[Mux.scala 27:72]
  wire  _T_5032 = _T_5031 | _T_4905; // @[Mux.scala 27:72]
  wire  _T_4778 = ifu_ic_rw_int_addr_ff == 7'h6b; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_107; // @[Reg.scala 27:20]
  wire  _T_4906 = _T_4778 & way_status_out_107; // @[Mux.scala 27:72]
  wire  _T_5033 = _T_5032 | _T_4906; // @[Mux.scala 27:72]
  wire  _T_4779 = ifu_ic_rw_int_addr_ff == 7'h6c; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_108; // @[Reg.scala 27:20]
  wire  _T_4907 = _T_4779 & way_status_out_108; // @[Mux.scala 27:72]
  wire  _T_5034 = _T_5033 | _T_4907; // @[Mux.scala 27:72]
  wire  _T_4780 = ifu_ic_rw_int_addr_ff == 7'h6d; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_109; // @[Reg.scala 27:20]
  wire  _T_4908 = _T_4780 & way_status_out_109; // @[Mux.scala 27:72]
  wire  _T_5035 = _T_5034 | _T_4908; // @[Mux.scala 27:72]
  wire  _T_4781 = ifu_ic_rw_int_addr_ff == 7'h6e; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_110; // @[Reg.scala 27:20]
  wire  _T_4909 = _T_4781 & way_status_out_110; // @[Mux.scala 27:72]
  wire  _T_5036 = _T_5035 | _T_4909; // @[Mux.scala 27:72]
  wire  _T_4782 = ifu_ic_rw_int_addr_ff == 7'h6f; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_111; // @[Reg.scala 27:20]
  wire  _T_4910 = _T_4782 & way_status_out_111; // @[Mux.scala 27:72]
  wire  _T_5037 = _T_5036 | _T_4910; // @[Mux.scala 27:72]
  wire  _T_4783 = ifu_ic_rw_int_addr_ff == 7'h70; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_112; // @[Reg.scala 27:20]
  wire  _T_4911 = _T_4783 & way_status_out_112; // @[Mux.scala 27:72]
  wire  _T_5038 = _T_5037 | _T_4911; // @[Mux.scala 27:72]
  wire  _T_4784 = ifu_ic_rw_int_addr_ff == 7'h71; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_113; // @[Reg.scala 27:20]
  wire  _T_4912 = _T_4784 & way_status_out_113; // @[Mux.scala 27:72]
  wire  _T_5039 = _T_5038 | _T_4912; // @[Mux.scala 27:72]
  wire  _T_4785 = ifu_ic_rw_int_addr_ff == 7'h72; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_114; // @[Reg.scala 27:20]
  wire  _T_4913 = _T_4785 & way_status_out_114; // @[Mux.scala 27:72]
  wire  _T_5040 = _T_5039 | _T_4913; // @[Mux.scala 27:72]
  wire  _T_4786 = ifu_ic_rw_int_addr_ff == 7'h73; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_115; // @[Reg.scala 27:20]
  wire  _T_4914 = _T_4786 & way_status_out_115; // @[Mux.scala 27:72]
  wire  _T_5041 = _T_5040 | _T_4914; // @[Mux.scala 27:72]
  wire  _T_4787 = ifu_ic_rw_int_addr_ff == 7'h74; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_116; // @[Reg.scala 27:20]
  wire  _T_4915 = _T_4787 & way_status_out_116; // @[Mux.scala 27:72]
  wire  _T_5042 = _T_5041 | _T_4915; // @[Mux.scala 27:72]
  wire  _T_4788 = ifu_ic_rw_int_addr_ff == 7'h75; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_117; // @[Reg.scala 27:20]
  wire  _T_4916 = _T_4788 & way_status_out_117; // @[Mux.scala 27:72]
  wire  _T_5043 = _T_5042 | _T_4916; // @[Mux.scala 27:72]
  wire  _T_4789 = ifu_ic_rw_int_addr_ff == 7'h76; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_118; // @[Reg.scala 27:20]
  wire  _T_4917 = _T_4789 & way_status_out_118; // @[Mux.scala 27:72]
  wire  _T_5044 = _T_5043 | _T_4917; // @[Mux.scala 27:72]
  wire  _T_4790 = ifu_ic_rw_int_addr_ff == 7'h77; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_119; // @[Reg.scala 27:20]
  wire  _T_4918 = _T_4790 & way_status_out_119; // @[Mux.scala 27:72]
  wire  _T_5045 = _T_5044 | _T_4918; // @[Mux.scala 27:72]
  wire  _T_4791 = ifu_ic_rw_int_addr_ff == 7'h78; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_120; // @[Reg.scala 27:20]
  wire  _T_4919 = _T_4791 & way_status_out_120; // @[Mux.scala 27:72]
  wire  _T_5046 = _T_5045 | _T_4919; // @[Mux.scala 27:72]
  wire  _T_4792 = ifu_ic_rw_int_addr_ff == 7'h79; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_121; // @[Reg.scala 27:20]
  wire  _T_4920 = _T_4792 & way_status_out_121; // @[Mux.scala 27:72]
  wire  _T_5047 = _T_5046 | _T_4920; // @[Mux.scala 27:72]
  wire  _T_4793 = ifu_ic_rw_int_addr_ff == 7'h7a; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_122; // @[Reg.scala 27:20]
  wire  _T_4921 = _T_4793 & way_status_out_122; // @[Mux.scala 27:72]
  wire  _T_5048 = _T_5047 | _T_4921; // @[Mux.scala 27:72]
  wire  _T_4794 = ifu_ic_rw_int_addr_ff == 7'h7b; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_123; // @[Reg.scala 27:20]
  wire  _T_4922 = _T_4794 & way_status_out_123; // @[Mux.scala 27:72]
  wire  _T_5049 = _T_5048 | _T_4922; // @[Mux.scala 27:72]
  wire  _T_4795 = ifu_ic_rw_int_addr_ff == 7'h7c; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_124; // @[Reg.scala 27:20]
  wire  _T_4923 = _T_4795 & way_status_out_124; // @[Mux.scala 27:72]
  wire  _T_5050 = _T_5049 | _T_4923; // @[Mux.scala 27:72]
  wire  _T_4796 = ifu_ic_rw_int_addr_ff == 7'h7d; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_125; // @[Reg.scala 27:20]
  wire  _T_4924 = _T_4796 & way_status_out_125; // @[Mux.scala 27:72]
  wire  _T_5051 = _T_5050 | _T_4924; // @[Mux.scala 27:72]
  wire  _T_4797 = ifu_ic_rw_int_addr_ff == 7'h7e; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_126; // @[Reg.scala 27:20]
  wire  _T_4925 = _T_4797 & way_status_out_126; // @[Mux.scala 27:72]
  wire  _T_5052 = _T_5051 | _T_4925; // @[Mux.scala 27:72]
  wire  _T_4798 = ifu_ic_rw_int_addr_ff == 7'h7f; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_127; // @[Reg.scala 27:20]
  wire  _T_4926 = _T_4798 & way_status_out_127; // @[Mux.scala 27:72]
  wire  way_status = _T_5052 | _T_4926; // @[Mux.scala 27:72]
  wire  _T_195 = ~reset_all_tags; // @[ifu_mem_ctl.scala 168:96]
  wire [1:0] _T_197 = _T_195 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire  _T_212 = _T_231 | _T_239; // @[ifu_mem_ctl.scala 182:59]
  wire  _T_214 = _T_212 | _T_2268; // @[ifu_mem_ctl.scala 182:91]
  wire  ic_iccm_hit_f = fetch_req_iccm_f & _T_214; // @[ifu_mem_ctl.scala 182:41]
  wire  _T_219 = _T_227 & fetch_req_icache_f; // @[ifu_mem_ctl.scala 188:39]
  wire  _T_221 = _T_219 & _T_195; // @[ifu_mem_ctl.scala 188:60]
  wire  _T_225 = _T_221 & _T_212; // @[ifu_mem_ctl.scala 188:78]
  wire  ic_act_hit_f = _T_225 & _T_247; // @[ifu_mem_ctl.scala 188:126]
  wire  _T_262 = ic_act_hit_f | ic_byp_hit_f; // @[ifu_mem_ctl.scala 195:31]
  wire  _T_263 = _T_262 | ic_iccm_hit_f; // @[ifu_mem_ctl.scala 195:46]
  wire  _T_264 = ifc_region_acc_fault_final_f & ifc_fetch_req_f; // @[ifu_mem_ctl.scala 195:94]
  reg  way_status_mb_ff; // @[ifu_mem_ctl.scala 223:59]
  wire  _T_9756 = ~way_status_mb_ff; // @[ifu_mem_ctl.scala 720:33]
  reg [1:0] tagv_mb_ff; // @[ifu_mem_ctl.scala 224:53]
  wire  _T_9758 = _T_9756 & tagv_mb_ff[0]; // @[ifu_mem_ctl.scala 720:51]
  wire  _T_9760 = _T_9758 & tagv_mb_ff[1]; // @[ifu_mem_ctl.scala 720:67]
  wire  _T_9762 = ~tagv_mb_ff[0]; // @[ifu_mem_ctl.scala 720:86]
  wire  replace_way_mb_any_0 = _T_9760 | _T_9762; // @[ifu_mem_ctl.scala 720:84]
  wire  _T_9765 = way_status_mb_ff & tagv_mb_ff[0]; // @[ifu_mem_ctl.scala 721:50]
  wire  _T_9767 = _T_9765 & tagv_mb_ff[1]; // @[ifu_mem_ctl.scala 721:66]
  wire  _T_9769 = ~tagv_mb_ff[1]; // @[ifu_mem_ctl.scala 721:85]
  wire  _T_9771 = _T_9769 & tagv_mb_ff[0]; // @[ifu_mem_ctl.scala 721:100]
  wire  replace_way_mb_any_1 = _T_9767 | _T_9771; // @[ifu_mem_ctl.scala 721:83]
  wire [1:0] _T_295 = io_ic_tag_valid & _T_197; // @[ifu_mem_ctl.scala 208:56]
  reg  reset_ic_ff; // @[ifu_mem_ctl.scala 212:48]
  wire  _T_299 = reset_all_tags | reset_ic_ff; // @[ifu_mem_ctl.scala 211:72]
  wire  reset_ic_in = miss_pending & _T_299; // @[ifu_mem_ctl.scala 211:53]
  reg  fetch_uncacheable_ff; // @[ifu_mem_ctl.scala 213:62]
  reg [25:0] miss_addr; // @[ifu_mem_ctl.scala 222:48]
  wire  _T_309 = io_ifu_bus_clk_en | ic_act_miss_f; // @[ifu_mem_ctl.scala 221:57]
  wire  _T_315 = _T_2283 & flush_final_f; // @[ifu_mem_ctl.scala 226:87]
  wire  _T_316 = ~_T_315; // @[ifu_mem_ctl.scala 226:55]
  wire  _T_317 = io_ifc_fetch_req_bf & _T_316; // @[ifu_mem_ctl.scala 226:53]
  wire  _T_2275 = ~_T_2270; // @[ifu_mem_ctl.scala 373:46]
  wire  _T_2276 = _T_2268 & _T_2275; // @[ifu_mem_ctl.scala 373:44]
  wire  stream_miss_f = _T_2276 & ifc_fetch_req_f; // @[ifu_mem_ctl.scala 373:84]
  wire  _T_318 = ~stream_miss_f; // @[ifu_mem_ctl.scala 226:106]
  reg  ifc_region_acc_fault_f; // @[ifu_mem_ctl.scala 232:68]
  reg [2:0] bus_rd_addr_count; // @[ifu_mem_ctl.scala 540:55]
  wire  _T_325 = _T_239 | _T_2268; // @[ifu_mem_ctl.scala 234:55]
  reg  ic_act_miss_f_delayed; // @[ifu_mem_ctl.scala 555:61]
  wire  _T_2687 = ic_act_miss_f_delayed & _T_2284; // @[ifu_mem_ctl.scala 556:53]
  wire  reset_tag_valid_for_miss = _T_2687 & _T_17; // @[ifu_mem_ctl.scala 556:84]
  wire [30:0] _T_338 = {imb_ff[30:5],3'h0,imb_ff[1:0]}; // @[Cat.scala 29:58]
  wire  _T_339 = ~reset_tag_valid_for_miss; // @[ifu_mem_ctl.scala 240:37]
  wire [30:0] _T_340 = reset_tag_valid_for_miss ? _T_338 : 31'h0; // @[Mux.scala 27:72]
  wire [30:0] _T_341 = _T_339 ? io_ifc_fetch_addr_bf : 31'h0; // @[Mux.scala 27:72]
  wire [30:0] ifu_ic_rw_int_addr = _T_340 | _T_341; // @[Mux.scala 27:72]
  wire [30:0] ifu_status_wr_addr = reset_tag_valid_for_miss ? _T_338 : ifu_fetch_addr_int_f; // @[ifu_mem_ctl.scala 243:31]
  wire  _T_1199 = |io_ic_eccerr; // @[ifu_mem_ctl.scala 256:73]
  wire  _T_1200 = _T_1199 & ic_act_hit_f; // @[ifu_mem_ctl.scala 256:100]
  wire [4:0] bypass_index = imb_ff[4:0]; // @[ifu_mem_ctl.scala 328:28]
  wire  _T_1404 = bypass_index[4:2] == 3'h0; // @[ifu_mem_ctl.scala 330:114]
  wire  _T_1330 = ~ic_act_miss_f; // @[ifu_mem_ctl.scala 319:118]
  wire  ic_miss_buff_data_valid_in_0 = ic_miss_buff_data_valid[0] & _T_1330; // @[ifu_mem_ctl.scala 319:116]
  wire  _T_1427 = _T_1404 & ic_miss_buff_data_valid_in_0; // @[Mux.scala 27:72]
  wire  _T_1407 = bypass_index[4:2] == 3'h1; // @[ifu_mem_ctl.scala 330:114]
  wire  ic_miss_buff_data_valid_in_1 = ic_miss_buff_data_valid[1] & _T_1330; // @[ifu_mem_ctl.scala 319:116]
  wire  _T_1428 = _T_1407 & ic_miss_buff_data_valid_in_1; // @[Mux.scala 27:72]
  wire  _T_1435 = _T_1427 | _T_1428; // @[Mux.scala 27:72]
  wire  _T_1410 = bypass_index[4:2] == 3'h2; // @[ifu_mem_ctl.scala 330:114]
  wire  ic_miss_buff_data_valid_in_2 = ic_miss_buff_data_valid[2] & _T_1330; // @[ifu_mem_ctl.scala 319:116]
  wire  _T_1429 = _T_1410 & ic_miss_buff_data_valid_in_2; // @[Mux.scala 27:72]
  wire  _T_1436 = _T_1435 | _T_1429; // @[Mux.scala 27:72]
  wire  _T_1413 = bypass_index[4:2] == 3'h3; // @[ifu_mem_ctl.scala 330:114]
  wire  ic_miss_buff_data_valid_in_3 = ic_miss_buff_data_valid[3] & _T_1330; // @[ifu_mem_ctl.scala 319:116]
  wire  _T_1430 = _T_1413 & ic_miss_buff_data_valid_in_3; // @[Mux.scala 27:72]
  wire  _T_1437 = _T_1436 | _T_1430; // @[Mux.scala 27:72]
  wire  _T_1416 = bypass_index[4:2] == 3'h4; // @[ifu_mem_ctl.scala 330:114]
  wire  ic_miss_buff_data_valid_in_4 = ic_miss_buff_data_valid[4] & _T_1330; // @[ifu_mem_ctl.scala 319:116]
  wire  _T_1431 = _T_1416 & ic_miss_buff_data_valid_in_4; // @[Mux.scala 27:72]
  wire  _T_1438 = _T_1437 | _T_1431; // @[Mux.scala 27:72]
  wire  _T_1419 = bypass_index[4:2] == 3'h5; // @[ifu_mem_ctl.scala 330:114]
  wire  ic_miss_buff_data_valid_in_5 = ic_miss_buff_data_valid[5] & _T_1330; // @[ifu_mem_ctl.scala 319:116]
  wire  _T_1432 = _T_1419 & ic_miss_buff_data_valid_in_5; // @[Mux.scala 27:72]
  wire  _T_1439 = _T_1438 | _T_1432; // @[Mux.scala 27:72]
  wire  _T_1422 = bypass_index[4:2] == 3'h6; // @[ifu_mem_ctl.scala 330:114]
  wire  ic_miss_buff_data_valid_in_6 = ic_miss_buff_data_valid[6] & _T_1330; // @[ifu_mem_ctl.scala 319:116]
  wire  _T_1433 = _T_1422 & ic_miss_buff_data_valid_in_6; // @[Mux.scala 27:72]
  wire  _T_1440 = _T_1439 | _T_1433; // @[Mux.scala 27:72]
  wire  _T_1425 = bypass_index[4:2] == 3'h7; // @[ifu_mem_ctl.scala 330:114]
  wire  ic_miss_buff_data_valid_in_7 = ic_miss_buff_data_valid[7] & _T_1330; // @[ifu_mem_ctl.scala 319:116]
  wire  _T_1434 = _T_1425 & ic_miss_buff_data_valid_in_7; // @[Mux.scala 27:72]
  wire  bypass_valid_value_check = _T_1440 | _T_1434; // @[Mux.scala 27:72]
  wire  _T_1443 = ~bypass_index[1]; // @[ifu_mem_ctl.scala 331:58]
  wire  _T_1444 = bypass_valid_value_check & _T_1443; // @[ifu_mem_ctl.scala 331:56]
  wire  _T_1446 = ~bypass_index[0]; // @[ifu_mem_ctl.scala 331:77]
  wire  _T_1447 = _T_1444 & _T_1446; // @[ifu_mem_ctl.scala 331:75]
  wire  _T_1452 = _T_1444 & bypass_index[0]; // @[ifu_mem_ctl.scala 332:75]
  wire  _T_1453 = _T_1447 | _T_1452; // @[ifu_mem_ctl.scala 331:95]
  wire  _T_1455 = bypass_valid_value_check & bypass_index[1]; // @[ifu_mem_ctl.scala 333:56]
  wire  _T_1458 = _T_1455 & _T_1446; // @[ifu_mem_ctl.scala 333:74]
  wire  _T_1459 = _T_1453 | _T_1458; // @[ifu_mem_ctl.scala 332:94]
  wire  _T_1463 = _T_1455 & bypass_index[0]; // @[ifu_mem_ctl.scala 334:51]
  wire [2:0] bypass_index_5_3_inc = bypass_index[4:2] + 3'h1; // @[ifu_mem_ctl.scala 329:70]
  wire  _T_1464 = bypass_index_5_3_inc == 3'h0; // @[ifu_mem_ctl.scala 334:132]
  wire  _T_1480 = _T_1464 & ic_miss_buff_data_valid_in_0; // @[Mux.scala 27:72]
  wire  _T_1466 = bypass_index_5_3_inc == 3'h1; // @[ifu_mem_ctl.scala 334:132]
  wire  _T_1481 = _T_1466 & ic_miss_buff_data_valid_in_1; // @[Mux.scala 27:72]
  wire  _T_1488 = _T_1480 | _T_1481; // @[Mux.scala 27:72]
  wire  _T_1468 = bypass_index_5_3_inc == 3'h2; // @[ifu_mem_ctl.scala 334:132]
  wire  _T_1482 = _T_1468 & ic_miss_buff_data_valid_in_2; // @[Mux.scala 27:72]
  wire  _T_1489 = _T_1488 | _T_1482; // @[Mux.scala 27:72]
  wire  _T_1470 = bypass_index_5_3_inc == 3'h3; // @[ifu_mem_ctl.scala 334:132]
  wire  _T_1483 = _T_1470 & ic_miss_buff_data_valid_in_3; // @[Mux.scala 27:72]
  wire  _T_1490 = _T_1489 | _T_1483; // @[Mux.scala 27:72]
  wire  _T_1472 = bypass_index_5_3_inc == 3'h4; // @[ifu_mem_ctl.scala 334:132]
  wire  _T_1484 = _T_1472 & ic_miss_buff_data_valid_in_4; // @[Mux.scala 27:72]
  wire  _T_1491 = _T_1490 | _T_1484; // @[Mux.scala 27:72]
  wire  _T_1474 = bypass_index_5_3_inc == 3'h5; // @[ifu_mem_ctl.scala 334:132]
  wire  _T_1485 = _T_1474 & ic_miss_buff_data_valid_in_5; // @[Mux.scala 27:72]
  wire  _T_1492 = _T_1491 | _T_1485; // @[Mux.scala 27:72]
  wire  _T_1476 = bypass_index_5_3_inc == 3'h6; // @[ifu_mem_ctl.scala 334:132]
  wire  _T_1486 = _T_1476 & ic_miss_buff_data_valid_in_6; // @[Mux.scala 27:72]
  wire  _T_1493 = _T_1492 | _T_1486; // @[Mux.scala 27:72]
  wire  _T_1478 = bypass_index_5_3_inc == 3'h7; // @[ifu_mem_ctl.scala 334:132]
  wire  _T_1487 = _T_1478 & ic_miss_buff_data_valid_in_7; // @[Mux.scala 27:72]
  wire  _T_1494 = _T_1493 | _T_1487; // @[Mux.scala 27:72]
  wire  _T_1496 = _T_1463 & _T_1494; // @[ifu_mem_ctl.scala 334:69]
  wire  _T_1497 = _T_1459 | _T_1496; // @[ifu_mem_ctl.scala 333:94]
  wire [4:0] _GEN_436 = {{2'd0}, bypass_index[4:2]}; // @[ifu_mem_ctl.scala 335:95]
  wire  _T_1500 = _GEN_436 == 5'h1f; // @[ifu_mem_ctl.scala 335:95]
  wire  _T_1501 = bypass_valid_value_check & _T_1500; // @[ifu_mem_ctl.scala 335:56]
  wire  bypass_data_ready_in = _T_1497 | _T_1501; // @[ifu_mem_ctl.scala 334:181]
  wire  _T_1502 = bypass_data_ready_in & crit_wd_byp_ok_ff; // @[ifu_mem_ctl.scala 339:53]
  wire  _T_1503 = _T_1502 & uncacheable_miss_ff; // @[ifu_mem_ctl.scala 339:73]
  wire  _T_1505 = _T_1503 & _T_319; // @[ifu_mem_ctl.scala 339:96]
  wire  _T_1507 = _T_1505 & _T_58; // @[ifu_mem_ctl.scala 339:118]
  wire  _T_1509 = crit_wd_byp_ok_ff & _T_17; // @[ifu_mem_ctl.scala 340:73]
  wire  _T_1511 = _T_1509 & _T_319; // @[ifu_mem_ctl.scala 340:96]
  wire  _T_1513 = _T_1511 & _T_58; // @[ifu_mem_ctl.scala 340:118]
  wire  _T_1514 = _T_1507 | _T_1513; // @[ifu_mem_ctl.scala 339:143]
  reg  ic_crit_wd_rdy_new_ff; // @[ifu_mem_ctl.scala 342:58]
  wire  _T_1515 = ic_crit_wd_rdy_new_ff & crit_wd_byp_ok_ff; // @[ifu_mem_ctl.scala 341:54]
  wire  _T_1516 = ~fetch_req_icache_f; // @[ifu_mem_ctl.scala 341:76]
  wire  _T_1517 = _T_1515 & _T_1516; // @[ifu_mem_ctl.scala 341:74]
  wire  _T_1519 = _T_1517 & _T_319; // @[ifu_mem_ctl.scala 341:96]
  wire  ic_crit_wd_rdy_new_in = _T_1514 | _T_1519; // @[ifu_mem_ctl.scala 340:143]
  wire  ic_crit_wd_rdy = ic_crit_wd_rdy_new_in | ic_crit_wd_rdy_new_ff; // @[ifu_mem_ctl.scala 561:43]
  wire  _T_1252 = ic_crit_wd_rdy | _T_2268; // @[ifu_mem_ctl.scala 280:38]
  wire  _T_1254 = _T_1252 | _T_2284; // @[ifu_mem_ctl.scala 280:64]
  wire  _T_1255 = ~_T_1254; // @[ifu_mem_ctl.scala 280:21]
  wire  _T_1256 = ~fetch_req_iccm_f; // @[ifu_mem_ctl.scala 280:98]
  wire  sel_ic_data = _T_1255 & _T_1256; // @[ifu_mem_ctl.scala 280:96]
  wire  _T_2491 = io_ic_tag_perr & sel_ic_data; // @[ifu_mem_ctl.scala 385:44]
  wire  _T_1612 = ~ifu_fetch_addr_int_f[1]; // @[ifu_mem_ctl.scala 351:30]
  wire  _T_1614 = ~ifu_fetch_addr_int_f[0]; // @[ifu_mem_ctl.scala 351:57]
  wire  _T_1615 = _T_1612 & _T_1614; // @[ifu_mem_ctl.scala 351:55]
  reg [7:0] ic_miss_buff_data_error; // @[ifu_mem_ctl.scala 325:60]
  wire [7:0] _T_1617 = ic_miss_buff_data_error >> byp_fetch_index[4:2]; // @[ifu_mem_ctl.scala 351:107]
  wire  _T_1619 = _T_1615 & _T_1617[0]; // @[ifu_mem_ctl.scala 351:82]
  wire  _T_1623 = _T_1612 & ifu_fetch_addr_int_f[0]; // @[ifu_mem_ctl.scala 352:33]
  wire  _T_1627 = _T_1623 & _T_1617[0]; // @[ifu_mem_ctl.scala 352:60]
  wire  _T_1628 = _T_1619 | _T_1627; // @[ifu_mem_ctl.scala 351:151]
  wire  _T_1637 = _T_1628 | _T_1627; // @[ifu_mem_ctl.scala 352:129]
  wire  _T_1641 = ifu_fetch_addr_int_f[1] & _T_1614; // @[ifu_mem_ctl.scala 354:33]
  wire  _T_1645 = _T_1641 & _T_1617[0]; // @[ifu_mem_ctl.scala 354:60]
  wire  _T_1646 = _T_1637 | _T_1645; // @[ifu_mem_ctl.scala 353:129]
  wire  _T_1649 = ifu_fetch_addr_int_f[1] & ifu_fetch_addr_int_f[0]; // @[ifu_mem_ctl.scala 355:32]
  wire [7:0] _T_1654 = ic_miss_buff_data_error >> byp_fetch_index_inc; // @[ifu_mem_ctl.scala 356:32]
  wire  _T_1656 = _T_1617[0] | _T_1654[0]; // @[ifu_mem_ctl.scala 355:127]
  wire  _T_1657 = _T_1649 & _T_1656; // @[ifu_mem_ctl.scala 355:58]
  wire  ifu_byp_data_err_new = _T_1646 | _T_1657; // @[ifu_mem_ctl.scala 354:129]
  wire  ifc_bus_acc_fault_f = ic_byp_hit_f & ifu_byp_data_err_new; // @[ifu_mem_ctl.scala 297:42]
  wire  _T_2492 = ifc_region_acc_fault_final_f | ifc_bus_acc_fault_f; // @[ifu_mem_ctl.scala 385:91]
  wire  _T_2493 = ~_T_2492; // @[ifu_mem_ctl.scala 385:60]
  wire  ic_rd_parity_final_err = _T_2491 & _T_2493; // @[ifu_mem_ctl.scala 385:58]
  reg  ic_debug_ict_array_sel_ff; // @[ifu_mem_ctl.scala 768:63]
  reg  ic_tag_valid_out_1_0; // @[Reg.scala 27:20]
  wire  _T_9374 = _T_4671 & ic_tag_valid_out_1_0; // @[ifu_mem_ctl.scala 696:10]
  reg  ic_tag_valid_out_1_1; // @[Reg.scala 27:20]
  wire  _T_9376 = _T_4672 & ic_tag_valid_out_1_1; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9629 = _T_9374 | _T_9376; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_2; // @[Reg.scala 27:20]
  wire  _T_9378 = _T_4673 & ic_tag_valid_out_1_2; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9630 = _T_9629 | _T_9378; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_3; // @[Reg.scala 27:20]
  wire  _T_9380 = _T_4674 & ic_tag_valid_out_1_3; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9631 = _T_9630 | _T_9380; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_4; // @[Reg.scala 27:20]
  wire  _T_9382 = _T_4675 & ic_tag_valid_out_1_4; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9632 = _T_9631 | _T_9382; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_5; // @[Reg.scala 27:20]
  wire  _T_9384 = _T_4676 & ic_tag_valid_out_1_5; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9633 = _T_9632 | _T_9384; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_6; // @[Reg.scala 27:20]
  wire  _T_9386 = _T_4677 & ic_tag_valid_out_1_6; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9634 = _T_9633 | _T_9386; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_7; // @[Reg.scala 27:20]
  wire  _T_9388 = _T_4678 & ic_tag_valid_out_1_7; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9635 = _T_9634 | _T_9388; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_8; // @[Reg.scala 27:20]
  wire  _T_9390 = _T_4679 & ic_tag_valid_out_1_8; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9636 = _T_9635 | _T_9390; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_9; // @[Reg.scala 27:20]
  wire  _T_9392 = _T_4680 & ic_tag_valid_out_1_9; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9637 = _T_9636 | _T_9392; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_10; // @[Reg.scala 27:20]
  wire  _T_9394 = _T_4681 & ic_tag_valid_out_1_10; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9638 = _T_9637 | _T_9394; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_11; // @[Reg.scala 27:20]
  wire  _T_9396 = _T_4682 & ic_tag_valid_out_1_11; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9639 = _T_9638 | _T_9396; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_12; // @[Reg.scala 27:20]
  wire  _T_9398 = _T_4683 & ic_tag_valid_out_1_12; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9640 = _T_9639 | _T_9398; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_13; // @[Reg.scala 27:20]
  wire  _T_9400 = _T_4684 & ic_tag_valid_out_1_13; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9641 = _T_9640 | _T_9400; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_14; // @[Reg.scala 27:20]
  wire  _T_9402 = _T_4685 & ic_tag_valid_out_1_14; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9642 = _T_9641 | _T_9402; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_15; // @[Reg.scala 27:20]
  wire  _T_9404 = _T_4686 & ic_tag_valid_out_1_15; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9643 = _T_9642 | _T_9404; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_16; // @[Reg.scala 27:20]
  wire  _T_9406 = _T_4687 & ic_tag_valid_out_1_16; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9644 = _T_9643 | _T_9406; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_17; // @[Reg.scala 27:20]
  wire  _T_9408 = _T_4688 & ic_tag_valid_out_1_17; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9645 = _T_9644 | _T_9408; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_18; // @[Reg.scala 27:20]
  wire  _T_9410 = _T_4689 & ic_tag_valid_out_1_18; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9646 = _T_9645 | _T_9410; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_19; // @[Reg.scala 27:20]
  wire  _T_9412 = _T_4690 & ic_tag_valid_out_1_19; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9647 = _T_9646 | _T_9412; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_20; // @[Reg.scala 27:20]
  wire  _T_9414 = _T_4691 & ic_tag_valid_out_1_20; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9648 = _T_9647 | _T_9414; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_21; // @[Reg.scala 27:20]
  wire  _T_9416 = _T_4692 & ic_tag_valid_out_1_21; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9649 = _T_9648 | _T_9416; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_22; // @[Reg.scala 27:20]
  wire  _T_9418 = _T_4693 & ic_tag_valid_out_1_22; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9650 = _T_9649 | _T_9418; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_23; // @[Reg.scala 27:20]
  wire  _T_9420 = _T_4694 & ic_tag_valid_out_1_23; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9651 = _T_9650 | _T_9420; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_24; // @[Reg.scala 27:20]
  wire  _T_9422 = _T_4695 & ic_tag_valid_out_1_24; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9652 = _T_9651 | _T_9422; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_25; // @[Reg.scala 27:20]
  wire  _T_9424 = _T_4696 & ic_tag_valid_out_1_25; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9653 = _T_9652 | _T_9424; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_26; // @[Reg.scala 27:20]
  wire  _T_9426 = _T_4697 & ic_tag_valid_out_1_26; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9654 = _T_9653 | _T_9426; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_27; // @[Reg.scala 27:20]
  wire  _T_9428 = _T_4698 & ic_tag_valid_out_1_27; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9655 = _T_9654 | _T_9428; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_28; // @[Reg.scala 27:20]
  wire  _T_9430 = _T_4699 & ic_tag_valid_out_1_28; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9656 = _T_9655 | _T_9430; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_29; // @[Reg.scala 27:20]
  wire  _T_9432 = _T_4700 & ic_tag_valid_out_1_29; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9657 = _T_9656 | _T_9432; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_30; // @[Reg.scala 27:20]
  wire  _T_9434 = _T_4701 & ic_tag_valid_out_1_30; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9658 = _T_9657 | _T_9434; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_31; // @[Reg.scala 27:20]
  wire  _T_9436 = _T_4702 & ic_tag_valid_out_1_31; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9659 = _T_9658 | _T_9436; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_32; // @[Reg.scala 27:20]
  wire  _T_9438 = _T_4703 & ic_tag_valid_out_1_32; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9660 = _T_9659 | _T_9438; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_33; // @[Reg.scala 27:20]
  wire  _T_9440 = _T_4704 & ic_tag_valid_out_1_33; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9661 = _T_9660 | _T_9440; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_34; // @[Reg.scala 27:20]
  wire  _T_9442 = _T_4705 & ic_tag_valid_out_1_34; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9662 = _T_9661 | _T_9442; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_35; // @[Reg.scala 27:20]
  wire  _T_9444 = _T_4706 & ic_tag_valid_out_1_35; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9663 = _T_9662 | _T_9444; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_36; // @[Reg.scala 27:20]
  wire  _T_9446 = _T_4707 & ic_tag_valid_out_1_36; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9664 = _T_9663 | _T_9446; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_37; // @[Reg.scala 27:20]
  wire  _T_9448 = _T_4708 & ic_tag_valid_out_1_37; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9665 = _T_9664 | _T_9448; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_38; // @[Reg.scala 27:20]
  wire  _T_9450 = _T_4709 & ic_tag_valid_out_1_38; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9666 = _T_9665 | _T_9450; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_39; // @[Reg.scala 27:20]
  wire  _T_9452 = _T_4710 & ic_tag_valid_out_1_39; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9667 = _T_9666 | _T_9452; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_40; // @[Reg.scala 27:20]
  wire  _T_9454 = _T_4711 & ic_tag_valid_out_1_40; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9668 = _T_9667 | _T_9454; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_41; // @[Reg.scala 27:20]
  wire  _T_9456 = _T_4712 & ic_tag_valid_out_1_41; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9669 = _T_9668 | _T_9456; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_42; // @[Reg.scala 27:20]
  wire  _T_9458 = _T_4713 & ic_tag_valid_out_1_42; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9670 = _T_9669 | _T_9458; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_43; // @[Reg.scala 27:20]
  wire  _T_9460 = _T_4714 & ic_tag_valid_out_1_43; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9671 = _T_9670 | _T_9460; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_44; // @[Reg.scala 27:20]
  wire  _T_9462 = _T_4715 & ic_tag_valid_out_1_44; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9672 = _T_9671 | _T_9462; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_45; // @[Reg.scala 27:20]
  wire  _T_9464 = _T_4716 & ic_tag_valid_out_1_45; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9673 = _T_9672 | _T_9464; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_46; // @[Reg.scala 27:20]
  wire  _T_9466 = _T_4717 & ic_tag_valid_out_1_46; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9674 = _T_9673 | _T_9466; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_47; // @[Reg.scala 27:20]
  wire  _T_9468 = _T_4718 & ic_tag_valid_out_1_47; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9675 = _T_9674 | _T_9468; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_48; // @[Reg.scala 27:20]
  wire  _T_9470 = _T_4719 & ic_tag_valid_out_1_48; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9676 = _T_9675 | _T_9470; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_49; // @[Reg.scala 27:20]
  wire  _T_9472 = _T_4720 & ic_tag_valid_out_1_49; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9677 = _T_9676 | _T_9472; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_50; // @[Reg.scala 27:20]
  wire  _T_9474 = _T_4721 & ic_tag_valid_out_1_50; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9678 = _T_9677 | _T_9474; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_51; // @[Reg.scala 27:20]
  wire  _T_9476 = _T_4722 & ic_tag_valid_out_1_51; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9679 = _T_9678 | _T_9476; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_52; // @[Reg.scala 27:20]
  wire  _T_9478 = _T_4723 & ic_tag_valid_out_1_52; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9680 = _T_9679 | _T_9478; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_53; // @[Reg.scala 27:20]
  wire  _T_9480 = _T_4724 & ic_tag_valid_out_1_53; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9681 = _T_9680 | _T_9480; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_54; // @[Reg.scala 27:20]
  wire  _T_9482 = _T_4725 & ic_tag_valid_out_1_54; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9682 = _T_9681 | _T_9482; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_55; // @[Reg.scala 27:20]
  wire  _T_9484 = _T_4726 & ic_tag_valid_out_1_55; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9683 = _T_9682 | _T_9484; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_56; // @[Reg.scala 27:20]
  wire  _T_9486 = _T_4727 & ic_tag_valid_out_1_56; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9684 = _T_9683 | _T_9486; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_57; // @[Reg.scala 27:20]
  wire  _T_9488 = _T_4728 & ic_tag_valid_out_1_57; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9685 = _T_9684 | _T_9488; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_58; // @[Reg.scala 27:20]
  wire  _T_9490 = _T_4729 & ic_tag_valid_out_1_58; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9686 = _T_9685 | _T_9490; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_59; // @[Reg.scala 27:20]
  wire  _T_9492 = _T_4730 & ic_tag_valid_out_1_59; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9687 = _T_9686 | _T_9492; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_60; // @[Reg.scala 27:20]
  wire  _T_9494 = _T_4731 & ic_tag_valid_out_1_60; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9688 = _T_9687 | _T_9494; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_61; // @[Reg.scala 27:20]
  wire  _T_9496 = _T_4732 & ic_tag_valid_out_1_61; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9689 = _T_9688 | _T_9496; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_62; // @[Reg.scala 27:20]
  wire  _T_9498 = _T_4733 & ic_tag_valid_out_1_62; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9690 = _T_9689 | _T_9498; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_63; // @[Reg.scala 27:20]
  wire  _T_9500 = _T_4734 & ic_tag_valid_out_1_63; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9691 = _T_9690 | _T_9500; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_64; // @[Reg.scala 27:20]
  wire  _T_9502 = _T_4735 & ic_tag_valid_out_1_64; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9692 = _T_9691 | _T_9502; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_65; // @[Reg.scala 27:20]
  wire  _T_9504 = _T_4736 & ic_tag_valid_out_1_65; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9693 = _T_9692 | _T_9504; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_66; // @[Reg.scala 27:20]
  wire  _T_9506 = _T_4737 & ic_tag_valid_out_1_66; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9694 = _T_9693 | _T_9506; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_67; // @[Reg.scala 27:20]
  wire  _T_9508 = _T_4738 & ic_tag_valid_out_1_67; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9695 = _T_9694 | _T_9508; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_68; // @[Reg.scala 27:20]
  wire  _T_9510 = _T_4739 & ic_tag_valid_out_1_68; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9696 = _T_9695 | _T_9510; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_69; // @[Reg.scala 27:20]
  wire  _T_9512 = _T_4740 & ic_tag_valid_out_1_69; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9697 = _T_9696 | _T_9512; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_70; // @[Reg.scala 27:20]
  wire  _T_9514 = _T_4741 & ic_tag_valid_out_1_70; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9698 = _T_9697 | _T_9514; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_71; // @[Reg.scala 27:20]
  wire  _T_9516 = _T_4742 & ic_tag_valid_out_1_71; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9699 = _T_9698 | _T_9516; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_72; // @[Reg.scala 27:20]
  wire  _T_9518 = _T_4743 & ic_tag_valid_out_1_72; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9700 = _T_9699 | _T_9518; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_73; // @[Reg.scala 27:20]
  wire  _T_9520 = _T_4744 & ic_tag_valid_out_1_73; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9701 = _T_9700 | _T_9520; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_74; // @[Reg.scala 27:20]
  wire  _T_9522 = _T_4745 & ic_tag_valid_out_1_74; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9702 = _T_9701 | _T_9522; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_75; // @[Reg.scala 27:20]
  wire  _T_9524 = _T_4746 & ic_tag_valid_out_1_75; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9703 = _T_9702 | _T_9524; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_76; // @[Reg.scala 27:20]
  wire  _T_9526 = _T_4747 & ic_tag_valid_out_1_76; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9704 = _T_9703 | _T_9526; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_77; // @[Reg.scala 27:20]
  wire  _T_9528 = _T_4748 & ic_tag_valid_out_1_77; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9705 = _T_9704 | _T_9528; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_78; // @[Reg.scala 27:20]
  wire  _T_9530 = _T_4749 & ic_tag_valid_out_1_78; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9706 = _T_9705 | _T_9530; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_79; // @[Reg.scala 27:20]
  wire  _T_9532 = _T_4750 & ic_tag_valid_out_1_79; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9707 = _T_9706 | _T_9532; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_80; // @[Reg.scala 27:20]
  wire  _T_9534 = _T_4751 & ic_tag_valid_out_1_80; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9708 = _T_9707 | _T_9534; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_81; // @[Reg.scala 27:20]
  wire  _T_9536 = _T_4752 & ic_tag_valid_out_1_81; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9709 = _T_9708 | _T_9536; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_82; // @[Reg.scala 27:20]
  wire  _T_9538 = _T_4753 & ic_tag_valid_out_1_82; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9710 = _T_9709 | _T_9538; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_83; // @[Reg.scala 27:20]
  wire  _T_9540 = _T_4754 & ic_tag_valid_out_1_83; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9711 = _T_9710 | _T_9540; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_84; // @[Reg.scala 27:20]
  wire  _T_9542 = _T_4755 & ic_tag_valid_out_1_84; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9712 = _T_9711 | _T_9542; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_85; // @[Reg.scala 27:20]
  wire  _T_9544 = _T_4756 & ic_tag_valid_out_1_85; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9713 = _T_9712 | _T_9544; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_86; // @[Reg.scala 27:20]
  wire  _T_9546 = _T_4757 & ic_tag_valid_out_1_86; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9714 = _T_9713 | _T_9546; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_87; // @[Reg.scala 27:20]
  wire  _T_9548 = _T_4758 & ic_tag_valid_out_1_87; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9715 = _T_9714 | _T_9548; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_88; // @[Reg.scala 27:20]
  wire  _T_9550 = _T_4759 & ic_tag_valid_out_1_88; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9716 = _T_9715 | _T_9550; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_89; // @[Reg.scala 27:20]
  wire  _T_9552 = _T_4760 & ic_tag_valid_out_1_89; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9717 = _T_9716 | _T_9552; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_90; // @[Reg.scala 27:20]
  wire  _T_9554 = _T_4761 & ic_tag_valid_out_1_90; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9718 = _T_9717 | _T_9554; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_91; // @[Reg.scala 27:20]
  wire  _T_9556 = _T_4762 & ic_tag_valid_out_1_91; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9719 = _T_9718 | _T_9556; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_92; // @[Reg.scala 27:20]
  wire  _T_9558 = _T_4763 & ic_tag_valid_out_1_92; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9720 = _T_9719 | _T_9558; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_93; // @[Reg.scala 27:20]
  wire  _T_9560 = _T_4764 & ic_tag_valid_out_1_93; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9721 = _T_9720 | _T_9560; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_94; // @[Reg.scala 27:20]
  wire  _T_9562 = _T_4765 & ic_tag_valid_out_1_94; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9722 = _T_9721 | _T_9562; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_95; // @[Reg.scala 27:20]
  wire  _T_9564 = _T_4766 & ic_tag_valid_out_1_95; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9723 = _T_9722 | _T_9564; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_96; // @[Reg.scala 27:20]
  wire  _T_9566 = _T_4767 & ic_tag_valid_out_1_96; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9724 = _T_9723 | _T_9566; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_97; // @[Reg.scala 27:20]
  wire  _T_9568 = _T_4768 & ic_tag_valid_out_1_97; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9725 = _T_9724 | _T_9568; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_98; // @[Reg.scala 27:20]
  wire  _T_9570 = _T_4769 & ic_tag_valid_out_1_98; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9726 = _T_9725 | _T_9570; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_99; // @[Reg.scala 27:20]
  wire  _T_9572 = _T_4770 & ic_tag_valid_out_1_99; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9727 = _T_9726 | _T_9572; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_100; // @[Reg.scala 27:20]
  wire  _T_9574 = _T_4771 & ic_tag_valid_out_1_100; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9728 = _T_9727 | _T_9574; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_101; // @[Reg.scala 27:20]
  wire  _T_9576 = _T_4772 & ic_tag_valid_out_1_101; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9729 = _T_9728 | _T_9576; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_102; // @[Reg.scala 27:20]
  wire  _T_9578 = _T_4773 & ic_tag_valid_out_1_102; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9730 = _T_9729 | _T_9578; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_103; // @[Reg.scala 27:20]
  wire  _T_9580 = _T_4774 & ic_tag_valid_out_1_103; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9731 = _T_9730 | _T_9580; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_104; // @[Reg.scala 27:20]
  wire  _T_9582 = _T_4775 & ic_tag_valid_out_1_104; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9732 = _T_9731 | _T_9582; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_105; // @[Reg.scala 27:20]
  wire  _T_9584 = _T_4776 & ic_tag_valid_out_1_105; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9733 = _T_9732 | _T_9584; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_106; // @[Reg.scala 27:20]
  wire  _T_9586 = _T_4777 & ic_tag_valid_out_1_106; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9734 = _T_9733 | _T_9586; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_107; // @[Reg.scala 27:20]
  wire  _T_9588 = _T_4778 & ic_tag_valid_out_1_107; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9735 = _T_9734 | _T_9588; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_108; // @[Reg.scala 27:20]
  wire  _T_9590 = _T_4779 & ic_tag_valid_out_1_108; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9736 = _T_9735 | _T_9590; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_109; // @[Reg.scala 27:20]
  wire  _T_9592 = _T_4780 & ic_tag_valid_out_1_109; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9737 = _T_9736 | _T_9592; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_110; // @[Reg.scala 27:20]
  wire  _T_9594 = _T_4781 & ic_tag_valid_out_1_110; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9738 = _T_9737 | _T_9594; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_111; // @[Reg.scala 27:20]
  wire  _T_9596 = _T_4782 & ic_tag_valid_out_1_111; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9739 = _T_9738 | _T_9596; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_112; // @[Reg.scala 27:20]
  wire  _T_9598 = _T_4783 & ic_tag_valid_out_1_112; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9740 = _T_9739 | _T_9598; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_113; // @[Reg.scala 27:20]
  wire  _T_9600 = _T_4784 & ic_tag_valid_out_1_113; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9741 = _T_9740 | _T_9600; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_114; // @[Reg.scala 27:20]
  wire  _T_9602 = _T_4785 & ic_tag_valid_out_1_114; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9742 = _T_9741 | _T_9602; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_115; // @[Reg.scala 27:20]
  wire  _T_9604 = _T_4786 & ic_tag_valid_out_1_115; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9743 = _T_9742 | _T_9604; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_116; // @[Reg.scala 27:20]
  wire  _T_9606 = _T_4787 & ic_tag_valid_out_1_116; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9744 = _T_9743 | _T_9606; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_117; // @[Reg.scala 27:20]
  wire  _T_9608 = _T_4788 & ic_tag_valid_out_1_117; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9745 = _T_9744 | _T_9608; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_118; // @[Reg.scala 27:20]
  wire  _T_9610 = _T_4789 & ic_tag_valid_out_1_118; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9746 = _T_9745 | _T_9610; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_119; // @[Reg.scala 27:20]
  wire  _T_9612 = _T_4790 & ic_tag_valid_out_1_119; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9747 = _T_9746 | _T_9612; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_120; // @[Reg.scala 27:20]
  wire  _T_9614 = _T_4791 & ic_tag_valid_out_1_120; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9748 = _T_9747 | _T_9614; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_121; // @[Reg.scala 27:20]
  wire  _T_9616 = _T_4792 & ic_tag_valid_out_1_121; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9749 = _T_9748 | _T_9616; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_122; // @[Reg.scala 27:20]
  wire  _T_9618 = _T_4793 & ic_tag_valid_out_1_122; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9750 = _T_9749 | _T_9618; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_123; // @[Reg.scala 27:20]
  wire  _T_9620 = _T_4794 & ic_tag_valid_out_1_123; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9751 = _T_9750 | _T_9620; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_124; // @[Reg.scala 27:20]
  wire  _T_9622 = _T_4795 & ic_tag_valid_out_1_124; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9752 = _T_9751 | _T_9622; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_125; // @[Reg.scala 27:20]
  wire  _T_9624 = _T_4796 & ic_tag_valid_out_1_125; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9753 = _T_9752 | _T_9624; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_126; // @[Reg.scala 27:20]
  wire  _T_9626 = _T_4797 & ic_tag_valid_out_1_126; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9754 = _T_9753 | _T_9626; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_127; // @[Reg.scala 27:20]
  wire  _T_9628 = _T_4798 & ic_tag_valid_out_1_127; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9755 = _T_9754 | _T_9628; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_0; // @[Reg.scala 27:20]
  wire  _T_8991 = _T_4671 & ic_tag_valid_out_0_0; // @[ifu_mem_ctl.scala 696:10]
  reg  ic_tag_valid_out_0_1; // @[Reg.scala 27:20]
  wire  _T_8993 = _T_4672 & ic_tag_valid_out_0_1; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9246 = _T_8991 | _T_8993; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_2; // @[Reg.scala 27:20]
  wire  _T_8995 = _T_4673 & ic_tag_valid_out_0_2; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9247 = _T_9246 | _T_8995; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_3; // @[Reg.scala 27:20]
  wire  _T_8997 = _T_4674 & ic_tag_valid_out_0_3; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9248 = _T_9247 | _T_8997; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_4; // @[Reg.scala 27:20]
  wire  _T_8999 = _T_4675 & ic_tag_valid_out_0_4; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9249 = _T_9248 | _T_8999; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_5; // @[Reg.scala 27:20]
  wire  _T_9001 = _T_4676 & ic_tag_valid_out_0_5; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9250 = _T_9249 | _T_9001; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_6; // @[Reg.scala 27:20]
  wire  _T_9003 = _T_4677 & ic_tag_valid_out_0_6; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9251 = _T_9250 | _T_9003; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_7; // @[Reg.scala 27:20]
  wire  _T_9005 = _T_4678 & ic_tag_valid_out_0_7; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9252 = _T_9251 | _T_9005; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_8; // @[Reg.scala 27:20]
  wire  _T_9007 = _T_4679 & ic_tag_valid_out_0_8; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9253 = _T_9252 | _T_9007; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_9; // @[Reg.scala 27:20]
  wire  _T_9009 = _T_4680 & ic_tag_valid_out_0_9; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9254 = _T_9253 | _T_9009; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_10; // @[Reg.scala 27:20]
  wire  _T_9011 = _T_4681 & ic_tag_valid_out_0_10; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9255 = _T_9254 | _T_9011; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_11; // @[Reg.scala 27:20]
  wire  _T_9013 = _T_4682 & ic_tag_valid_out_0_11; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9256 = _T_9255 | _T_9013; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_12; // @[Reg.scala 27:20]
  wire  _T_9015 = _T_4683 & ic_tag_valid_out_0_12; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9257 = _T_9256 | _T_9015; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_13; // @[Reg.scala 27:20]
  wire  _T_9017 = _T_4684 & ic_tag_valid_out_0_13; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9258 = _T_9257 | _T_9017; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_14; // @[Reg.scala 27:20]
  wire  _T_9019 = _T_4685 & ic_tag_valid_out_0_14; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9259 = _T_9258 | _T_9019; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_15; // @[Reg.scala 27:20]
  wire  _T_9021 = _T_4686 & ic_tag_valid_out_0_15; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9260 = _T_9259 | _T_9021; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_16; // @[Reg.scala 27:20]
  wire  _T_9023 = _T_4687 & ic_tag_valid_out_0_16; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9261 = _T_9260 | _T_9023; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_17; // @[Reg.scala 27:20]
  wire  _T_9025 = _T_4688 & ic_tag_valid_out_0_17; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9262 = _T_9261 | _T_9025; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_18; // @[Reg.scala 27:20]
  wire  _T_9027 = _T_4689 & ic_tag_valid_out_0_18; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9263 = _T_9262 | _T_9027; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_19; // @[Reg.scala 27:20]
  wire  _T_9029 = _T_4690 & ic_tag_valid_out_0_19; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9264 = _T_9263 | _T_9029; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_20; // @[Reg.scala 27:20]
  wire  _T_9031 = _T_4691 & ic_tag_valid_out_0_20; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9265 = _T_9264 | _T_9031; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_21; // @[Reg.scala 27:20]
  wire  _T_9033 = _T_4692 & ic_tag_valid_out_0_21; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9266 = _T_9265 | _T_9033; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_22; // @[Reg.scala 27:20]
  wire  _T_9035 = _T_4693 & ic_tag_valid_out_0_22; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9267 = _T_9266 | _T_9035; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_23; // @[Reg.scala 27:20]
  wire  _T_9037 = _T_4694 & ic_tag_valid_out_0_23; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9268 = _T_9267 | _T_9037; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_24; // @[Reg.scala 27:20]
  wire  _T_9039 = _T_4695 & ic_tag_valid_out_0_24; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9269 = _T_9268 | _T_9039; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_25; // @[Reg.scala 27:20]
  wire  _T_9041 = _T_4696 & ic_tag_valid_out_0_25; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9270 = _T_9269 | _T_9041; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_26; // @[Reg.scala 27:20]
  wire  _T_9043 = _T_4697 & ic_tag_valid_out_0_26; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9271 = _T_9270 | _T_9043; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_27; // @[Reg.scala 27:20]
  wire  _T_9045 = _T_4698 & ic_tag_valid_out_0_27; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9272 = _T_9271 | _T_9045; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_28; // @[Reg.scala 27:20]
  wire  _T_9047 = _T_4699 & ic_tag_valid_out_0_28; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9273 = _T_9272 | _T_9047; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_29; // @[Reg.scala 27:20]
  wire  _T_9049 = _T_4700 & ic_tag_valid_out_0_29; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9274 = _T_9273 | _T_9049; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_30; // @[Reg.scala 27:20]
  wire  _T_9051 = _T_4701 & ic_tag_valid_out_0_30; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9275 = _T_9274 | _T_9051; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_31; // @[Reg.scala 27:20]
  wire  _T_9053 = _T_4702 & ic_tag_valid_out_0_31; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9276 = _T_9275 | _T_9053; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_32; // @[Reg.scala 27:20]
  wire  _T_9055 = _T_4703 & ic_tag_valid_out_0_32; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9277 = _T_9276 | _T_9055; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_33; // @[Reg.scala 27:20]
  wire  _T_9057 = _T_4704 & ic_tag_valid_out_0_33; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9278 = _T_9277 | _T_9057; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_34; // @[Reg.scala 27:20]
  wire  _T_9059 = _T_4705 & ic_tag_valid_out_0_34; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9279 = _T_9278 | _T_9059; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_35; // @[Reg.scala 27:20]
  wire  _T_9061 = _T_4706 & ic_tag_valid_out_0_35; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9280 = _T_9279 | _T_9061; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_36; // @[Reg.scala 27:20]
  wire  _T_9063 = _T_4707 & ic_tag_valid_out_0_36; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9281 = _T_9280 | _T_9063; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_37; // @[Reg.scala 27:20]
  wire  _T_9065 = _T_4708 & ic_tag_valid_out_0_37; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9282 = _T_9281 | _T_9065; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_38; // @[Reg.scala 27:20]
  wire  _T_9067 = _T_4709 & ic_tag_valid_out_0_38; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9283 = _T_9282 | _T_9067; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_39; // @[Reg.scala 27:20]
  wire  _T_9069 = _T_4710 & ic_tag_valid_out_0_39; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9284 = _T_9283 | _T_9069; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_40; // @[Reg.scala 27:20]
  wire  _T_9071 = _T_4711 & ic_tag_valid_out_0_40; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9285 = _T_9284 | _T_9071; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_41; // @[Reg.scala 27:20]
  wire  _T_9073 = _T_4712 & ic_tag_valid_out_0_41; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9286 = _T_9285 | _T_9073; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_42; // @[Reg.scala 27:20]
  wire  _T_9075 = _T_4713 & ic_tag_valid_out_0_42; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9287 = _T_9286 | _T_9075; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_43; // @[Reg.scala 27:20]
  wire  _T_9077 = _T_4714 & ic_tag_valid_out_0_43; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9288 = _T_9287 | _T_9077; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_44; // @[Reg.scala 27:20]
  wire  _T_9079 = _T_4715 & ic_tag_valid_out_0_44; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9289 = _T_9288 | _T_9079; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_45; // @[Reg.scala 27:20]
  wire  _T_9081 = _T_4716 & ic_tag_valid_out_0_45; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9290 = _T_9289 | _T_9081; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_46; // @[Reg.scala 27:20]
  wire  _T_9083 = _T_4717 & ic_tag_valid_out_0_46; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9291 = _T_9290 | _T_9083; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_47; // @[Reg.scala 27:20]
  wire  _T_9085 = _T_4718 & ic_tag_valid_out_0_47; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9292 = _T_9291 | _T_9085; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_48; // @[Reg.scala 27:20]
  wire  _T_9087 = _T_4719 & ic_tag_valid_out_0_48; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9293 = _T_9292 | _T_9087; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_49; // @[Reg.scala 27:20]
  wire  _T_9089 = _T_4720 & ic_tag_valid_out_0_49; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9294 = _T_9293 | _T_9089; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_50; // @[Reg.scala 27:20]
  wire  _T_9091 = _T_4721 & ic_tag_valid_out_0_50; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9295 = _T_9294 | _T_9091; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_51; // @[Reg.scala 27:20]
  wire  _T_9093 = _T_4722 & ic_tag_valid_out_0_51; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9296 = _T_9295 | _T_9093; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_52; // @[Reg.scala 27:20]
  wire  _T_9095 = _T_4723 & ic_tag_valid_out_0_52; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9297 = _T_9296 | _T_9095; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_53; // @[Reg.scala 27:20]
  wire  _T_9097 = _T_4724 & ic_tag_valid_out_0_53; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9298 = _T_9297 | _T_9097; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_54; // @[Reg.scala 27:20]
  wire  _T_9099 = _T_4725 & ic_tag_valid_out_0_54; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9299 = _T_9298 | _T_9099; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_55; // @[Reg.scala 27:20]
  wire  _T_9101 = _T_4726 & ic_tag_valid_out_0_55; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9300 = _T_9299 | _T_9101; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_56; // @[Reg.scala 27:20]
  wire  _T_9103 = _T_4727 & ic_tag_valid_out_0_56; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9301 = _T_9300 | _T_9103; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_57; // @[Reg.scala 27:20]
  wire  _T_9105 = _T_4728 & ic_tag_valid_out_0_57; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9302 = _T_9301 | _T_9105; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_58; // @[Reg.scala 27:20]
  wire  _T_9107 = _T_4729 & ic_tag_valid_out_0_58; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9303 = _T_9302 | _T_9107; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_59; // @[Reg.scala 27:20]
  wire  _T_9109 = _T_4730 & ic_tag_valid_out_0_59; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9304 = _T_9303 | _T_9109; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_60; // @[Reg.scala 27:20]
  wire  _T_9111 = _T_4731 & ic_tag_valid_out_0_60; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9305 = _T_9304 | _T_9111; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_61; // @[Reg.scala 27:20]
  wire  _T_9113 = _T_4732 & ic_tag_valid_out_0_61; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9306 = _T_9305 | _T_9113; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_62; // @[Reg.scala 27:20]
  wire  _T_9115 = _T_4733 & ic_tag_valid_out_0_62; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9307 = _T_9306 | _T_9115; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_63; // @[Reg.scala 27:20]
  wire  _T_9117 = _T_4734 & ic_tag_valid_out_0_63; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9308 = _T_9307 | _T_9117; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_64; // @[Reg.scala 27:20]
  wire  _T_9119 = _T_4735 & ic_tag_valid_out_0_64; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9309 = _T_9308 | _T_9119; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_65; // @[Reg.scala 27:20]
  wire  _T_9121 = _T_4736 & ic_tag_valid_out_0_65; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9310 = _T_9309 | _T_9121; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_66; // @[Reg.scala 27:20]
  wire  _T_9123 = _T_4737 & ic_tag_valid_out_0_66; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9311 = _T_9310 | _T_9123; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_67; // @[Reg.scala 27:20]
  wire  _T_9125 = _T_4738 & ic_tag_valid_out_0_67; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9312 = _T_9311 | _T_9125; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_68; // @[Reg.scala 27:20]
  wire  _T_9127 = _T_4739 & ic_tag_valid_out_0_68; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9313 = _T_9312 | _T_9127; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_69; // @[Reg.scala 27:20]
  wire  _T_9129 = _T_4740 & ic_tag_valid_out_0_69; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9314 = _T_9313 | _T_9129; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_70; // @[Reg.scala 27:20]
  wire  _T_9131 = _T_4741 & ic_tag_valid_out_0_70; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9315 = _T_9314 | _T_9131; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_71; // @[Reg.scala 27:20]
  wire  _T_9133 = _T_4742 & ic_tag_valid_out_0_71; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9316 = _T_9315 | _T_9133; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_72; // @[Reg.scala 27:20]
  wire  _T_9135 = _T_4743 & ic_tag_valid_out_0_72; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9317 = _T_9316 | _T_9135; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_73; // @[Reg.scala 27:20]
  wire  _T_9137 = _T_4744 & ic_tag_valid_out_0_73; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9318 = _T_9317 | _T_9137; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_74; // @[Reg.scala 27:20]
  wire  _T_9139 = _T_4745 & ic_tag_valid_out_0_74; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9319 = _T_9318 | _T_9139; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_75; // @[Reg.scala 27:20]
  wire  _T_9141 = _T_4746 & ic_tag_valid_out_0_75; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9320 = _T_9319 | _T_9141; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_76; // @[Reg.scala 27:20]
  wire  _T_9143 = _T_4747 & ic_tag_valid_out_0_76; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9321 = _T_9320 | _T_9143; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_77; // @[Reg.scala 27:20]
  wire  _T_9145 = _T_4748 & ic_tag_valid_out_0_77; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9322 = _T_9321 | _T_9145; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_78; // @[Reg.scala 27:20]
  wire  _T_9147 = _T_4749 & ic_tag_valid_out_0_78; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9323 = _T_9322 | _T_9147; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_79; // @[Reg.scala 27:20]
  wire  _T_9149 = _T_4750 & ic_tag_valid_out_0_79; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9324 = _T_9323 | _T_9149; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_80; // @[Reg.scala 27:20]
  wire  _T_9151 = _T_4751 & ic_tag_valid_out_0_80; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9325 = _T_9324 | _T_9151; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_81; // @[Reg.scala 27:20]
  wire  _T_9153 = _T_4752 & ic_tag_valid_out_0_81; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9326 = _T_9325 | _T_9153; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_82; // @[Reg.scala 27:20]
  wire  _T_9155 = _T_4753 & ic_tag_valid_out_0_82; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9327 = _T_9326 | _T_9155; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_83; // @[Reg.scala 27:20]
  wire  _T_9157 = _T_4754 & ic_tag_valid_out_0_83; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9328 = _T_9327 | _T_9157; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_84; // @[Reg.scala 27:20]
  wire  _T_9159 = _T_4755 & ic_tag_valid_out_0_84; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9329 = _T_9328 | _T_9159; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_85; // @[Reg.scala 27:20]
  wire  _T_9161 = _T_4756 & ic_tag_valid_out_0_85; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9330 = _T_9329 | _T_9161; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_86; // @[Reg.scala 27:20]
  wire  _T_9163 = _T_4757 & ic_tag_valid_out_0_86; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9331 = _T_9330 | _T_9163; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_87; // @[Reg.scala 27:20]
  wire  _T_9165 = _T_4758 & ic_tag_valid_out_0_87; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9332 = _T_9331 | _T_9165; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_88; // @[Reg.scala 27:20]
  wire  _T_9167 = _T_4759 & ic_tag_valid_out_0_88; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9333 = _T_9332 | _T_9167; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_89; // @[Reg.scala 27:20]
  wire  _T_9169 = _T_4760 & ic_tag_valid_out_0_89; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9334 = _T_9333 | _T_9169; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_90; // @[Reg.scala 27:20]
  wire  _T_9171 = _T_4761 & ic_tag_valid_out_0_90; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9335 = _T_9334 | _T_9171; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_91; // @[Reg.scala 27:20]
  wire  _T_9173 = _T_4762 & ic_tag_valid_out_0_91; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9336 = _T_9335 | _T_9173; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_92; // @[Reg.scala 27:20]
  wire  _T_9175 = _T_4763 & ic_tag_valid_out_0_92; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9337 = _T_9336 | _T_9175; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_93; // @[Reg.scala 27:20]
  wire  _T_9177 = _T_4764 & ic_tag_valid_out_0_93; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9338 = _T_9337 | _T_9177; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_94; // @[Reg.scala 27:20]
  wire  _T_9179 = _T_4765 & ic_tag_valid_out_0_94; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9339 = _T_9338 | _T_9179; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_95; // @[Reg.scala 27:20]
  wire  _T_9181 = _T_4766 & ic_tag_valid_out_0_95; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9340 = _T_9339 | _T_9181; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_96; // @[Reg.scala 27:20]
  wire  _T_9183 = _T_4767 & ic_tag_valid_out_0_96; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9341 = _T_9340 | _T_9183; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_97; // @[Reg.scala 27:20]
  wire  _T_9185 = _T_4768 & ic_tag_valid_out_0_97; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9342 = _T_9341 | _T_9185; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_98; // @[Reg.scala 27:20]
  wire  _T_9187 = _T_4769 & ic_tag_valid_out_0_98; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9343 = _T_9342 | _T_9187; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_99; // @[Reg.scala 27:20]
  wire  _T_9189 = _T_4770 & ic_tag_valid_out_0_99; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9344 = _T_9343 | _T_9189; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_100; // @[Reg.scala 27:20]
  wire  _T_9191 = _T_4771 & ic_tag_valid_out_0_100; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9345 = _T_9344 | _T_9191; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_101; // @[Reg.scala 27:20]
  wire  _T_9193 = _T_4772 & ic_tag_valid_out_0_101; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9346 = _T_9345 | _T_9193; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_102; // @[Reg.scala 27:20]
  wire  _T_9195 = _T_4773 & ic_tag_valid_out_0_102; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9347 = _T_9346 | _T_9195; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_103; // @[Reg.scala 27:20]
  wire  _T_9197 = _T_4774 & ic_tag_valid_out_0_103; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9348 = _T_9347 | _T_9197; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_104; // @[Reg.scala 27:20]
  wire  _T_9199 = _T_4775 & ic_tag_valid_out_0_104; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9349 = _T_9348 | _T_9199; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_105; // @[Reg.scala 27:20]
  wire  _T_9201 = _T_4776 & ic_tag_valid_out_0_105; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9350 = _T_9349 | _T_9201; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_106; // @[Reg.scala 27:20]
  wire  _T_9203 = _T_4777 & ic_tag_valid_out_0_106; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9351 = _T_9350 | _T_9203; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_107; // @[Reg.scala 27:20]
  wire  _T_9205 = _T_4778 & ic_tag_valid_out_0_107; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9352 = _T_9351 | _T_9205; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_108; // @[Reg.scala 27:20]
  wire  _T_9207 = _T_4779 & ic_tag_valid_out_0_108; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9353 = _T_9352 | _T_9207; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_109; // @[Reg.scala 27:20]
  wire  _T_9209 = _T_4780 & ic_tag_valid_out_0_109; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9354 = _T_9353 | _T_9209; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_110; // @[Reg.scala 27:20]
  wire  _T_9211 = _T_4781 & ic_tag_valid_out_0_110; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9355 = _T_9354 | _T_9211; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_111; // @[Reg.scala 27:20]
  wire  _T_9213 = _T_4782 & ic_tag_valid_out_0_111; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9356 = _T_9355 | _T_9213; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_112; // @[Reg.scala 27:20]
  wire  _T_9215 = _T_4783 & ic_tag_valid_out_0_112; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9357 = _T_9356 | _T_9215; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_113; // @[Reg.scala 27:20]
  wire  _T_9217 = _T_4784 & ic_tag_valid_out_0_113; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9358 = _T_9357 | _T_9217; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_114; // @[Reg.scala 27:20]
  wire  _T_9219 = _T_4785 & ic_tag_valid_out_0_114; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9359 = _T_9358 | _T_9219; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_115; // @[Reg.scala 27:20]
  wire  _T_9221 = _T_4786 & ic_tag_valid_out_0_115; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9360 = _T_9359 | _T_9221; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_116; // @[Reg.scala 27:20]
  wire  _T_9223 = _T_4787 & ic_tag_valid_out_0_116; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9361 = _T_9360 | _T_9223; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_117; // @[Reg.scala 27:20]
  wire  _T_9225 = _T_4788 & ic_tag_valid_out_0_117; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9362 = _T_9361 | _T_9225; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_118; // @[Reg.scala 27:20]
  wire  _T_9227 = _T_4789 & ic_tag_valid_out_0_118; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9363 = _T_9362 | _T_9227; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_119; // @[Reg.scala 27:20]
  wire  _T_9229 = _T_4790 & ic_tag_valid_out_0_119; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9364 = _T_9363 | _T_9229; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_120; // @[Reg.scala 27:20]
  wire  _T_9231 = _T_4791 & ic_tag_valid_out_0_120; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9365 = _T_9364 | _T_9231; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_121; // @[Reg.scala 27:20]
  wire  _T_9233 = _T_4792 & ic_tag_valid_out_0_121; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9366 = _T_9365 | _T_9233; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_122; // @[Reg.scala 27:20]
  wire  _T_9235 = _T_4793 & ic_tag_valid_out_0_122; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9367 = _T_9366 | _T_9235; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_123; // @[Reg.scala 27:20]
  wire  _T_9237 = _T_4794 & ic_tag_valid_out_0_123; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9368 = _T_9367 | _T_9237; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_124; // @[Reg.scala 27:20]
  wire  _T_9239 = _T_4795 & ic_tag_valid_out_0_124; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9369 = _T_9368 | _T_9239; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_125; // @[Reg.scala 27:20]
  wire  _T_9241 = _T_4796 & ic_tag_valid_out_0_125; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9370 = _T_9369 | _T_9241; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_126; // @[Reg.scala 27:20]
  wire  _T_9243 = _T_4797 & ic_tag_valid_out_0_126; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9371 = _T_9370 | _T_9243; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_127; // @[Reg.scala 27:20]
  wire  _T_9245 = _T_4798 & ic_tag_valid_out_0_127; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9372 = _T_9371 | _T_9245; // @[ifu_mem_ctl.scala 696:91]
  wire [1:0] ic_tag_valid_unq = {_T_9755,_T_9372}; // @[Cat.scala 29:58]
  reg [1:0] ic_debug_way_ff; // @[ifu_mem_ctl.scala 767:53]
  reg  ic_debug_rd_en_ff; // @[ifu_mem_ctl.scala 769:54]
  wire [1:0] _T_9795 = ic_debug_rd_en_ff ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [1:0] _T_9796 = ic_debug_way_ff & _T_9795; // @[ifu_mem_ctl.scala 750:67]
  wire [1:0] _T_9797 = ic_tag_valid_unq & _T_9796; // @[ifu_mem_ctl.scala 750:48]
  wire  ic_debug_tag_val_rd_out = |_T_9797; // @[ifu_mem_ctl.scala 750:115]
  wire [70:0] _T_1211 = {2'h0,io_ic_tag_debug_rd_data[25:21],32'h0,io_ic_tag_debug_rd_data[20:0],6'h0,way_status,3'h0,ic_debug_tag_val_rd_out}; // @[Cat.scala 29:58]
  reg [70:0] _T_1212; // @[ifu_mem_ctl.scala 263:76]
  wire  _T_1250 = ~ifu_byp_data_err_new; // @[ifu_mem_ctl.scala 279:98]
  wire  sel_byp_data = _T_1254 & _T_1250; // @[ifu_mem_ctl.scala 279:96]
  wire  _T_1257 = sel_byp_data | fetch_req_iccm_f; // @[ifu_mem_ctl.scala 284:46]
  wire  final_data_sel1_0 = _T_1257 | sel_ic_data; // @[ifu_mem_ctl.scala 284:62]
  wire [63:0] _T_1263 = final_data_sel1_0 ? 64'hffffffffffffffff : 64'h0; // @[Bitwise.scala 72:12]
  wire [63:0] ic_final_data = _T_1263 & io_ic_rd_data; // @[ifu_mem_ctl.scala 288:92]
  wire [63:0] _T_1265 = fetch_req_iccm_f ? 64'hffffffffffffffff : 64'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_1266 = _T_1265 & io_iccm_rd_data; // @[ifu_mem_ctl.scala 292:69]
  wire [79:0] ic_premux_data_temp = {{16'd0}, _T_1266}; // @[ifu_mem_ctl.scala 292:88]
  wire  fetch_req_f_qual = io_ic_hit_f & _T_319; // @[ifu_mem_ctl.scala 299:38]
  reg  ifc_region_acc_fault_memory_f; // @[ifu_mem_ctl.scala 783:66]
  wire [1:0] _T_1277 = ifc_region_acc_fault_memory_f ? 2'h3 : 2'h0; // @[ifu_mem_ctl.scala 304:10]
  wire [1:0] _T_1278 = ifc_region_acc_fault_f ? 2'h2 : _T_1277; // @[ifu_mem_ctl.scala 303:8]
  wire  _T_1280 = fetch_req_f_qual & io_ifu_bp_inst_mask_f; // @[ifu_mem_ctl.scala 305:45]
  wire  _T_1282 = byp_fetch_index == 5'h1f; // @[ifu_mem_ctl.scala 305:80]
  wire  _T_1283 = ~_T_1282; // @[ifu_mem_ctl.scala 305:71]
  wire  _T_1284 = _T_1280 & _T_1283; // @[ifu_mem_ctl.scala 305:69]
  wire  _T_1285 = err_stop_state != 2'h2; // @[ifu_mem_ctl.scala 305:131]
  wire  _T_1286 = _T_1284 & _T_1285; // @[ifu_mem_ctl.scala 305:114]
  wire [6:0] _T_1358 = {ic_miss_buff_data_valid_in_7,ic_miss_buff_data_valid_in_6,ic_miss_buff_data_valid_in_5,ic_miss_buff_data_valid_in_4,ic_miss_buff_data_valid_in_3,ic_miss_buff_data_valid_in_2,ic_miss_buff_data_valid_in_1}; // @[Cat.scala 29:58]
  wire  ic_miss_buff_data_error_in_0 = ic_miss_buff_data_error[0] & _T_1330; // @[ifu_mem_ctl.scala 324:32]
  wire  ic_miss_buff_data_error_in_1 = ic_miss_buff_data_error[1] & _T_1330; // @[ifu_mem_ctl.scala 324:32]
  wire  ic_miss_buff_data_error_in_2 = ic_miss_buff_data_error[2] & _T_1330; // @[ifu_mem_ctl.scala 324:32]
  wire  ic_miss_buff_data_error_in_3 = ic_miss_buff_data_error[3] & _T_1330; // @[ifu_mem_ctl.scala 324:32]
  wire  ic_miss_buff_data_error_in_4 = ic_miss_buff_data_error[4] & _T_1330; // @[ifu_mem_ctl.scala 324:32]
  wire  ic_miss_buff_data_error_in_5 = ic_miss_buff_data_error[5] & _T_1330; // @[ifu_mem_ctl.scala 324:32]
  wire  ic_miss_buff_data_error_in_6 = ic_miss_buff_data_error[6] & _T_1330; // @[ifu_mem_ctl.scala 324:32]
  wire  ic_miss_buff_data_error_in_7 = ic_miss_buff_data_error[7] & _T_1330; // @[ifu_mem_ctl.scala 324:32]
  wire [6:0] _T_1398 = {ic_miss_buff_data_error_in_7,ic_miss_buff_data_error_in_6,ic_miss_buff_data_error_in_5,ic_miss_buff_data_error_in_4,ic_miss_buff_data_error_in_3,ic_miss_buff_data_error_in_2,ic_miss_buff_data_error_in_1}; // @[Cat.scala 29:58]
  reg [6:0] perr_ic_index_ff; // @[Reg.scala 27:20]
  wire  _T_2500 = 3'h0 == perr_state; // @[Conditional.scala 37:30]
  wire  _T_2508 = _T_6 & _T_319; // @[ifu_mem_ctl.scala 405:82]
  wire  _T_2509 = _T_2508 | io_iccm_dma_sb_error; // @[ifu_mem_ctl.scala 405:105]
  wire  _T_2511 = _T_2509 & _T_2623; // @[ifu_mem_ctl.scala 405:129]
  wire  _T_2512 = 3'h1 == perr_state; // @[Conditional.scala 37:30]
  wire  _T_2513 = io_dec_tlu_flush_lower_wb | io_dec_mem_ctrl_dec_tlu_force_halt; // @[ifu_mem_ctl.scala 410:50]
  wire  _T_2515 = 3'h2 == perr_state; // @[Conditional.scala 37:30]
  wire  _T_2522 = 3'h4 == perr_state; // @[Conditional.scala 37:30]
  wire  _T_2524 = 3'h3 == perr_state; // @[Conditional.scala 37:30]
  wire  _GEN_21 = _T_2522 | _T_2524; // @[Conditional.scala 39:67]
  wire  _GEN_23 = _T_2515 ? _T_2513 : _GEN_21; // @[Conditional.scala 39:67]
  wire  _GEN_25 = _T_2512 ? _T_2513 : _GEN_23; // @[Conditional.scala 39:67]
  wire  perr_state_en = _T_2500 ? _T_2511 : _GEN_25; // @[Conditional.scala 40:58]
  wire  perr_sb_write_status = _T_2500 & perr_state_en; // @[Conditional.scala 40:58]
  wire  _T_2514 = io_dec_tlu_flush_lower_wb & io_dec_mem_ctrl_dec_tlu_flush_err_wb; // @[ifu_mem_ctl.scala 411:56]
  wire  _GEN_26 = _T_2512 & _T_2514; // @[Conditional.scala 39:67]
  wire  perr_sel_invalidate = _T_2500 ? 1'h0 : _GEN_26; // @[Conditional.scala 40:58]
  wire [1:0] perr_err_inv_way = perr_sel_invalidate ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  reg  dma_sb_err_state_ff; // @[ifu_mem_ctl.scala 396:58]
  wire  _T_2497 = ~dma_sb_err_state_ff; // @[ifu_mem_ctl.scala 395:49]
  wire  _T_2502 = io_dec_mem_ctrl_ifu_ic_error_start & _T_319; // @[ifu_mem_ctl.scala 404:104]
  wire  _T_2516 = ~io_dec_mem_ctrl_dec_tlu_flush_err_wb; // @[ifu_mem_ctl.scala 414:30]
  wire  _T_2517 = _T_2516 & io_dec_tlu_flush_lower_wb; // @[ifu_mem_ctl.scala 414:68]
  wire  _T_2518 = _T_2517 | io_dec_mem_ctrl_dec_tlu_force_halt; // @[ifu_mem_ctl.scala 414:98]
  wire  _T_2527 = perr_state == 3'h2; // @[ifu_mem_ctl.scala 434:79]
  wire  _T_2528 = io_dec_mem_ctrl_dec_tlu_flush_err_wb & _T_2527; // @[ifu_mem_ctl.scala 434:65]
  wire  _T_2530 = _T_2528 & _T_2623; // @[ifu_mem_ctl.scala 434:94]
  wire  _T_2532 = io_dec_tlu_flush_lower_wb | io_dec_mem_ctrl_dec_tlu_i0_commit_cmt; // @[ifu_mem_ctl.scala 437:59]
  wire  _T_2533 = _T_2532 | io_dec_mem_ctrl_dec_tlu_force_halt; // @[ifu_mem_ctl.scala 437:99]
  wire  _T_2547 = _T_2532 | io_ifu_fetch_val[0]; // @[ifu_mem_ctl.scala 440:94]
  wire  _T_2548 = _T_2547 | ifu_bp_hit_taken_q_f; // @[ifu_mem_ctl.scala 440:116]
  wire  _T_2549 = _T_2548 | io_dec_mem_ctrl_dec_tlu_force_halt; // @[ifu_mem_ctl.scala 440:139]
  wire  _T_2569 = _T_2547 | io_dec_mem_ctrl_dec_tlu_force_halt; // @[ifu_mem_ctl.scala 447:116]
  wire  _T_2577 = io_dec_tlu_flush_lower_wb & _T_2516; // @[ifu_mem_ctl.scala 452:60]
  wire  _T_2578 = _T_2577 | io_dec_mem_ctrl_dec_tlu_i0_commit_cmt; // @[ifu_mem_ctl.scala 452:101]
  wire  _T_2579 = _T_2578 | io_dec_mem_ctrl_dec_tlu_force_halt; // @[ifu_mem_ctl.scala 452:141]
  wire  _GEN_33 = _T_2575 & _T_2533; // @[Conditional.scala 39:67]
  wire  _GEN_36 = _T_2558 ? _T_2569 : _GEN_33; // @[Conditional.scala 39:67]
  wire  _GEN_38 = _T_2558 | _T_2575; // @[Conditional.scala 39:67]
  wire  _GEN_40 = _T_2531 ? _T_2549 : _GEN_36; // @[Conditional.scala 39:67]
  wire  _GEN_42 = _T_2531 | _GEN_38; // @[Conditional.scala 39:67]
  wire  err_stop_state_en = _T_2526 ? _T_2530 : _GEN_40; // @[Conditional.scala 40:58]
  reg  bus_cmd_req_hold; // @[ifu_mem_ctl.scala 475:53]
  wire  _T_2591 = ic_act_miss_f | bus_cmd_req_hold; // @[ifu_mem_ctl.scala 471:45]
  reg  ifu_bus_cmd_valid; // @[ifu_mem_ctl.scala 472:55]
  wire  _T_2592 = _T_2591 | ifu_bus_cmd_valid; // @[ifu_mem_ctl.scala 471:64]
  wire [31:0] _T_2610 = {miss_addr,bus_rd_addr_count,3'h0}; // @[Cat.scala 29:58]
  wire [31:0] _T_2612 = ifu_bus_cmd_valid ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  reg  ifu_bus_arvalid_ff; // @[ifu_mem_ctl.scala 511:53]
  reg  ifc_dma_access_ok_prev; // @[ifu_mem_ctl.scala 560:62]
  wire  _T_2698 = ~iccm_correct_ecc; // @[ifu_mem_ctl.scala 565:50]
  wire  _T_2699 = io_ifc_dma_access_ok & _T_2698; // @[ifu_mem_ctl.scala 565:47]
  wire  _T_2700 = ~io_iccm_dma_sb_error; // @[ifu_mem_ctl.scala 565:70]
  wire  _T_2704 = _T_2699 & ifc_dma_access_ok_prev; // @[ifu_mem_ctl.scala 566:72]
  wire  _T_2705 = perr_state == 3'h0; // @[ifu_mem_ctl.scala 566:111]
  wire  _T_2706 = _T_2704 & _T_2705; // @[ifu_mem_ctl.scala 566:97]
  wire  ifc_dma_access_q_ok = _T_2706 & _T_2700; // @[ifu_mem_ctl.scala 566:127]
  wire  _T_2709 = ifc_dma_access_q_ok & io_dma_mem_ctl_dma_iccm_req; // @[ifu_mem_ctl.scala 569:40]
  wire  _T_2710 = _T_2709 & io_dma_mem_ctl_dma_mem_write; // @[ifu_mem_ctl.scala 569:70]
  wire  _T_2713 = ~io_dma_mem_ctl_dma_mem_write; // @[ifu_mem_ctl.scala 570:72]
  wire  _T_2714 = _T_2709 & _T_2713; // @[ifu_mem_ctl.scala 570:70]
  wire  _T_2715 = io_ifc_iccm_access_bf & io_ifc_fetch_req_bf; // @[ifu_mem_ctl.scala 570:128]
  wire [2:0] _T_2720 = io_dma_mem_ctl_dma_iccm_req ? 3'h7 : 3'h0; // @[Bitwise.scala 72:12]
  wire  _T_2741 = io_dma_mem_ctl_dma_mem_wdata[32] ^ io_dma_mem_ctl_dma_mem_wdata[33]; // @[lib.scala 119:74]
  wire  _T_2742 = _T_2741 ^ io_dma_mem_ctl_dma_mem_wdata[35]; // @[lib.scala 119:74]
  wire  _T_2743 = _T_2742 ^ io_dma_mem_ctl_dma_mem_wdata[36]; // @[lib.scala 119:74]
  wire  _T_2744 = _T_2743 ^ io_dma_mem_ctl_dma_mem_wdata[38]; // @[lib.scala 119:74]
  wire  _T_2745 = _T_2744 ^ io_dma_mem_ctl_dma_mem_wdata[40]; // @[lib.scala 119:74]
  wire  _T_2746 = _T_2745 ^ io_dma_mem_ctl_dma_mem_wdata[42]; // @[lib.scala 119:74]
  wire  _T_2747 = _T_2746 ^ io_dma_mem_ctl_dma_mem_wdata[43]; // @[lib.scala 119:74]
  wire  _T_2748 = _T_2747 ^ io_dma_mem_ctl_dma_mem_wdata[45]; // @[lib.scala 119:74]
  wire  _T_2749 = _T_2748 ^ io_dma_mem_ctl_dma_mem_wdata[47]; // @[lib.scala 119:74]
  wire  _T_2750 = _T_2749 ^ io_dma_mem_ctl_dma_mem_wdata[49]; // @[lib.scala 119:74]
  wire  _T_2751 = _T_2750 ^ io_dma_mem_ctl_dma_mem_wdata[51]; // @[lib.scala 119:74]
  wire  _T_2752 = _T_2751 ^ io_dma_mem_ctl_dma_mem_wdata[53]; // @[lib.scala 119:74]
  wire  _T_2753 = _T_2752 ^ io_dma_mem_ctl_dma_mem_wdata[55]; // @[lib.scala 119:74]
  wire  _T_2754 = _T_2753 ^ io_dma_mem_ctl_dma_mem_wdata[57]; // @[lib.scala 119:74]
  wire  _T_2755 = _T_2754 ^ io_dma_mem_ctl_dma_mem_wdata[58]; // @[lib.scala 119:74]
  wire  _T_2756 = _T_2755 ^ io_dma_mem_ctl_dma_mem_wdata[60]; // @[lib.scala 119:74]
  wire  _T_2757 = _T_2756 ^ io_dma_mem_ctl_dma_mem_wdata[62]; // @[lib.scala 119:74]
  wire  _T_2776 = io_dma_mem_ctl_dma_mem_wdata[32] ^ io_dma_mem_ctl_dma_mem_wdata[34]; // @[lib.scala 119:74]
  wire  _T_2777 = _T_2776 ^ io_dma_mem_ctl_dma_mem_wdata[35]; // @[lib.scala 119:74]
  wire  _T_2778 = _T_2777 ^ io_dma_mem_ctl_dma_mem_wdata[37]; // @[lib.scala 119:74]
  wire  _T_2779 = _T_2778 ^ io_dma_mem_ctl_dma_mem_wdata[38]; // @[lib.scala 119:74]
  wire  _T_2780 = _T_2779 ^ io_dma_mem_ctl_dma_mem_wdata[41]; // @[lib.scala 119:74]
  wire  _T_2781 = _T_2780 ^ io_dma_mem_ctl_dma_mem_wdata[42]; // @[lib.scala 119:74]
  wire  _T_2782 = _T_2781 ^ io_dma_mem_ctl_dma_mem_wdata[44]; // @[lib.scala 119:74]
  wire  _T_2783 = _T_2782 ^ io_dma_mem_ctl_dma_mem_wdata[45]; // @[lib.scala 119:74]
  wire  _T_2784 = _T_2783 ^ io_dma_mem_ctl_dma_mem_wdata[48]; // @[lib.scala 119:74]
  wire  _T_2785 = _T_2784 ^ io_dma_mem_ctl_dma_mem_wdata[49]; // @[lib.scala 119:74]
  wire  _T_2786 = _T_2785 ^ io_dma_mem_ctl_dma_mem_wdata[52]; // @[lib.scala 119:74]
  wire  _T_2787 = _T_2786 ^ io_dma_mem_ctl_dma_mem_wdata[53]; // @[lib.scala 119:74]
  wire  _T_2788 = _T_2787 ^ io_dma_mem_ctl_dma_mem_wdata[56]; // @[lib.scala 119:74]
  wire  _T_2789 = _T_2788 ^ io_dma_mem_ctl_dma_mem_wdata[57]; // @[lib.scala 119:74]
  wire  _T_2790 = _T_2789 ^ io_dma_mem_ctl_dma_mem_wdata[59]; // @[lib.scala 119:74]
  wire  _T_2791 = _T_2790 ^ io_dma_mem_ctl_dma_mem_wdata[60]; // @[lib.scala 119:74]
  wire  _T_2792 = _T_2791 ^ io_dma_mem_ctl_dma_mem_wdata[63]; // @[lib.scala 119:74]
  wire  _T_2811 = io_dma_mem_ctl_dma_mem_wdata[33] ^ io_dma_mem_ctl_dma_mem_wdata[34]; // @[lib.scala 119:74]
  wire  _T_2812 = _T_2811 ^ io_dma_mem_ctl_dma_mem_wdata[35]; // @[lib.scala 119:74]
  wire  _T_2813 = _T_2812 ^ io_dma_mem_ctl_dma_mem_wdata[39]; // @[lib.scala 119:74]
  wire  _T_2814 = _T_2813 ^ io_dma_mem_ctl_dma_mem_wdata[40]; // @[lib.scala 119:74]
  wire  _T_2815 = _T_2814 ^ io_dma_mem_ctl_dma_mem_wdata[41]; // @[lib.scala 119:74]
  wire  _T_2816 = _T_2815 ^ io_dma_mem_ctl_dma_mem_wdata[42]; // @[lib.scala 119:74]
  wire  _T_2817 = _T_2816 ^ io_dma_mem_ctl_dma_mem_wdata[46]; // @[lib.scala 119:74]
  wire  _T_2818 = _T_2817 ^ io_dma_mem_ctl_dma_mem_wdata[47]; // @[lib.scala 119:74]
  wire  _T_2819 = _T_2818 ^ io_dma_mem_ctl_dma_mem_wdata[48]; // @[lib.scala 119:74]
  wire  _T_2820 = _T_2819 ^ io_dma_mem_ctl_dma_mem_wdata[49]; // @[lib.scala 119:74]
  wire  _T_2821 = _T_2820 ^ io_dma_mem_ctl_dma_mem_wdata[54]; // @[lib.scala 119:74]
  wire  _T_2822 = _T_2821 ^ io_dma_mem_ctl_dma_mem_wdata[55]; // @[lib.scala 119:74]
  wire  _T_2823 = _T_2822 ^ io_dma_mem_ctl_dma_mem_wdata[56]; // @[lib.scala 119:74]
  wire  _T_2824 = _T_2823 ^ io_dma_mem_ctl_dma_mem_wdata[57]; // @[lib.scala 119:74]
  wire  _T_2825 = _T_2824 ^ io_dma_mem_ctl_dma_mem_wdata[61]; // @[lib.scala 119:74]
  wire  _T_2826 = _T_2825 ^ io_dma_mem_ctl_dma_mem_wdata[62]; // @[lib.scala 119:74]
  wire  _T_2827 = _T_2826 ^ io_dma_mem_ctl_dma_mem_wdata[63]; // @[lib.scala 119:74]
  wire  _T_2843 = io_dma_mem_ctl_dma_mem_wdata[36] ^ io_dma_mem_ctl_dma_mem_wdata[37]; // @[lib.scala 119:74]
  wire  _T_2844 = _T_2843 ^ io_dma_mem_ctl_dma_mem_wdata[38]; // @[lib.scala 119:74]
  wire  _T_2845 = _T_2844 ^ io_dma_mem_ctl_dma_mem_wdata[39]; // @[lib.scala 119:74]
  wire  _T_2846 = _T_2845 ^ io_dma_mem_ctl_dma_mem_wdata[40]; // @[lib.scala 119:74]
  wire  _T_2847 = _T_2846 ^ io_dma_mem_ctl_dma_mem_wdata[41]; // @[lib.scala 119:74]
  wire  _T_2848 = _T_2847 ^ io_dma_mem_ctl_dma_mem_wdata[42]; // @[lib.scala 119:74]
  wire  _T_2849 = _T_2848 ^ io_dma_mem_ctl_dma_mem_wdata[50]; // @[lib.scala 119:74]
  wire  _T_2850 = _T_2849 ^ io_dma_mem_ctl_dma_mem_wdata[51]; // @[lib.scala 119:74]
  wire  _T_2851 = _T_2850 ^ io_dma_mem_ctl_dma_mem_wdata[52]; // @[lib.scala 119:74]
  wire  _T_2852 = _T_2851 ^ io_dma_mem_ctl_dma_mem_wdata[53]; // @[lib.scala 119:74]
  wire  _T_2853 = _T_2852 ^ io_dma_mem_ctl_dma_mem_wdata[54]; // @[lib.scala 119:74]
  wire  _T_2854 = _T_2853 ^ io_dma_mem_ctl_dma_mem_wdata[55]; // @[lib.scala 119:74]
  wire  _T_2855 = _T_2854 ^ io_dma_mem_ctl_dma_mem_wdata[56]; // @[lib.scala 119:74]
  wire  _T_2856 = _T_2855 ^ io_dma_mem_ctl_dma_mem_wdata[57]; // @[lib.scala 119:74]
  wire  _T_2872 = io_dma_mem_ctl_dma_mem_wdata[43] ^ io_dma_mem_ctl_dma_mem_wdata[44]; // @[lib.scala 119:74]
  wire  _T_2873 = _T_2872 ^ io_dma_mem_ctl_dma_mem_wdata[45]; // @[lib.scala 119:74]
  wire  _T_2874 = _T_2873 ^ io_dma_mem_ctl_dma_mem_wdata[46]; // @[lib.scala 119:74]
  wire  _T_2875 = _T_2874 ^ io_dma_mem_ctl_dma_mem_wdata[47]; // @[lib.scala 119:74]
  wire  _T_2876 = _T_2875 ^ io_dma_mem_ctl_dma_mem_wdata[48]; // @[lib.scala 119:74]
  wire  _T_2877 = _T_2876 ^ io_dma_mem_ctl_dma_mem_wdata[49]; // @[lib.scala 119:74]
  wire  _T_2878 = _T_2877 ^ io_dma_mem_ctl_dma_mem_wdata[50]; // @[lib.scala 119:74]
  wire  _T_2879 = _T_2878 ^ io_dma_mem_ctl_dma_mem_wdata[51]; // @[lib.scala 119:74]
  wire  _T_2880 = _T_2879 ^ io_dma_mem_ctl_dma_mem_wdata[52]; // @[lib.scala 119:74]
  wire  _T_2881 = _T_2880 ^ io_dma_mem_ctl_dma_mem_wdata[53]; // @[lib.scala 119:74]
  wire  _T_2882 = _T_2881 ^ io_dma_mem_ctl_dma_mem_wdata[54]; // @[lib.scala 119:74]
  wire  _T_2883 = _T_2882 ^ io_dma_mem_ctl_dma_mem_wdata[55]; // @[lib.scala 119:74]
  wire  _T_2884 = _T_2883 ^ io_dma_mem_ctl_dma_mem_wdata[56]; // @[lib.scala 119:74]
  wire  _T_2885 = _T_2884 ^ io_dma_mem_ctl_dma_mem_wdata[57]; // @[lib.scala 119:74]
  wire  _T_2892 = io_dma_mem_ctl_dma_mem_wdata[58] ^ io_dma_mem_ctl_dma_mem_wdata[59]; // @[lib.scala 119:74]
  wire  _T_2893 = _T_2892 ^ io_dma_mem_ctl_dma_mem_wdata[60]; // @[lib.scala 119:74]
  wire  _T_2894 = _T_2893 ^ io_dma_mem_ctl_dma_mem_wdata[61]; // @[lib.scala 119:74]
  wire  _T_2895 = _T_2894 ^ io_dma_mem_ctl_dma_mem_wdata[62]; // @[lib.scala 119:74]
  wire  _T_2896 = _T_2895 ^ io_dma_mem_ctl_dma_mem_wdata[63]; // @[lib.scala 119:74]
  wire [5:0] _T_2901 = {_T_2896,_T_2885,_T_2856,_T_2827,_T_2792,_T_2757}; // @[Cat.scala 29:58]
  wire  _T_2902 = ^io_dma_mem_ctl_dma_mem_wdata[63:32]; // @[lib.scala 127:13]
  wire  _T_2903 = ^_T_2901; // @[lib.scala 127:23]
  wire  _T_2904 = _T_2902 ^ _T_2903; // @[lib.scala 127:18]
  wire  _T_2925 = io_dma_mem_ctl_dma_mem_wdata[0] ^ io_dma_mem_ctl_dma_mem_wdata[1]; // @[lib.scala 119:74]
  wire  _T_2926 = _T_2925 ^ io_dma_mem_ctl_dma_mem_wdata[3]; // @[lib.scala 119:74]
  wire  _T_2927 = _T_2926 ^ io_dma_mem_ctl_dma_mem_wdata[4]; // @[lib.scala 119:74]
  wire  _T_2928 = _T_2927 ^ io_dma_mem_ctl_dma_mem_wdata[6]; // @[lib.scala 119:74]
  wire  _T_2929 = _T_2928 ^ io_dma_mem_ctl_dma_mem_wdata[8]; // @[lib.scala 119:74]
  wire  _T_2930 = _T_2929 ^ io_dma_mem_ctl_dma_mem_wdata[10]; // @[lib.scala 119:74]
  wire  _T_2931 = _T_2930 ^ io_dma_mem_ctl_dma_mem_wdata[11]; // @[lib.scala 119:74]
  wire  _T_2932 = _T_2931 ^ io_dma_mem_ctl_dma_mem_wdata[13]; // @[lib.scala 119:74]
  wire  _T_2933 = _T_2932 ^ io_dma_mem_ctl_dma_mem_wdata[15]; // @[lib.scala 119:74]
  wire  _T_2934 = _T_2933 ^ io_dma_mem_ctl_dma_mem_wdata[17]; // @[lib.scala 119:74]
  wire  _T_2935 = _T_2934 ^ io_dma_mem_ctl_dma_mem_wdata[19]; // @[lib.scala 119:74]
  wire  _T_2936 = _T_2935 ^ io_dma_mem_ctl_dma_mem_wdata[21]; // @[lib.scala 119:74]
  wire  _T_2937 = _T_2936 ^ io_dma_mem_ctl_dma_mem_wdata[23]; // @[lib.scala 119:74]
  wire  _T_2938 = _T_2937 ^ io_dma_mem_ctl_dma_mem_wdata[25]; // @[lib.scala 119:74]
  wire  _T_2939 = _T_2938 ^ io_dma_mem_ctl_dma_mem_wdata[26]; // @[lib.scala 119:74]
  wire  _T_2940 = _T_2939 ^ io_dma_mem_ctl_dma_mem_wdata[28]; // @[lib.scala 119:74]
  wire  _T_2941 = _T_2940 ^ io_dma_mem_ctl_dma_mem_wdata[30]; // @[lib.scala 119:74]
  wire  _T_2960 = io_dma_mem_ctl_dma_mem_wdata[0] ^ io_dma_mem_ctl_dma_mem_wdata[2]; // @[lib.scala 119:74]
  wire  _T_2961 = _T_2960 ^ io_dma_mem_ctl_dma_mem_wdata[3]; // @[lib.scala 119:74]
  wire  _T_2962 = _T_2961 ^ io_dma_mem_ctl_dma_mem_wdata[5]; // @[lib.scala 119:74]
  wire  _T_2963 = _T_2962 ^ io_dma_mem_ctl_dma_mem_wdata[6]; // @[lib.scala 119:74]
  wire  _T_2964 = _T_2963 ^ io_dma_mem_ctl_dma_mem_wdata[9]; // @[lib.scala 119:74]
  wire  _T_2965 = _T_2964 ^ io_dma_mem_ctl_dma_mem_wdata[10]; // @[lib.scala 119:74]
  wire  _T_2966 = _T_2965 ^ io_dma_mem_ctl_dma_mem_wdata[12]; // @[lib.scala 119:74]
  wire  _T_2967 = _T_2966 ^ io_dma_mem_ctl_dma_mem_wdata[13]; // @[lib.scala 119:74]
  wire  _T_2968 = _T_2967 ^ io_dma_mem_ctl_dma_mem_wdata[16]; // @[lib.scala 119:74]
  wire  _T_2969 = _T_2968 ^ io_dma_mem_ctl_dma_mem_wdata[17]; // @[lib.scala 119:74]
  wire  _T_2970 = _T_2969 ^ io_dma_mem_ctl_dma_mem_wdata[20]; // @[lib.scala 119:74]
  wire  _T_2971 = _T_2970 ^ io_dma_mem_ctl_dma_mem_wdata[21]; // @[lib.scala 119:74]
  wire  _T_2972 = _T_2971 ^ io_dma_mem_ctl_dma_mem_wdata[24]; // @[lib.scala 119:74]
  wire  _T_2973 = _T_2972 ^ io_dma_mem_ctl_dma_mem_wdata[25]; // @[lib.scala 119:74]
  wire  _T_2974 = _T_2973 ^ io_dma_mem_ctl_dma_mem_wdata[27]; // @[lib.scala 119:74]
  wire  _T_2975 = _T_2974 ^ io_dma_mem_ctl_dma_mem_wdata[28]; // @[lib.scala 119:74]
  wire  _T_2976 = _T_2975 ^ io_dma_mem_ctl_dma_mem_wdata[31]; // @[lib.scala 119:74]
  wire  _T_2995 = io_dma_mem_ctl_dma_mem_wdata[1] ^ io_dma_mem_ctl_dma_mem_wdata[2]; // @[lib.scala 119:74]
  wire  _T_2996 = _T_2995 ^ io_dma_mem_ctl_dma_mem_wdata[3]; // @[lib.scala 119:74]
  wire  _T_2997 = _T_2996 ^ io_dma_mem_ctl_dma_mem_wdata[7]; // @[lib.scala 119:74]
  wire  _T_2998 = _T_2997 ^ io_dma_mem_ctl_dma_mem_wdata[8]; // @[lib.scala 119:74]
  wire  _T_2999 = _T_2998 ^ io_dma_mem_ctl_dma_mem_wdata[9]; // @[lib.scala 119:74]
  wire  _T_3000 = _T_2999 ^ io_dma_mem_ctl_dma_mem_wdata[10]; // @[lib.scala 119:74]
  wire  _T_3001 = _T_3000 ^ io_dma_mem_ctl_dma_mem_wdata[14]; // @[lib.scala 119:74]
  wire  _T_3002 = _T_3001 ^ io_dma_mem_ctl_dma_mem_wdata[15]; // @[lib.scala 119:74]
  wire  _T_3003 = _T_3002 ^ io_dma_mem_ctl_dma_mem_wdata[16]; // @[lib.scala 119:74]
  wire  _T_3004 = _T_3003 ^ io_dma_mem_ctl_dma_mem_wdata[17]; // @[lib.scala 119:74]
  wire  _T_3005 = _T_3004 ^ io_dma_mem_ctl_dma_mem_wdata[22]; // @[lib.scala 119:74]
  wire  _T_3006 = _T_3005 ^ io_dma_mem_ctl_dma_mem_wdata[23]; // @[lib.scala 119:74]
  wire  _T_3007 = _T_3006 ^ io_dma_mem_ctl_dma_mem_wdata[24]; // @[lib.scala 119:74]
  wire  _T_3008 = _T_3007 ^ io_dma_mem_ctl_dma_mem_wdata[25]; // @[lib.scala 119:74]
  wire  _T_3009 = _T_3008 ^ io_dma_mem_ctl_dma_mem_wdata[29]; // @[lib.scala 119:74]
  wire  _T_3010 = _T_3009 ^ io_dma_mem_ctl_dma_mem_wdata[30]; // @[lib.scala 119:74]
  wire  _T_3011 = _T_3010 ^ io_dma_mem_ctl_dma_mem_wdata[31]; // @[lib.scala 119:74]
  wire  _T_3027 = io_dma_mem_ctl_dma_mem_wdata[4] ^ io_dma_mem_ctl_dma_mem_wdata[5]; // @[lib.scala 119:74]
  wire  _T_3028 = _T_3027 ^ io_dma_mem_ctl_dma_mem_wdata[6]; // @[lib.scala 119:74]
  wire  _T_3029 = _T_3028 ^ io_dma_mem_ctl_dma_mem_wdata[7]; // @[lib.scala 119:74]
  wire  _T_3030 = _T_3029 ^ io_dma_mem_ctl_dma_mem_wdata[8]; // @[lib.scala 119:74]
  wire  _T_3031 = _T_3030 ^ io_dma_mem_ctl_dma_mem_wdata[9]; // @[lib.scala 119:74]
  wire  _T_3032 = _T_3031 ^ io_dma_mem_ctl_dma_mem_wdata[10]; // @[lib.scala 119:74]
  wire  _T_3033 = _T_3032 ^ io_dma_mem_ctl_dma_mem_wdata[18]; // @[lib.scala 119:74]
  wire  _T_3034 = _T_3033 ^ io_dma_mem_ctl_dma_mem_wdata[19]; // @[lib.scala 119:74]
  wire  _T_3035 = _T_3034 ^ io_dma_mem_ctl_dma_mem_wdata[20]; // @[lib.scala 119:74]
  wire  _T_3036 = _T_3035 ^ io_dma_mem_ctl_dma_mem_wdata[21]; // @[lib.scala 119:74]
  wire  _T_3037 = _T_3036 ^ io_dma_mem_ctl_dma_mem_wdata[22]; // @[lib.scala 119:74]
  wire  _T_3038 = _T_3037 ^ io_dma_mem_ctl_dma_mem_wdata[23]; // @[lib.scala 119:74]
  wire  _T_3039 = _T_3038 ^ io_dma_mem_ctl_dma_mem_wdata[24]; // @[lib.scala 119:74]
  wire  _T_3040 = _T_3039 ^ io_dma_mem_ctl_dma_mem_wdata[25]; // @[lib.scala 119:74]
  wire  _T_3056 = io_dma_mem_ctl_dma_mem_wdata[11] ^ io_dma_mem_ctl_dma_mem_wdata[12]; // @[lib.scala 119:74]
  wire  _T_3057 = _T_3056 ^ io_dma_mem_ctl_dma_mem_wdata[13]; // @[lib.scala 119:74]
  wire  _T_3058 = _T_3057 ^ io_dma_mem_ctl_dma_mem_wdata[14]; // @[lib.scala 119:74]
  wire  _T_3059 = _T_3058 ^ io_dma_mem_ctl_dma_mem_wdata[15]; // @[lib.scala 119:74]
  wire  _T_3060 = _T_3059 ^ io_dma_mem_ctl_dma_mem_wdata[16]; // @[lib.scala 119:74]
  wire  _T_3061 = _T_3060 ^ io_dma_mem_ctl_dma_mem_wdata[17]; // @[lib.scala 119:74]
  wire  _T_3062 = _T_3061 ^ io_dma_mem_ctl_dma_mem_wdata[18]; // @[lib.scala 119:74]
  wire  _T_3063 = _T_3062 ^ io_dma_mem_ctl_dma_mem_wdata[19]; // @[lib.scala 119:74]
  wire  _T_3064 = _T_3063 ^ io_dma_mem_ctl_dma_mem_wdata[20]; // @[lib.scala 119:74]
  wire  _T_3065 = _T_3064 ^ io_dma_mem_ctl_dma_mem_wdata[21]; // @[lib.scala 119:74]
  wire  _T_3066 = _T_3065 ^ io_dma_mem_ctl_dma_mem_wdata[22]; // @[lib.scala 119:74]
  wire  _T_3067 = _T_3066 ^ io_dma_mem_ctl_dma_mem_wdata[23]; // @[lib.scala 119:74]
  wire  _T_3068 = _T_3067 ^ io_dma_mem_ctl_dma_mem_wdata[24]; // @[lib.scala 119:74]
  wire  _T_3069 = _T_3068 ^ io_dma_mem_ctl_dma_mem_wdata[25]; // @[lib.scala 119:74]
  wire  _T_3076 = io_dma_mem_ctl_dma_mem_wdata[26] ^ io_dma_mem_ctl_dma_mem_wdata[27]; // @[lib.scala 119:74]
  wire  _T_3077 = _T_3076 ^ io_dma_mem_ctl_dma_mem_wdata[28]; // @[lib.scala 119:74]
  wire  _T_3078 = _T_3077 ^ io_dma_mem_ctl_dma_mem_wdata[29]; // @[lib.scala 119:74]
  wire  _T_3079 = _T_3078 ^ io_dma_mem_ctl_dma_mem_wdata[30]; // @[lib.scala 119:74]
  wire  _T_3080 = _T_3079 ^ io_dma_mem_ctl_dma_mem_wdata[31]; // @[lib.scala 119:74]
  wire [5:0] _T_3085 = {_T_3080,_T_3069,_T_3040,_T_3011,_T_2976,_T_2941}; // @[Cat.scala 29:58]
  wire  _T_3086 = ^io_dma_mem_ctl_dma_mem_wdata[31:0]; // @[lib.scala 127:13]
  wire  _T_3087 = ^_T_3085; // @[lib.scala 127:23]
  wire  _T_3088 = _T_3086 ^ _T_3087; // @[lib.scala 127:18]
  wire [6:0] _T_3089 = {_T_3088,_T_3080,_T_3069,_T_3040,_T_3011,_T_2976,_T_2941}; // @[Cat.scala 29:58]
  wire [13:0] dma_mem_ecc = {_T_2904,_T_2896,_T_2885,_T_2856,_T_2827,_T_2792,_T_2757,_T_3089}; // @[Cat.scala 29:58]
  wire  _T_3091 = ~_T_2709; // @[ifu_mem_ctl.scala 576:45]
  wire  _T_3092 = iccm_correct_ecc & _T_3091; // @[ifu_mem_ctl.scala 576:43]
  reg [38:0] iccm_ecc_corr_data_ff; // @[Reg.scala 27:20]
  wire [77:0] _T_3093 = {iccm_ecc_corr_data_ff,iccm_ecc_corr_data_ff}; // @[Cat.scala 29:58]
  wire [77:0] _T_3100 = {dma_mem_ecc[13:7],io_dma_mem_ctl_dma_mem_wdata[63:32],dma_mem_ecc[6:0],io_dma_mem_ctl_dma_mem_wdata[31:0]}; // @[Cat.scala 29:58]
  reg [1:0] dma_mem_addr_ff; // @[ifu_mem_ctl.scala 590:53]
  wire  _T_3435 = _T_3347[5:0] == 6'h27; // @[lib.scala 199:41]
  wire  _T_3433 = _T_3347[5:0] == 6'h26; // @[lib.scala 199:41]
  wire  _T_3431 = _T_3347[5:0] == 6'h25; // @[lib.scala 199:41]
  wire  _T_3429 = _T_3347[5:0] == 6'h24; // @[lib.scala 199:41]
  wire  _T_3427 = _T_3347[5:0] == 6'h23; // @[lib.scala 199:41]
  wire  _T_3425 = _T_3347[5:0] == 6'h22; // @[lib.scala 199:41]
  wire  _T_3423 = _T_3347[5:0] == 6'h21; // @[lib.scala 199:41]
  wire  _T_3421 = _T_3347[5:0] == 6'h20; // @[lib.scala 199:41]
  wire  _T_3419 = _T_3347[5:0] == 6'h1f; // @[lib.scala 199:41]
  wire  _T_3417 = _T_3347[5:0] == 6'h1e; // @[lib.scala 199:41]
  wire [9:0] _T_3493 = {_T_3435,_T_3433,_T_3431,_T_3429,_T_3427,_T_3425,_T_3423,_T_3421,_T_3419,_T_3417}; // @[lib.scala 202:69]
  wire  _T_3415 = _T_3347[5:0] == 6'h1d; // @[lib.scala 199:41]
  wire  _T_3413 = _T_3347[5:0] == 6'h1c; // @[lib.scala 199:41]
  wire  _T_3411 = _T_3347[5:0] == 6'h1b; // @[lib.scala 199:41]
  wire  _T_3409 = _T_3347[5:0] == 6'h1a; // @[lib.scala 199:41]
  wire  _T_3407 = _T_3347[5:0] == 6'h19; // @[lib.scala 199:41]
  wire  _T_3405 = _T_3347[5:0] == 6'h18; // @[lib.scala 199:41]
  wire  _T_3403 = _T_3347[5:0] == 6'h17; // @[lib.scala 199:41]
  wire  _T_3401 = _T_3347[5:0] == 6'h16; // @[lib.scala 199:41]
  wire  _T_3399 = _T_3347[5:0] == 6'h15; // @[lib.scala 199:41]
  wire  _T_3397 = _T_3347[5:0] == 6'h14; // @[lib.scala 199:41]
  wire [9:0] _T_3484 = {_T_3415,_T_3413,_T_3411,_T_3409,_T_3407,_T_3405,_T_3403,_T_3401,_T_3399,_T_3397}; // @[lib.scala 202:69]
  wire  _T_3395 = _T_3347[5:0] == 6'h13; // @[lib.scala 199:41]
  wire  _T_3393 = _T_3347[5:0] == 6'h12; // @[lib.scala 199:41]
  wire  _T_3391 = _T_3347[5:0] == 6'h11; // @[lib.scala 199:41]
  wire  _T_3389 = _T_3347[5:0] == 6'h10; // @[lib.scala 199:41]
  wire  _T_3387 = _T_3347[5:0] == 6'hf; // @[lib.scala 199:41]
  wire  _T_3385 = _T_3347[5:0] == 6'he; // @[lib.scala 199:41]
  wire  _T_3383 = _T_3347[5:0] == 6'hd; // @[lib.scala 199:41]
  wire  _T_3381 = _T_3347[5:0] == 6'hc; // @[lib.scala 199:41]
  wire  _T_3379 = _T_3347[5:0] == 6'hb; // @[lib.scala 199:41]
  wire  _T_3377 = _T_3347[5:0] == 6'ha; // @[lib.scala 199:41]
  wire [9:0] _T_3474 = {_T_3395,_T_3393,_T_3391,_T_3389,_T_3387,_T_3385,_T_3383,_T_3381,_T_3379,_T_3377}; // @[lib.scala 202:69]
  wire  _T_3375 = _T_3347[5:0] == 6'h9; // @[lib.scala 199:41]
  wire  _T_3373 = _T_3347[5:0] == 6'h8; // @[lib.scala 199:41]
  wire  _T_3371 = _T_3347[5:0] == 6'h7; // @[lib.scala 199:41]
  wire  _T_3369 = _T_3347[5:0] == 6'h6; // @[lib.scala 199:41]
  wire  _T_3367 = _T_3347[5:0] == 6'h5; // @[lib.scala 199:41]
  wire  _T_3365 = _T_3347[5:0] == 6'h4; // @[lib.scala 199:41]
  wire  _T_3363 = _T_3347[5:0] == 6'h3; // @[lib.scala 199:41]
  wire  _T_3361 = _T_3347[5:0] == 6'h2; // @[lib.scala 199:41]
  wire  _T_3359 = _T_3347[5:0] == 6'h1; // @[lib.scala 199:41]
  wire [18:0] _T_3475 = {_T_3474,_T_3375,_T_3373,_T_3371,_T_3369,_T_3367,_T_3365,_T_3363,_T_3361,_T_3359}; // @[lib.scala 202:69]
  wire [38:0] _T_3495 = {_T_3493,_T_3484,_T_3475}; // @[lib.scala 202:69]
  wire [7:0] _T_3450 = {io_iccm_rd_data_ecc[35],io_iccm_rd_data_ecc[3:1],io_iccm_rd_data_ecc[34],io_iccm_rd_data_ecc[0],io_iccm_rd_data_ecc[33:32]}; // @[Cat.scala 29:58]
  wire [38:0] _T_3456 = {io_iccm_rd_data_ecc[38],io_iccm_rd_data_ecc[31:26],io_iccm_rd_data_ecc[37],io_iccm_rd_data_ecc[25:11],io_iccm_rd_data_ecc[36],io_iccm_rd_data_ecc[10:4],_T_3450}; // @[Cat.scala 29:58]
  wire [38:0] _T_3496 = _T_3495 ^ _T_3456; // @[lib.scala 202:76]
  wire [38:0] _T_3497 = _T_3351 ? _T_3496 : _T_3456; // @[lib.scala 202:31]
  wire [31:0] iccm_corrected_data_0 = {_T_3497[37:32],_T_3497[30:16],_T_3497[14:8],_T_3497[6:4],_T_3497[2]}; // @[Cat.scala 29:58]
  wire  _T_3820 = _T_3732[5:0] == 6'h27; // @[lib.scala 199:41]
  wire  _T_3818 = _T_3732[5:0] == 6'h26; // @[lib.scala 199:41]
  wire  _T_3816 = _T_3732[5:0] == 6'h25; // @[lib.scala 199:41]
  wire  _T_3814 = _T_3732[5:0] == 6'h24; // @[lib.scala 199:41]
  wire  _T_3812 = _T_3732[5:0] == 6'h23; // @[lib.scala 199:41]
  wire  _T_3810 = _T_3732[5:0] == 6'h22; // @[lib.scala 199:41]
  wire  _T_3808 = _T_3732[5:0] == 6'h21; // @[lib.scala 199:41]
  wire  _T_3806 = _T_3732[5:0] == 6'h20; // @[lib.scala 199:41]
  wire  _T_3804 = _T_3732[5:0] == 6'h1f; // @[lib.scala 199:41]
  wire  _T_3802 = _T_3732[5:0] == 6'h1e; // @[lib.scala 199:41]
  wire [9:0] _T_3878 = {_T_3820,_T_3818,_T_3816,_T_3814,_T_3812,_T_3810,_T_3808,_T_3806,_T_3804,_T_3802}; // @[lib.scala 202:69]
  wire  _T_3800 = _T_3732[5:0] == 6'h1d; // @[lib.scala 199:41]
  wire  _T_3798 = _T_3732[5:0] == 6'h1c; // @[lib.scala 199:41]
  wire  _T_3796 = _T_3732[5:0] == 6'h1b; // @[lib.scala 199:41]
  wire  _T_3794 = _T_3732[5:0] == 6'h1a; // @[lib.scala 199:41]
  wire  _T_3792 = _T_3732[5:0] == 6'h19; // @[lib.scala 199:41]
  wire  _T_3790 = _T_3732[5:0] == 6'h18; // @[lib.scala 199:41]
  wire  _T_3788 = _T_3732[5:0] == 6'h17; // @[lib.scala 199:41]
  wire  _T_3786 = _T_3732[5:0] == 6'h16; // @[lib.scala 199:41]
  wire  _T_3784 = _T_3732[5:0] == 6'h15; // @[lib.scala 199:41]
  wire  _T_3782 = _T_3732[5:0] == 6'h14; // @[lib.scala 199:41]
  wire [9:0] _T_3869 = {_T_3800,_T_3798,_T_3796,_T_3794,_T_3792,_T_3790,_T_3788,_T_3786,_T_3784,_T_3782}; // @[lib.scala 202:69]
  wire  _T_3780 = _T_3732[5:0] == 6'h13; // @[lib.scala 199:41]
  wire  _T_3778 = _T_3732[5:0] == 6'h12; // @[lib.scala 199:41]
  wire  _T_3776 = _T_3732[5:0] == 6'h11; // @[lib.scala 199:41]
  wire  _T_3774 = _T_3732[5:0] == 6'h10; // @[lib.scala 199:41]
  wire  _T_3772 = _T_3732[5:0] == 6'hf; // @[lib.scala 199:41]
  wire  _T_3770 = _T_3732[5:0] == 6'he; // @[lib.scala 199:41]
  wire  _T_3768 = _T_3732[5:0] == 6'hd; // @[lib.scala 199:41]
  wire  _T_3766 = _T_3732[5:0] == 6'hc; // @[lib.scala 199:41]
  wire  _T_3764 = _T_3732[5:0] == 6'hb; // @[lib.scala 199:41]
  wire  _T_3762 = _T_3732[5:0] == 6'ha; // @[lib.scala 199:41]
  wire [9:0] _T_3859 = {_T_3780,_T_3778,_T_3776,_T_3774,_T_3772,_T_3770,_T_3768,_T_3766,_T_3764,_T_3762}; // @[lib.scala 202:69]
  wire  _T_3760 = _T_3732[5:0] == 6'h9; // @[lib.scala 199:41]
  wire  _T_3758 = _T_3732[5:0] == 6'h8; // @[lib.scala 199:41]
  wire  _T_3756 = _T_3732[5:0] == 6'h7; // @[lib.scala 199:41]
  wire  _T_3754 = _T_3732[5:0] == 6'h6; // @[lib.scala 199:41]
  wire  _T_3752 = _T_3732[5:0] == 6'h5; // @[lib.scala 199:41]
  wire  _T_3750 = _T_3732[5:0] == 6'h4; // @[lib.scala 199:41]
  wire  _T_3748 = _T_3732[5:0] == 6'h3; // @[lib.scala 199:41]
  wire  _T_3746 = _T_3732[5:0] == 6'h2; // @[lib.scala 199:41]
  wire  _T_3744 = _T_3732[5:0] == 6'h1; // @[lib.scala 199:41]
  wire [18:0] _T_3860 = {_T_3859,_T_3760,_T_3758,_T_3756,_T_3754,_T_3752,_T_3750,_T_3748,_T_3746,_T_3744}; // @[lib.scala 202:69]
  wire [38:0] _T_3880 = {_T_3878,_T_3869,_T_3860}; // @[lib.scala 202:69]
  wire [7:0] _T_3835 = {io_iccm_rd_data_ecc[74],io_iccm_rd_data_ecc[42:40],io_iccm_rd_data_ecc[73],io_iccm_rd_data_ecc[39],io_iccm_rd_data_ecc[72:71]}; // @[Cat.scala 29:58]
  wire [38:0] _T_3841 = {io_iccm_rd_data_ecc[77],io_iccm_rd_data_ecc[70:65],io_iccm_rd_data_ecc[76],io_iccm_rd_data_ecc[64:50],io_iccm_rd_data_ecc[75],io_iccm_rd_data_ecc[49:43],_T_3835}; // @[Cat.scala 29:58]
  wire [38:0] _T_3881 = _T_3880 ^ _T_3841; // @[lib.scala 202:76]
  wire [38:0] _T_3882 = _T_3736 ? _T_3881 : _T_3841; // @[lib.scala 202:31]
  wire [31:0] iccm_corrected_data_1 = {_T_3882[37:32],_T_3882[30:16],_T_3882[14:8],_T_3882[6:4],_T_3882[2]}; // @[Cat.scala 29:58]
  wire [31:0] iccm_dma_rdata_1_muxed = dma_mem_addr_ff[0] ? iccm_corrected_data_0 : iccm_corrected_data_1; // @[ifu_mem_ctl.scala 582:35]
  wire  _T_3740 = ~_T_3732[6]; // @[lib.scala 195:55]
  wire  _T_3741 = _T_3734 & _T_3740; // @[lib.scala 195:53]
  wire  _T_3355 = ~_T_3347[6]; // @[lib.scala 195:55]
  wire  _T_3356 = _T_3349 & _T_3355; // @[lib.scala 195:53]
  wire [1:0] iccm_double_ecc_error = {_T_3741,_T_3356}; // @[Cat.scala 29:58]
  wire  iccm_dma_ecc_error_in = |iccm_double_ecc_error; // @[ifu_mem_ctl.scala 584:53]
  wire [63:0] _T_3104 = {io_dma_mem_ctl_dma_mem_addr,io_dma_mem_ctl_dma_mem_addr}; // @[Cat.scala 29:58]
  wire [63:0] _T_3105 = {iccm_dma_rdata_1_muxed,_T_3497[37:32],_T_3497[30:16],_T_3497[14:8],_T_3497[6:4],_T_3497[2]}; // @[Cat.scala 29:58]
  reg [2:0] dma_mem_tag_ff; // @[ifu_mem_ctl.scala 586:54]
  reg [2:0] iccm_dma_rtag_temp; // @[ifu_mem_ctl.scala 587:74]
  reg  iccm_dma_rvalid_temp; // @[ifu_mem_ctl.scala 592:76]
  reg  iccm_dma_ecc_error; // @[ifu_mem_ctl.scala 594:74]
  reg [63:0] iccm_dma_rdata_temp; // @[ifu_mem_ctl.scala 596:75]
  wire  _T_3110 = _T_2709 & _T_2698; // @[ifu_mem_ctl.scala 599:77]
  wire  _T_3114 = _T_3091 & iccm_correct_ecc; // @[ifu_mem_ctl.scala 600:62]
  reg [13:0] iccm_ecc_corr_index_ff; // @[Reg.scala 27:20]
  wire [14:0] _T_3115 = {iccm_ecc_corr_index_ff,1'h0}; // @[Cat.scala 29:58]
  wire [14:0] _T_3117 = _T_3114 ? _T_3115 : io_ifc_fetch_addr_bf[14:0]; // @[ifu_mem_ctl.scala 600:8]
  wire  _T_3509 = _T_3347 == 7'h40; // @[lib.scala 205:62]
  wire  _T_3510 = _T_3497[38] ^ _T_3509; // @[lib.scala 205:44]
  wire [6:0] iccm_corrected_ecc_0 = {_T_3510,_T_3497[31],_T_3497[15],_T_3497[7],_T_3497[3],_T_3497[1:0]}; // @[Cat.scala 29:58]
  wire  _T_3894 = _T_3732 == 7'h40; // @[lib.scala 205:62]
  wire  _T_3895 = _T_3882[38] ^ _T_3894; // @[lib.scala 205:44]
  wire [6:0] iccm_corrected_ecc_1 = {_T_3895,_T_3882[31],_T_3882[15],_T_3882[7],_T_3882[3],_T_3882[1:0]}; // @[Cat.scala 29:58]
  wire  _T_3911 = _T_3 & ifc_iccm_access_f; // @[ifu_mem_ctl.scala 612:75]
  wire [31:0] iccm_corrected_data_f_mux = iccm_single_ecc_error[0] ? iccm_corrected_data_0 : iccm_corrected_data_1; // @[ifu_mem_ctl.scala 614:38]
  wire [6:0] iccm_corrected_ecc_f_mux = iccm_single_ecc_error[0] ? iccm_corrected_ecc_0 : iccm_corrected_ecc_1; // @[ifu_mem_ctl.scala 615:37]
  reg  iccm_rd_ecc_single_err_ff; // @[ifu_mem_ctl.scala 623:62]
  wire  _T_3919 = ~iccm_rd_ecc_single_err_ff; // @[ifu_mem_ctl.scala 617:93]
  wire  _T_3920 = io_dec_mem_ctrl_ifu_iccm_rd_ecc_single_err & _T_3919; // @[ifu_mem_ctl.scala 617:91]
  wire  _T_3922 = _T_3920 & _T_319; // @[ifu_mem_ctl.scala 617:121]
  wire  iccm_ecc_write_status = _T_3922 | io_iccm_dma_sb_error; // @[ifu_mem_ctl.scala 617:144]
  wire  _T_3923 = io_dec_mem_ctrl_ifu_iccm_rd_ecc_single_err | iccm_rd_ecc_single_err_ff; // @[ifu_mem_ctl.scala 618:84]
  reg [13:0] iccm_rw_addr_f; // @[ifu_mem_ctl.scala 622:51]
  wire [13:0] _T_3928 = iccm_rw_addr_f + 14'h1; // @[ifu_mem_ctl.scala 621:102]
  wire [38:0] _T_3932 = {iccm_corrected_ecc_f_mux,iccm_corrected_data_f_mux}; // @[Cat.scala 29:58]
  wire  _T_3937 = ~io_ifc_fetch_uncacheable_bf; // @[ifu_mem_ctl.scala 626:41]
  wire  _T_3938 = io_ifc_fetch_req_bf & _T_3937; // @[ifu_mem_ctl.scala 626:39]
  wire  _T_3939 = ~io_ifc_iccm_access_bf; // @[ifu_mem_ctl.scala 626:72]
  wire  _T_3940 = _T_3938 & _T_3939; // @[ifu_mem_ctl.scala 626:70]
  wire  _T_3942 = ~miss_state_en; // @[ifu_mem_ctl.scala 627:34]
  wire  _T_3943 = _T_2268 & _T_3942; // @[ifu_mem_ctl.scala 627:32]
  wire  _T_3946 = _T_2284 & _T_3942; // @[ifu_mem_ctl.scala 628:37]
  wire  _T_3947 = _T_3943 | _T_3946; // @[ifu_mem_ctl.scala 627:88]
  wire  _T_3948 = miss_state == 3'h7; // @[ifu_mem_ctl.scala 629:19]
  wire  _T_3950 = _T_3948 & _T_3942; // @[ifu_mem_ctl.scala 629:41]
  wire  _T_3951 = _T_3947 | _T_3950; // @[ifu_mem_ctl.scala 628:88]
  wire  _T_3952 = miss_state == 3'h3; // @[ifu_mem_ctl.scala 630:19]
  wire  _T_3954 = _T_3952 & _T_3942; // @[ifu_mem_ctl.scala 630:35]
  wire  _T_3955 = _T_3951 | _T_3954; // @[ifu_mem_ctl.scala 629:88]
  wire  _T_3958 = _T_2283 & _T_3942; // @[ifu_mem_ctl.scala 631:38]
  wire  _T_3959 = _T_3955 | _T_3958; // @[ifu_mem_ctl.scala 630:88]
  wire  _T_3961 = _T_2284 & miss_state_en; // @[ifu_mem_ctl.scala 632:37]
  wire  _T_3962 = miss_nxtstate == 3'h3; // @[ifu_mem_ctl.scala 632:71]
  wire  _T_3963 = _T_3961 & _T_3962; // @[ifu_mem_ctl.scala 632:54]
  wire  _T_3964 = _T_3959 | _T_3963; // @[ifu_mem_ctl.scala 631:57]
  wire  _T_3965 = ~_T_3964; // @[ifu_mem_ctl.scala 627:5]
  wire  _T_3966 = _T_3940 & _T_3965; // @[ifu_mem_ctl.scala 626:96]
  wire  _T_3967 = io_ifc_fetch_req_bf & io_exu_flush_final; // @[ifu_mem_ctl.scala 633:28]
  wire  _T_3969 = _T_3967 & _T_3937; // @[ifu_mem_ctl.scala 633:50]
  wire  _T_3971 = _T_3969 & _T_3939; // @[ifu_mem_ctl.scala 633:81]
  wire  _T_3992 = reset_ic_in | reset_ic_ff; // @[ifu_mem_ctl.scala 639:64]
  wire  _T_3993 = ~_T_3992; // @[ifu_mem_ctl.scala 639:50]
  wire  ic_valid = _T_3993 & _T_339; // @[ifu_mem_ctl.scala 639:79]
  wire  _T_3997 = debug_c1_clken & io_ic_debug_tag_array; // @[ifu_mem_ctl.scala 640:82]
  reg [6:0] ifu_status_wr_addr_ff; // @[ifu_mem_ctl.scala 643:14]
  wire  _T_4000 = io_ic_debug_wr_en & io_ic_debug_tag_array; // @[ifu_mem_ctl.scala 646:74]
  reg  way_status_wr_en_ff; // @[ifu_mem_ctl.scala 648:14]
  wire  way_status_hit_new = io_ic_rd_hit[0]; // @[ifu_mem_ctl.scala 722:41]
  reg  way_status_new_ff; // @[ifu_mem_ctl.scala 654:14]
  wire  _T_4020 = ifu_status_wr_addr_ff[2:0] == 3'h0; // @[ifu_mem_ctl.scala 660:128]
  wire  _T_4021 = _T_4020 & way_status_wr_en_ff; // @[ifu_mem_ctl.scala 660:136]
  wire  _T_4024 = ifu_status_wr_addr_ff[2:0] == 3'h1; // @[ifu_mem_ctl.scala 660:128]
  wire  _T_4025 = _T_4024 & way_status_wr_en_ff; // @[ifu_mem_ctl.scala 660:136]
  wire  _T_4028 = ifu_status_wr_addr_ff[2:0] == 3'h2; // @[ifu_mem_ctl.scala 660:128]
  wire  _T_4029 = _T_4028 & way_status_wr_en_ff; // @[ifu_mem_ctl.scala 660:136]
  wire  _T_4032 = ifu_status_wr_addr_ff[2:0] == 3'h3; // @[ifu_mem_ctl.scala 660:128]
  wire  _T_4033 = _T_4032 & way_status_wr_en_ff; // @[ifu_mem_ctl.scala 660:136]
  wire  _T_4036 = ifu_status_wr_addr_ff[2:0] == 3'h4; // @[ifu_mem_ctl.scala 660:128]
  wire  _T_4037 = _T_4036 & way_status_wr_en_ff; // @[ifu_mem_ctl.scala 660:136]
  wire  _T_4040 = ifu_status_wr_addr_ff[2:0] == 3'h5; // @[ifu_mem_ctl.scala 660:128]
  wire  _T_4041 = _T_4040 & way_status_wr_en_ff; // @[ifu_mem_ctl.scala 660:136]
  wire  _T_4044 = ifu_status_wr_addr_ff[2:0] == 3'h6; // @[ifu_mem_ctl.scala 660:128]
  wire  _T_4045 = _T_4044 & way_status_wr_en_ff; // @[ifu_mem_ctl.scala 660:136]
  wire  _T_4048 = ifu_status_wr_addr_ff[2:0] == 3'h7; // @[ifu_mem_ctl.scala 660:128]
  wire  _T_4049 = _T_4048 & way_status_wr_en_ff; // @[ifu_mem_ctl.scala 660:136]
  wire  wren_reset_miss_1 = replace_way_mb_any_1 & reset_tag_valid_for_miss; // @[ifu_mem_ctl.scala 730:84]
  wire  wren_reset_miss_0 = replace_way_mb_any_0 & reset_tag_valid_for_miss; // @[ifu_mem_ctl.scala 730:84]
  wire [1:0] ifu_tag_wren = {wren_reset_miss_1,wren_reset_miss_0}; // @[Cat.scala 29:58]
  wire [1:0] _T_9821 = _T_4000 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [1:0] ic_debug_tag_wr_en = _T_9821 & io_ic_debug_way; // @[ifu_mem_ctl.scala 765:90]
  reg [1:0] ifu_tag_wren_ff; // @[ifu_mem_ctl.scala 675:14]
  reg  ic_valid_ff; // @[ifu_mem_ctl.scala 679:14]
  wire  _T_5063 = ifu_ic_rw_int_addr_ff[6:5] == 2'h0; // @[ifu_mem_ctl.scala 683:78]
  wire  _T_5065 = _T_5063 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 683:87]
  wire  _T_5067 = perr_ic_index_ff[6:5] == 2'h0; // @[ifu_mem_ctl.scala 684:70]
  wire  _T_5069 = _T_5067 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 684:79]
  wire  _T_5070 = _T_5065 | _T_5069; // @[ifu_mem_ctl.scala 683:109]
  wire  _T_5071 = _T_5070 | reset_all_tags; // @[ifu_mem_ctl.scala 684:102]
  wire  _T_5075 = _T_5063 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 683:87]
  wire  _T_5079 = _T_5067 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 684:79]
  wire  _T_5080 = _T_5075 | _T_5079; // @[ifu_mem_ctl.scala 683:109]
  wire  _T_5081 = _T_5080 | reset_all_tags; // @[ifu_mem_ctl.scala 684:102]
  wire [1:0] tag_valid_clken_0 = {_T_5081,_T_5071}; // @[Cat.scala 29:58]
  wire  _T_5083 = ifu_ic_rw_int_addr_ff[6:5] == 2'h1; // @[ifu_mem_ctl.scala 683:78]
  wire  _T_5085 = _T_5083 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 683:87]
  wire  _T_5087 = perr_ic_index_ff[6:5] == 2'h1; // @[ifu_mem_ctl.scala 684:70]
  wire  _T_5089 = _T_5087 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 684:79]
  wire  _T_5090 = _T_5085 | _T_5089; // @[ifu_mem_ctl.scala 683:109]
  wire  _T_5091 = _T_5090 | reset_all_tags; // @[ifu_mem_ctl.scala 684:102]
  wire  _T_5095 = _T_5083 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 683:87]
  wire  _T_5099 = _T_5087 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 684:79]
  wire  _T_5100 = _T_5095 | _T_5099; // @[ifu_mem_ctl.scala 683:109]
  wire  _T_5101 = _T_5100 | reset_all_tags; // @[ifu_mem_ctl.scala 684:102]
  wire [1:0] tag_valid_clken_1 = {_T_5101,_T_5091}; // @[Cat.scala 29:58]
  wire  _T_5103 = ifu_ic_rw_int_addr_ff[6:5] == 2'h2; // @[ifu_mem_ctl.scala 683:78]
  wire  _T_5105 = _T_5103 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 683:87]
  wire  _T_5107 = perr_ic_index_ff[6:5] == 2'h2; // @[ifu_mem_ctl.scala 684:70]
  wire  _T_5109 = _T_5107 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 684:79]
  wire  _T_5110 = _T_5105 | _T_5109; // @[ifu_mem_ctl.scala 683:109]
  wire  _T_5111 = _T_5110 | reset_all_tags; // @[ifu_mem_ctl.scala 684:102]
  wire  _T_5115 = _T_5103 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 683:87]
  wire  _T_5119 = _T_5107 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 684:79]
  wire  _T_5120 = _T_5115 | _T_5119; // @[ifu_mem_ctl.scala 683:109]
  wire  _T_5121 = _T_5120 | reset_all_tags; // @[ifu_mem_ctl.scala 684:102]
  wire [1:0] tag_valid_clken_2 = {_T_5121,_T_5111}; // @[Cat.scala 29:58]
  wire  _T_5123 = ifu_ic_rw_int_addr_ff[6:5] == 2'h3; // @[ifu_mem_ctl.scala 683:78]
  wire  _T_5125 = _T_5123 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 683:87]
  wire  _T_5127 = perr_ic_index_ff[6:5] == 2'h3; // @[ifu_mem_ctl.scala 684:70]
  wire  _T_5129 = _T_5127 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 684:79]
  wire  _T_5130 = _T_5125 | _T_5129; // @[ifu_mem_ctl.scala 683:109]
  wire  _T_5131 = _T_5130 | reset_all_tags; // @[ifu_mem_ctl.scala 684:102]
  wire  _T_5135 = _T_5123 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 683:87]
  wire  _T_5139 = _T_5127 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 684:79]
  wire  _T_5140 = _T_5135 | _T_5139; // @[ifu_mem_ctl.scala 683:109]
  wire  _T_5141 = _T_5140 | reset_all_tags; // @[ifu_mem_ctl.scala 684:102]
  wire [1:0] tag_valid_clken_3 = {_T_5141,_T_5131}; // @[Cat.scala 29:58]
  wire  _T_5152 = ic_valid_ff & _T_195; // @[ifu_mem_ctl.scala 692:97]
  wire  _T_5153 = ~perr_sel_invalidate; // @[ifu_mem_ctl.scala 692:124]
  wire  _T_5154 = _T_5152 & _T_5153; // @[ifu_mem_ctl.scala 692:122]
  wire  _T_5157 = _T_4671 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_5158 = perr_ic_index_ff == 7'h0; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_5160 = _T_5158 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_5161 = _T_5157 | _T_5160; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_5162 = _T_5161 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_5172 = _T_4672 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_5173 = perr_ic_index_ff == 7'h1; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_5175 = _T_5173 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_5176 = _T_5172 | _T_5175; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_5177 = _T_5176 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_5187 = _T_4673 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_5188 = perr_ic_index_ff == 7'h2; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_5190 = _T_5188 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_5191 = _T_5187 | _T_5190; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_5192 = _T_5191 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_5202 = _T_4674 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_5203 = perr_ic_index_ff == 7'h3; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_5205 = _T_5203 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_5206 = _T_5202 | _T_5205; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_5207 = _T_5206 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_5217 = _T_4675 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_5218 = perr_ic_index_ff == 7'h4; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_5220 = _T_5218 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_5221 = _T_5217 | _T_5220; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_5222 = _T_5221 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_5232 = _T_4676 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_5233 = perr_ic_index_ff == 7'h5; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_5235 = _T_5233 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_5236 = _T_5232 | _T_5235; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_5237 = _T_5236 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_5247 = _T_4677 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_5248 = perr_ic_index_ff == 7'h6; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_5250 = _T_5248 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_5251 = _T_5247 | _T_5250; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_5252 = _T_5251 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_5262 = _T_4678 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_5263 = perr_ic_index_ff == 7'h7; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_5265 = _T_5263 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_5266 = _T_5262 | _T_5265; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_5267 = _T_5266 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_5277 = _T_4679 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_5278 = perr_ic_index_ff == 7'h8; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_5280 = _T_5278 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_5281 = _T_5277 | _T_5280; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_5282 = _T_5281 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_5292 = _T_4680 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_5293 = perr_ic_index_ff == 7'h9; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_5295 = _T_5293 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_5296 = _T_5292 | _T_5295; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_5297 = _T_5296 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_5307 = _T_4681 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_5308 = perr_ic_index_ff == 7'ha; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_5310 = _T_5308 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_5311 = _T_5307 | _T_5310; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_5312 = _T_5311 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_5322 = _T_4682 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_5323 = perr_ic_index_ff == 7'hb; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_5325 = _T_5323 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_5326 = _T_5322 | _T_5325; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_5327 = _T_5326 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_5337 = _T_4683 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_5338 = perr_ic_index_ff == 7'hc; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_5340 = _T_5338 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_5341 = _T_5337 | _T_5340; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_5342 = _T_5341 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_5352 = _T_4684 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_5353 = perr_ic_index_ff == 7'hd; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_5355 = _T_5353 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_5356 = _T_5352 | _T_5355; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_5357 = _T_5356 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_5367 = _T_4685 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_5368 = perr_ic_index_ff == 7'he; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_5370 = _T_5368 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_5371 = _T_5367 | _T_5370; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_5372 = _T_5371 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_5382 = _T_4686 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_5383 = perr_ic_index_ff == 7'hf; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_5385 = _T_5383 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_5386 = _T_5382 | _T_5385; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_5387 = _T_5386 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_5397 = _T_4687 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_5398 = perr_ic_index_ff == 7'h10; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_5400 = _T_5398 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_5401 = _T_5397 | _T_5400; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_5402 = _T_5401 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_5412 = _T_4688 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_5413 = perr_ic_index_ff == 7'h11; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_5415 = _T_5413 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_5416 = _T_5412 | _T_5415; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_5417 = _T_5416 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_5427 = _T_4689 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_5428 = perr_ic_index_ff == 7'h12; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_5430 = _T_5428 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_5431 = _T_5427 | _T_5430; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_5432 = _T_5431 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_5442 = _T_4690 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_5443 = perr_ic_index_ff == 7'h13; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_5445 = _T_5443 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_5446 = _T_5442 | _T_5445; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_5447 = _T_5446 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_5457 = _T_4691 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_5458 = perr_ic_index_ff == 7'h14; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_5460 = _T_5458 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_5461 = _T_5457 | _T_5460; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_5462 = _T_5461 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_5472 = _T_4692 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_5473 = perr_ic_index_ff == 7'h15; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_5475 = _T_5473 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_5476 = _T_5472 | _T_5475; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_5477 = _T_5476 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_5487 = _T_4693 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_5488 = perr_ic_index_ff == 7'h16; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_5490 = _T_5488 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_5491 = _T_5487 | _T_5490; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_5492 = _T_5491 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_5502 = _T_4694 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_5503 = perr_ic_index_ff == 7'h17; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_5505 = _T_5503 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_5506 = _T_5502 | _T_5505; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_5507 = _T_5506 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_5517 = _T_4695 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_5518 = perr_ic_index_ff == 7'h18; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_5520 = _T_5518 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_5521 = _T_5517 | _T_5520; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_5522 = _T_5521 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_5532 = _T_4696 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_5533 = perr_ic_index_ff == 7'h19; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_5535 = _T_5533 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_5536 = _T_5532 | _T_5535; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_5537 = _T_5536 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_5547 = _T_4697 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_5548 = perr_ic_index_ff == 7'h1a; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_5550 = _T_5548 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_5551 = _T_5547 | _T_5550; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_5552 = _T_5551 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_5562 = _T_4698 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_5563 = perr_ic_index_ff == 7'h1b; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_5565 = _T_5563 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_5566 = _T_5562 | _T_5565; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_5567 = _T_5566 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_5577 = _T_4699 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_5578 = perr_ic_index_ff == 7'h1c; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_5580 = _T_5578 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_5581 = _T_5577 | _T_5580; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_5582 = _T_5581 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_5592 = _T_4700 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_5593 = perr_ic_index_ff == 7'h1d; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_5595 = _T_5593 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_5596 = _T_5592 | _T_5595; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_5597 = _T_5596 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_5607 = _T_4701 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_5608 = perr_ic_index_ff == 7'h1e; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_5610 = _T_5608 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_5611 = _T_5607 | _T_5610; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_5612 = _T_5611 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_5622 = _T_4702 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_5623 = perr_ic_index_ff == 7'h1f; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_5625 = _T_5623 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_5626 = _T_5622 | _T_5625; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_5627 = _T_5626 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_5637 = _T_4671 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_5640 = _T_5158 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_5641 = _T_5637 | _T_5640; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_5642 = _T_5641 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_5652 = _T_4672 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_5655 = _T_5173 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_5656 = _T_5652 | _T_5655; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_5657 = _T_5656 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_5667 = _T_4673 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_5670 = _T_5188 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_5671 = _T_5667 | _T_5670; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_5672 = _T_5671 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_5682 = _T_4674 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_5685 = _T_5203 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_5686 = _T_5682 | _T_5685; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_5687 = _T_5686 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_5697 = _T_4675 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_5700 = _T_5218 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_5701 = _T_5697 | _T_5700; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_5702 = _T_5701 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_5712 = _T_4676 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_5715 = _T_5233 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_5716 = _T_5712 | _T_5715; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_5717 = _T_5716 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_5727 = _T_4677 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_5730 = _T_5248 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_5731 = _T_5727 | _T_5730; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_5732 = _T_5731 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_5742 = _T_4678 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_5745 = _T_5263 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_5746 = _T_5742 | _T_5745; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_5747 = _T_5746 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_5757 = _T_4679 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_5760 = _T_5278 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_5761 = _T_5757 | _T_5760; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_5762 = _T_5761 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_5772 = _T_4680 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_5775 = _T_5293 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_5776 = _T_5772 | _T_5775; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_5777 = _T_5776 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_5787 = _T_4681 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_5790 = _T_5308 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_5791 = _T_5787 | _T_5790; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_5792 = _T_5791 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_5802 = _T_4682 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_5805 = _T_5323 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_5806 = _T_5802 | _T_5805; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_5807 = _T_5806 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_5817 = _T_4683 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_5820 = _T_5338 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_5821 = _T_5817 | _T_5820; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_5822 = _T_5821 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_5832 = _T_4684 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_5835 = _T_5353 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_5836 = _T_5832 | _T_5835; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_5837 = _T_5836 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_5847 = _T_4685 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_5850 = _T_5368 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_5851 = _T_5847 | _T_5850; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_5852 = _T_5851 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_5862 = _T_4686 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_5865 = _T_5383 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_5866 = _T_5862 | _T_5865; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_5867 = _T_5866 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_5877 = _T_4687 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_5880 = _T_5398 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_5881 = _T_5877 | _T_5880; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_5882 = _T_5881 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_5892 = _T_4688 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_5895 = _T_5413 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_5896 = _T_5892 | _T_5895; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_5897 = _T_5896 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_5907 = _T_4689 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_5910 = _T_5428 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_5911 = _T_5907 | _T_5910; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_5912 = _T_5911 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_5922 = _T_4690 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_5925 = _T_5443 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_5926 = _T_5922 | _T_5925; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_5927 = _T_5926 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_5937 = _T_4691 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_5940 = _T_5458 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_5941 = _T_5937 | _T_5940; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_5942 = _T_5941 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_5952 = _T_4692 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_5955 = _T_5473 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_5956 = _T_5952 | _T_5955; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_5957 = _T_5956 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_5967 = _T_4693 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_5970 = _T_5488 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_5971 = _T_5967 | _T_5970; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_5972 = _T_5971 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_5982 = _T_4694 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_5985 = _T_5503 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_5986 = _T_5982 | _T_5985; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_5987 = _T_5986 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_5997 = _T_4695 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6000 = _T_5518 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6001 = _T_5997 | _T_6000; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6002 = _T_6001 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6012 = _T_4696 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6015 = _T_5533 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6016 = _T_6012 | _T_6015; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6017 = _T_6016 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6027 = _T_4697 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6030 = _T_5548 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6031 = _T_6027 | _T_6030; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6032 = _T_6031 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6042 = _T_4698 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6045 = _T_5563 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6046 = _T_6042 | _T_6045; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6047 = _T_6046 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6057 = _T_4699 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6060 = _T_5578 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6061 = _T_6057 | _T_6060; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6062 = _T_6061 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6072 = _T_4700 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6075 = _T_5593 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6076 = _T_6072 | _T_6075; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6077 = _T_6076 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6087 = _T_4701 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6090 = _T_5608 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6091 = _T_6087 | _T_6090; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6092 = _T_6091 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6102 = _T_4702 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6105 = _T_5623 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6106 = _T_6102 | _T_6105; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6107 = _T_6106 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6117 = _T_4703 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6118 = perr_ic_index_ff == 7'h20; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_6120 = _T_6118 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6121 = _T_6117 | _T_6120; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6122 = _T_6121 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6132 = _T_4704 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6133 = perr_ic_index_ff == 7'h21; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_6135 = _T_6133 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6136 = _T_6132 | _T_6135; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6137 = _T_6136 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6147 = _T_4705 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6148 = perr_ic_index_ff == 7'h22; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_6150 = _T_6148 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6151 = _T_6147 | _T_6150; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6152 = _T_6151 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6162 = _T_4706 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6163 = perr_ic_index_ff == 7'h23; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_6165 = _T_6163 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6166 = _T_6162 | _T_6165; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6167 = _T_6166 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6177 = _T_4707 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6178 = perr_ic_index_ff == 7'h24; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_6180 = _T_6178 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6181 = _T_6177 | _T_6180; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6182 = _T_6181 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6192 = _T_4708 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6193 = perr_ic_index_ff == 7'h25; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_6195 = _T_6193 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6196 = _T_6192 | _T_6195; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6197 = _T_6196 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6207 = _T_4709 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6208 = perr_ic_index_ff == 7'h26; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_6210 = _T_6208 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6211 = _T_6207 | _T_6210; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6212 = _T_6211 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6222 = _T_4710 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6223 = perr_ic_index_ff == 7'h27; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_6225 = _T_6223 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6226 = _T_6222 | _T_6225; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6227 = _T_6226 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6237 = _T_4711 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6238 = perr_ic_index_ff == 7'h28; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_6240 = _T_6238 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6241 = _T_6237 | _T_6240; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6242 = _T_6241 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6252 = _T_4712 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6253 = perr_ic_index_ff == 7'h29; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_6255 = _T_6253 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6256 = _T_6252 | _T_6255; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6257 = _T_6256 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6267 = _T_4713 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6268 = perr_ic_index_ff == 7'h2a; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_6270 = _T_6268 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6271 = _T_6267 | _T_6270; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6272 = _T_6271 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6282 = _T_4714 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6283 = perr_ic_index_ff == 7'h2b; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_6285 = _T_6283 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6286 = _T_6282 | _T_6285; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6287 = _T_6286 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6297 = _T_4715 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6298 = perr_ic_index_ff == 7'h2c; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_6300 = _T_6298 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6301 = _T_6297 | _T_6300; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6302 = _T_6301 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6312 = _T_4716 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6313 = perr_ic_index_ff == 7'h2d; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_6315 = _T_6313 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6316 = _T_6312 | _T_6315; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6317 = _T_6316 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6327 = _T_4717 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6328 = perr_ic_index_ff == 7'h2e; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_6330 = _T_6328 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6331 = _T_6327 | _T_6330; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6332 = _T_6331 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6342 = _T_4718 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6343 = perr_ic_index_ff == 7'h2f; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_6345 = _T_6343 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6346 = _T_6342 | _T_6345; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6347 = _T_6346 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6357 = _T_4719 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6358 = perr_ic_index_ff == 7'h30; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_6360 = _T_6358 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6361 = _T_6357 | _T_6360; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6362 = _T_6361 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6372 = _T_4720 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6373 = perr_ic_index_ff == 7'h31; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_6375 = _T_6373 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6376 = _T_6372 | _T_6375; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6377 = _T_6376 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6387 = _T_4721 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6388 = perr_ic_index_ff == 7'h32; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_6390 = _T_6388 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6391 = _T_6387 | _T_6390; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6392 = _T_6391 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6402 = _T_4722 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6403 = perr_ic_index_ff == 7'h33; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_6405 = _T_6403 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6406 = _T_6402 | _T_6405; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6407 = _T_6406 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6417 = _T_4723 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6418 = perr_ic_index_ff == 7'h34; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_6420 = _T_6418 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6421 = _T_6417 | _T_6420; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6422 = _T_6421 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6432 = _T_4724 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6433 = perr_ic_index_ff == 7'h35; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_6435 = _T_6433 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6436 = _T_6432 | _T_6435; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6437 = _T_6436 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6447 = _T_4725 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6448 = perr_ic_index_ff == 7'h36; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_6450 = _T_6448 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6451 = _T_6447 | _T_6450; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6452 = _T_6451 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6462 = _T_4726 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6463 = perr_ic_index_ff == 7'h37; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_6465 = _T_6463 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6466 = _T_6462 | _T_6465; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6467 = _T_6466 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6477 = _T_4727 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6478 = perr_ic_index_ff == 7'h38; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_6480 = _T_6478 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6481 = _T_6477 | _T_6480; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6482 = _T_6481 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6492 = _T_4728 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6493 = perr_ic_index_ff == 7'h39; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_6495 = _T_6493 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6496 = _T_6492 | _T_6495; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6497 = _T_6496 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6507 = _T_4729 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6508 = perr_ic_index_ff == 7'h3a; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_6510 = _T_6508 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6511 = _T_6507 | _T_6510; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6512 = _T_6511 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6522 = _T_4730 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6523 = perr_ic_index_ff == 7'h3b; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_6525 = _T_6523 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6526 = _T_6522 | _T_6525; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6527 = _T_6526 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6537 = _T_4731 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6538 = perr_ic_index_ff == 7'h3c; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_6540 = _T_6538 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6541 = _T_6537 | _T_6540; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6542 = _T_6541 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6552 = _T_4732 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6553 = perr_ic_index_ff == 7'h3d; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_6555 = _T_6553 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6556 = _T_6552 | _T_6555; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6557 = _T_6556 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6567 = _T_4733 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6568 = perr_ic_index_ff == 7'h3e; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_6570 = _T_6568 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6571 = _T_6567 | _T_6570; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6572 = _T_6571 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6582 = _T_4734 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6583 = perr_ic_index_ff == 7'h3f; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_6585 = _T_6583 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6586 = _T_6582 | _T_6585; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6587 = _T_6586 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6597 = _T_4703 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6600 = _T_6118 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6601 = _T_6597 | _T_6600; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6602 = _T_6601 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6612 = _T_4704 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6615 = _T_6133 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6616 = _T_6612 | _T_6615; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6617 = _T_6616 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6627 = _T_4705 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6630 = _T_6148 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6631 = _T_6627 | _T_6630; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6632 = _T_6631 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6642 = _T_4706 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6645 = _T_6163 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6646 = _T_6642 | _T_6645; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6647 = _T_6646 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6657 = _T_4707 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6660 = _T_6178 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6661 = _T_6657 | _T_6660; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6662 = _T_6661 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6672 = _T_4708 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6675 = _T_6193 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6676 = _T_6672 | _T_6675; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6677 = _T_6676 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6687 = _T_4709 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6690 = _T_6208 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6691 = _T_6687 | _T_6690; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6692 = _T_6691 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6702 = _T_4710 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6705 = _T_6223 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6706 = _T_6702 | _T_6705; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6707 = _T_6706 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6717 = _T_4711 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6720 = _T_6238 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6721 = _T_6717 | _T_6720; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6722 = _T_6721 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6732 = _T_4712 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6735 = _T_6253 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6736 = _T_6732 | _T_6735; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6737 = _T_6736 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6747 = _T_4713 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6750 = _T_6268 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6751 = _T_6747 | _T_6750; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6752 = _T_6751 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6762 = _T_4714 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6765 = _T_6283 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6766 = _T_6762 | _T_6765; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6767 = _T_6766 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6777 = _T_4715 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6780 = _T_6298 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6781 = _T_6777 | _T_6780; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6782 = _T_6781 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6792 = _T_4716 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6795 = _T_6313 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6796 = _T_6792 | _T_6795; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6797 = _T_6796 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6807 = _T_4717 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6810 = _T_6328 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6811 = _T_6807 | _T_6810; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6812 = _T_6811 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6822 = _T_4718 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6825 = _T_6343 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6826 = _T_6822 | _T_6825; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6827 = _T_6826 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6837 = _T_4719 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6840 = _T_6358 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6841 = _T_6837 | _T_6840; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6842 = _T_6841 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6852 = _T_4720 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6855 = _T_6373 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6856 = _T_6852 | _T_6855; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6857 = _T_6856 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6867 = _T_4721 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6870 = _T_6388 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6871 = _T_6867 | _T_6870; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6872 = _T_6871 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6882 = _T_4722 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6885 = _T_6403 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6886 = _T_6882 | _T_6885; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6887 = _T_6886 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6897 = _T_4723 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6900 = _T_6418 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6901 = _T_6897 | _T_6900; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6902 = _T_6901 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6912 = _T_4724 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6915 = _T_6433 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6916 = _T_6912 | _T_6915; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6917 = _T_6916 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6927 = _T_4725 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6930 = _T_6448 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6931 = _T_6927 | _T_6930; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6932 = _T_6931 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6942 = _T_4726 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6945 = _T_6463 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6946 = _T_6942 | _T_6945; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6947 = _T_6946 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6957 = _T_4727 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6960 = _T_6478 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6961 = _T_6957 | _T_6960; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6962 = _T_6961 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6972 = _T_4728 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6975 = _T_6493 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6976 = _T_6972 | _T_6975; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6977 = _T_6976 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6987 = _T_4729 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6990 = _T_6508 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6991 = _T_6987 | _T_6990; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6992 = _T_6991 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7002 = _T_4730 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7005 = _T_6523 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7006 = _T_7002 | _T_7005; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7007 = _T_7006 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7017 = _T_4731 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7020 = _T_6538 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7021 = _T_7017 | _T_7020; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7022 = _T_7021 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7032 = _T_4732 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7035 = _T_6553 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7036 = _T_7032 | _T_7035; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7037 = _T_7036 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7047 = _T_4733 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7050 = _T_6568 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7051 = _T_7047 | _T_7050; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7052 = _T_7051 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7062 = _T_4734 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7065 = _T_6583 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7066 = _T_7062 | _T_7065; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7067 = _T_7066 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7077 = _T_4735 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7078 = perr_ic_index_ff == 7'h40; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_7080 = _T_7078 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7081 = _T_7077 | _T_7080; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7082 = _T_7081 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7092 = _T_4736 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7093 = perr_ic_index_ff == 7'h41; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_7095 = _T_7093 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7096 = _T_7092 | _T_7095; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7097 = _T_7096 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7107 = _T_4737 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7108 = perr_ic_index_ff == 7'h42; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_7110 = _T_7108 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7111 = _T_7107 | _T_7110; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7112 = _T_7111 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7122 = _T_4738 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7123 = perr_ic_index_ff == 7'h43; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_7125 = _T_7123 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7126 = _T_7122 | _T_7125; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7127 = _T_7126 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7137 = _T_4739 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7138 = perr_ic_index_ff == 7'h44; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_7140 = _T_7138 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7141 = _T_7137 | _T_7140; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7142 = _T_7141 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7152 = _T_4740 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7153 = perr_ic_index_ff == 7'h45; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_7155 = _T_7153 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7156 = _T_7152 | _T_7155; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7157 = _T_7156 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7167 = _T_4741 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7168 = perr_ic_index_ff == 7'h46; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_7170 = _T_7168 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7171 = _T_7167 | _T_7170; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7172 = _T_7171 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7182 = _T_4742 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7183 = perr_ic_index_ff == 7'h47; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_7185 = _T_7183 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7186 = _T_7182 | _T_7185; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7187 = _T_7186 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7197 = _T_4743 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7198 = perr_ic_index_ff == 7'h48; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_7200 = _T_7198 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7201 = _T_7197 | _T_7200; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7202 = _T_7201 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7212 = _T_4744 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7213 = perr_ic_index_ff == 7'h49; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_7215 = _T_7213 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7216 = _T_7212 | _T_7215; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7217 = _T_7216 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7227 = _T_4745 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7228 = perr_ic_index_ff == 7'h4a; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_7230 = _T_7228 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7231 = _T_7227 | _T_7230; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7232 = _T_7231 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7242 = _T_4746 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7243 = perr_ic_index_ff == 7'h4b; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_7245 = _T_7243 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7246 = _T_7242 | _T_7245; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7247 = _T_7246 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7257 = _T_4747 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7258 = perr_ic_index_ff == 7'h4c; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_7260 = _T_7258 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7261 = _T_7257 | _T_7260; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7262 = _T_7261 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7272 = _T_4748 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7273 = perr_ic_index_ff == 7'h4d; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_7275 = _T_7273 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7276 = _T_7272 | _T_7275; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7277 = _T_7276 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7287 = _T_4749 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7288 = perr_ic_index_ff == 7'h4e; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_7290 = _T_7288 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7291 = _T_7287 | _T_7290; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7292 = _T_7291 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7302 = _T_4750 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7303 = perr_ic_index_ff == 7'h4f; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_7305 = _T_7303 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7306 = _T_7302 | _T_7305; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7307 = _T_7306 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7317 = _T_4751 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7318 = perr_ic_index_ff == 7'h50; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_7320 = _T_7318 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7321 = _T_7317 | _T_7320; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7322 = _T_7321 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7332 = _T_4752 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7333 = perr_ic_index_ff == 7'h51; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_7335 = _T_7333 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7336 = _T_7332 | _T_7335; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7337 = _T_7336 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7347 = _T_4753 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7348 = perr_ic_index_ff == 7'h52; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_7350 = _T_7348 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7351 = _T_7347 | _T_7350; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7352 = _T_7351 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7362 = _T_4754 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7363 = perr_ic_index_ff == 7'h53; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_7365 = _T_7363 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7366 = _T_7362 | _T_7365; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7367 = _T_7366 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7377 = _T_4755 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7378 = perr_ic_index_ff == 7'h54; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_7380 = _T_7378 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7381 = _T_7377 | _T_7380; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7382 = _T_7381 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7392 = _T_4756 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7393 = perr_ic_index_ff == 7'h55; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_7395 = _T_7393 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7396 = _T_7392 | _T_7395; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7397 = _T_7396 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7407 = _T_4757 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7408 = perr_ic_index_ff == 7'h56; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_7410 = _T_7408 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7411 = _T_7407 | _T_7410; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7412 = _T_7411 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7422 = _T_4758 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7423 = perr_ic_index_ff == 7'h57; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_7425 = _T_7423 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7426 = _T_7422 | _T_7425; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7427 = _T_7426 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7437 = _T_4759 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7438 = perr_ic_index_ff == 7'h58; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_7440 = _T_7438 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7441 = _T_7437 | _T_7440; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7442 = _T_7441 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7452 = _T_4760 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7453 = perr_ic_index_ff == 7'h59; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_7455 = _T_7453 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7456 = _T_7452 | _T_7455; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7457 = _T_7456 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7467 = _T_4761 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7468 = perr_ic_index_ff == 7'h5a; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_7470 = _T_7468 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7471 = _T_7467 | _T_7470; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7472 = _T_7471 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7482 = _T_4762 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7483 = perr_ic_index_ff == 7'h5b; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_7485 = _T_7483 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7486 = _T_7482 | _T_7485; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7487 = _T_7486 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7497 = _T_4763 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7498 = perr_ic_index_ff == 7'h5c; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_7500 = _T_7498 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7501 = _T_7497 | _T_7500; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7502 = _T_7501 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7512 = _T_4764 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7513 = perr_ic_index_ff == 7'h5d; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_7515 = _T_7513 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7516 = _T_7512 | _T_7515; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7517 = _T_7516 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7527 = _T_4765 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7528 = perr_ic_index_ff == 7'h5e; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_7530 = _T_7528 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7531 = _T_7527 | _T_7530; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7532 = _T_7531 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7542 = _T_4766 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7543 = perr_ic_index_ff == 7'h5f; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_7545 = _T_7543 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7546 = _T_7542 | _T_7545; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7547 = _T_7546 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7557 = _T_4735 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7560 = _T_7078 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7561 = _T_7557 | _T_7560; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7562 = _T_7561 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7572 = _T_4736 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7575 = _T_7093 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7576 = _T_7572 | _T_7575; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7577 = _T_7576 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7587 = _T_4737 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7590 = _T_7108 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7591 = _T_7587 | _T_7590; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7592 = _T_7591 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7602 = _T_4738 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7605 = _T_7123 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7606 = _T_7602 | _T_7605; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7607 = _T_7606 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7617 = _T_4739 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7620 = _T_7138 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7621 = _T_7617 | _T_7620; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7622 = _T_7621 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7632 = _T_4740 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7635 = _T_7153 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7636 = _T_7632 | _T_7635; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7637 = _T_7636 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7647 = _T_4741 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7650 = _T_7168 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7651 = _T_7647 | _T_7650; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7652 = _T_7651 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7662 = _T_4742 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7665 = _T_7183 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7666 = _T_7662 | _T_7665; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7667 = _T_7666 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7677 = _T_4743 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7680 = _T_7198 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7681 = _T_7677 | _T_7680; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7682 = _T_7681 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7692 = _T_4744 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7695 = _T_7213 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7696 = _T_7692 | _T_7695; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7697 = _T_7696 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7707 = _T_4745 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7710 = _T_7228 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7711 = _T_7707 | _T_7710; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7712 = _T_7711 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7722 = _T_4746 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7725 = _T_7243 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7726 = _T_7722 | _T_7725; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7727 = _T_7726 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7737 = _T_4747 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7740 = _T_7258 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7741 = _T_7737 | _T_7740; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7742 = _T_7741 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7752 = _T_4748 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7755 = _T_7273 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7756 = _T_7752 | _T_7755; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7757 = _T_7756 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7767 = _T_4749 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7770 = _T_7288 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7771 = _T_7767 | _T_7770; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7772 = _T_7771 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7782 = _T_4750 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7785 = _T_7303 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7786 = _T_7782 | _T_7785; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7787 = _T_7786 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7797 = _T_4751 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7800 = _T_7318 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7801 = _T_7797 | _T_7800; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7802 = _T_7801 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7812 = _T_4752 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7815 = _T_7333 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7816 = _T_7812 | _T_7815; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7817 = _T_7816 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7827 = _T_4753 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7830 = _T_7348 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7831 = _T_7827 | _T_7830; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7832 = _T_7831 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7842 = _T_4754 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7845 = _T_7363 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7846 = _T_7842 | _T_7845; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7847 = _T_7846 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7857 = _T_4755 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7860 = _T_7378 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7861 = _T_7857 | _T_7860; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7862 = _T_7861 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7872 = _T_4756 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7875 = _T_7393 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7876 = _T_7872 | _T_7875; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7877 = _T_7876 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7887 = _T_4757 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7890 = _T_7408 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7891 = _T_7887 | _T_7890; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7892 = _T_7891 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7902 = _T_4758 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7905 = _T_7423 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7906 = _T_7902 | _T_7905; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7907 = _T_7906 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7917 = _T_4759 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7920 = _T_7438 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7921 = _T_7917 | _T_7920; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7922 = _T_7921 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7932 = _T_4760 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7935 = _T_7453 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7936 = _T_7932 | _T_7935; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7937 = _T_7936 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7947 = _T_4761 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7950 = _T_7468 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7951 = _T_7947 | _T_7950; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7952 = _T_7951 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7962 = _T_4762 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7965 = _T_7483 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7966 = _T_7962 | _T_7965; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7967 = _T_7966 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7977 = _T_4763 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7980 = _T_7498 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7981 = _T_7977 | _T_7980; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7982 = _T_7981 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7992 = _T_4764 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7995 = _T_7513 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7996 = _T_7992 | _T_7995; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7997 = _T_7996 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8007 = _T_4765 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8010 = _T_7528 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8011 = _T_8007 | _T_8010; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8012 = _T_8011 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8022 = _T_4766 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8025 = _T_7543 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8026 = _T_8022 | _T_8025; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8027 = _T_8026 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8037 = _T_4767 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8038 = perr_ic_index_ff == 7'h60; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_8040 = _T_8038 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8041 = _T_8037 | _T_8040; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8042 = _T_8041 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8052 = _T_4768 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8053 = perr_ic_index_ff == 7'h61; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_8055 = _T_8053 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8056 = _T_8052 | _T_8055; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8057 = _T_8056 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8067 = _T_4769 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8068 = perr_ic_index_ff == 7'h62; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_8070 = _T_8068 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8071 = _T_8067 | _T_8070; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8072 = _T_8071 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8082 = _T_4770 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8083 = perr_ic_index_ff == 7'h63; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_8085 = _T_8083 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8086 = _T_8082 | _T_8085; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8087 = _T_8086 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8097 = _T_4771 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8098 = perr_ic_index_ff == 7'h64; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_8100 = _T_8098 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8101 = _T_8097 | _T_8100; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8102 = _T_8101 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8112 = _T_4772 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8113 = perr_ic_index_ff == 7'h65; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_8115 = _T_8113 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8116 = _T_8112 | _T_8115; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8117 = _T_8116 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8127 = _T_4773 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8128 = perr_ic_index_ff == 7'h66; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_8130 = _T_8128 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8131 = _T_8127 | _T_8130; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8132 = _T_8131 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8142 = _T_4774 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8143 = perr_ic_index_ff == 7'h67; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_8145 = _T_8143 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8146 = _T_8142 | _T_8145; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8147 = _T_8146 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8157 = _T_4775 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8158 = perr_ic_index_ff == 7'h68; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_8160 = _T_8158 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8161 = _T_8157 | _T_8160; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8162 = _T_8161 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8172 = _T_4776 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8173 = perr_ic_index_ff == 7'h69; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_8175 = _T_8173 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8176 = _T_8172 | _T_8175; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8177 = _T_8176 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8187 = _T_4777 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8188 = perr_ic_index_ff == 7'h6a; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_8190 = _T_8188 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8191 = _T_8187 | _T_8190; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8192 = _T_8191 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8202 = _T_4778 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8203 = perr_ic_index_ff == 7'h6b; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_8205 = _T_8203 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8206 = _T_8202 | _T_8205; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8207 = _T_8206 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8217 = _T_4779 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8218 = perr_ic_index_ff == 7'h6c; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_8220 = _T_8218 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8221 = _T_8217 | _T_8220; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8222 = _T_8221 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8232 = _T_4780 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8233 = perr_ic_index_ff == 7'h6d; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_8235 = _T_8233 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8236 = _T_8232 | _T_8235; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8237 = _T_8236 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8247 = _T_4781 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8248 = perr_ic_index_ff == 7'h6e; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_8250 = _T_8248 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8251 = _T_8247 | _T_8250; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8252 = _T_8251 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8262 = _T_4782 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8263 = perr_ic_index_ff == 7'h6f; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_8265 = _T_8263 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8266 = _T_8262 | _T_8265; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8267 = _T_8266 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8277 = _T_4783 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8278 = perr_ic_index_ff == 7'h70; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_8280 = _T_8278 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8281 = _T_8277 | _T_8280; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8282 = _T_8281 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8292 = _T_4784 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8293 = perr_ic_index_ff == 7'h71; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_8295 = _T_8293 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8296 = _T_8292 | _T_8295; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8297 = _T_8296 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8307 = _T_4785 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8308 = perr_ic_index_ff == 7'h72; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_8310 = _T_8308 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8311 = _T_8307 | _T_8310; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8312 = _T_8311 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8322 = _T_4786 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8323 = perr_ic_index_ff == 7'h73; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_8325 = _T_8323 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8326 = _T_8322 | _T_8325; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8327 = _T_8326 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8337 = _T_4787 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8338 = perr_ic_index_ff == 7'h74; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_8340 = _T_8338 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8341 = _T_8337 | _T_8340; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8342 = _T_8341 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8352 = _T_4788 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8353 = perr_ic_index_ff == 7'h75; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_8355 = _T_8353 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8356 = _T_8352 | _T_8355; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8357 = _T_8356 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8367 = _T_4789 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8368 = perr_ic_index_ff == 7'h76; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_8370 = _T_8368 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8371 = _T_8367 | _T_8370; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8372 = _T_8371 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8382 = _T_4790 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8383 = perr_ic_index_ff == 7'h77; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_8385 = _T_8383 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8386 = _T_8382 | _T_8385; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8387 = _T_8386 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8397 = _T_4791 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8398 = perr_ic_index_ff == 7'h78; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_8400 = _T_8398 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8401 = _T_8397 | _T_8400; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8402 = _T_8401 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8412 = _T_4792 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8413 = perr_ic_index_ff == 7'h79; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_8415 = _T_8413 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8416 = _T_8412 | _T_8415; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8417 = _T_8416 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8427 = _T_4793 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8428 = perr_ic_index_ff == 7'h7a; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_8430 = _T_8428 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8431 = _T_8427 | _T_8430; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8432 = _T_8431 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8442 = _T_4794 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8443 = perr_ic_index_ff == 7'h7b; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_8445 = _T_8443 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8446 = _T_8442 | _T_8445; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8447 = _T_8446 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8457 = _T_4795 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8458 = perr_ic_index_ff == 7'h7c; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_8460 = _T_8458 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8461 = _T_8457 | _T_8460; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8462 = _T_8461 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8472 = _T_4796 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8473 = perr_ic_index_ff == 7'h7d; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_8475 = _T_8473 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8476 = _T_8472 | _T_8475; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8477 = _T_8476 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8487 = _T_4797 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8488 = perr_ic_index_ff == 7'h7e; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_8490 = _T_8488 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8491 = _T_8487 | _T_8490; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8492 = _T_8491 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8502 = _T_4798 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8503 = perr_ic_index_ff == 7'h7f; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_8505 = _T_8503 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8506 = _T_8502 | _T_8505; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8507 = _T_8506 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8517 = _T_4767 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8520 = _T_8038 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8521 = _T_8517 | _T_8520; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8522 = _T_8521 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8532 = _T_4768 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8535 = _T_8053 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8536 = _T_8532 | _T_8535; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8537 = _T_8536 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8547 = _T_4769 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8550 = _T_8068 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8551 = _T_8547 | _T_8550; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8552 = _T_8551 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8562 = _T_4770 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8565 = _T_8083 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8566 = _T_8562 | _T_8565; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8567 = _T_8566 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8577 = _T_4771 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8580 = _T_8098 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8581 = _T_8577 | _T_8580; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8582 = _T_8581 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8592 = _T_4772 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8595 = _T_8113 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8596 = _T_8592 | _T_8595; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8597 = _T_8596 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8607 = _T_4773 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8610 = _T_8128 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8611 = _T_8607 | _T_8610; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8612 = _T_8611 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8622 = _T_4774 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8625 = _T_8143 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8626 = _T_8622 | _T_8625; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8627 = _T_8626 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8637 = _T_4775 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8640 = _T_8158 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8641 = _T_8637 | _T_8640; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8642 = _T_8641 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8652 = _T_4776 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8655 = _T_8173 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8656 = _T_8652 | _T_8655; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8657 = _T_8656 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8667 = _T_4777 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8670 = _T_8188 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8671 = _T_8667 | _T_8670; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8672 = _T_8671 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8682 = _T_4778 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8685 = _T_8203 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8686 = _T_8682 | _T_8685; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8687 = _T_8686 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8697 = _T_4779 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8700 = _T_8218 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8701 = _T_8697 | _T_8700; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8702 = _T_8701 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8712 = _T_4780 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8715 = _T_8233 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8716 = _T_8712 | _T_8715; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8717 = _T_8716 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8727 = _T_4781 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8730 = _T_8248 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8731 = _T_8727 | _T_8730; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8732 = _T_8731 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8742 = _T_4782 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8745 = _T_8263 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8746 = _T_8742 | _T_8745; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8747 = _T_8746 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8757 = _T_4783 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8760 = _T_8278 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8761 = _T_8757 | _T_8760; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8762 = _T_8761 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8772 = _T_4784 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8775 = _T_8293 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8776 = _T_8772 | _T_8775; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8777 = _T_8776 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8787 = _T_4785 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8790 = _T_8308 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8791 = _T_8787 | _T_8790; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8792 = _T_8791 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8802 = _T_4786 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8805 = _T_8323 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8806 = _T_8802 | _T_8805; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8807 = _T_8806 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8817 = _T_4787 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8820 = _T_8338 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8821 = _T_8817 | _T_8820; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8822 = _T_8821 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8832 = _T_4788 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8835 = _T_8353 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8836 = _T_8832 | _T_8835; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8837 = _T_8836 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8847 = _T_4789 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8850 = _T_8368 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8851 = _T_8847 | _T_8850; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8852 = _T_8851 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8862 = _T_4790 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8865 = _T_8383 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8866 = _T_8862 | _T_8865; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8867 = _T_8866 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8877 = _T_4791 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8880 = _T_8398 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8881 = _T_8877 | _T_8880; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8882 = _T_8881 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8892 = _T_4792 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8895 = _T_8413 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8896 = _T_8892 | _T_8895; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8897 = _T_8896 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8907 = _T_4793 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8910 = _T_8428 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8911 = _T_8907 | _T_8910; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8912 = _T_8911 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8922 = _T_4794 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8925 = _T_8443 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8926 = _T_8922 | _T_8925; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8927 = _T_8926 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8937 = _T_4795 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8940 = _T_8458 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8941 = _T_8937 | _T_8940; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8942 = _T_8941 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8952 = _T_4796 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8955 = _T_8473 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8956 = _T_8952 | _T_8955; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8957 = _T_8956 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8967 = _T_4797 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8970 = _T_8488 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8971 = _T_8967 | _T_8970; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8972 = _T_8971 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8982 = _T_4798 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8985 = _T_8503 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8986 = _T_8982 | _T_8985; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8987 = _T_8986 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_9789 = ~fetch_uncacheable_ff; // @[ifu_mem_ctl.scala 747:63]
  wire  _T_9790 = _T_9789 & ifc_fetch_req_f; // @[ifu_mem_ctl.scala 747:85]
  wire [1:0] _T_9792 = _T_9790 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  reg  _T_9799; // @[ifu_mem_ctl.scala 752:70]
  reg  _T_9800; // @[ifu_mem_ctl.scala 753:69]
  reg  _T_9801; // @[ifu_mem_ctl.scala 754:72]
  reg  _T_9805; // @[ifu_mem_ctl.scala 755:71]
  wire  _T_9809 = io_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_dicawics[15:14] == 2'h3; // @[ifu_mem_ctl.scala 763:84]
  wire  _T_9811 = io_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_dicawics[15:14] == 2'h2; // @[ifu_mem_ctl.scala 763:150]
  wire  _T_9813 = io_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_dicawics[15:14] == 2'h1; // @[ifu_mem_ctl.scala 764:63]
  wire  _T_9815 = io_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_dicawics[15:14] == 2'h0; // @[ifu_mem_ctl.scala 764:129]
  wire [3:0] _T_9818 = {_T_9809,_T_9811,_T_9813,_T_9815}; // @[Cat.scala 29:58]
  reg  _T_9826; // @[ifu_mem_ctl.scala 770:79]
  wire [31:0] _T_9836 = {io_ifc_fetch_addr_bf,1'h0}; // @[Cat.scala 29:58]
  wire [31:0] _T_9837 = _T_9836 | 32'h7fffffff; // @[ifu_mem_ctl.scala 773:65]
  wire  _T_9839 = _T_9837 == 32'h7fffffff; // @[ifu_mem_ctl.scala 773:96]
  wire [31:0] _T_9843 = _T_9836 | 32'h3fffffff; // @[ifu_mem_ctl.scala 774:65]
  wire  _T_9845 = _T_9843 == 32'hffffffff; // @[ifu_mem_ctl.scala 774:96]
  wire  _T_9847 = _T_9839 | _T_9845; // @[ifu_mem_ctl.scala 773:162]
  wire [31:0] _T_9849 = _T_9836 | 32'h1fffffff; // @[ifu_mem_ctl.scala 775:65]
  wire  _T_9851 = _T_9849 == 32'hbfffffff; // @[ifu_mem_ctl.scala 775:96]
  wire  _T_9853 = _T_9847 | _T_9851; // @[ifu_mem_ctl.scala 774:162]
  wire [31:0] _T_9855 = _T_9836 | 32'hfffffff; // @[ifu_mem_ctl.scala 776:65]
  wire  _T_9857 = _T_9855 == 32'h8fffffff; // @[ifu_mem_ctl.scala 776:96]
  wire  ifc_region_acc_okay = _T_9853 | _T_9857; // @[ifu_mem_ctl.scala 775:162]
  wire  _T_9884 = ~ifc_region_acc_okay; // @[ifu_mem_ctl.scala 781:65]
  wire  _T_9885 = _T_3939 & _T_9884; // @[ifu_mem_ctl.scala 781:63]
  wire  ifc_region_acc_fault_memory_bf = _T_9885 & io_ifc_fetch_req_bf; // @[ifu_mem_ctl.scala 781:86]
  rvclkhdr rvclkhdr ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_io_l1clk),
    .io_clk(rvclkhdr_io_clk),
    .io_en(rvclkhdr_io_en),
    .io_scan_mode(rvclkhdr_io_scan_mode)
  );
  rvclkhdr rvclkhdr_1 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_1_io_l1clk),
    .io_clk(rvclkhdr_1_io_clk),
    .io_en(rvclkhdr_1_io_en),
    .io_scan_mode(rvclkhdr_1_io_scan_mode)
  );
  rvclkhdr rvclkhdr_2 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_2_io_l1clk),
    .io_clk(rvclkhdr_2_io_clk),
    .io_en(rvclkhdr_2_io_en),
    .io_scan_mode(rvclkhdr_2_io_scan_mode)
  );
  rvclkhdr rvclkhdr_3 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_3_io_l1clk),
    .io_clk(rvclkhdr_3_io_clk),
    .io_en(rvclkhdr_3_io_en),
    .io_scan_mode(rvclkhdr_3_io_scan_mode)
  );
  rvclkhdr rvclkhdr_4 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_4_io_l1clk),
    .io_clk(rvclkhdr_4_io_clk),
    .io_en(rvclkhdr_4_io_en),
    .io_scan_mode(rvclkhdr_4_io_scan_mode)
  );
  rvclkhdr rvclkhdr_5 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_5_io_l1clk),
    .io_clk(rvclkhdr_5_io_clk),
    .io_en(rvclkhdr_5_io_en),
    .io_scan_mode(rvclkhdr_5_io_scan_mode)
  );
  rvclkhdr rvclkhdr_6 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_6_io_l1clk),
    .io_clk(rvclkhdr_6_io_clk),
    .io_en(rvclkhdr_6_io_en),
    .io_scan_mode(rvclkhdr_6_io_scan_mode)
  );
  rvclkhdr rvclkhdr_7 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_7_io_l1clk),
    .io_clk(rvclkhdr_7_io_clk),
    .io_en(rvclkhdr_7_io_en),
    .io_scan_mode(rvclkhdr_7_io_scan_mode)
  );
  rvclkhdr rvclkhdr_8 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_8_io_l1clk),
    .io_clk(rvclkhdr_8_io_clk),
    .io_en(rvclkhdr_8_io_en),
    .io_scan_mode(rvclkhdr_8_io_scan_mode)
  );
  rvclkhdr rvclkhdr_9 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_9_io_l1clk),
    .io_clk(rvclkhdr_9_io_clk),
    .io_en(rvclkhdr_9_io_en),
    .io_scan_mode(rvclkhdr_9_io_scan_mode)
  );
  rvclkhdr rvclkhdr_10 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_10_io_l1clk),
    .io_clk(rvclkhdr_10_io_clk),
    .io_en(rvclkhdr_10_io_en),
    .io_scan_mode(rvclkhdr_10_io_scan_mode)
  );
  rvclkhdr rvclkhdr_11 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_11_io_l1clk),
    .io_clk(rvclkhdr_11_io_clk),
    .io_en(rvclkhdr_11_io_en),
    .io_scan_mode(rvclkhdr_11_io_scan_mode)
  );
  rvclkhdr rvclkhdr_12 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_12_io_l1clk),
    .io_clk(rvclkhdr_12_io_clk),
    .io_en(rvclkhdr_12_io_en),
    .io_scan_mode(rvclkhdr_12_io_scan_mode)
  );
  rvclkhdr rvclkhdr_13 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_13_io_l1clk),
    .io_clk(rvclkhdr_13_io_clk),
    .io_en(rvclkhdr_13_io_en),
    .io_scan_mode(rvclkhdr_13_io_scan_mode)
  );
  rvclkhdr rvclkhdr_14 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_14_io_l1clk),
    .io_clk(rvclkhdr_14_io_clk),
    .io_en(rvclkhdr_14_io_en),
    .io_scan_mode(rvclkhdr_14_io_scan_mode)
  );
  rvclkhdr rvclkhdr_15 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_15_io_l1clk),
    .io_clk(rvclkhdr_15_io_clk),
    .io_en(rvclkhdr_15_io_en),
    .io_scan_mode(rvclkhdr_15_io_scan_mode)
  );
  rvclkhdr rvclkhdr_16 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_16_io_l1clk),
    .io_clk(rvclkhdr_16_io_clk),
    .io_en(rvclkhdr_16_io_en),
    .io_scan_mode(rvclkhdr_16_io_scan_mode)
  );
  rvclkhdr rvclkhdr_17 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_17_io_l1clk),
    .io_clk(rvclkhdr_17_io_clk),
    .io_en(rvclkhdr_17_io_en),
    .io_scan_mode(rvclkhdr_17_io_scan_mode)
  );
  rvclkhdr rvclkhdr_18 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_18_io_l1clk),
    .io_clk(rvclkhdr_18_io_clk),
    .io_en(rvclkhdr_18_io_en),
    .io_scan_mode(rvclkhdr_18_io_scan_mode)
  );
  rvclkhdr rvclkhdr_19 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_19_io_l1clk),
    .io_clk(rvclkhdr_19_io_clk),
    .io_en(rvclkhdr_19_io_en),
    .io_scan_mode(rvclkhdr_19_io_scan_mode)
  );
  rvclkhdr rvclkhdr_20 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_20_io_l1clk),
    .io_clk(rvclkhdr_20_io_clk),
    .io_en(rvclkhdr_20_io_en),
    .io_scan_mode(rvclkhdr_20_io_scan_mode)
  );
  rvclkhdr rvclkhdr_21 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_21_io_l1clk),
    .io_clk(rvclkhdr_21_io_clk),
    .io_en(rvclkhdr_21_io_en),
    .io_scan_mode(rvclkhdr_21_io_scan_mode)
  );
  rvclkhdr rvclkhdr_22 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_22_io_l1clk),
    .io_clk(rvclkhdr_22_io_clk),
    .io_en(rvclkhdr_22_io_en),
    .io_scan_mode(rvclkhdr_22_io_scan_mode)
  );
  rvclkhdr rvclkhdr_23 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_23_io_l1clk),
    .io_clk(rvclkhdr_23_io_clk),
    .io_en(rvclkhdr_23_io_en),
    .io_scan_mode(rvclkhdr_23_io_scan_mode)
  );
  rvclkhdr rvclkhdr_24 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_24_io_l1clk),
    .io_clk(rvclkhdr_24_io_clk),
    .io_en(rvclkhdr_24_io_en),
    .io_scan_mode(rvclkhdr_24_io_scan_mode)
  );
  rvclkhdr rvclkhdr_25 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_25_io_l1clk),
    .io_clk(rvclkhdr_25_io_clk),
    .io_en(rvclkhdr_25_io_en),
    .io_scan_mode(rvclkhdr_25_io_scan_mode)
  );
  rvclkhdr rvclkhdr_26 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_26_io_l1clk),
    .io_clk(rvclkhdr_26_io_clk),
    .io_en(rvclkhdr_26_io_en),
    .io_scan_mode(rvclkhdr_26_io_scan_mode)
  );
  rvclkhdr rvclkhdr_27 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_27_io_l1clk),
    .io_clk(rvclkhdr_27_io_clk),
    .io_en(rvclkhdr_27_io_en),
    .io_scan_mode(rvclkhdr_27_io_scan_mode)
  );
  rvclkhdr rvclkhdr_28 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_28_io_l1clk),
    .io_clk(rvclkhdr_28_io_clk),
    .io_en(rvclkhdr_28_io_en),
    .io_scan_mode(rvclkhdr_28_io_scan_mode)
  );
  rvclkhdr rvclkhdr_29 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_29_io_l1clk),
    .io_clk(rvclkhdr_29_io_clk),
    .io_en(rvclkhdr_29_io_en),
    .io_scan_mode(rvclkhdr_29_io_scan_mode)
  );
  rvclkhdr rvclkhdr_30 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_30_io_l1clk),
    .io_clk(rvclkhdr_30_io_clk),
    .io_en(rvclkhdr_30_io_en),
    .io_scan_mode(rvclkhdr_30_io_scan_mode)
  );
  rvclkhdr rvclkhdr_31 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_31_io_l1clk),
    .io_clk(rvclkhdr_31_io_clk),
    .io_en(rvclkhdr_31_io_en),
    .io_scan_mode(rvclkhdr_31_io_scan_mode)
  );
  rvclkhdr rvclkhdr_32 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_32_io_l1clk),
    .io_clk(rvclkhdr_32_io_clk),
    .io_en(rvclkhdr_32_io_en),
    .io_scan_mode(rvclkhdr_32_io_scan_mode)
  );
  rvclkhdr rvclkhdr_33 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_33_io_l1clk),
    .io_clk(rvclkhdr_33_io_clk),
    .io_en(rvclkhdr_33_io_en),
    .io_scan_mode(rvclkhdr_33_io_scan_mode)
  );
  rvclkhdr rvclkhdr_34 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_34_io_l1clk),
    .io_clk(rvclkhdr_34_io_clk),
    .io_en(rvclkhdr_34_io_en),
    .io_scan_mode(rvclkhdr_34_io_scan_mode)
  );
  rvclkhdr rvclkhdr_35 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_35_io_l1clk),
    .io_clk(rvclkhdr_35_io_clk),
    .io_en(rvclkhdr_35_io_en),
    .io_scan_mode(rvclkhdr_35_io_scan_mode)
  );
  rvclkhdr rvclkhdr_36 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_36_io_l1clk),
    .io_clk(rvclkhdr_36_io_clk),
    .io_en(rvclkhdr_36_io_en),
    .io_scan_mode(rvclkhdr_36_io_scan_mode)
  );
  rvclkhdr rvclkhdr_37 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_37_io_l1clk),
    .io_clk(rvclkhdr_37_io_clk),
    .io_en(rvclkhdr_37_io_en),
    .io_scan_mode(rvclkhdr_37_io_scan_mode)
  );
  rvclkhdr rvclkhdr_38 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_38_io_l1clk),
    .io_clk(rvclkhdr_38_io_clk),
    .io_en(rvclkhdr_38_io_en),
    .io_scan_mode(rvclkhdr_38_io_scan_mode)
  );
  rvclkhdr rvclkhdr_39 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_39_io_l1clk),
    .io_clk(rvclkhdr_39_io_clk),
    .io_en(rvclkhdr_39_io_en),
    .io_scan_mode(rvclkhdr_39_io_scan_mode)
  );
  rvclkhdr rvclkhdr_40 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_40_io_l1clk),
    .io_clk(rvclkhdr_40_io_clk),
    .io_en(rvclkhdr_40_io_en),
    .io_scan_mode(rvclkhdr_40_io_scan_mode)
  );
  rvclkhdr rvclkhdr_41 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_41_io_l1clk),
    .io_clk(rvclkhdr_41_io_clk),
    .io_en(rvclkhdr_41_io_en),
    .io_scan_mode(rvclkhdr_41_io_scan_mode)
  );
  rvclkhdr rvclkhdr_42 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_42_io_l1clk),
    .io_clk(rvclkhdr_42_io_clk),
    .io_en(rvclkhdr_42_io_en),
    .io_scan_mode(rvclkhdr_42_io_scan_mode)
  );
  rvclkhdr rvclkhdr_43 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_43_io_l1clk),
    .io_clk(rvclkhdr_43_io_clk),
    .io_en(rvclkhdr_43_io_en),
    .io_scan_mode(rvclkhdr_43_io_scan_mode)
  );
  rvclkhdr rvclkhdr_44 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_44_io_l1clk),
    .io_clk(rvclkhdr_44_io_clk),
    .io_en(rvclkhdr_44_io_en),
    .io_scan_mode(rvclkhdr_44_io_scan_mode)
  );
  rvclkhdr rvclkhdr_45 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_45_io_l1clk),
    .io_clk(rvclkhdr_45_io_clk),
    .io_en(rvclkhdr_45_io_en),
    .io_scan_mode(rvclkhdr_45_io_scan_mode)
  );
  rvclkhdr rvclkhdr_46 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_46_io_l1clk),
    .io_clk(rvclkhdr_46_io_clk),
    .io_en(rvclkhdr_46_io_en),
    .io_scan_mode(rvclkhdr_46_io_scan_mode)
  );
  rvclkhdr rvclkhdr_47 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_47_io_l1clk),
    .io_clk(rvclkhdr_47_io_clk),
    .io_en(rvclkhdr_47_io_en),
    .io_scan_mode(rvclkhdr_47_io_scan_mode)
  );
  rvclkhdr rvclkhdr_48 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_48_io_l1clk),
    .io_clk(rvclkhdr_48_io_clk),
    .io_en(rvclkhdr_48_io_en),
    .io_scan_mode(rvclkhdr_48_io_scan_mode)
  );
  rvclkhdr rvclkhdr_49 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_49_io_l1clk),
    .io_clk(rvclkhdr_49_io_clk),
    .io_en(rvclkhdr_49_io_en),
    .io_scan_mode(rvclkhdr_49_io_scan_mode)
  );
  rvclkhdr rvclkhdr_50 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_50_io_l1clk),
    .io_clk(rvclkhdr_50_io_clk),
    .io_en(rvclkhdr_50_io_en),
    .io_scan_mode(rvclkhdr_50_io_scan_mode)
  );
  rvclkhdr rvclkhdr_51 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_51_io_l1clk),
    .io_clk(rvclkhdr_51_io_clk),
    .io_en(rvclkhdr_51_io_en),
    .io_scan_mode(rvclkhdr_51_io_scan_mode)
  );
  rvclkhdr rvclkhdr_52 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_52_io_l1clk),
    .io_clk(rvclkhdr_52_io_clk),
    .io_en(rvclkhdr_52_io_en),
    .io_scan_mode(rvclkhdr_52_io_scan_mode)
  );
  rvclkhdr rvclkhdr_53 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_53_io_l1clk),
    .io_clk(rvclkhdr_53_io_clk),
    .io_en(rvclkhdr_53_io_en),
    .io_scan_mode(rvclkhdr_53_io_scan_mode)
  );
  rvclkhdr rvclkhdr_54 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_54_io_l1clk),
    .io_clk(rvclkhdr_54_io_clk),
    .io_en(rvclkhdr_54_io_en),
    .io_scan_mode(rvclkhdr_54_io_scan_mode)
  );
  rvclkhdr rvclkhdr_55 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_55_io_l1clk),
    .io_clk(rvclkhdr_55_io_clk),
    .io_en(rvclkhdr_55_io_en),
    .io_scan_mode(rvclkhdr_55_io_scan_mode)
  );
  rvclkhdr rvclkhdr_56 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_56_io_l1clk),
    .io_clk(rvclkhdr_56_io_clk),
    .io_en(rvclkhdr_56_io_en),
    .io_scan_mode(rvclkhdr_56_io_scan_mode)
  );
  rvclkhdr rvclkhdr_57 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_57_io_l1clk),
    .io_clk(rvclkhdr_57_io_clk),
    .io_en(rvclkhdr_57_io_en),
    .io_scan_mode(rvclkhdr_57_io_scan_mode)
  );
  rvclkhdr rvclkhdr_58 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_58_io_l1clk),
    .io_clk(rvclkhdr_58_io_clk),
    .io_en(rvclkhdr_58_io_en),
    .io_scan_mode(rvclkhdr_58_io_scan_mode)
  );
  rvclkhdr rvclkhdr_59 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_59_io_l1clk),
    .io_clk(rvclkhdr_59_io_clk),
    .io_en(rvclkhdr_59_io_en),
    .io_scan_mode(rvclkhdr_59_io_scan_mode)
  );
  rvclkhdr rvclkhdr_60 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_60_io_l1clk),
    .io_clk(rvclkhdr_60_io_clk),
    .io_en(rvclkhdr_60_io_en),
    .io_scan_mode(rvclkhdr_60_io_scan_mode)
  );
  rvclkhdr rvclkhdr_61 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_61_io_l1clk),
    .io_clk(rvclkhdr_61_io_clk),
    .io_en(rvclkhdr_61_io_en),
    .io_scan_mode(rvclkhdr_61_io_scan_mode)
  );
  rvclkhdr rvclkhdr_62 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_62_io_l1clk),
    .io_clk(rvclkhdr_62_io_clk),
    .io_en(rvclkhdr_62_io_en),
    .io_scan_mode(rvclkhdr_62_io_scan_mode)
  );
  rvclkhdr rvclkhdr_63 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_63_io_l1clk),
    .io_clk(rvclkhdr_63_io_clk),
    .io_en(rvclkhdr_63_io_en),
    .io_scan_mode(rvclkhdr_63_io_scan_mode)
  );
  rvclkhdr rvclkhdr_64 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_64_io_l1clk),
    .io_clk(rvclkhdr_64_io_clk),
    .io_en(rvclkhdr_64_io_en),
    .io_scan_mode(rvclkhdr_64_io_scan_mode)
  );
  rvclkhdr rvclkhdr_65 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_65_io_l1clk),
    .io_clk(rvclkhdr_65_io_clk),
    .io_en(rvclkhdr_65_io_en),
    .io_scan_mode(rvclkhdr_65_io_scan_mode)
  );
  rvclkhdr rvclkhdr_66 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_66_io_l1clk),
    .io_clk(rvclkhdr_66_io_clk),
    .io_en(rvclkhdr_66_io_en),
    .io_scan_mode(rvclkhdr_66_io_scan_mode)
  );
  rvclkhdr rvclkhdr_67 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_67_io_l1clk),
    .io_clk(rvclkhdr_67_io_clk),
    .io_en(rvclkhdr_67_io_en),
    .io_scan_mode(rvclkhdr_67_io_scan_mode)
  );
  rvclkhdr rvclkhdr_68 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_68_io_l1clk),
    .io_clk(rvclkhdr_68_io_clk),
    .io_en(rvclkhdr_68_io_en),
    .io_scan_mode(rvclkhdr_68_io_scan_mode)
  );
  rvclkhdr rvclkhdr_69 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_69_io_l1clk),
    .io_clk(rvclkhdr_69_io_clk),
    .io_en(rvclkhdr_69_io_en),
    .io_scan_mode(rvclkhdr_69_io_scan_mode)
  );
  rvclkhdr rvclkhdr_70 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_70_io_l1clk),
    .io_clk(rvclkhdr_70_io_clk),
    .io_en(rvclkhdr_70_io_en),
    .io_scan_mode(rvclkhdr_70_io_scan_mode)
  );
  rvclkhdr rvclkhdr_71 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_71_io_l1clk),
    .io_clk(rvclkhdr_71_io_clk),
    .io_en(rvclkhdr_71_io_en),
    .io_scan_mode(rvclkhdr_71_io_scan_mode)
  );
  rvclkhdr rvclkhdr_72 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_72_io_l1clk),
    .io_clk(rvclkhdr_72_io_clk),
    .io_en(rvclkhdr_72_io_en),
    .io_scan_mode(rvclkhdr_72_io_scan_mode)
  );
  rvclkhdr rvclkhdr_73 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_73_io_l1clk),
    .io_clk(rvclkhdr_73_io_clk),
    .io_en(rvclkhdr_73_io_en),
    .io_scan_mode(rvclkhdr_73_io_scan_mode)
  );
  rvclkhdr rvclkhdr_74 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_74_io_l1clk),
    .io_clk(rvclkhdr_74_io_clk),
    .io_en(rvclkhdr_74_io_en),
    .io_scan_mode(rvclkhdr_74_io_scan_mode)
  );
  rvclkhdr rvclkhdr_75 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_75_io_l1clk),
    .io_clk(rvclkhdr_75_io_clk),
    .io_en(rvclkhdr_75_io_en),
    .io_scan_mode(rvclkhdr_75_io_scan_mode)
  );
  rvclkhdr rvclkhdr_76 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_76_io_l1clk),
    .io_clk(rvclkhdr_76_io_clk),
    .io_en(rvclkhdr_76_io_en),
    .io_scan_mode(rvclkhdr_76_io_scan_mode)
  );
  rvclkhdr rvclkhdr_77 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_77_io_l1clk),
    .io_clk(rvclkhdr_77_io_clk),
    .io_en(rvclkhdr_77_io_en),
    .io_scan_mode(rvclkhdr_77_io_scan_mode)
  );
  rvclkhdr rvclkhdr_78 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_78_io_l1clk),
    .io_clk(rvclkhdr_78_io_clk),
    .io_en(rvclkhdr_78_io_en),
    .io_scan_mode(rvclkhdr_78_io_scan_mode)
  );
  rvclkhdr rvclkhdr_79 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_79_io_l1clk),
    .io_clk(rvclkhdr_79_io_clk),
    .io_en(rvclkhdr_79_io_en),
    .io_scan_mode(rvclkhdr_79_io_scan_mode)
  );
  rvclkhdr rvclkhdr_80 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_80_io_l1clk),
    .io_clk(rvclkhdr_80_io_clk),
    .io_en(rvclkhdr_80_io_en),
    .io_scan_mode(rvclkhdr_80_io_scan_mode)
  );
  rvclkhdr rvclkhdr_81 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_81_io_l1clk),
    .io_clk(rvclkhdr_81_io_clk),
    .io_en(rvclkhdr_81_io_en),
    .io_scan_mode(rvclkhdr_81_io_scan_mode)
  );
  rvclkhdr rvclkhdr_82 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_82_io_l1clk),
    .io_clk(rvclkhdr_82_io_clk),
    .io_en(rvclkhdr_82_io_en),
    .io_scan_mode(rvclkhdr_82_io_scan_mode)
  );
  rvclkhdr rvclkhdr_83 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_83_io_l1clk),
    .io_clk(rvclkhdr_83_io_clk),
    .io_en(rvclkhdr_83_io_en),
    .io_scan_mode(rvclkhdr_83_io_scan_mode)
  );
  rvclkhdr rvclkhdr_84 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_84_io_l1clk),
    .io_clk(rvclkhdr_84_io_clk),
    .io_en(rvclkhdr_84_io_en),
    .io_scan_mode(rvclkhdr_84_io_scan_mode)
  );
  rvclkhdr rvclkhdr_85 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_85_io_l1clk),
    .io_clk(rvclkhdr_85_io_clk),
    .io_en(rvclkhdr_85_io_en),
    .io_scan_mode(rvclkhdr_85_io_scan_mode)
  );
  rvclkhdr rvclkhdr_86 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_86_io_l1clk),
    .io_clk(rvclkhdr_86_io_clk),
    .io_en(rvclkhdr_86_io_en),
    .io_scan_mode(rvclkhdr_86_io_scan_mode)
  );
  rvclkhdr rvclkhdr_87 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_87_io_l1clk),
    .io_clk(rvclkhdr_87_io_clk),
    .io_en(rvclkhdr_87_io_en),
    .io_scan_mode(rvclkhdr_87_io_scan_mode)
  );
  rvclkhdr rvclkhdr_88 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_88_io_l1clk),
    .io_clk(rvclkhdr_88_io_clk),
    .io_en(rvclkhdr_88_io_en),
    .io_scan_mode(rvclkhdr_88_io_scan_mode)
  );
  rvclkhdr rvclkhdr_89 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_89_io_l1clk),
    .io_clk(rvclkhdr_89_io_clk),
    .io_en(rvclkhdr_89_io_en),
    .io_scan_mode(rvclkhdr_89_io_scan_mode)
  );
  rvclkhdr rvclkhdr_90 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_90_io_l1clk),
    .io_clk(rvclkhdr_90_io_clk),
    .io_en(rvclkhdr_90_io_en),
    .io_scan_mode(rvclkhdr_90_io_scan_mode)
  );
  rvclkhdr rvclkhdr_91 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_91_io_l1clk),
    .io_clk(rvclkhdr_91_io_clk),
    .io_en(rvclkhdr_91_io_en),
    .io_scan_mode(rvclkhdr_91_io_scan_mode)
  );
  rvclkhdr rvclkhdr_92 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_92_io_l1clk),
    .io_clk(rvclkhdr_92_io_clk),
    .io_en(rvclkhdr_92_io_en),
    .io_scan_mode(rvclkhdr_92_io_scan_mode)
  );
  rvclkhdr rvclkhdr_93 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_93_io_l1clk),
    .io_clk(rvclkhdr_93_io_clk),
    .io_en(rvclkhdr_93_io_en),
    .io_scan_mode(rvclkhdr_93_io_scan_mode)
  );
  assign io_dec_mem_ctrl_ifu_pmu_ic_miss = _T_9799; // @[ifu_mem_ctl.scala 752:35]
  assign io_dec_mem_ctrl_ifu_pmu_ic_hit = _T_9800; // @[ifu_mem_ctl.scala 753:34]
  assign io_dec_mem_ctrl_ifu_pmu_bus_error = _T_9801; // @[ifu_mem_ctl.scala 754:37]
  assign io_dec_mem_ctrl_ifu_pmu_bus_busy = _T_9805; // @[ifu_mem_ctl.scala 755:36]
  assign io_dec_mem_ctrl_ifu_ic_error_start = _T_1200 | ic_rd_parity_final_err; // @[ifu_mem_ctl.scala 256:38]
  assign io_dec_mem_ctrl_ifu_iccm_rd_ecc_single_err = _T_3911 & ifc_fetch_req_f; // @[ifu_mem_ctl.scala 612:46]
  assign io_dec_mem_ctrl_ifu_ic_debug_rd_data = _T_1212; // @[ifu_mem_ctl.scala 263:40]
  assign io_dec_mem_ctrl_ifu_ic_debug_rd_data_valid = _T_9826; // @[ifu_mem_ctl.scala 770:46]
  assign io_dec_mem_ctrl_ifu_miss_state_idle = miss_state == 3'h0; // @[ifu_mem_ctl.scala 235:39]
  assign io_ifu_axi_ar_valid = ifu_bus_cmd_valid; // @[ifu_mem_ctl.scala 497:23]
  assign io_ifu_axi_ar_bits_addr = _T_2610 & _T_2612; // @[ifu_mem_ctl.scala 499:27]
  assign io_iccm_rw_addr = _T_3110 ? io_dma_mem_ctl_dma_mem_addr[15:1] : _T_3117; // @[ifu_mem_ctl.scala 599:19]
  assign io_iccm_buf_correct_ecc = iccm_correct_ecc & _T_2497; // @[ifu_mem_ctl.scala 395:27]
  assign io_iccm_correction_state = _T_2526 ? 1'h0 : _GEN_42; // @[ifu_mem_ctl.scala 430:28 ifu_mem_ctl.scala 442:32 ifu_mem_ctl.scala 449:32 ifu_mem_ctl.scala 456:32]
  assign io_iccm_wren = _T_2710 | iccm_correct_ecc; // @[ifu_mem_ctl.scala 569:16]
  assign io_iccm_rden = _T_2714 | _T_2715; // @[ifu_mem_ctl.scala 570:16]
  assign io_iccm_wr_size = _T_2720 & io_dma_mem_ctl_dma_mem_sz; // @[ifu_mem_ctl.scala 572:19]
  assign io_iccm_wr_data = _T_3092 ? _T_3093 : _T_3100; // @[ifu_mem_ctl.scala 576:19]
  assign io_ic_rw_addr = _T_340 | _T_341; // @[ifu_mem_ctl.scala 244:17]
  assign io_ic_tag_valid = ic_tag_valid_unq & _T_9792; // @[ifu_mem_ctl.scala 747:19]
  assign io_ic_rd_en = _T_3966 | _T_3971; // @[ifu_mem_ctl.scala 626:15]
  assign io_ic_debug_wr_data = io_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_wrdata; // @[ifu_mem_ctl.scala 254:23]
  assign io_ic_debug_addr = io_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_dicawics[9:0]; // @[ifu_mem_ctl.scala 759:20]
  assign io_ic_debug_rd_en = io_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_rd_valid; // @[ifu_mem_ctl.scala 761:21]
  assign io_ic_debug_wr_en = io_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_wr_valid; // @[ifu_mem_ctl.scala 762:21]
  assign io_ic_debug_tag_array = io_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_dicawics[16]; // @[ifu_mem_ctl.scala 760:25]
  assign io_ic_debug_way = _T_9818[1:0]; // @[ifu_mem_ctl.scala 763:19]
  assign io_ic_premux_data = ic_premux_data_temp[63:0]; // @[ifu_mem_ctl.scala 295:21]
  assign io_ic_sel_premux_data = fetch_req_iccm_f | sel_byp_data; // @[ifu_mem_ctl.scala 296:25]
  assign io_ifu_ic_mb_empty = _T_325 | _T_231; // @[ifu_mem_ctl.scala 234:22]
  assign io_ic_dma_active = _T_11 | io_dec_mem_ctrl_dec_tlu_flush_err_wb; // @[ifu_mem_ctl.scala 97:20]
  assign io_iccm_dma_ecc_error = iccm_dma_ecc_error; // @[ifu_mem_ctl.scala 595:25]
  assign io_iccm_dma_rvalid = iccm_dma_rvalid_temp; // @[ifu_mem_ctl.scala 593:22]
  assign io_iccm_dma_rdata = iccm_dma_rdata_temp; // @[ifu_mem_ctl.scala 597:21]
  assign io_iccm_dma_rtag = iccm_dma_rtag_temp; // @[ifu_mem_ctl.scala 588:20]
  assign io_iccm_ready = _T_2706 & _T_2700; // @[ifu_mem_ctl.scala 567:17]
  assign io_iccm_rd_ecc_double_err = iccm_dma_ecc_error_in & ifc_iccm_access_f; // @[ifu_mem_ctl.scala 613:29]
  assign io_iccm_dma_sb_error = _T_3 & dma_iccm_req_f; // @[ifu_mem_ctl.scala 95:24]
  assign io_ic_hit_f = _T_263 | _T_264; // @[ifu_mem_ctl.scala 195:15]
  assign io_ic_access_fault_f = _T_2492 & _T_319; // @[ifu_mem_ctl.scala 301:24]
  assign io_ic_access_fault_type_f = io_iccm_rd_ecc_double_err ? 2'h1 : _T_1278; // @[ifu_mem_ctl.scala 302:29]
  assign io_ifu_async_error_start = io_dec_mem_ctrl_ifu_iccm_rd_ecc_single_err | io_dec_mem_ctrl_ifu_ic_error_start; // @[ifu_mem_ctl.scala 96:28]
  assign io_ic_fetch_val_f = {_T_1286,fetch_req_f_qual}; // @[ifu_mem_ctl.scala 305:21]
  assign io_ic_data_f = ic_final_data[31:0]; // @[ifu_mem_ctl.scala 298:16]
  assign rvclkhdr_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_io_en = ic_debug_rd_en_ff; // @[lib.scala 345:16]
  assign rvclkhdr_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_1_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_1_io_en = io_ic_debug_rd_en | io_ic_debug_wr_en; // @[lib.scala 345:16]
  assign rvclkhdr_1_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_2_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_2_io_en = _T_1 | io_exu_flush_final; // @[lib.scala 345:16]
  assign rvclkhdr_2_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_3_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_3_io_en = _T_309 | io_dec_mem_ctrl_dec_tlu_force_halt; // @[lib.scala 345:16]
  assign rvclkhdr_3_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_4_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_4_io_en = 1'h0; // @[lib.scala 345:16]
  assign rvclkhdr_4_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_5_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_5_io_en = 1'h0; // @[lib.scala 345:16]
  assign rvclkhdr_5_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_6_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_6_io_en = 1'h0; // @[lib.scala 345:16]
  assign rvclkhdr_6_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_7_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_7_io_en = 1'h0; // @[lib.scala 345:16]
  assign rvclkhdr_7_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_8_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_8_io_en = 1'h0; // @[lib.scala 345:16]
  assign rvclkhdr_8_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_9_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_9_io_en = 1'h0; // @[lib.scala 345:16]
  assign rvclkhdr_9_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_10_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_10_io_en = 1'h0; // @[lib.scala 345:16]
  assign rvclkhdr_10_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_11_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_11_io_en = 1'h0; // @[lib.scala 345:16]
  assign rvclkhdr_11_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_12_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_12_io_en = 1'h0; // @[lib.scala 345:16]
  assign rvclkhdr_12_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_13_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_13_io_en = 1'h0; // @[lib.scala 345:16]
  assign rvclkhdr_13_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_14_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_14_io_en = 1'h0; // @[lib.scala 345:16]
  assign rvclkhdr_14_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_15_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_15_io_en = 1'h0; // @[lib.scala 345:16]
  assign rvclkhdr_15_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_16_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_16_io_en = 1'h0; // @[lib.scala 345:16]
  assign rvclkhdr_16_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_17_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_17_io_en = 1'h0; // @[lib.scala 345:16]
  assign rvclkhdr_17_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_18_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_18_io_en = 1'h0; // @[lib.scala 345:16]
  assign rvclkhdr_18_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_19_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_19_io_en = 1'h0; // @[lib.scala 345:16]
  assign rvclkhdr_19_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_20_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_20_io_en = 1'h0; // @[lib.scala 345:16]
  assign rvclkhdr_20_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_21_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_21_io_en = 1'h0; // @[lib.scala 345:16]
  assign rvclkhdr_21_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_22_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_22_io_en = 1'h0; // @[lib.scala 345:16]
  assign rvclkhdr_22_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_23_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_23_io_en = 1'h0; // @[lib.scala 345:16]
  assign rvclkhdr_23_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_24_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_24_io_en = 1'h0; // @[lib.scala 345:16]
  assign rvclkhdr_24_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_25_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_25_io_en = 1'h0; // @[lib.scala 345:16]
  assign rvclkhdr_25_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_26_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_26_io_en = 1'h0; // @[lib.scala 345:16]
  assign rvclkhdr_26_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_27_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_27_io_en = 1'h0; // @[lib.scala 345:16]
  assign rvclkhdr_27_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_28_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_28_io_en = 1'h0; // @[lib.scala 345:16]
  assign rvclkhdr_28_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_29_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_29_io_en = 1'h0; // @[lib.scala 345:16]
  assign rvclkhdr_29_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_30_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_30_io_en = 1'h0; // @[lib.scala 345:16]
  assign rvclkhdr_30_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_31_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_31_io_en = 1'h0; // @[lib.scala 345:16]
  assign rvclkhdr_31_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_32_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_32_io_en = 1'h0; // @[lib.scala 345:16]
  assign rvclkhdr_32_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_33_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_33_io_en = 1'h0; // @[lib.scala 345:16]
  assign rvclkhdr_33_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_34_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_34_io_en = 1'h0; // @[lib.scala 345:16]
  assign rvclkhdr_34_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_35_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_35_io_en = 1'h0; // @[lib.scala 345:16]
  assign rvclkhdr_35_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_36_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_36_io_en = 1'h0; // @[lib.scala 345:16]
  assign rvclkhdr_36_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_37_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_37_io_en = 1'h0; // @[lib.scala 345:16]
  assign rvclkhdr_37_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_38_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_38_io_en = 1'h0; // @[lib.scala 345:16]
  assign rvclkhdr_38_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_39_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_39_io_en = 1'h0; // @[lib.scala 345:16]
  assign rvclkhdr_39_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_40_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_40_io_en = 1'h0; // @[lib.scala 345:16]
  assign rvclkhdr_40_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_41_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_41_io_en = 1'h0; // @[lib.scala 345:16]
  assign rvclkhdr_41_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_42_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_42_io_en = 1'h0; // @[lib.scala 345:16]
  assign rvclkhdr_42_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_43_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_43_io_en = 1'h0; // @[lib.scala 345:16]
  assign rvclkhdr_43_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_44_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_44_io_en = 1'h0; // @[lib.scala 345:16]
  assign rvclkhdr_44_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_45_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_45_io_en = 1'h0; // @[lib.scala 345:16]
  assign rvclkhdr_45_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_46_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_46_io_en = 1'h0; // @[lib.scala 345:16]
  assign rvclkhdr_46_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_47_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_47_io_en = 1'h0; // @[lib.scala 345:16]
  assign rvclkhdr_47_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_48_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_48_io_en = 1'h0; // @[lib.scala 345:16]
  assign rvclkhdr_48_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_49_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_49_io_en = 1'h0; // @[lib.scala 345:16]
  assign rvclkhdr_49_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_50_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_50_io_en = 1'h0; // @[lib.scala 345:16]
  assign rvclkhdr_50_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_51_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_51_io_en = 1'h0; // @[lib.scala 345:16]
  assign rvclkhdr_51_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_52_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_52_io_en = 1'h0; // @[lib.scala 345:16]
  assign rvclkhdr_52_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_53_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_53_io_en = 1'h0; // @[lib.scala 345:16]
  assign rvclkhdr_53_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_54_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_54_io_en = 1'h0; // @[lib.scala 345:16]
  assign rvclkhdr_54_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_55_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_55_io_en = 1'h0; // @[lib.scala 345:16]
  assign rvclkhdr_55_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_56_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_56_io_en = 1'h0; // @[lib.scala 345:16]
  assign rvclkhdr_56_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_57_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_57_io_en = 1'h0; // @[lib.scala 345:16]
  assign rvclkhdr_57_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_58_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_58_io_en = 1'h0; // @[lib.scala 345:16]
  assign rvclkhdr_58_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_59_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_59_io_en = 1'h0; // @[lib.scala 345:16]
  assign rvclkhdr_59_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_60_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_60_io_en = 1'h0; // @[lib.scala 345:16]
  assign rvclkhdr_60_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_61_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_61_io_en = 1'h0; // @[lib.scala 345:16]
  assign rvclkhdr_61_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_62_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_62_io_en = 1'h0; // @[lib.scala 345:16]
  assign rvclkhdr_62_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_63_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_63_io_en = 1'h0; // @[lib.scala 345:16]
  assign rvclkhdr_63_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_64_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_64_io_en = 1'h0; // @[lib.scala 345:16]
  assign rvclkhdr_64_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_65_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_65_io_en = 1'h0; // @[lib.scala 345:16]
  assign rvclkhdr_65_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_66_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_66_io_en = 1'h0; // @[lib.scala 345:16]
  assign rvclkhdr_66_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_67_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_67_io_en = 1'h0; // @[lib.scala 345:16]
  assign rvclkhdr_67_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_68_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_68_io_en = io_ifu_bus_clk_en; // @[lib.scala 345:16]
  assign rvclkhdr_68_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_69_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_69_io_en = io_ifu_bus_clk_en | io_dec_mem_ctrl_dec_tlu_force_halt; // @[lib.scala 345:16]
  assign rvclkhdr_69_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_70_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_70_io_en = ifu_status_wr_addr_ff[6:3] == 4'h0; // @[lib.scala 345:16]
  assign rvclkhdr_70_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_71_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_71_io_en = ifu_status_wr_addr_ff[6:3] == 4'h1; // @[lib.scala 345:16]
  assign rvclkhdr_71_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_72_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_72_io_en = ifu_status_wr_addr_ff[6:3] == 4'h2; // @[lib.scala 345:16]
  assign rvclkhdr_72_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_73_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_73_io_en = ifu_status_wr_addr_ff[6:3] == 4'h3; // @[lib.scala 345:16]
  assign rvclkhdr_73_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_74_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_74_io_en = ifu_status_wr_addr_ff[6:3] == 4'h4; // @[lib.scala 345:16]
  assign rvclkhdr_74_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_75_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_75_io_en = ifu_status_wr_addr_ff[6:3] == 4'h5; // @[lib.scala 345:16]
  assign rvclkhdr_75_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_76_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_76_io_en = ifu_status_wr_addr_ff[6:3] == 4'h6; // @[lib.scala 345:16]
  assign rvclkhdr_76_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_77_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_77_io_en = ifu_status_wr_addr_ff[6:3] == 4'h7; // @[lib.scala 345:16]
  assign rvclkhdr_77_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_78_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_78_io_en = ifu_status_wr_addr_ff[6:3] == 4'h8; // @[lib.scala 345:16]
  assign rvclkhdr_78_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_79_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_79_io_en = ifu_status_wr_addr_ff[6:3] == 4'h9; // @[lib.scala 345:16]
  assign rvclkhdr_79_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_80_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_80_io_en = ifu_status_wr_addr_ff[6:3] == 4'ha; // @[lib.scala 345:16]
  assign rvclkhdr_80_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_81_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_81_io_en = ifu_status_wr_addr_ff[6:3] == 4'hb; // @[lib.scala 345:16]
  assign rvclkhdr_81_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_82_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_82_io_en = ifu_status_wr_addr_ff[6:3] == 4'hc; // @[lib.scala 345:16]
  assign rvclkhdr_82_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_83_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_83_io_en = ifu_status_wr_addr_ff[6:3] == 4'hd; // @[lib.scala 345:16]
  assign rvclkhdr_83_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_84_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_84_io_en = ifu_status_wr_addr_ff[6:3] == 4'he; // @[lib.scala 345:16]
  assign rvclkhdr_84_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_85_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_85_io_en = ifu_status_wr_addr_ff[6:3] == 4'hf; // @[lib.scala 345:16]
  assign rvclkhdr_85_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_86_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_86_io_en = tag_valid_clken_0[0]; // @[lib.scala 345:16]
  assign rvclkhdr_86_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_87_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_87_io_en = tag_valid_clken_0[1]; // @[lib.scala 345:16]
  assign rvclkhdr_87_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_88_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_88_io_en = tag_valid_clken_1[0]; // @[lib.scala 345:16]
  assign rvclkhdr_88_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_89_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_89_io_en = tag_valid_clken_1[1]; // @[lib.scala 345:16]
  assign rvclkhdr_89_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_90_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_90_io_en = tag_valid_clken_2[0]; // @[lib.scala 345:16]
  assign rvclkhdr_90_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_91_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_91_io_en = tag_valid_clken_2[1]; // @[lib.scala 345:16]
  assign rvclkhdr_91_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_92_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_92_io_en = tag_valid_clken_3[0]; // @[lib.scala 345:16]
  assign rvclkhdr_92_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_93_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_93_io_en = tag_valid_clken_3[1]; // @[lib.scala 345:16]
  assign rvclkhdr_93_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  flush_final_f = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  ifc_fetch_req_f_raw = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  miss_state = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  ifu_fetch_addr_int_f = _RAND_3[30:0];
  _RAND_4 = {1{`RANDOM}};
  ifc_iccm_access_f = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  iccm_dma_rvalid_in = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  dma_iccm_req_f = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  perr_state = _RAND_7[2:0];
  _RAND_8 = {1{`RANDOM}};
  err_stop_state = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  reset_all_tags = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  ifc_region_acc_fault_final_f = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  uncacheable_miss_ff = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  ic_miss_buff_data_valid = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  imb_ff = _RAND_13[30:0];
  _RAND_14 = {1{`RANDOM}};
  sel_mb_addr_ff = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  ifu_ic_rw_int_addr_ff = _RAND_15[6:0];
  _RAND_16 = {1{`RANDOM}};
  way_status_out_0 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  way_status_out_1 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  way_status_out_2 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  way_status_out_3 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  way_status_out_4 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  way_status_out_5 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  way_status_out_6 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  way_status_out_7 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  way_status_out_8 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  way_status_out_9 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  way_status_out_10 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  way_status_out_11 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  way_status_out_12 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  way_status_out_13 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  way_status_out_14 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  way_status_out_15 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  way_status_out_16 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  way_status_out_17 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  way_status_out_18 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  way_status_out_19 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  way_status_out_20 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  way_status_out_21 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  way_status_out_22 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  way_status_out_23 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  way_status_out_24 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  way_status_out_25 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  way_status_out_26 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  way_status_out_27 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  way_status_out_28 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  way_status_out_29 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  way_status_out_30 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  way_status_out_31 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  way_status_out_32 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  way_status_out_33 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  way_status_out_34 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  way_status_out_35 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  way_status_out_36 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  way_status_out_37 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  way_status_out_38 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  way_status_out_39 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  way_status_out_40 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  way_status_out_41 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  way_status_out_42 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  way_status_out_43 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  way_status_out_44 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  way_status_out_45 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  way_status_out_46 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  way_status_out_47 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  way_status_out_48 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  way_status_out_49 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  way_status_out_50 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  way_status_out_51 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  way_status_out_52 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  way_status_out_53 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  way_status_out_54 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  way_status_out_55 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  way_status_out_56 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  way_status_out_57 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  way_status_out_58 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  way_status_out_59 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  way_status_out_60 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  way_status_out_61 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  way_status_out_62 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  way_status_out_63 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  way_status_out_64 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  way_status_out_65 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  way_status_out_66 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  way_status_out_67 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  way_status_out_68 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  way_status_out_69 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  way_status_out_70 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  way_status_out_71 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  way_status_out_72 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  way_status_out_73 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  way_status_out_74 = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  way_status_out_75 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  way_status_out_76 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  way_status_out_77 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  way_status_out_78 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  way_status_out_79 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  way_status_out_80 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  way_status_out_81 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  way_status_out_82 = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  way_status_out_83 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  way_status_out_84 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  way_status_out_85 = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  way_status_out_86 = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  way_status_out_87 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  way_status_out_88 = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  way_status_out_89 = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  way_status_out_90 = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  way_status_out_91 = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  way_status_out_92 = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  way_status_out_93 = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  way_status_out_94 = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  way_status_out_95 = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  way_status_out_96 = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  way_status_out_97 = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  way_status_out_98 = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  way_status_out_99 = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  way_status_out_100 = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  way_status_out_101 = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  way_status_out_102 = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  way_status_out_103 = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  way_status_out_104 = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  way_status_out_105 = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  way_status_out_106 = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  way_status_out_107 = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  way_status_out_108 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  way_status_out_109 = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  way_status_out_110 = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  way_status_out_111 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  way_status_out_112 = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  way_status_out_113 = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  way_status_out_114 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  way_status_out_115 = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  way_status_out_116 = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  way_status_out_117 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  way_status_out_118 = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  way_status_out_119 = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  way_status_out_120 = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  way_status_out_121 = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  way_status_out_122 = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  way_status_out_123 = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  way_status_out_124 = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  way_status_out_125 = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  way_status_out_126 = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  way_status_out_127 = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  way_status_mb_ff = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  tagv_mb_ff = _RAND_145[1:0];
  _RAND_146 = {1{`RANDOM}};
  reset_ic_ff = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  fetch_uncacheable_ff = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  miss_addr = _RAND_148[25:0];
  _RAND_149 = {1{`RANDOM}};
  ifc_region_acc_fault_f = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  bus_rd_addr_count = _RAND_150[2:0];
  _RAND_151 = {1{`RANDOM}};
  ic_act_miss_f_delayed = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  ic_crit_wd_rdy_new_ff = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  ic_miss_buff_data_error = _RAND_153[7:0];
  _RAND_154 = {1{`RANDOM}};
  ic_debug_ict_array_sel_ff = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  ic_tag_valid_out_1_0 = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  ic_tag_valid_out_1_1 = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  ic_tag_valid_out_1_2 = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  ic_tag_valid_out_1_3 = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  ic_tag_valid_out_1_4 = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  ic_tag_valid_out_1_5 = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  ic_tag_valid_out_1_6 = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  ic_tag_valid_out_1_7 = _RAND_162[0:0];
  _RAND_163 = {1{`RANDOM}};
  ic_tag_valid_out_1_8 = _RAND_163[0:0];
  _RAND_164 = {1{`RANDOM}};
  ic_tag_valid_out_1_9 = _RAND_164[0:0];
  _RAND_165 = {1{`RANDOM}};
  ic_tag_valid_out_1_10 = _RAND_165[0:0];
  _RAND_166 = {1{`RANDOM}};
  ic_tag_valid_out_1_11 = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  ic_tag_valid_out_1_12 = _RAND_167[0:0];
  _RAND_168 = {1{`RANDOM}};
  ic_tag_valid_out_1_13 = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  ic_tag_valid_out_1_14 = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  ic_tag_valid_out_1_15 = _RAND_170[0:0];
  _RAND_171 = {1{`RANDOM}};
  ic_tag_valid_out_1_16 = _RAND_171[0:0];
  _RAND_172 = {1{`RANDOM}};
  ic_tag_valid_out_1_17 = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  ic_tag_valid_out_1_18 = _RAND_173[0:0];
  _RAND_174 = {1{`RANDOM}};
  ic_tag_valid_out_1_19 = _RAND_174[0:0];
  _RAND_175 = {1{`RANDOM}};
  ic_tag_valid_out_1_20 = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  ic_tag_valid_out_1_21 = _RAND_176[0:0];
  _RAND_177 = {1{`RANDOM}};
  ic_tag_valid_out_1_22 = _RAND_177[0:0];
  _RAND_178 = {1{`RANDOM}};
  ic_tag_valid_out_1_23 = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  ic_tag_valid_out_1_24 = _RAND_179[0:0];
  _RAND_180 = {1{`RANDOM}};
  ic_tag_valid_out_1_25 = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  ic_tag_valid_out_1_26 = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  ic_tag_valid_out_1_27 = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  ic_tag_valid_out_1_28 = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  ic_tag_valid_out_1_29 = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  ic_tag_valid_out_1_30 = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  ic_tag_valid_out_1_31 = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  ic_tag_valid_out_1_32 = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  ic_tag_valid_out_1_33 = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  ic_tag_valid_out_1_34 = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  ic_tag_valid_out_1_35 = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  ic_tag_valid_out_1_36 = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  ic_tag_valid_out_1_37 = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  ic_tag_valid_out_1_38 = _RAND_193[0:0];
  _RAND_194 = {1{`RANDOM}};
  ic_tag_valid_out_1_39 = _RAND_194[0:0];
  _RAND_195 = {1{`RANDOM}};
  ic_tag_valid_out_1_40 = _RAND_195[0:0];
  _RAND_196 = {1{`RANDOM}};
  ic_tag_valid_out_1_41 = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  ic_tag_valid_out_1_42 = _RAND_197[0:0];
  _RAND_198 = {1{`RANDOM}};
  ic_tag_valid_out_1_43 = _RAND_198[0:0];
  _RAND_199 = {1{`RANDOM}};
  ic_tag_valid_out_1_44 = _RAND_199[0:0];
  _RAND_200 = {1{`RANDOM}};
  ic_tag_valid_out_1_45 = _RAND_200[0:0];
  _RAND_201 = {1{`RANDOM}};
  ic_tag_valid_out_1_46 = _RAND_201[0:0];
  _RAND_202 = {1{`RANDOM}};
  ic_tag_valid_out_1_47 = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  ic_tag_valid_out_1_48 = _RAND_203[0:0];
  _RAND_204 = {1{`RANDOM}};
  ic_tag_valid_out_1_49 = _RAND_204[0:0];
  _RAND_205 = {1{`RANDOM}};
  ic_tag_valid_out_1_50 = _RAND_205[0:0];
  _RAND_206 = {1{`RANDOM}};
  ic_tag_valid_out_1_51 = _RAND_206[0:0];
  _RAND_207 = {1{`RANDOM}};
  ic_tag_valid_out_1_52 = _RAND_207[0:0];
  _RAND_208 = {1{`RANDOM}};
  ic_tag_valid_out_1_53 = _RAND_208[0:0];
  _RAND_209 = {1{`RANDOM}};
  ic_tag_valid_out_1_54 = _RAND_209[0:0];
  _RAND_210 = {1{`RANDOM}};
  ic_tag_valid_out_1_55 = _RAND_210[0:0];
  _RAND_211 = {1{`RANDOM}};
  ic_tag_valid_out_1_56 = _RAND_211[0:0];
  _RAND_212 = {1{`RANDOM}};
  ic_tag_valid_out_1_57 = _RAND_212[0:0];
  _RAND_213 = {1{`RANDOM}};
  ic_tag_valid_out_1_58 = _RAND_213[0:0];
  _RAND_214 = {1{`RANDOM}};
  ic_tag_valid_out_1_59 = _RAND_214[0:0];
  _RAND_215 = {1{`RANDOM}};
  ic_tag_valid_out_1_60 = _RAND_215[0:0];
  _RAND_216 = {1{`RANDOM}};
  ic_tag_valid_out_1_61 = _RAND_216[0:0];
  _RAND_217 = {1{`RANDOM}};
  ic_tag_valid_out_1_62 = _RAND_217[0:0];
  _RAND_218 = {1{`RANDOM}};
  ic_tag_valid_out_1_63 = _RAND_218[0:0];
  _RAND_219 = {1{`RANDOM}};
  ic_tag_valid_out_1_64 = _RAND_219[0:0];
  _RAND_220 = {1{`RANDOM}};
  ic_tag_valid_out_1_65 = _RAND_220[0:0];
  _RAND_221 = {1{`RANDOM}};
  ic_tag_valid_out_1_66 = _RAND_221[0:0];
  _RAND_222 = {1{`RANDOM}};
  ic_tag_valid_out_1_67 = _RAND_222[0:0];
  _RAND_223 = {1{`RANDOM}};
  ic_tag_valid_out_1_68 = _RAND_223[0:0];
  _RAND_224 = {1{`RANDOM}};
  ic_tag_valid_out_1_69 = _RAND_224[0:0];
  _RAND_225 = {1{`RANDOM}};
  ic_tag_valid_out_1_70 = _RAND_225[0:0];
  _RAND_226 = {1{`RANDOM}};
  ic_tag_valid_out_1_71 = _RAND_226[0:0];
  _RAND_227 = {1{`RANDOM}};
  ic_tag_valid_out_1_72 = _RAND_227[0:0];
  _RAND_228 = {1{`RANDOM}};
  ic_tag_valid_out_1_73 = _RAND_228[0:0];
  _RAND_229 = {1{`RANDOM}};
  ic_tag_valid_out_1_74 = _RAND_229[0:0];
  _RAND_230 = {1{`RANDOM}};
  ic_tag_valid_out_1_75 = _RAND_230[0:0];
  _RAND_231 = {1{`RANDOM}};
  ic_tag_valid_out_1_76 = _RAND_231[0:0];
  _RAND_232 = {1{`RANDOM}};
  ic_tag_valid_out_1_77 = _RAND_232[0:0];
  _RAND_233 = {1{`RANDOM}};
  ic_tag_valid_out_1_78 = _RAND_233[0:0];
  _RAND_234 = {1{`RANDOM}};
  ic_tag_valid_out_1_79 = _RAND_234[0:0];
  _RAND_235 = {1{`RANDOM}};
  ic_tag_valid_out_1_80 = _RAND_235[0:0];
  _RAND_236 = {1{`RANDOM}};
  ic_tag_valid_out_1_81 = _RAND_236[0:0];
  _RAND_237 = {1{`RANDOM}};
  ic_tag_valid_out_1_82 = _RAND_237[0:0];
  _RAND_238 = {1{`RANDOM}};
  ic_tag_valid_out_1_83 = _RAND_238[0:0];
  _RAND_239 = {1{`RANDOM}};
  ic_tag_valid_out_1_84 = _RAND_239[0:0];
  _RAND_240 = {1{`RANDOM}};
  ic_tag_valid_out_1_85 = _RAND_240[0:0];
  _RAND_241 = {1{`RANDOM}};
  ic_tag_valid_out_1_86 = _RAND_241[0:0];
  _RAND_242 = {1{`RANDOM}};
  ic_tag_valid_out_1_87 = _RAND_242[0:0];
  _RAND_243 = {1{`RANDOM}};
  ic_tag_valid_out_1_88 = _RAND_243[0:0];
  _RAND_244 = {1{`RANDOM}};
  ic_tag_valid_out_1_89 = _RAND_244[0:0];
  _RAND_245 = {1{`RANDOM}};
  ic_tag_valid_out_1_90 = _RAND_245[0:0];
  _RAND_246 = {1{`RANDOM}};
  ic_tag_valid_out_1_91 = _RAND_246[0:0];
  _RAND_247 = {1{`RANDOM}};
  ic_tag_valid_out_1_92 = _RAND_247[0:0];
  _RAND_248 = {1{`RANDOM}};
  ic_tag_valid_out_1_93 = _RAND_248[0:0];
  _RAND_249 = {1{`RANDOM}};
  ic_tag_valid_out_1_94 = _RAND_249[0:0];
  _RAND_250 = {1{`RANDOM}};
  ic_tag_valid_out_1_95 = _RAND_250[0:0];
  _RAND_251 = {1{`RANDOM}};
  ic_tag_valid_out_1_96 = _RAND_251[0:0];
  _RAND_252 = {1{`RANDOM}};
  ic_tag_valid_out_1_97 = _RAND_252[0:0];
  _RAND_253 = {1{`RANDOM}};
  ic_tag_valid_out_1_98 = _RAND_253[0:0];
  _RAND_254 = {1{`RANDOM}};
  ic_tag_valid_out_1_99 = _RAND_254[0:0];
  _RAND_255 = {1{`RANDOM}};
  ic_tag_valid_out_1_100 = _RAND_255[0:0];
  _RAND_256 = {1{`RANDOM}};
  ic_tag_valid_out_1_101 = _RAND_256[0:0];
  _RAND_257 = {1{`RANDOM}};
  ic_tag_valid_out_1_102 = _RAND_257[0:0];
  _RAND_258 = {1{`RANDOM}};
  ic_tag_valid_out_1_103 = _RAND_258[0:0];
  _RAND_259 = {1{`RANDOM}};
  ic_tag_valid_out_1_104 = _RAND_259[0:0];
  _RAND_260 = {1{`RANDOM}};
  ic_tag_valid_out_1_105 = _RAND_260[0:0];
  _RAND_261 = {1{`RANDOM}};
  ic_tag_valid_out_1_106 = _RAND_261[0:0];
  _RAND_262 = {1{`RANDOM}};
  ic_tag_valid_out_1_107 = _RAND_262[0:0];
  _RAND_263 = {1{`RANDOM}};
  ic_tag_valid_out_1_108 = _RAND_263[0:0];
  _RAND_264 = {1{`RANDOM}};
  ic_tag_valid_out_1_109 = _RAND_264[0:0];
  _RAND_265 = {1{`RANDOM}};
  ic_tag_valid_out_1_110 = _RAND_265[0:0];
  _RAND_266 = {1{`RANDOM}};
  ic_tag_valid_out_1_111 = _RAND_266[0:0];
  _RAND_267 = {1{`RANDOM}};
  ic_tag_valid_out_1_112 = _RAND_267[0:0];
  _RAND_268 = {1{`RANDOM}};
  ic_tag_valid_out_1_113 = _RAND_268[0:0];
  _RAND_269 = {1{`RANDOM}};
  ic_tag_valid_out_1_114 = _RAND_269[0:0];
  _RAND_270 = {1{`RANDOM}};
  ic_tag_valid_out_1_115 = _RAND_270[0:0];
  _RAND_271 = {1{`RANDOM}};
  ic_tag_valid_out_1_116 = _RAND_271[0:0];
  _RAND_272 = {1{`RANDOM}};
  ic_tag_valid_out_1_117 = _RAND_272[0:0];
  _RAND_273 = {1{`RANDOM}};
  ic_tag_valid_out_1_118 = _RAND_273[0:0];
  _RAND_274 = {1{`RANDOM}};
  ic_tag_valid_out_1_119 = _RAND_274[0:0];
  _RAND_275 = {1{`RANDOM}};
  ic_tag_valid_out_1_120 = _RAND_275[0:0];
  _RAND_276 = {1{`RANDOM}};
  ic_tag_valid_out_1_121 = _RAND_276[0:0];
  _RAND_277 = {1{`RANDOM}};
  ic_tag_valid_out_1_122 = _RAND_277[0:0];
  _RAND_278 = {1{`RANDOM}};
  ic_tag_valid_out_1_123 = _RAND_278[0:0];
  _RAND_279 = {1{`RANDOM}};
  ic_tag_valid_out_1_124 = _RAND_279[0:0];
  _RAND_280 = {1{`RANDOM}};
  ic_tag_valid_out_1_125 = _RAND_280[0:0];
  _RAND_281 = {1{`RANDOM}};
  ic_tag_valid_out_1_126 = _RAND_281[0:0];
  _RAND_282 = {1{`RANDOM}};
  ic_tag_valid_out_1_127 = _RAND_282[0:0];
  _RAND_283 = {1{`RANDOM}};
  ic_tag_valid_out_0_0 = _RAND_283[0:0];
  _RAND_284 = {1{`RANDOM}};
  ic_tag_valid_out_0_1 = _RAND_284[0:0];
  _RAND_285 = {1{`RANDOM}};
  ic_tag_valid_out_0_2 = _RAND_285[0:0];
  _RAND_286 = {1{`RANDOM}};
  ic_tag_valid_out_0_3 = _RAND_286[0:0];
  _RAND_287 = {1{`RANDOM}};
  ic_tag_valid_out_0_4 = _RAND_287[0:0];
  _RAND_288 = {1{`RANDOM}};
  ic_tag_valid_out_0_5 = _RAND_288[0:0];
  _RAND_289 = {1{`RANDOM}};
  ic_tag_valid_out_0_6 = _RAND_289[0:0];
  _RAND_290 = {1{`RANDOM}};
  ic_tag_valid_out_0_7 = _RAND_290[0:0];
  _RAND_291 = {1{`RANDOM}};
  ic_tag_valid_out_0_8 = _RAND_291[0:0];
  _RAND_292 = {1{`RANDOM}};
  ic_tag_valid_out_0_9 = _RAND_292[0:0];
  _RAND_293 = {1{`RANDOM}};
  ic_tag_valid_out_0_10 = _RAND_293[0:0];
  _RAND_294 = {1{`RANDOM}};
  ic_tag_valid_out_0_11 = _RAND_294[0:0];
  _RAND_295 = {1{`RANDOM}};
  ic_tag_valid_out_0_12 = _RAND_295[0:0];
  _RAND_296 = {1{`RANDOM}};
  ic_tag_valid_out_0_13 = _RAND_296[0:0];
  _RAND_297 = {1{`RANDOM}};
  ic_tag_valid_out_0_14 = _RAND_297[0:0];
  _RAND_298 = {1{`RANDOM}};
  ic_tag_valid_out_0_15 = _RAND_298[0:0];
  _RAND_299 = {1{`RANDOM}};
  ic_tag_valid_out_0_16 = _RAND_299[0:0];
  _RAND_300 = {1{`RANDOM}};
  ic_tag_valid_out_0_17 = _RAND_300[0:0];
  _RAND_301 = {1{`RANDOM}};
  ic_tag_valid_out_0_18 = _RAND_301[0:0];
  _RAND_302 = {1{`RANDOM}};
  ic_tag_valid_out_0_19 = _RAND_302[0:0];
  _RAND_303 = {1{`RANDOM}};
  ic_tag_valid_out_0_20 = _RAND_303[0:0];
  _RAND_304 = {1{`RANDOM}};
  ic_tag_valid_out_0_21 = _RAND_304[0:0];
  _RAND_305 = {1{`RANDOM}};
  ic_tag_valid_out_0_22 = _RAND_305[0:0];
  _RAND_306 = {1{`RANDOM}};
  ic_tag_valid_out_0_23 = _RAND_306[0:0];
  _RAND_307 = {1{`RANDOM}};
  ic_tag_valid_out_0_24 = _RAND_307[0:0];
  _RAND_308 = {1{`RANDOM}};
  ic_tag_valid_out_0_25 = _RAND_308[0:0];
  _RAND_309 = {1{`RANDOM}};
  ic_tag_valid_out_0_26 = _RAND_309[0:0];
  _RAND_310 = {1{`RANDOM}};
  ic_tag_valid_out_0_27 = _RAND_310[0:0];
  _RAND_311 = {1{`RANDOM}};
  ic_tag_valid_out_0_28 = _RAND_311[0:0];
  _RAND_312 = {1{`RANDOM}};
  ic_tag_valid_out_0_29 = _RAND_312[0:0];
  _RAND_313 = {1{`RANDOM}};
  ic_tag_valid_out_0_30 = _RAND_313[0:0];
  _RAND_314 = {1{`RANDOM}};
  ic_tag_valid_out_0_31 = _RAND_314[0:0];
  _RAND_315 = {1{`RANDOM}};
  ic_tag_valid_out_0_32 = _RAND_315[0:0];
  _RAND_316 = {1{`RANDOM}};
  ic_tag_valid_out_0_33 = _RAND_316[0:0];
  _RAND_317 = {1{`RANDOM}};
  ic_tag_valid_out_0_34 = _RAND_317[0:0];
  _RAND_318 = {1{`RANDOM}};
  ic_tag_valid_out_0_35 = _RAND_318[0:0];
  _RAND_319 = {1{`RANDOM}};
  ic_tag_valid_out_0_36 = _RAND_319[0:0];
  _RAND_320 = {1{`RANDOM}};
  ic_tag_valid_out_0_37 = _RAND_320[0:0];
  _RAND_321 = {1{`RANDOM}};
  ic_tag_valid_out_0_38 = _RAND_321[0:0];
  _RAND_322 = {1{`RANDOM}};
  ic_tag_valid_out_0_39 = _RAND_322[0:0];
  _RAND_323 = {1{`RANDOM}};
  ic_tag_valid_out_0_40 = _RAND_323[0:0];
  _RAND_324 = {1{`RANDOM}};
  ic_tag_valid_out_0_41 = _RAND_324[0:0];
  _RAND_325 = {1{`RANDOM}};
  ic_tag_valid_out_0_42 = _RAND_325[0:0];
  _RAND_326 = {1{`RANDOM}};
  ic_tag_valid_out_0_43 = _RAND_326[0:0];
  _RAND_327 = {1{`RANDOM}};
  ic_tag_valid_out_0_44 = _RAND_327[0:0];
  _RAND_328 = {1{`RANDOM}};
  ic_tag_valid_out_0_45 = _RAND_328[0:0];
  _RAND_329 = {1{`RANDOM}};
  ic_tag_valid_out_0_46 = _RAND_329[0:0];
  _RAND_330 = {1{`RANDOM}};
  ic_tag_valid_out_0_47 = _RAND_330[0:0];
  _RAND_331 = {1{`RANDOM}};
  ic_tag_valid_out_0_48 = _RAND_331[0:0];
  _RAND_332 = {1{`RANDOM}};
  ic_tag_valid_out_0_49 = _RAND_332[0:0];
  _RAND_333 = {1{`RANDOM}};
  ic_tag_valid_out_0_50 = _RAND_333[0:0];
  _RAND_334 = {1{`RANDOM}};
  ic_tag_valid_out_0_51 = _RAND_334[0:0];
  _RAND_335 = {1{`RANDOM}};
  ic_tag_valid_out_0_52 = _RAND_335[0:0];
  _RAND_336 = {1{`RANDOM}};
  ic_tag_valid_out_0_53 = _RAND_336[0:0];
  _RAND_337 = {1{`RANDOM}};
  ic_tag_valid_out_0_54 = _RAND_337[0:0];
  _RAND_338 = {1{`RANDOM}};
  ic_tag_valid_out_0_55 = _RAND_338[0:0];
  _RAND_339 = {1{`RANDOM}};
  ic_tag_valid_out_0_56 = _RAND_339[0:0];
  _RAND_340 = {1{`RANDOM}};
  ic_tag_valid_out_0_57 = _RAND_340[0:0];
  _RAND_341 = {1{`RANDOM}};
  ic_tag_valid_out_0_58 = _RAND_341[0:0];
  _RAND_342 = {1{`RANDOM}};
  ic_tag_valid_out_0_59 = _RAND_342[0:0];
  _RAND_343 = {1{`RANDOM}};
  ic_tag_valid_out_0_60 = _RAND_343[0:0];
  _RAND_344 = {1{`RANDOM}};
  ic_tag_valid_out_0_61 = _RAND_344[0:0];
  _RAND_345 = {1{`RANDOM}};
  ic_tag_valid_out_0_62 = _RAND_345[0:0];
  _RAND_346 = {1{`RANDOM}};
  ic_tag_valid_out_0_63 = _RAND_346[0:0];
  _RAND_347 = {1{`RANDOM}};
  ic_tag_valid_out_0_64 = _RAND_347[0:0];
  _RAND_348 = {1{`RANDOM}};
  ic_tag_valid_out_0_65 = _RAND_348[0:0];
  _RAND_349 = {1{`RANDOM}};
  ic_tag_valid_out_0_66 = _RAND_349[0:0];
  _RAND_350 = {1{`RANDOM}};
  ic_tag_valid_out_0_67 = _RAND_350[0:0];
  _RAND_351 = {1{`RANDOM}};
  ic_tag_valid_out_0_68 = _RAND_351[0:0];
  _RAND_352 = {1{`RANDOM}};
  ic_tag_valid_out_0_69 = _RAND_352[0:0];
  _RAND_353 = {1{`RANDOM}};
  ic_tag_valid_out_0_70 = _RAND_353[0:0];
  _RAND_354 = {1{`RANDOM}};
  ic_tag_valid_out_0_71 = _RAND_354[0:0];
  _RAND_355 = {1{`RANDOM}};
  ic_tag_valid_out_0_72 = _RAND_355[0:0];
  _RAND_356 = {1{`RANDOM}};
  ic_tag_valid_out_0_73 = _RAND_356[0:0];
  _RAND_357 = {1{`RANDOM}};
  ic_tag_valid_out_0_74 = _RAND_357[0:0];
  _RAND_358 = {1{`RANDOM}};
  ic_tag_valid_out_0_75 = _RAND_358[0:0];
  _RAND_359 = {1{`RANDOM}};
  ic_tag_valid_out_0_76 = _RAND_359[0:0];
  _RAND_360 = {1{`RANDOM}};
  ic_tag_valid_out_0_77 = _RAND_360[0:0];
  _RAND_361 = {1{`RANDOM}};
  ic_tag_valid_out_0_78 = _RAND_361[0:0];
  _RAND_362 = {1{`RANDOM}};
  ic_tag_valid_out_0_79 = _RAND_362[0:0];
  _RAND_363 = {1{`RANDOM}};
  ic_tag_valid_out_0_80 = _RAND_363[0:0];
  _RAND_364 = {1{`RANDOM}};
  ic_tag_valid_out_0_81 = _RAND_364[0:0];
  _RAND_365 = {1{`RANDOM}};
  ic_tag_valid_out_0_82 = _RAND_365[0:0];
  _RAND_366 = {1{`RANDOM}};
  ic_tag_valid_out_0_83 = _RAND_366[0:0];
  _RAND_367 = {1{`RANDOM}};
  ic_tag_valid_out_0_84 = _RAND_367[0:0];
  _RAND_368 = {1{`RANDOM}};
  ic_tag_valid_out_0_85 = _RAND_368[0:0];
  _RAND_369 = {1{`RANDOM}};
  ic_tag_valid_out_0_86 = _RAND_369[0:0];
  _RAND_370 = {1{`RANDOM}};
  ic_tag_valid_out_0_87 = _RAND_370[0:0];
  _RAND_371 = {1{`RANDOM}};
  ic_tag_valid_out_0_88 = _RAND_371[0:0];
  _RAND_372 = {1{`RANDOM}};
  ic_tag_valid_out_0_89 = _RAND_372[0:0];
  _RAND_373 = {1{`RANDOM}};
  ic_tag_valid_out_0_90 = _RAND_373[0:0];
  _RAND_374 = {1{`RANDOM}};
  ic_tag_valid_out_0_91 = _RAND_374[0:0];
  _RAND_375 = {1{`RANDOM}};
  ic_tag_valid_out_0_92 = _RAND_375[0:0];
  _RAND_376 = {1{`RANDOM}};
  ic_tag_valid_out_0_93 = _RAND_376[0:0];
  _RAND_377 = {1{`RANDOM}};
  ic_tag_valid_out_0_94 = _RAND_377[0:0];
  _RAND_378 = {1{`RANDOM}};
  ic_tag_valid_out_0_95 = _RAND_378[0:0];
  _RAND_379 = {1{`RANDOM}};
  ic_tag_valid_out_0_96 = _RAND_379[0:0];
  _RAND_380 = {1{`RANDOM}};
  ic_tag_valid_out_0_97 = _RAND_380[0:0];
  _RAND_381 = {1{`RANDOM}};
  ic_tag_valid_out_0_98 = _RAND_381[0:0];
  _RAND_382 = {1{`RANDOM}};
  ic_tag_valid_out_0_99 = _RAND_382[0:0];
  _RAND_383 = {1{`RANDOM}};
  ic_tag_valid_out_0_100 = _RAND_383[0:0];
  _RAND_384 = {1{`RANDOM}};
  ic_tag_valid_out_0_101 = _RAND_384[0:0];
  _RAND_385 = {1{`RANDOM}};
  ic_tag_valid_out_0_102 = _RAND_385[0:0];
  _RAND_386 = {1{`RANDOM}};
  ic_tag_valid_out_0_103 = _RAND_386[0:0];
  _RAND_387 = {1{`RANDOM}};
  ic_tag_valid_out_0_104 = _RAND_387[0:0];
  _RAND_388 = {1{`RANDOM}};
  ic_tag_valid_out_0_105 = _RAND_388[0:0];
  _RAND_389 = {1{`RANDOM}};
  ic_tag_valid_out_0_106 = _RAND_389[0:0];
  _RAND_390 = {1{`RANDOM}};
  ic_tag_valid_out_0_107 = _RAND_390[0:0];
  _RAND_391 = {1{`RANDOM}};
  ic_tag_valid_out_0_108 = _RAND_391[0:0];
  _RAND_392 = {1{`RANDOM}};
  ic_tag_valid_out_0_109 = _RAND_392[0:0];
  _RAND_393 = {1{`RANDOM}};
  ic_tag_valid_out_0_110 = _RAND_393[0:0];
  _RAND_394 = {1{`RANDOM}};
  ic_tag_valid_out_0_111 = _RAND_394[0:0];
  _RAND_395 = {1{`RANDOM}};
  ic_tag_valid_out_0_112 = _RAND_395[0:0];
  _RAND_396 = {1{`RANDOM}};
  ic_tag_valid_out_0_113 = _RAND_396[0:0];
  _RAND_397 = {1{`RANDOM}};
  ic_tag_valid_out_0_114 = _RAND_397[0:0];
  _RAND_398 = {1{`RANDOM}};
  ic_tag_valid_out_0_115 = _RAND_398[0:0];
  _RAND_399 = {1{`RANDOM}};
  ic_tag_valid_out_0_116 = _RAND_399[0:0];
  _RAND_400 = {1{`RANDOM}};
  ic_tag_valid_out_0_117 = _RAND_400[0:0];
  _RAND_401 = {1{`RANDOM}};
  ic_tag_valid_out_0_118 = _RAND_401[0:0];
  _RAND_402 = {1{`RANDOM}};
  ic_tag_valid_out_0_119 = _RAND_402[0:0];
  _RAND_403 = {1{`RANDOM}};
  ic_tag_valid_out_0_120 = _RAND_403[0:0];
  _RAND_404 = {1{`RANDOM}};
  ic_tag_valid_out_0_121 = _RAND_404[0:0];
  _RAND_405 = {1{`RANDOM}};
  ic_tag_valid_out_0_122 = _RAND_405[0:0];
  _RAND_406 = {1{`RANDOM}};
  ic_tag_valid_out_0_123 = _RAND_406[0:0];
  _RAND_407 = {1{`RANDOM}};
  ic_tag_valid_out_0_124 = _RAND_407[0:0];
  _RAND_408 = {1{`RANDOM}};
  ic_tag_valid_out_0_125 = _RAND_408[0:0];
  _RAND_409 = {1{`RANDOM}};
  ic_tag_valid_out_0_126 = _RAND_409[0:0];
  _RAND_410 = {1{`RANDOM}};
  ic_tag_valid_out_0_127 = _RAND_410[0:0];
  _RAND_411 = {1{`RANDOM}};
  ic_debug_way_ff = _RAND_411[1:0];
  _RAND_412 = {1{`RANDOM}};
  ic_debug_rd_en_ff = _RAND_412[0:0];
  _RAND_413 = {3{`RANDOM}};
  _T_1212 = _RAND_413[70:0];
  _RAND_414 = {1{`RANDOM}};
  ifc_region_acc_fault_memory_f = _RAND_414[0:0];
  _RAND_415 = {1{`RANDOM}};
  perr_ic_index_ff = _RAND_415[6:0];
  _RAND_416 = {1{`RANDOM}};
  dma_sb_err_state_ff = _RAND_416[0:0];
  _RAND_417 = {1{`RANDOM}};
  bus_cmd_req_hold = _RAND_417[0:0];
  _RAND_418 = {1{`RANDOM}};
  ifu_bus_cmd_valid = _RAND_418[0:0];
  _RAND_419 = {1{`RANDOM}};
  ifu_bus_arvalid_ff = _RAND_419[0:0];
  _RAND_420 = {1{`RANDOM}};
  ifc_dma_access_ok_prev = _RAND_420[0:0];
  _RAND_421 = {2{`RANDOM}};
  iccm_ecc_corr_data_ff = _RAND_421[38:0];
  _RAND_422 = {1{`RANDOM}};
  dma_mem_addr_ff = _RAND_422[1:0];
  _RAND_423 = {1{`RANDOM}};
  dma_mem_tag_ff = _RAND_423[2:0];
  _RAND_424 = {1{`RANDOM}};
  iccm_dma_rtag_temp = _RAND_424[2:0];
  _RAND_425 = {1{`RANDOM}};
  iccm_dma_rvalid_temp = _RAND_425[0:0];
  _RAND_426 = {1{`RANDOM}};
  iccm_dma_ecc_error = _RAND_426[0:0];
  _RAND_427 = {2{`RANDOM}};
  iccm_dma_rdata_temp = _RAND_427[63:0];
  _RAND_428 = {1{`RANDOM}};
  iccm_ecc_corr_index_ff = _RAND_428[13:0];
  _RAND_429 = {1{`RANDOM}};
  iccm_rd_ecc_single_err_ff = _RAND_429[0:0];
  _RAND_430 = {1{`RANDOM}};
  iccm_rw_addr_f = _RAND_430[13:0];
  _RAND_431 = {1{`RANDOM}};
  ifu_status_wr_addr_ff = _RAND_431[6:0];
  _RAND_432 = {1{`RANDOM}};
  way_status_wr_en_ff = _RAND_432[0:0];
  _RAND_433 = {1{`RANDOM}};
  way_status_new_ff = _RAND_433[0:0];
  _RAND_434 = {1{`RANDOM}};
  ifu_tag_wren_ff = _RAND_434[1:0];
  _RAND_435 = {1{`RANDOM}};
  ic_valid_ff = _RAND_435[0:0];
  _RAND_436 = {1{`RANDOM}};
  _T_9799 = _RAND_436[0:0];
  _RAND_437 = {1{`RANDOM}};
  _T_9800 = _RAND_437[0:0];
  _RAND_438 = {1{`RANDOM}};
  _T_9801 = _RAND_438[0:0];
  _RAND_439 = {1{`RANDOM}};
  _T_9805 = _RAND_439[0:0];
  _RAND_440 = {1{`RANDOM}};
  _T_9826 = _RAND_440[0:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    flush_final_f = 1'h0;
  end
  if (reset) begin
    ifc_fetch_req_f_raw = 1'h0;
  end
  if (reset) begin
    miss_state = 3'h0;
  end
  if (reset) begin
    ifu_fetch_addr_int_f = 31'h0;
  end
  if (reset) begin
    ifc_iccm_access_f = 1'h0;
  end
  if (reset) begin
    iccm_dma_rvalid_in = 1'h0;
  end
  if (reset) begin
    dma_iccm_req_f = 1'h0;
  end
  if (reset) begin
    perr_state = 3'h0;
  end
  if (reset) begin
    err_stop_state = 2'h0;
  end
  if (reset) begin
    reset_all_tags = 1'h0;
  end
  if (reset) begin
    ifc_region_acc_fault_final_f = 1'h0;
  end
  if (reset) begin
    uncacheable_miss_ff = 1'h0;
  end
  if (reset) begin
    ic_miss_buff_data_valid = 8'h0;
  end
  if (reset) begin
    imb_ff = 31'h0;
  end
  if (reset) begin
    sel_mb_addr_ff = 1'h0;
  end
  if (reset) begin
    ifu_ic_rw_int_addr_ff = 7'h0;
  end
  if (reset) begin
    way_status_out_0 = 1'h0;
  end
  if (reset) begin
    way_status_out_1 = 1'h0;
  end
  if (reset) begin
    way_status_out_2 = 1'h0;
  end
  if (reset) begin
    way_status_out_3 = 1'h0;
  end
  if (reset) begin
    way_status_out_4 = 1'h0;
  end
  if (reset) begin
    way_status_out_5 = 1'h0;
  end
  if (reset) begin
    way_status_out_6 = 1'h0;
  end
  if (reset) begin
    way_status_out_7 = 1'h0;
  end
  if (reset) begin
    way_status_out_8 = 1'h0;
  end
  if (reset) begin
    way_status_out_9 = 1'h0;
  end
  if (reset) begin
    way_status_out_10 = 1'h0;
  end
  if (reset) begin
    way_status_out_11 = 1'h0;
  end
  if (reset) begin
    way_status_out_12 = 1'h0;
  end
  if (reset) begin
    way_status_out_13 = 1'h0;
  end
  if (reset) begin
    way_status_out_14 = 1'h0;
  end
  if (reset) begin
    way_status_out_15 = 1'h0;
  end
  if (reset) begin
    way_status_out_16 = 1'h0;
  end
  if (reset) begin
    way_status_out_17 = 1'h0;
  end
  if (reset) begin
    way_status_out_18 = 1'h0;
  end
  if (reset) begin
    way_status_out_19 = 1'h0;
  end
  if (reset) begin
    way_status_out_20 = 1'h0;
  end
  if (reset) begin
    way_status_out_21 = 1'h0;
  end
  if (reset) begin
    way_status_out_22 = 1'h0;
  end
  if (reset) begin
    way_status_out_23 = 1'h0;
  end
  if (reset) begin
    way_status_out_24 = 1'h0;
  end
  if (reset) begin
    way_status_out_25 = 1'h0;
  end
  if (reset) begin
    way_status_out_26 = 1'h0;
  end
  if (reset) begin
    way_status_out_27 = 1'h0;
  end
  if (reset) begin
    way_status_out_28 = 1'h0;
  end
  if (reset) begin
    way_status_out_29 = 1'h0;
  end
  if (reset) begin
    way_status_out_30 = 1'h0;
  end
  if (reset) begin
    way_status_out_31 = 1'h0;
  end
  if (reset) begin
    way_status_out_32 = 1'h0;
  end
  if (reset) begin
    way_status_out_33 = 1'h0;
  end
  if (reset) begin
    way_status_out_34 = 1'h0;
  end
  if (reset) begin
    way_status_out_35 = 1'h0;
  end
  if (reset) begin
    way_status_out_36 = 1'h0;
  end
  if (reset) begin
    way_status_out_37 = 1'h0;
  end
  if (reset) begin
    way_status_out_38 = 1'h0;
  end
  if (reset) begin
    way_status_out_39 = 1'h0;
  end
  if (reset) begin
    way_status_out_40 = 1'h0;
  end
  if (reset) begin
    way_status_out_41 = 1'h0;
  end
  if (reset) begin
    way_status_out_42 = 1'h0;
  end
  if (reset) begin
    way_status_out_43 = 1'h0;
  end
  if (reset) begin
    way_status_out_44 = 1'h0;
  end
  if (reset) begin
    way_status_out_45 = 1'h0;
  end
  if (reset) begin
    way_status_out_46 = 1'h0;
  end
  if (reset) begin
    way_status_out_47 = 1'h0;
  end
  if (reset) begin
    way_status_out_48 = 1'h0;
  end
  if (reset) begin
    way_status_out_49 = 1'h0;
  end
  if (reset) begin
    way_status_out_50 = 1'h0;
  end
  if (reset) begin
    way_status_out_51 = 1'h0;
  end
  if (reset) begin
    way_status_out_52 = 1'h0;
  end
  if (reset) begin
    way_status_out_53 = 1'h0;
  end
  if (reset) begin
    way_status_out_54 = 1'h0;
  end
  if (reset) begin
    way_status_out_55 = 1'h0;
  end
  if (reset) begin
    way_status_out_56 = 1'h0;
  end
  if (reset) begin
    way_status_out_57 = 1'h0;
  end
  if (reset) begin
    way_status_out_58 = 1'h0;
  end
  if (reset) begin
    way_status_out_59 = 1'h0;
  end
  if (reset) begin
    way_status_out_60 = 1'h0;
  end
  if (reset) begin
    way_status_out_61 = 1'h0;
  end
  if (reset) begin
    way_status_out_62 = 1'h0;
  end
  if (reset) begin
    way_status_out_63 = 1'h0;
  end
  if (reset) begin
    way_status_out_64 = 1'h0;
  end
  if (reset) begin
    way_status_out_65 = 1'h0;
  end
  if (reset) begin
    way_status_out_66 = 1'h0;
  end
  if (reset) begin
    way_status_out_67 = 1'h0;
  end
  if (reset) begin
    way_status_out_68 = 1'h0;
  end
  if (reset) begin
    way_status_out_69 = 1'h0;
  end
  if (reset) begin
    way_status_out_70 = 1'h0;
  end
  if (reset) begin
    way_status_out_71 = 1'h0;
  end
  if (reset) begin
    way_status_out_72 = 1'h0;
  end
  if (reset) begin
    way_status_out_73 = 1'h0;
  end
  if (reset) begin
    way_status_out_74 = 1'h0;
  end
  if (reset) begin
    way_status_out_75 = 1'h0;
  end
  if (reset) begin
    way_status_out_76 = 1'h0;
  end
  if (reset) begin
    way_status_out_77 = 1'h0;
  end
  if (reset) begin
    way_status_out_78 = 1'h0;
  end
  if (reset) begin
    way_status_out_79 = 1'h0;
  end
  if (reset) begin
    way_status_out_80 = 1'h0;
  end
  if (reset) begin
    way_status_out_81 = 1'h0;
  end
  if (reset) begin
    way_status_out_82 = 1'h0;
  end
  if (reset) begin
    way_status_out_83 = 1'h0;
  end
  if (reset) begin
    way_status_out_84 = 1'h0;
  end
  if (reset) begin
    way_status_out_85 = 1'h0;
  end
  if (reset) begin
    way_status_out_86 = 1'h0;
  end
  if (reset) begin
    way_status_out_87 = 1'h0;
  end
  if (reset) begin
    way_status_out_88 = 1'h0;
  end
  if (reset) begin
    way_status_out_89 = 1'h0;
  end
  if (reset) begin
    way_status_out_90 = 1'h0;
  end
  if (reset) begin
    way_status_out_91 = 1'h0;
  end
  if (reset) begin
    way_status_out_92 = 1'h0;
  end
  if (reset) begin
    way_status_out_93 = 1'h0;
  end
  if (reset) begin
    way_status_out_94 = 1'h0;
  end
  if (reset) begin
    way_status_out_95 = 1'h0;
  end
  if (reset) begin
    way_status_out_96 = 1'h0;
  end
  if (reset) begin
    way_status_out_97 = 1'h0;
  end
  if (reset) begin
    way_status_out_98 = 1'h0;
  end
  if (reset) begin
    way_status_out_99 = 1'h0;
  end
  if (reset) begin
    way_status_out_100 = 1'h0;
  end
  if (reset) begin
    way_status_out_101 = 1'h0;
  end
  if (reset) begin
    way_status_out_102 = 1'h0;
  end
  if (reset) begin
    way_status_out_103 = 1'h0;
  end
  if (reset) begin
    way_status_out_104 = 1'h0;
  end
  if (reset) begin
    way_status_out_105 = 1'h0;
  end
  if (reset) begin
    way_status_out_106 = 1'h0;
  end
  if (reset) begin
    way_status_out_107 = 1'h0;
  end
  if (reset) begin
    way_status_out_108 = 1'h0;
  end
  if (reset) begin
    way_status_out_109 = 1'h0;
  end
  if (reset) begin
    way_status_out_110 = 1'h0;
  end
  if (reset) begin
    way_status_out_111 = 1'h0;
  end
  if (reset) begin
    way_status_out_112 = 1'h0;
  end
  if (reset) begin
    way_status_out_113 = 1'h0;
  end
  if (reset) begin
    way_status_out_114 = 1'h0;
  end
  if (reset) begin
    way_status_out_115 = 1'h0;
  end
  if (reset) begin
    way_status_out_116 = 1'h0;
  end
  if (reset) begin
    way_status_out_117 = 1'h0;
  end
  if (reset) begin
    way_status_out_118 = 1'h0;
  end
  if (reset) begin
    way_status_out_119 = 1'h0;
  end
  if (reset) begin
    way_status_out_120 = 1'h0;
  end
  if (reset) begin
    way_status_out_121 = 1'h0;
  end
  if (reset) begin
    way_status_out_122 = 1'h0;
  end
  if (reset) begin
    way_status_out_123 = 1'h0;
  end
  if (reset) begin
    way_status_out_124 = 1'h0;
  end
  if (reset) begin
    way_status_out_125 = 1'h0;
  end
  if (reset) begin
    way_status_out_126 = 1'h0;
  end
  if (reset) begin
    way_status_out_127 = 1'h0;
  end
  if (reset) begin
    way_status_mb_ff = 1'h0;
  end
  if (reset) begin
    tagv_mb_ff = 2'h0;
  end
  if (reset) begin
    reset_ic_ff = 1'h0;
  end
  if (reset) begin
    fetch_uncacheable_ff = 1'h0;
  end
  if (reset) begin
    miss_addr = 26'h0;
  end
  if (reset) begin
    ifc_region_acc_fault_f = 1'h0;
  end
  if (reset) begin
    bus_rd_addr_count = 3'h0;
  end
  if (reset) begin
    ic_act_miss_f_delayed = 1'h0;
  end
  if (reset) begin
    ic_crit_wd_rdy_new_ff = 1'h0;
  end
  if (reset) begin
    ic_miss_buff_data_error = 8'h0;
  end
  if (reset) begin
    ic_debug_ict_array_sel_ff = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_0 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_1 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_2 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_3 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_4 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_5 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_6 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_7 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_8 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_9 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_10 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_11 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_12 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_13 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_14 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_15 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_16 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_17 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_18 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_19 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_20 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_21 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_22 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_23 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_24 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_25 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_26 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_27 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_28 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_29 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_30 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_31 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_32 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_33 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_34 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_35 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_36 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_37 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_38 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_39 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_40 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_41 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_42 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_43 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_44 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_45 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_46 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_47 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_48 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_49 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_50 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_51 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_52 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_53 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_54 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_55 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_56 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_57 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_58 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_59 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_60 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_61 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_62 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_63 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_64 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_65 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_66 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_67 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_68 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_69 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_70 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_71 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_72 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_73 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_74 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_75 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_76 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_77 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_78 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_79 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_80 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_81 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_82 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_83 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_84 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_85 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_86 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_87 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_88 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_89 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_90 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_91 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_92 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_93 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_94 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_95 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_96 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_97 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_98 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_99 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_100 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_101 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_102 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_103 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_104 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_105 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_106 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_107 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_108 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_109 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_110 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_111 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_112 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_113 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_114 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_115 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_116 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_117 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_118 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_119 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_120 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_121 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_122 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_123 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_124 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_125 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_126 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_127 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_0 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_1 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_2 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_3 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_4 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_5 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_6 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_7 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_8 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_9 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_10 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_11 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_12 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_13 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_14 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_15 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_16 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_17 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_18 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_19 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_20 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_21 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_22 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_23 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_24 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_25 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_26 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_27 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_28 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_29 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_30 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_31 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_32 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_33 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_34 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_35 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_36 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_37 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_38 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_39 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_40 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_41 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_42 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_43 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_44 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_45 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_46 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_47 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_48 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_49 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_50 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_51 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_52 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_53 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_54 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_55 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_56 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_57 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_58 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_59 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_60 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_61 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_62 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_63 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_64 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_65 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_66 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_67 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_68 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_69 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_70 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_71 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_72 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_73 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_74 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_75 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_76 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_77 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_78 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_79 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_80 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_81 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_82 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_83 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_84 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_85 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_86 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_87 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_88 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_89 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_90 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_91 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_92 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_93 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_94 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_95 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_96 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_97 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_98 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_99 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_100 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_101 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_102 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_103 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_104 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_105 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_106 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_107 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_108 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_109 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_110 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_111 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_112 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_113 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_114 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_115 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_116 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_117 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_118 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_119 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_120 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_121 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_122 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_123 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_124 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_125 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_126 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_127 = 1'h0;
  end
  if (reset) begin
    ic_debug_way_ff = 2'h0;
  end
  if (reset) begin
    ic_debug_rd_en_ff = 1'h0;
  end
  if (reset) begin
    _T_1212 = 71'h0;
  end
  if (reset) begin
    ifc_region_acc_fault_memory_f = 1'h0;
  end
  if (reset) begin
    perr_ic_index_ff = 7'h0;
  end
  if (reset) begin
    dma_sb_err_state_ff = 1'h0;
  end
  if (reset) begin
    bus_cmd_req_hold = 1'h0;
  end
  if (reset) begin
    ifu_bus_cmd_valid = 1'h0;
  end
  if (reset) begin
    ifu_bus_arvalid_ff = 1'h0;
  end
  if (reset) begin
    ifc_dma_access_ok_prev = 1'h0;
  end
  if (reset) begin
    iccm_ecc_corr_data_ff = 39'h0;
  end
  if (reset) begin
    dma_mem_addr_ff = 2'h0;
  end
  if (reset) begin
    dma_mem_tag_ff = 3'h0;
  end
  if (reset) begin
    iccm_dma_rtag_temp = 3'h0;
  end
  if (reset) begin
    iccm_dma_rvalid_temp = 1'h0;
  end
  if (reset) begin
    iccm_dma_ecc_error = 1'h0;
  end
  if (reset) begin
    iccm_dma_rdata_temp = 64'h0;
  end
  if (reset) begin
    iccm_ecc_corr_index_ff = 14'h0;
  end
  if (reset) begin
    iccm_rd_ecc_single_err_ff = 1'h0;
  end
  if (reset) begin
    iccm_rw_addr_f = 14'h0;
  end
  if (reset) begin
    ifu_status_wr_addr_ff = 7'h0;
  end
  if (reset) begin
    way_status_wr_en_ff = 1'h0;
  end
  if (reset) begin
    way_status_new_ff = 1'h0;
  end
  if (reset) begin
    ifu_tag_wren_ff = 2'h0;
  end
  if (reset) begin
    ic_valid_ff = 1'h0;
  end
  if (reset) begin
    _T_9799 = 1'h0;
  end
  if (reset) begin
    _T_9800 = 1'h0;
  end
  if (reset) begin
    _T_9801 = 1'h0;
  end
  if (reset) begin
    _T_9805 = 1'h0;
  end
  if (reset) begin
    _T_9826 = 1'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      flush_final_f <= 1'h0;
    end else begin
      flush_final_f <= io_exu_flush_final;
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      ifc_fetch_req_f_raw <= 1'h0;
    end else begin
      ifc_fetch_req_f_raw <= _T_317 & _T_318;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      miss_state <= 3'h0;
    end else if (miss_state_en) begin
      if (_T_24) begin
        if (_T_26) begin
          miss_state <= 3'h1;
        end else begin
          miss_state <= 3'h2;
        end
      end else if (_T_31) begin
        if (io_dec_mem_ctrl_dec_tlu_force_halt) begin
          miss_state <= 3'h0;
        end else if (_T_40) begin
          miss_state <= 3'h3;
        end else if (_T_61) begin
          miss_state <= 3'h6;
        end else if (_T_81) begin
          miss_state <= 3'h2;
        end else begin
          miss_state <= 3'h0;
        end
      end else if (_T_102) begin
        miss_state <= 3'h0;
      end else if (_T_106) begin
        if (_T_113) begin
          miss_state <= 3'h2;
        end else begin
          miss_state <= 3'h0;
        end
      end else if (_T_121) begin
        if (_T_126) begin
          miss_state <= 3'h2;
        end else begin
          miss_state <= 3'h0;
        end
      end else if (_T_132) begin
        if (_T_137) begin
          miss_state <= 3'h5;
        end else if (_T_143) begin
          miss_state <= 3'h7;
        end else begin
          miss_state <= 3'h0;
        end
      end else if (_T_151) begin
        if (io_dec_mem_ctrl_dec_tlu_force_halt) begin
          miss_state <= 3'h0;
        end else if (io_exu_flush_final) begin
          miss_state <= 3'h2;
        end else begin
          miss_state <= 3'h1;
        end
      end else if (_T_160) begin
        if (io_dec_mem_ctrl_dec_tlu_force_halt) begin
          miss_state <= 3'h0;
        end else if (io_exu_flush_final) begin
          miss_state <= 3'h2;
        end else begin
          miss_state <= 3'h0;
        end
      end else begin
        miss_state <= 3'h0;
      end
    end
  end
  always @(posedge rvclkhdr_2_io_l1clk or posedge reset) begin
    if (reset) begin
      ifu_fetch_addr_int_f <= 31'h0;
    end else begin
      ifu_fetch_addr_int_f <= io_ifc_fetch_addr_bf;
    end
  end
  always @(posedge rvclkhdr_2_io_l1clk or posedge reset) begin
    if (reset) begin
      ifc_iccm_access_f <= 1'h0;
    end else begin
      ifc_iccm_access_f <= io_ifc_iccm_access_bf;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      iccm_dma_rvalid_in <= 1'h0;
    end else begin
      iccm_dma_rvalid_in <= _T_2709 & _T_2713;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      dma_iccm_req_f <= 1'h0;
    end else begin
      dma_iccm_req_f <= io_dma_mem_ctl_dma_iccm_req;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      perr_state <= 3'h0;
    end else if (perr_state_en) begin
      if (_T_2500) begin
        if (io_iccm_dma_sb_error) begin
          perr_state <= 3'h4;
        end else if (_T_2502) begin
          perr_state <= 3'h1;
        end else begin
          perr_state <= 3'h2;
        end
      end else if (_T_2512) begin
        perr_state <= 3'h0;
      end else if (_T_2515) begin
        if (_T_2518) begin
          perr_state <= 3'h0;
        end else begin
          perr_state <= 3'h3;
        end
      end else if (_T_2522) begin
        if (io_dec_mem_ctrl_dec_tlu_force_halt) begin
          perr_state <= 3'h0;
        end else begin
          perr_state <= 3'h3;
        end
      end else begin
        perr_state <= 3'h0;
      end
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      err_stop_state <= 2'h0;
    end else if (err_stop_state_en) begin
      if (_T_2526) begin
        err_stop_state <= 2'h1;
      end else if (_T_2531) begin
        if (_T_2533) begin
          err_stop_state <= 2'h0;
        end else if (_T_2554) begin
          err_stop_state <= 2'h3;
        end else if (io_ifu_fetch_val[0]) begin
          err_stop_state <= 2'h2;
        end else begin
          err_stop_state <= 2'h1;
        end
      end else if (_T_2558) begin
        if (_T_2533) begin
          err_stop_state <= 2'h0;
        end else if (io_ifu_fetch_val[0]) begin
          err_stop_state <= 2'h3;
        end else begin
          err_stop_state <= 2'h2;
        end
      end else if (_T_2575) begin
        if (_T_2579) begin
          err_stop_state <= 2'h0;
        end else if (io_dec_mem_ctrl_dec_tlu_flush_err_wb) begin
          err_stop_state <= 2'h1;
        end else begin
          err_stop_state <= 2'h3;
        end
      end else begin
        err_stop_state <= 2'h0;
      end
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      reset_all_tags <= 1'h0;
    end else begin
      reset_all_tags <= io_dec_mem_ctrl_dec_tlu_fence_i_wb;
    end
  end
  always @(posedge rvclkhdr_2_io_l1clk or posedge reset) begin
    if (reset) begin
      ifc_region_acc_fault_final_f <= 1'h0;
    end else begin
      ifc_region_acc_fault_final_f <= io_ifc_region_acc_fault_bf | ifc_region_acc_fault_memory_bf;
    end
  end
  always @(posedge rvclkhdr_2_io_l1clk or posedge reset) begin
    if (reset) begin
      uncacheable_miss_ff <= 1'h0;
    end else if (!(sel_hold_imb)) begin
      uncacheable_miss_ff <= io_ifc_fetch_uncacheable_bf;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      ic_miss_buff_data_valid <= 8'h0;
    end else begin
      ic_miss_buff_data_valid <= {_T_1358,ic_miss_buff_data_valid_in_0};
    end
  end
  always @(posedge rvclkhdr_2_io_l1clk or posedge reset) begin
    if (reset) begin
      imb_ff <= 31'h0;
    end else if (!(sel_hold_imb)) begin
      imb_ff <= io_ifc_fetch_addr_bf;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      sel_mb_addr_ff <= 1'h0;
    end else begin
      sel_mb_addr_ff <= _T_2687 & _T_17;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      ifu_ic_rw_int_addr_ff <= 7'h0;
    end else if (_T_3997) begin
      ifu_ic_rw_int_addr_ff <= io_ic_debug_addr[9:3];
    end else begin
      ifu_ic_rw_int_addr_ff <= ifu_ic_rw_int_addr[11:5];
    end
  end
  always @(posedge rvclkhdr_70_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_0 <= 1'h0;
    end else if (_T_4021) begin
      way_status_out_0 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_70_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_1 <= 1'h0;
    end else if (_T_4025) begin
      way_status_out_1 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_70_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_2 <= 1'h0;
    end else if (_T_4029) begin
      way_status_out_2 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_70_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_3 <= 1'h0;
    end else if (_T_4033) begin
      way_status_out_3 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_70_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_4 <= 1'h0;
    end else if (_T_4037) begin
      way_status_out_4 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_70_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_5 <= 1'h0;
    end else if (_T_4041) begin
      way_status_out_5 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_70_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_6 <= 1'h0;
    end else if (_T_4045) begin
      way_status_out_6 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_70_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_7 <= 1'h0;
    end else if (_T_4049) begin
      way_status_out_7 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_71_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_8 <= 1'h0;
    end else if (_T_4021) begin
      way_status_out_8 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_71_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_9 <= 1'h0;
    end else if (_T_4025) begin
      way_status_out_9 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_71_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_10 <= 1'h0;
    end else if (_T_4029) begin
      way_status_out_10 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_71_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_11 <= 1'h0;
    end else if (_T_4033) begin
      way_status_out_11 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_71_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_12 <= 1'h0;
    end else if (_T_4037) begin
      way_status_out_12 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_71_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_13 <= 1'h0;
    end else if (_T_4041) begin
      way_status_out_13 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_71_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_14 <= 1'h0;
    end else if (_T_4045) begin
      way_status_out_14 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_71_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_15 <= 1'h0;
    end else if (_T_4049) begin
      way_status_out_15 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_72_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_16 <= 1'h0;
    end else if (_T_4021) begin
      way_status_out_16 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_72_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_17 <= 1'h0;
    end else if (_T_4025) begin
      way_status_out_17 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_72_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_18 <= 1'h0;
    end else if (_T_4029) begin
      way_status_out_18 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_72_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_19 <= 1'h0;
    end else if (_T_4033) begin
      way_status_out_19 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_72_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_20 <= 1'h0;
    end else if (_T_4037) begin
      way_status_out_20 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_72_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_21 <= 1'h0;
    end else if (_T_4041) begin
      way_status_out_21 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_72_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_22 <= 1'h0;
    end else if (_T_4045) begin
      way_status_out_22 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_72_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_23 <= 1'h0;
    end else if (_T_4049) begin
      way_status_out_23 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_73_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_24 <= 1'h0;
    end else if (_T_4021) begin
      way_status_out_24 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_73_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_25 <= 1'h0;
    end else if (_T_4025) begin
      way_status_out_25 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_73_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_26 <= 1'h0;
    end else if (_T_4029) begin
      way_status_out_26 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_73_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_27 <= 1'h0;
    end else if (_T_4033) begin
      way_status_out_27 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_73_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_28 <= 1'h0;
    end else if (_T_4037) begin
      way_status_out_28 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_73_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_29 <= 1'h0;
    end else if (_T_4041) begin
      way_status_out_29 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_73_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_30 <= 1'h0;
    end else if (_T_4045) begin
      way_status_out_30 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_73_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_31 <= 1'h0;
    end else if (_T_4049) begin
      way_status_out_31 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_74_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_32 <= 1'h0;
    end else if (_T_4021) begin
      way_status_out_32 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_74_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_33 <= 1'h0;
    end else if (_T_4025) begin
      way_status_out_33 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_74_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_34 <= 1'h0;
    end else if (_T_4029) begin
      way_status_out_34 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_74_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_35 <= 1'h0;
    end else if (_T_4033) begin
      way_status_out_35 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_74_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_36 <= 1'h0;
    end else if (_T_4037) begin
      way_status_out_36 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_74_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_37 <= 1'h0;
    end else if (_T_4041) begin
      way_status_out_37 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_74_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_38 <= 1'h0;
    end else if (_T_4045) begin
      way_status_out_38 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_74_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_39 <= 1'h0;
    end else if (_T_4049) begin
      way_status_out_39 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_75_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_40 <= 1'h0;
    end else if (_T_4021) begin
      way_status_out_40 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_75_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_41 <= 1'h0;
    end else if (_T_4025) begin
      way_status_out_41 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_75_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_42 <= 1'h0;
    end else if (_T_4029) begin
      way_status_out_42 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_75_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_43 <= 1'h0;
    end else if (_T_4033) begin
      way_status_out_43 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_75_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_44 <= 1'h0;
    end else if (_T_4037) begin
      way_status_out_44 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_75_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_45 <= 1'h0;
    end else if (_T_4041) begin
      way_status_out_45 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_75_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_46 <= 1'h0;
    end else if (_T_4045) begin
      way_status_out_46 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_75_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_47 <= 1'h0;
    end else if (_T_4049) begin
      way_status_out_47 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_76_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_48 <= 1'h0;
    end else if (_T_4021) begin
      way_status_out_48 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_76_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_49 <= 1'h0;
    end else if (_T_4025) begin
      way_status_out_49 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_76_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_50 <= 1'h0;
    end else if (_T_4029) begin
      way_status_out_50 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_76_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_51 <= 1'h0;
    end else if (_T_4033) begin
      way_status_out_51 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_76_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_52 <= 1'h0;
    end else if (_T_4037) begin
      way_status_out_52 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_76_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_53 <= 1'h0;
    end else if (_T_4041) begin
      way_status_out_53 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_76_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_54 <= 1'h0;
    end else if (_T_4045) begin
      way_status_out_54 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_76_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_55 <= 1'h0;
    end else if (_T_4049) begin
      way_status_out_55 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_77_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_56 <= 1'h0;
    end else if (_T_4021) begin
      way_status_out_56 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_77_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_57 <= 1'h0;
    end else if (_T_4025) begin
      way_status_out_57 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_77_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_58 <= 1'h0;
    end else if (_T_4029) begin
      way_status_out_58 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_77_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_59 <= 1'h0;
    end else if (_T_4033) begin
      way_status_out_59 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_77_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_60 <= 1'h0;
    end else if (_T_4037) begin
      way_status_out_60 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_77_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_61 <= 1'h0;
    end else if (_T_4041) begin
      way_status_out_61 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_77_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_62 <= 1'h0;
    end else if (_T_4045) begin
      way_status_out_62 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_77_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_63 <= 1'h0;
    end else if (_T_4049) begin
      way_status_out_63 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_78_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_64 <= 1'h0;
    end else if (_T_4021) begin
      way_status_out_64 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_78_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_65 <= 1'h0;
    end else if (_T_4025) begin
      way_status_out_65 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_78_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_66 <= 1'h0;
    end else if (_T_4029) begin
      way_status_out_66 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_78_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_67 <= 1'h0;
    end else if (_T_4033) begin
      way_status_out_67 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_78_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_68 <= 1'h0;
    end else if (_T_4037) begin
      way_status_out_68 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_78_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_69 <= 1'h0;
    end else if (_T_4041) begin
      way_status_out_69 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_78_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_70 <= 1'h0;
    end else if (_T_4045) begin
      way_status_out_70 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_78_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_71 <= 1'h0;
    end else if (_T_4049) begin
      way_status_out_71 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_79_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_72 <= 1'h0;
    end else if (_T_4021) begin
      way_status_out_72 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_79_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_73 <= 1'h0;
    end else if (_T_4025) begin
      way_status_out_73 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_79_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_74 <= 1'h0;
    end else if (_T_4029) begin
      way_status_out_74 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_79_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_75 <= 1'h0;
    end else if (_T_4033) begin
      way_status_out_75 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_79_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_76 <= 1'h0;
    end else if (_T_4037) begin
      way_status_out_76 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_79_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_77 <= 1'h0;
    end else if (_T_4041) begin
      way_status_out_77 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_79_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_78 <= 1'h0;
    end else if (_T_4045) begin
      way_status_out_78 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_79_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_79 <= 1'h0;
    end else if (_T_4049) begin
      way_status_out_79 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_80_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_80 <= 1'h0;
    end else if (_T_4021) begin
      way_status_out_80 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_80_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_81 <= 1'h0;
    end else if (_T_4025) begin
      way_status_out_81 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_80_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_82 <= 1'h0;
    end else if (_T_4029) begin
      way_status_out_82 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_80_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_83 <= 1'h0;
    end else if (_T_4033) begin
      way_status_out_83 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_80_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_84 <= 1'h0;
    end else if (_T_4037) begin
      way_status_out_84 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_80_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_85 <= 1'h0;
    end else if (_T_4041) begin
      way_status_out_85 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_80_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_86 <= 1'h0;
    end else if (_T_4045) begin
      way_status_out_86 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_80_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_87 <= 1'h0;
    end else if (_T_4049) begin
      way_status_out_87 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_81_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_88 <= 1'h0;
    end else if (_T_4021) begin
      way_status_out_88 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_81_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_89 <= 1'h0;
    end else if (_T_4025) begin
      way_status_out_89 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_81_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_90 <= 1'h0;
    end else if (_T_4029) begin
      way_status_out_90 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_81_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_91 <= 1'h0;
    end else if (_T_4033) begin
      way_status_out_91 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_81_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_92 <= 1'h0;
    end else if (_T_4037) begin
      way_status_out_92 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_81_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_93 <= 1'h0;
    end else if (_T_4041) begin
      way_status_out_93 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_81_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_94 <= 1'h0;
    end else if (_T_4045) begin
      way_status_out_94 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_81_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_95 <= 1'h0;
    end else if (_T_4049) begin
      way_status_out_95 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_82_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_96 <= 1'h0;
    end else if (_T_4021) begin
      way_status_out_96 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_82_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_97 <= 1'h0;
    end else if (_T_4025) begin
      way_status_out_97 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_82_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_98 <= 1'h0;
    end else if (_T_4029) begin
      way_status_out_98 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_82_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_99 <= 1'h0;
    end else if (_T_4033) begin
      way_status_out_99 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_82_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_100 <= 1'h0;
    end else if (_T_4037) begin
      way_status_out_100 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_82_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_101 <= 1'h0;
    end else if (_T_4041) begin
      way_status_out_101 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_82_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_102 <= 1'h0;
    end else if (_T_4045) begin
      way_status_out_102 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_82_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_103 <= 1'h0;
    end else if (_T_4049) begin
      way_status_out_103 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_83_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_104 <= 1'h0;
    end else if (_T_4021) begin
      way_status_out_104 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_83_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_105 <= 1'h0;
    end else if (_T_4025) begin
      way_status_out_105 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_83_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_106 <= 1'h0;
    end else if (_T_4029) begin
      way_status_out_106 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_83_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_107 <= 1'h0;
    end else if (_T_4033) begin
      way_status_out_107 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_83_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_108 <= 1'h0;
    end else if (_T_4037) begin
      way_status_out_108 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_83_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_109 <= 1'h0;
    end else if (_T_4041) begin
      way_status_out_109 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_83_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_110 <= 1'h0;
    end else if (_T_4045) begin
      way_status_out_110 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_83_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_111 <= 1'h0;
    end else if (_T_4049) begin
      way_status_out_111 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_84_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_112 <= 1'h0;
    end else if (_T_4021) begin
      way_status_out_112 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_84_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_113 <= 1'h0;
    end else if (_T_4025) begin
      way_status_out_113 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_84_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_114 <= 1'h0;
    end else if (_T_4029) begin
      way_status_out_114 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_84_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_115 <= 1'h0;
    end else if (_T_4033) begin
      way_status_out_115 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_84_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_116 <= 1'h0;
    end else if (_T_4037) begin
      way_status_out_116 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_84_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_117 <= 1'h0;
    end else if (_T_4041) begin
      way_status_out_117 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_84_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_118 <= 1'h0;
    end else if (_T_4045) begin
      way_status_out_118 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_84_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_119 <= 1'h0;
    end else if (_T_4049) begin
      way_status_out_119 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_85_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_120 <= 1'h0;
    end else if (_T_4021) begin
      way_status_out_120 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_85_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_121 <= 1'h0;
    end else if (_T_4025) begin
      way_status_out_121 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_85_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_122 <= 1'h0;
    end else if (_T_4029) begin
      way_status_out_122 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_85_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_123 <= 1'h0;
    end else if (_T_4033) begin
      way_status_out_123 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_85_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_124 <= 1'h0;
    end else if (_T_4037) begin
      way_status_out_124 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_85_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_125 <= 1'h0;
    end else if (_T_4041) begin
      way_status_out_125 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_85_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_126 <= 1'h0;
    end else if (_T_4045) begin
      way_status_out_126 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_85_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_127 <= 1'h0;
    end else if (_T_4049) begin
      way_status_out_127 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_2_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_mb_ff <= 1'h0;
    end else if (!(miss_pending)) begin
      way_status_mb_ff <= way_status;
    end
  end
  always @(posedge rvclkhdr_2_io_l1clk or posedge reset) begin
    if (reset) begin
      tagv_mb_ff <= 2'h0;
    end else if (!(miss_pending)) begin
      tagv_mb_ff <= _T_295;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      reset_ic_ff <= 1'h0;
    end else begin
      reset_ic_ff <= miss_pending & _T_299;
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      fetch_uncacheable_ff <= 1'h0;
    end else begin
      fetch_uncacheable_ff <= io_ifc_fetch_uncacheable_bf;
    end
  end
  always @(posedge rvclkhdr_3_io_l1clk or posedge reset) begin
    if (reset) begin
      miss_addr <= 26'h0;
    end else if (_T_231) begin
      miss_addr <= imb_ff[30:5];
    end
  end
  always @(posedge rvclkhdr_2_io_l1clk or posedge reset) begin
    if (reset) begin
      ifc_region_acc_fault_f <= 1'h0;
    end else begin
      ifc_region_acc_fault_f <= io_ifc_region_acc_fault_bf;
    end
  end
  always @(posedge rvclkhdr_3_io_l1clk or posedge reset) begin
    if (reset) begin
      bus_rd_addr_count <= 3'h0;
    end else if (_T_231) begin
      bus_rd_addr_count <= imb_ff[4:2];
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      ic_act_miss_f_delayed <= 1'h0;
    end else begin
      ic_act_miss_f_delayed <= _T_232 & _T_209;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      ic_crit_wd_rdy_new_ff <= 1'h0;
    end else begin
      ic_crit_wd_rdy_new_ff <= _T_1514 | _T_1519;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      ic_miss_buff_data_error <= 8'h0;
    end else begin
      ic_miss_buff_data_error <= {_T_1398,ic_miss_buff_data_error_in_0};
    end
  end
  always @(posedge rvclkhdr_1_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_debug_ict_array_sel_ff <= 1'h0;
    end else begin
      ic_debug_ict_array_sel_ff <= io_ic_debug_rd_en & io_ic_debug_tag_array;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_0 <= 1'h0;
    end else if (_T_5642) begin
      ic_tag_valid_out_1_0 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_1 <= 1'h0;
    end else if (_T_5657) begin
      ic_tag_valid_out_1_1 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_2 <= 1'h0;
    end else if (_T_5672) begin
      ic_tag_valid_out_1_2 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_3 <= 1'h0;
    end else if (_T_5687) begin
      ic_tag_valid_out_1_3 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_4 <= 1'h0;
    end else if (_T_5702) begin
      ic_tag_valid_out_1_4 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_5 <= 1'h0;
    end else if (_T_5717) begin
      ic_tag_valid_out_1_5 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_6 <= 1'h0;
    end else if (_T_5732) begin
      ic_tag_valid_out_1_6 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_7 <= 1'h0;
    end else if (_T_5747) begin
      ic_tag_valid_out_1_7 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_8 <= 1'h0;
    end else if (_T_5762) begin
      ic_tag_valid_out_1_8 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_9 <= 1'h0;
    end else if (_T_5777) begin
      ic_tag_valid_out_1_9 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_10 <= 1'h0;
    end else if (_T_5792) begin
      ic_tag_valid_out_1_10 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_11 <= 1'h0;
    end else if (_T_5807) begin
      ic_tag_valid_out_1_11 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_12 <= 1'h0;
    end else if (_T_5822) begin
      ic_tag_valid_out_1_12 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_13 <= 1'h0;
    end else if (_T_5837) begin
      ic_tag_valid_out_1_13 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_14 <= 1'h0;
    end else if (_T_5852) begin
      ic_tag_valid_out_1_14 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_15 <= 1'h0;
    end else if (_T_5867) begin
      ic_tag_valid_out_1_15 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_16 <= 1'h0;
    end else if (_T_5882) begin
      ic_tag_valid_out_1_16 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_17 <= 1'h0;
    end else if (_T_5897) begin
      ic_tag_valid_out_1_17 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_18 <= 1'h0;
    end else if (_T_5912) begin
      ic_tag_valid_out_1_18 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_19 <= 1'h0;
    end else if (_T_5927) begin
      ic_tag_valid_out_1_19 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_20 <= 1'h0;
    end else if (_T_5942) begin
      ic_tag_valid_out_1_20 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_21 <= 1'h0;
    end else if (_T_5957) begin
      ic_tag_valid_out_1_21 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_22 <= 1'h0;
    end else if (_T_5972) begin
      ic_tag_valid_out_1_22 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_23 <= 1'h0;
    end else if (_T_5987) begin
      ic_tag_valid_out_1_23 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_24 <= 1'h0;
    end else if (_T_6002) begin
      ic_tag_valid_out_1_24 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_25 <= 1'h0;
    end else if (_T_6017) begin
      ic_tag_valid_out_1_25 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_26 <= 1'h0;
    end else if (_T_6032) begin
      ic_tag_valid_out_1_26 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_27 <= 1'h0;
    end else if (_T_6047) begin
      ic_tag_valid_out_1_27 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_28 <= 1'h0;
    end else if (_T_6062) begin
      ic_tag_valid_out_1_28 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_29 <= 1'h0;
    end else if (_T_6077) begin
      ic_tag_valid_out_1_29 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_30 <= 1'h0;
    end else if (_T_6092) begin
      ic_tag_valid_out_1_30 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_31 <= 1'h0;
    end else if (_T_6107) begin
      ic_tag_valid_out_1_31 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_32 <= 1'h0;
    end else if (_T_6602) begin
      ic_tag_valid_out_1_32 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_33 <= 1'h0;
    end else if (_T_6617) begin
      ic_tag_valid_out_1_33 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_34 <= 1'h0;
    end else if (_T_6632) begin
      ic_tag_valid_out_1_34 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_35 <= 1'h0;
    end else if (_T_6647) begin
      ic_tag_valid_out_1_35 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_36 <= 1'h0;
    end else if (_T_6662) begin
      ic_tag_valid_out_1_36 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_37 <= 1'h0;
    end else if (_T_6677) begin
      ic_tag_valid_out_1_37 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_38 <= 1'h0;
    end else if (_T_6692) begin
      ic_tag_valid_out_1_38 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_39 <= 1'h0;
    end else if (_T_6707) begin
      ic_tag_valid_out_1_39 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_40 <= 1'h0;
    end else if (_T_6722) begin
      ic_tag_valid_out_1_40 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_41 <= 1'h0;
    end else if (_T_6737) begin
      ic_tag_valid_out_1_41 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_42 <= 1'h0;
    end else if (_T_6752) begin
      ic_tag_valid_out_1_42 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_43 <= 1'h0;
    end else if (_T_6767) begin
      ic_tag_valid_out_1_43 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_44 <= 1'h0;
    end else if (_T_6782) begin
      ic_tag_valid_out_1_44 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_45 <= 1'h0;
    end else if (_T_6797) begin
      ic_tag_valid_out_1_45 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_46 <= 1'h0;
    end else if (_T_6812) begin
      ic_tag_valid_out_1_46 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_47 <= 1'h0;
    end else if (_T_6827) begin
      ic_tag_valid_out_1_47 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_48 <= 1'h0;
    end else if (_T_6842) begin
      ic_tag_valid_out_1_48 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_49 <= 1'h0;
    end else if (_T_6857) begin
      ic_tag_valid_out_1_49 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_50 <= 1'h0;
    end else if (_T_6872) begin
      ic_tag_valid_out_1_50 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_51 <= 1'h0;
    end else if (_T_6887) begin
      ic_tag_valid_out_1_51 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_52 <= 1'h0;
    end else if (_T_6902) begin
      ic_tag_valid_out_1_52 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_53 <= 1'h0;
    end else if (_T_6917) begin
      ic_tag_valid_out_1_53 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_54 <= 1'h0;
    end else if (_T_6932) begin
      ic_tag_valid_out_1_54 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_55 <= 1'h0;
    end else if (_T_6947) begin
      ic_tag_valid_out_1_55 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_56 <= 1'h0;
    end else if (_T_6962) begin
      ic_tag_valid_out_1_56 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_57 <= 1'h0;
    end else if (_T_6977) begin
      ic_tag_valid_out_1_57 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_58 <= 1'h0;
    end else if (_T_6992) begin
      ic_tag_valid_out_1_58 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_59 <= 1'h0;
    end else if (_T_7007) begin
      ic_tag_valid_out_1_59 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_60 <= 1'h0;
    end else if (_T_7022) begin
      ic_tag_valid_out_1_60 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_61 <= 1'h0;
    end else if (_T_7037) begin
      ic_tag_valid_out_1_61 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_62 <= 1'h0;
    end else if (_T_7052) begin
      ic_tag_valid_out_1_62 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_63 <= 1'h0;
    end else if (_T_7067) begin
      ic_tag_valid_out_1_63 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_64 <= 1'h0;
    end else if (_T_7562) begin
      ic_tag_valid_out_1_64 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_65 <= 1'h0;
    end else if (_T_7577) begin
      ic_tag_valid_out_1_65 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_66 <= 1'h0;
    end else if (_T_7592) begin
      ic_tag_valid_out_1_66 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_67 <= 1'h0;
    end else if (_T_7607) begin
      ic_tag_valid_out_1_67 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_68 <= 1'h0;
    end else if (_T_7622) begin
      ic_tag_valid_out_1_68 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_69 <= 1'h0;
    end else if (_T_7637) begin
      ic_tag_valid_out_1_69 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_70 <= 1'h0;
    end else if (_T_7652) begin
      ic_tag_valid_out_1_70 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_71 <= 1'h0;
    end else if (_T_7667) begin
      ic_tag_valid_out_1_71 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_72 <= 1'h0;
    end else if (_T_7682) begin
      ic_tag_valid_out_1_72 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_73 <= 1'h0;
    end else if (_T_7697) begin
      ic_tag_valid_out_1_73 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_74 <= 1'h0;
    end else if (_T_7712) begin
      ic_tag_valid_out_1_74 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_75 <= 1'h0;
    end else if (_T_7727) begin
      ic_tag_valid_out_1_75 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_76 <= 1'h0;
    end else if (_T_7742) begin
      ic_tag_valid_out_1_76 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_77 <= 1'h0;
    end else if (_T_7757) begin
      ic_tag_valid_out_1_77 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_78 <= 1'h0;
    end else if (_T_7772) begin
      ic_tag_valid_out_1_78 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_79 <= 1'h0;
    end else if (_T_7787) begin
      ic_tag_valid_out_1_79 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_80 <= 1'h0;
    end else if (_T_7802) begin
      ic_tag_valid_out_1_80 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_81 <= 1'h0;
    end else if (_T_7817) begin
      ic_tag_valid_out_1_81 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_82 <= 1'h0;
    end else if (_T_7832) begin
      ic_tag_valid_out_1_82 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_83 <= 1'h0;
    end else if (_T_7847) begin
      ic_tag_valid_out_1_83 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_84 <= 1'h0;
    end else if (_T_7862) begin
      ic_tag_valid_out_1_84 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_85 <= 1'h0;
    end else if (_T_7877) begin
      ic_tag_valid_out_1_85 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_86 <= 1'h0;
    end else if (_T_7892) begin
      ic_tag_valid_out_1_86 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_87 <= 1'h0;
    end else if (_T_7907) begin
      ic_tag_valid_out_1_87 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_88 <= 1'h0;
    end else if (_T_7922) begin
      ic_tag_valid_out_1_88 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_89 <= 1'h0;
    end else if (_T_7937) begin
      ic_tag_valid_out_1_89 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_90 <= 1'h0;
    end else if (_T_7952) begin
      ic_tag_valid_out_1_90 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_91 <= 1'h0;
    end else if (_T_7967) begin
      ic_tag_valid_out_1_91 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_92 <= 1'h0;
    end else if (_T_7982) begin
      ic_tag_valid_out_1_92 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_93 <= 1'h0;
    end else if (_T_7997) begin
      ic_tag_valid_out_1_93 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_94 <= 1'h0;
    end else if (_T_8012) begin
      ic_tag_valid_out_1_94 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_95 <= 1'h0;
    end else if (_T_8027) begin
      ic_tag_valid_out_1_95 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_96 <= 1'h0;
    end else if (_T_8522) begin
      ic_tag_valid_out_1_96 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_97 <= 1'h0;
    end else if (_T_8537) begin
      ic_tag_valid_out_1_97 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_98 <= 1'h0;
    end else if (_T_8552) begin
      ic_tag_valid_out_1_98 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_99 <= 1'h0;
    end else if (_T_8567) begin
      ic_tag_valid_out_1_99 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_100 <= 1'h0;
    end else if (_T_8582) begin
      ic_tag_valid_out_1_100 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_101 <= 1'h0;
    end else if (_T_8597) begin
      ic_tag_valid_out_1_101 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_102 <= 1'h0;
    end else if (_T_8612) begin
      ic_tag_valid_out_1_102 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_103 <= 1'h0;
    end else if (_T_8627) begin
      ic_tag_valid_out_1_103 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_104 <= 1'h0;
    end else if (_T_8642) begin
      ic_tag_valid_out_1_104 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_105 <= 1'h0;
    end else if (_T_8657) begin
      ic_tag_valid_out_1_105 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_106 <= 1'h0;
    end else if (_T_8672) begin
      ic_tag_valid_out_1_106 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_107 <= 1'h0;
    end else if (_T_8687) begin
      ic_tag_valid_out_1_107 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_108 <= 1'h0;
    end else if (_T_8702) begin
      ic_tag_valid_out_1_108 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_109 <= 1'h0;
    end else if (_T_8717) begin
      ic_tag_valid_out_1_109 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_110 <= 1'h0;
    end else if (_T_8732) begin
      ic_tag_valid_out_1_110 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_111 <= 1'h0;
    end else if (_T_8747) begin
      ic_tag_valid_out_1_111 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_112 <= 1'h0;
    end else if (_T_8762) begin
      ic_tag_valid_out_1_112 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_113 <= 1'h0;
    end else if (_T_8777) begin
      ic_tag_valid_out_1_113 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_114 <= 1'h0;
    end else if (_T_8792) begin
      ic_tag_valid_out_1_114 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_115 <= 1'h0;
    end else if (_T_8807) begin
      ic_tag_valid_out_1_115 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_116 <= 1'h0;
    end else if (_T_8822) begin
      ic_tag_valid_out_1_116 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_117 <= 1'h0;
    end else if (_T_8837) begin
      ic_tag_valid_out_1_117 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_118 <= 1'h0;
    end else if (_T_8852) begin
      ic_tag_valid_out_1_118 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_119 <= 1'h0;
    end else if (_T_8867) begin
      ic_tag_valid_out_1_119 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_120 <= 1'h0;
    end else if (_T_8882) begin
      ic_tag_valid_out_1_120 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_121 <= 1'h0;
    end else if (_T_8897) begin
      ic_tag_valid_out_1_121 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_122 <= 1'h0;
    end else if (_T_8912) begin
      ic_tag_valid_out_1_122 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_123 <= 1'h0;
    end else if (_T_8927) begin
      ic_tag_valid_out_1_123 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_124 <= 1'h0;
    end else if (_T_8942) begin
      ic_tag_valid_out_1_124 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_125 <= 1'h0;
    end else if (_T_8957) begin
      ic_tag_valid_out_1_125 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_126 <= 1'h0;
    end else if (_T_8972) begin
      ic_tag_valid_out_1_126 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_127 <= 1'h0;
    end else if (_T_8987) begin
      ic_tag_valid_out_1_127 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_0 <= 1'h0;
    end else if (_T_5162) begin
      ic_tag_valid_out_0_0 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_1 <= 1'h0;
    end else if (_T_5177) begin
      ic_tag_valid_out_0_1 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_2 <= 1'h0;
    end else if (_T_5192) begin
      ic_tag_valid_out_0_2 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_3 <= 1'h0;
    end else if (_T_5207) begin
      ic_tag_valid_out_0_3 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_4 <= 1'h0;
    end else if (_T_5222) begin
      ic_tag_valid_out_0_4 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_5 <= 1'h0;
    end else if (_T_5237) begin
      ic_tag_valid_out_0_5 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_6 <= 1'h0;
    end else if (_T_5252) begin
      ic_tag_valid_out_0_6 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_7 <= 1'h0;
    end else if (_T_5267) begin
      ic_tag_valid_out_0_7 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_8 <= 1'h0;
    end else if (_T_5282) begin
      ic_tag_valid_out_0_8 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_9 <= 1'h0;
    end else if (_T_5297) begin
      ic_tag_valid_out_0_9 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_10 <= 1'h0;
    end else if (_T_5312) begin
      ic_tag_valid_out_0_10 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_11 <= 1'h0;
    end else if (_T_5327) begin
      ic_tag_valid_out_0_11 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_12 <= 1'h0;
    end else if (_T_5342) begin
      ic_tag_valid_out_0_12 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_13 <= 1'h0;
    end else if (_T_5357) begin
      ic_tag_valid_out_0_13 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_14 <= 1'h0;
    end else if (_T_5372) begin
      ic_tag_valid_out_0_14 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_15 <= 1'h0;
    end else if (_T_5387) begin
      ic_tag_valid_out_0_15 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_16 <= 1'h0;
    end else if (_T_5402) begin
      ic_tag_valid_out_0_16 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_17 <= 1'h0;
    end else if (_T_5417) begin
      ic_tag_valid_out_0_17 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_18 <= 1'h0;
    end else if (_T_5432) begin
      ic_tag_valid_out_0_18 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_19 <= 1'h0;
    end else if (_T_5447) begin
      ic_tag_valid_out_0_19 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_20 <= 1'h0;
    end else if (_T_5462) begin
      ic_tag_valid_out_0_20 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_21 <= 1'h0;
    end else if (_T_5477) begin
      ic_tag_valid_out_0_21 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_22 <= 1'h0;
    end else if (_T_5492) begin
      ic_tag_valid_out_0_22 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_23 <= 1'h0;
    end else if (_T_5507) begin
      ic_tag_valid_out_0_23 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_24 <= 1'h0;
    end else if (_T_5522) begin
      ic_tag_valid_out_0_24 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_25 <= 1'h0;
    end else if (_T_5537) begin
      ic_tag_valid_out_0_25 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_26 <= 1'h0;
    end else if (_T_5552) begin
      ic_tag_valid_out_0_26 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_27 <= 1'h0;
    end else if (_T_5567) begin
      ic_tag_valid_out_0_27 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_28 <= 1'h0;
    end else if (_T_5582) begin
      ic_tag_valid_out_0_28 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_29 <= 1'h0;
    end else if (_T_5597) begin
      ic_tag_valid_out_0_29 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_30 <= 1'h0;
    end else if (_T_5612) begin
      ic_tag_valid_out_0_30 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_31 <= 1'h0;
    end else if (_T_5627) begin
      ic_tag_valid_out_0_31 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_32 <= 1'h0;
    end else if (_T_6122) begin
      ic_tag_valid_out_0_32 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_33 <= 1'h0;
    end else if (_T_6137) begin
      ic_tag_valid_out_0_33 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_34 <= 1'h0;
    end else if (_T_6152) begin
      ic_tag_valid_out_0_34 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_35 <= 1'h0;
    end else if (_T_6167) begin
      ic_tag_valid_out_0_35 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_36 <= 1'h0;
    end else if (_T_6182) begin
      ic_tag_valid_out_0_36 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_37 <= 1'h0;
    end else if (_T_6197) begin
      ic_tag_valid_out_0_37 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_38 <= 1'h0;
    end else if (_T_6212) begin
      ic_tag_valid_out_0_38 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_39 <= 1'h0;
    end else if (_T_6227) begin
      ic_tag_valid_out_0_39 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_40 <= 1'h0;
    end else if (_T_6242) begin
      ic_tag_valid_out_0_40 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_41 <= 1'h0;
    end else if (_T_6257) begin
      ic_tag_valid_out_0_41 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_42 <= 1'h0;
    end else if (_T_6272) begin
      ic_tag_valid_out_0_42 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_43 <= 1'h0;
    end else if (_T_6287) begin
      ic_tag_valid_out_0_43 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_44 <= 1'h0;
    end else if (_T_6302) begin
      ic_tag_valid_out_0_44 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_45 <= 1'h0;
    end else if (_T_6317) begin
      ic_tag_valid_out_0_45 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_46 <= 1'h0;
    end else if (_T_6332) begin
      ic_tag_valid_out_0_46 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_47 <= 1'h0;
    end else if (_T_6347) begin
      ic_tag_valid_out_0_47 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_48 <= 1'h0;
    end else if (_T_6362) begin
      ic_tag_valid_out_0_48 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_49 <= 1'h0;
    end else if (_T_6377) begin
      ic_tag_valid_out_0_49 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_50 <= 1'h0;
    end else if (_T_6392) begin
      ic_tag_valid_out_0_50 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_51 <= 1'h0;
    end else if (_T_6407) begin
      ic_tag_valid_out_0_51 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_52 <= 1'h0;
    end else if (_T_6422) begin
      ic_tag_valid_out_0_52 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_53 <= 1'h0;
    end else if (_T_6437) begin
      ic_tag_valid_out_0_53 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_54 <= 1'h0;
    end else if (_T_6452) begin
      ic_tag_valid_out_0_54 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_55 <= 1'h0;
    end else if (_T_6467) begin
      ic_tag_valid_out_0_55 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_56 <= 1'h0;
    end else if (_T_6482) begin
      ic_tag_valid_out_0_56 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_57 <= 1'h0;
    end else if (_T_6497) begin
      ic_tag_valid_out_0_57 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_58 <= 1'h0;
    end else if (_T_6512) begin
      ic_tag_valid_out_0_58 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_59 <= 1'h0;
    end else if (_T_6527) begin
      ic_tag_valid_out_0_59 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_60 <= 1'h0;
    end else if (_T_6542) begin
      ic_tag_valid_out_0_60 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_61 <= 1'h0;
    end else if (_T_6557) begin
      ic_tag_valid_out_0_61 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_62 <= 1'h0;
    end else if (_T_6572) begin
      ic_tag_valid_out_0_62 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_63 <= 1'h0;
    end else if (_T_6587) begin
      ic_tag_valid_out_0_63 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_64 <= 1'h0;
    end else if (_T_7082) begin
      ic_tag_valid_out_0_64 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_65 <= 1'h0;
    end else if (_T_7097) begin
      ic_tag_valid_out_0_65 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_66 <= 1'h0;
    end else if (_T_7112) begin
      ic_tag_valid_out_0_66 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_67 <= 1'h0;
    end else if (_T_7127) begin
      ic_tag_valid_out_0_67 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_68 <= 1'h0;
    end else if (_T_7142) begin
      ic_tag_valid_out_0_68 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_69 <= 1'h0;
    end else if (_T_7157) begin
      ic_tag_valid_out_0_69 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_70 <= 1'h0;
    end else if (_T_7172) begin
      ic_tag_valid_out_0_70 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_71 <= 1'h0;
    end else if (_T_7187) begin
      ic_tag_valid_out_0_71 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_72 <= 1'h0;
    end else if (_T_7202) begin
      ic_tag_valid_out_0_72 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_73 <= 1'h0;
    end else if (_T_7217) begin
      ic_tag_valid_out_0_73 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_74 <= 1'h0;
    end else if (_T_7232) begin
      ic_tag_valid_out_0_74 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_75 <= 1'h0;
    end else if (_T_7247) begin
      ic_tag_valid_out_0_75 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_76 <= 1'h0;
    end else if (_T_7262) begin
      ic_tag_valid_out_0_76 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_77 <= 1'h0;
    end else if (_T_7277) begin
      ic_tag_valid_out_0_77 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_78 <= 1'h0;
    end else if (_T_7292) begin
      ic_tag_valid_out_0_78 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_79 <= 1'h0;
    end else if (_T_7307) begin
      ic_tag_valid_out_0_79 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_80 <= 1'h0;
    end else if (_T_7322) begin
      ic_tag_valid_out_0_80 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_81 <= 1'h0;
    end else if (_T_7337) begin
      ic_tag_valid_out_0_81 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_82 <= 1'h0;
    end else if (_T_7352) begin
      ic_tag_valid_out_0_82 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_83 <= 1'h0;
    end else if (_T_7367) begin
      ic_tag_valid_out_0_83 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_84 <= 1'h0;
    end else if (_T_7382) begin
      ic_tag_valid_out_0_84 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_85 <= 1'h0;
    end else if (_T_7397) begin
      ic_tag_valid_out_0_85 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_86 <= 1'h0;
    end else if (_T_7412) begin
      ic_tag_valid_out_0_86 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_87 <= 1'h0;
    end else if (_T_7427) begin
      ic_tag_valid_out_0_87 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_88 <= 1'h0;
    end else if (_T_7442) begin
      ic_tag_valid_out_0_88 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_89 <= 1'h0;
    end else if (_T_7457) begin
      ic_tag_valid_out_0_89 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_90 <= 1'h0;
    end else if (_T_7472) begin
      ic_tag_valid_out_0_90 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_91 <= 1'h0;
    end else if (_T_7487) begin
      ic_tag_valid_out_0_91 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_92 <= 1'h0;
    end else if (_T_7502) begin
      ic_tag_valid_out_0_92 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_93 <= 1'h0;
    end else if (_T_7517) begin
      ic_tag_valid_out_0_93 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_94 <= 1'h0;
    end else if (_T_7532) begin
      ic_tag_valid_out_0_94 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_95 <= 1'h0;
    end else if (_T_7547) begin
      ic_tag_valid_out_0_95 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_96 <= 1'h0;
    end else if (_T_8042) begin
      ic_tag_valid_out_0_96 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_97 <= 1'h0;
    end else if (_T_8057) begin
      ic_tag_valid_out_0_97 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_98 <= 1'h0;
    end else if (_T_8072) begin
      ic_tag_valid_out_0_98 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_99 <= 1'h0;
    end else if (_T_8087) begin
      ic_tag_valid_out_0_99 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_100 <= 1'h0;
    end else if (_T_8102) begin
      ic_tag_valid_out_0_100 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_101 <= 1'h0;
    end else if (_T_8117) begin
      ic_tag_valid_out_0_101 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_102 <= 1'h0;
    end else if (_T_8132) begin
      ic_tag_valid_out_0_102 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_103 <= 1'h0;
    end else if (_T_8147) begin
      ic_tag_valid_out_0_103 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_104 <= 1'h0;
    end else if (_T_8162) begin
      ic_tag_valid_out_0_104 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_105 <= 1'h0;
    end else if (_T_8177) begin
      ic_tag_valid_out_0_105 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_106 <= 1'h0;
    end else if (_T_8192) begin
      ic_tag_valid_out_0_106 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_107 <= 1'h0;
    end else if (_T_8207) begin
      ic_tag_valid_out_0_107 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_108 <= 1'h0;
    end else if (_T_8222) begin
      ic_tag_valid_out_0_108 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_109 <= 1'h0;
    end else if (_T_8237) begin
      ic_tag_valid_out_0_109 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_110 <= 1'h0;
    end else if (_T_8252) begin
      ic_tag_valid_out_0_110 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_111 <= 1'h0;
    end else if (_T_8267) begin
      ic_tag_valid_out_0_111 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_112 <= 1'h0;
    end else if (_T_8282) begin
      ic_tag_valid_out_0_112 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_113 <= 1'h0;
    end else if (_T_8297) begin
      ic_tag_valid_out_0_113 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_114 <= 1'h0;
    end else if (_T_8312) begin
      ic_tag_valid_out_0_114 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_115 <= 1'h0;
    end else if (_T_8327) begin
      ic_tag_valid_out_0_115 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_116 <= 1'h0;
    end else if (_T_8342) begin
      ic_tag_valid_out_0_116 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_117 <= 1'h0;
    end else if (_T_8357) begin
      ic_tag_valid_out_0_117 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_118 <= 1'h0;
    end else if (_T_8372) begin
      ic_tag_valid_out_0_118 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_119 <= 1'h0;
    end else if (_T_8387) begin
      ic_tag_valid_out_0_119 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_120 <= 1'h0;
    end else if (_T_8402) begin
      ic_tag_valid_out_0_120 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_121 <= 1'h0;
    end else if (_T_8417) begin
      ic_tag_valid_out_0_121 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_122 <= 1'h0;
    end else if (_T_8432) begin
      ic_tag_valid_out_0_122 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_123 <= 1'h0;
    end else if (_T_8447) begin
      ic_tag_valid_out_0_123 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_124 <= 1'h0;
    end else if (_T_8462) begin
      ic_tag_valid_out_0_124 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_125 <= 1'h0;
    end else if (_T_8477) begin
      ic_tag_valid_out_0_125 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_126 <= 1'h0;
    end else if (_T_8492) begin
      ic_tag_valid_out_0_126 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_127 <= 1'h0;
    end else if (_T_8507) begin
      ic_tag_valid_out_0_127 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_1_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_debug_way_ff <= 2'h0;
    end else begin
      ic_debug_way_ff <= io_ic_debug_way;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      ic_debug_rd_en_ff <= 1'h0;
    end else begin
      ic_debug_rd_en_ff <= io_ic_debug_rd_en;
    end
  end
  always @(posedge rvclkhdr_io_l1clk or posedge reset) begin
    if (reset) begin
      _T_1212 <= 71'h0;
    end else if (ic_debug_ict_array_sel_ff) begin
      _T_1212 <= _T_1211;
    end else begin
      _T_1212 <= io_ic_debug_rd_data;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      ifc_region_acc_fault_memory_f <= 1'h0;
    end else begin
      ifc_region_acc_fault_memory_f <= _T_9885 & io_ifc_fetch_req_bf;
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      perr_ic_index_ff <= 7'h0;
    end else if (perr_sb_write_status) begin
      perr_ic_index_ff <= ifu_ic_rw_int_addr_ff;
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      dma_sb_err_state_ff <= 1'h0;
    end else begin
      dma_sb_err_state_ff <= perr_state == 3'h4;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      bus_cmd_req_hold <= 1'h0;
    end else begin
      bus_cmd_req_hold <= _T_2591 & _T_2623;
    end
  end
  always @(posedge rvclkhdr_69_io_l1clk or posedge reset) begin
    if (reset) begin
      ifu_bus_cmd_valid <= 1'h0;
    end else begin
      ifu_bus_cmd_valid <= _T_2592 & _T_2623;
    end
  end
  always @(posedge rvclkhdr_68_io_l1clk or posedge reset) begin
    if (reset) begin
      ifu_bus_arvalid_ff <= 1'h0;
    end else begin
      ifu_bus_arvalid_ff <= io_ifu_axi_ar_valid;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      ifc_dma_access_ok_prev <= 1'h0;
    end else begin
      ifc_dma_access_ok_prev <= _T_2699 & _T_2700;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      iccm_ecc_corr_data_ff <= 39'h0;
    end else if (iccm_ecc_write_status) begin
      iccm_ecc_corr_data_ff <= _T_3932;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      dma_mem_addr_ff <= 2'h0;
    end else begin
      dma_mem_addr_ff <= io_dma_mem_ctl_dma_mem_addr[3:2];
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      dma_mem_tag_ff <= 3'h0;
    end else begin
      dma_mem_tag_ff <= io_dma_mem_ctl_dma_mem_tag;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      iccm_dma_rtag_temp <= 3'h0;
    end else begin
      iccm_dma_rtag_temp <= dma_mem_tag_ff;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      iccm_dma_rvalid_temp <= 1'h0;
    end else begin
      iccm_dma_rvalid_temp <= iccm_dma_rvalid_in;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      iccm_dma_ecc_error <= 1'h0;
    end else begin
      iccm_dma_ecc_error <= |iccm_double_ecc_error;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      iccm_dma_rdata_temp <= 64'h0;
    end else if (iccm_dma_ecc_error_in) begin
      iccm_dma_rdata_temp <= _T_3104;
    end else begin
      iccm_dma_rdata_temp <= _T_3105;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      iccm_ecc_corr_index_ff <= 14'h0;
    end else if (iccm_ecc_write_status) begin
      if (iccm_single_ecc_error[0]) begin
        iccm_ecc_corr_index_ff <= iccm_rw_addr_f;
      end else begin
        iccm_ecc_corr_index_ff <= _T_3928;
      end
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      iccm_rd_ecc_single_err_ff <= 1'h0;
    end else begin
      iccm_rd_ecc_single_err_ff <= _T_3923 & _T_319;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      iccm_rw_addr_f <= 14'h0;
    end else begin
      iccm_rw_addr_f <= io_iccm_rw_addr[14:1];
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      ifu_status_wr_addr_ff <= 7'h0;
    end else if (_T_3997) begin
      ifu_status_wr_addr_ff <= io_ic_debug_addr[9:3];
    end else begin
      ifu_status_wr_addr_ff <= ifu_status_wr_addr[11:5];
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      way_status_wr_en_ff <= 1'h0;
    end else begin
      way_status_wr_en_ff <= ic_act_hit_f | _T_4000;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      way_status_new_ff <= 1'h0;
    end else if (_T_4000) begin
      way_status_new_ff <= io_ic_debug_wr_data[4];
    end else begin
      way_status_new_ff <= way_status_hit_new;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      ifu_tag_wren_ff <= 2'h0;
    end else begin
      ifu_tag_wren_ff <= ifu_tag_wren | ic_debug_tag_wr_en;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      ic_valid_ff <= 1'h0;
    end else if (_T_4000) begin
      ic_valid_ff <= io_ic_debug_wr_data[0];
    end else begin
      ic_valid_ff <= ic_valid;
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      _T_9799 <= 1'h0;
    end else begin
      _T_9799 <= _T_232 & _T_209;
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      _T_9800 <= 1'h0;
    end else begin
      _T_9800 <= _T_225 & _T_247;
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      _T_9801 <= 1'h0;
    end else begin
      _T_9801 <= ic_byp_hit_f & ifu_byp_data_err_new;
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      _T_9805 <= 1'h0;
    end else begin
      _T_9805 <= ifu_bus_arvalid_ff & miss_pending;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      _T_9826 <= 1'h0;
    end else begin
      _T_9826 <= ic_debug_rd_en_ff;
    end
  end
endmodule
module ifu_bp_ctl(
  input         clock,
  input         reset,
  input         io_active_clk,
  input         io_ic_hit_f,
  input         io_exu_flush_final,
  input  [30:0] io_ifc_fetch_addr_f,
  input         io_ifc_fetch_req_f,
  input         io_dec_bp_dec_tlu_br0_r_pkt_valid,
  input  [1:0]  io_dec_bp_dec_tlu_br0_r_pkt_bits_hist,
  input         io_dec_bp_dec_tlu_br0_r_pkt_bits_br_error,
  input         io_dec_bp_dec_tlu_br0_r_pkt_bits_br_start_error,
  input         io_dec_bp_dec_tlu_br0_r_pkt_bits_way,
  input         io_dec_bp_dec_tlu_br0_r_pkt_bits_middle,
  input         io_dec_bp_dec_tlu_flush_leak_one_wb,
  input         io_dec_bp_dec_tlu_bpred_disable,
  input         io_dec_tlu_flush_lower_wb,
  input  [7:0]  io_exu_bp_exu_i0_br_index_r,
  input  [7:0]  io_exu_bp_exu_i0_br_fghr_r,
  input         io_exu_bp_exu_mp_pkt_bits_misp,
  input         io_exu_bp_exu_mp_pkt_bits_ataken,
  input         io_exu_bp_exu_mp_pkt_bits_boffset,
  input         io_exu_bp_exu_mp_pkt_bits_pc4,
  input  [1:0]  io_exu_bp_exu_mp_pkt_bits_hist,
  input  [11:0] io_exu_bp_exu_mp_pkt_bits_toffset,
  input         io_exu_bp_exu_mp_pkt_bits_pcall,
  input         io_exu_bp_exu_mp_pkt_bits_pret,
  input         io_exu_bp_exu_mp_pkt_bits_pja,
  input         io_exu_bp_exu_mp_pkt_bits_way,
  input  [7:0]  io_exu_bp_exu_mp_eghr,
  input  [7:0]  io_exu_bp_exu_mp_fghr,
  input  [7:0]  io_exu_bp_exu_mp_index,
  input  [4:0]  io_exu_bp_exu_mp_btag,
  output        io_ifu_bp_hit_taken_f,
  output [30:0] io_ifu_bp_btb_target_f,
  output        io_ifu_bp_inst_mask_f,
  output [7:0]  io_ifu_bp_fghr_f,
  output [1:0]  io_ifu_bp_way_f,
  output [1:0]  io_ifu_bp_ret_f,
  output [1:0]  io_ifu_bp_hist1_f,
  output [1:0]  io_ifu_bp_hist0_f,
  output [1:0]  io_ifu_bp_pc4_f,
  output [1:0]  io_ifu_bp_valid_f,
  output [11:0] io_ifu_bp_poffset_f,
  input         io_scan_mode
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_576;
  reg [31:0] _RAND_577;
  reg [31:0] _RAND_578;
  reg [31:0] _RAND_579;
  reg [31:0] _RAND_580;
  reg [31:0] _RAND_581;
  reg [31:0] _RAND_582;
  reg [31:0] _RAND_583;
  reg [31:0] _RAND_584;
  reg [31:0] _RAND_585;
  reg [31:0] _RAND_586;
  reg [31:0] _RAND_587;
  reg [31:0] _RAND_588;
  reg [31:0] _RAND_589;
  reg [31:0] _RAND_590;
  reg [31:0] _RAND_591;
  reg [31:0] _RAND_592;
  reg [31:0] _RAND_593;
  reg [31:0] _RAND_594;
  reg [31:0] _RAND_595;
  reg [31:0] _RAND_596;
  reg [31:0] _RAND_597;
  reg [31:0] _RAND_598;
  reg [31:0] _RAND_599;
  reg [31:0] _RAND_600;
  reg [31:0] _RAND_601;
  reg [31:0] _RAND_602;
  reg [31:0] _RAND_603;
  reg [31:0] _RAND_604;
  reg [31:0] _RAND_605;
  reg [31:0] _RAND_606;
  reg [31:0] _RAND_607;
  reg [31:0] _RAND_608;
  reg [31:0] _RAND_609;
  reg [31:0] _RAND_610;
  reg [31:0] _RAND_611;
  reg [31:0] _RAND_612;
  reg [31:0] _RAND_613;
  reg [31:0] _RAND_614;
  reg [31:0] _RAND_615;
  reg [31:0] _RAND_616;
  reg [31:0] _RAND_617;
  reg [31:0] _RAND_618;
  reg [31:0] _RAND_619;
  reg [31:0] _RAND_620;
  reg [31:0] _RAND_621;
  reg [31:0] _RAND_622;
  reg [31:0] _RAND_623;
  reg [31:0] _RAND_624;
  reg [31:0] _RAND_625;
  reg [31:0] _RAND_626;
  reg [31:0] _RAND_627;
  reg [31:0] _RAND_628;
  reg [31:0] _RAND_629;
  reg [31:0] _RAND_630;
  reg [31:0] _RAND_631;
  reg [31:0] _RAND_632;
  reg [31:0] _RAND_633;
  reg [31:0] _RAND_634;
  reg [31:0] _RAND_635;
  reg [31:0] _RAND_636;
  reg [31:0] _RAND_637;
  reg [31:0] _RAND_638;
  reg [31:0] _RAND_639;
  reg [31:0] _RAND_640;
  reg [31:0] _RAND_641;
  reg [31:0] _RAND_642;
  reg [31:0] _RAND_643;
  reg [31:0] _RAND_644;
  reg [31:0] _RAND_645;
  reg [31:0] _RAND_646;
  reg [31:0] _RAND_647;
  reg [31:0] _RAND_648;
  reg [31:0] _RAND_649;
  reg [31:0] _RAND_650;
  reg [31:0] _RAND_651;
  reg [31:0] _RAND_652;
  reg [31:0] _RAND_653;
  reg [31:0] _RAND_654;
  reg [31:0] _RAND_655;
  reg [31:0] _RAND_656;
  reg [31:0] _RAND_657;
  reg [31:0] _RAND_658;
  reg [31:0] _RAND_659;
  reg [31:0] _RAND_660;
  reg [31:0] _RAND_661;
  reg [31:0] _RAND_662;
  reg [31:0] _RAND_663;
  reg [31:0] _RAND_664;
  reg [31:0] _RAND_665;
  reg [31:0] _RAND_666;
  reg [31:0] _RAND_667;
  reg [31:0] _RAND_668;
  reg [31:0] _RAND_669;
  reg [31:0] _RAND_670;
  reg [31:0] _RAND_671;
  reg [31:0] _RAND_672;
  reg [31:0] _RAND_673;
  reg [31:0] _RAND_674;
  reg [31:0] _RAND_675;
  reg [31:0] _RAND_676;
  reg [31:0] _RAND_677;
  reg [31:0] _RAND_678;
  reg [31:0] _RAND_679;
  reg [31:0] _RAND_680;
  reg [31:0] _RAND_681;
  reg [31:0] _RAND_682;
  reg [31:0] _RAND_683;
  reg [31:0] _RAND_684;
  reg [31:0] _RAND_685;
  reg [31:0] _RAND_686;
  reg [31:0] _RAND_687;
  reg [31:0] _RAND_688;
  reg [31:0] _RAND_689;
  reg [31:0] _RAND_690;
  reg [31:0] _RAND_691;
  reg [31:0] _RAND_692;
  reg [31:0] _RAND_693;
  reg [31:0] _RAND_694;
  reg [31:0] _RAND_695;
  reg [31:0] _RAND_696;
  reg [31:0] _RAND_697;
  reg [31:0] _RAND_698;
  reg [31:0] _RAND_699;
  reg [31:0] _RAND_700;
  reg [31:0] _RAND_701;
  reg [31:0] _RAND_702;
  reg [31:0] _RAND_703;
  reg [31:0] _RAND_704;
  reg [31:0] _RAND_705;
  reg [31:0] _RAND_706;
  reg [31:0] _RAND_707;
  reg [31:0] _RAND_708;
  reg [31:0] _RAND_709;
  reg [31:0] _RAND_710;
  reg [31:0] _RAND_711;
  reg [31:0] _RAND_712;
  reg [31:0] _RAND_713;
  reg [31:0] _RAND_714;
  reg [31:0] _RAND_715;
  reg [31:0] _RAND_716;
  reg [31:0] _RAND_717;
  reg [31:0] _RAND_718;
  reg [31:0] _RAND_719;
  reg [31:0] _RAND_720;
  reg [31:0] _RAND_721;
  reg [31:0] _RAND_722;
  reg [31:0] _RAND_723;
  reg [31:0] _RAND_724;
  reg [31:0] _RAND_725;
  reg [31:0] _RAND_726;
  reg [31:0] _RAND_727;
  reg [31:0] _RAND_728;
  reg [31:0] _RAND_729;
  reg [31:0] _RAND_730;
  reg [31:0] _RAND_731;
  reg [31:0] _RAND_732;
  reg [31:0] _RAND_733;
  reg [31:0] _RAND_734;
  reg [31:0] _RAND_735;
  reg [31:0] _RAND_736;
  reg [31:0] _RAND_737;
  reg [31:0] _RAND_738;
  reg [31:0] _RAND_739;
  reg [31:0] _RAND_740;
  reg [31:0] _RAND_741;
  reg [31:0] _RAND_742;
  reg [31:0] _RAND_743;
  reg [31:0] _RAND_744;
  reg [31:0] _RAND_745;
  reg [31:0] _RAND_746;
  reg [31:0] _RAND_747;
  reg [31:0] _RAND_748;
  reg [31:0] _RAND_749;
  reg [31:0] _RAND_750;
  reg [31:0] _RAND_751;
  reg [31:0] _RAND_752;
  reg [31:0] _RAND_753;
  reg [31:0] _RAND_754;
  reg [31:0] _RAND_755;
  reg [31:0] _RAND_756;
  reg [31:0] _RAND_757;
  reg [31:0] _RAND_758;
  reg [31:0] _RAND_759;
  reg [31:0] _RAND_760;
  reg [31:0] _RAND_761;
  reg [31:0] _RAND_762;
  reg [31:0] _RAND_763;
  reg [31:0] _RAND_764;
  reg [31:0] _RAND_765;
  reg [31:0] _RAND_766;
  reg [31:0] _RAND_767;
  reg [31:0] _RAND_768;
  reg [31:0] _RAND_769;
  reg [31:0] _RAND_770;
  reg [31:0] _RAND_771;
  reg [31:0] _RAND_772;
  reg [31:0] _RAND_773;
  reg [31:0] _RAND_774;
  reg [31:0] _RAND_775;
  reg [31:0] _RAND_776;
  reg [31:0] _RAND_777;
  reg [31:0] _RAND_778;
  reg [31:0] _RAND_779;
  reg [31:0] _RAND_780;
  reg [31:0] _RAND_781;
  reg [31:0] _RAND_782;
  reg [31:0] _RAND_783;
  reg [31:0] _RAND_784;
  reg [31:0] _RAND_785;
  reg [31:0] _RAND_786;
  reg [31:0] _RAND_787;
  reg [31:0] _RAND_788;
  reg [31:0] _RAND_789;
  reg [31:0] _RAND_790;
  reg [31:0] _RAND_791;
  reg [31:0] _RAND_792;
  reg [31:0] _RAND_793;
  reg [31:0] _RAND_794;
  reg [31:0] _RAND_795;
  reg [31:0] _RAND_796;
  reg [31:0] _RAND_797;
  reg [31:0] _RAND_798;
  reg [31:0] _RAND_799;
  reg [31:0] _RAND_800;
  reg [31:0] _RAND_801;
  reg [31:0] _RAND_802;
  reg [31:0] _RAND_803;
  reg [31:0] _RAND_804;
  reg [31:0] _RAND_805;
  reg [31:0] _RAND_806;
  reg [31:0] _RAND_807;
  reg [31:0] _RAND_808;
  reg [31:0] _RAND_809;
  reg [31:0] _RAND_810;
  reg [31:0] _RAND_811;
  reg [31:0] _RAND_812;
  reg [31:0] _RAND_813;
  reg [31:0] _RAND_814;
  reg [31:0] _RAND_815;
  reg [31:0] _RAND_816;
  reg [31:0] _RAND_817;
  reg [31:0] _RAND_818;
  reg [31:0] _RAND_819;
  reg [31:0] _RAND_820;
  reg [31:0] _RAND_821;
  reg [31:0] _RAND_822;
  reg [31:0] _RAND_823;
  reg [31:0] _RAND_824;
  reg [31:0] _RAND_825;
  reg [31:0] _RAND_826;
  reg [31:0] _RAND_827;
  reg [31:0] _RAND_828;
  reg [31:0] _RAND_829;
  reg [31:0] _RAND_830;
  reg [31:0] _RAND_831;
  reg [31:0] _RAND_832;
  reg [31:0] _RAND_833;
  reg [31:0] _RAND_834;
  reg [31:0] _RAND_835;
  reg [31:0] _RAND_836;
  reg [31:0] _RAND_837;
  reg [31:0] _RAND_838;
  reg [31:0] _RAND_839;
  reg [31:0] _RAND_840;
  reg [31:0] _RAND_841;
  reg [31:0] _RAND_842;
  reg [31:0] _RAND_843;
  reg [31:0] _RAND_844;
  reg [31:0] _RAND_845;
  reg [31:0] _RAND_846;
  reg [31:0] _RAND_847;
  reg [31:0] _RAND_848;
  reg [31:0] _RAND_849;
  reg [31:0] _RAND_850;
  reg [31:0] _RAND_851;
  reg [31:0] _RAND_852;
  reg [31:0] _RAND_853;
  reg [31:0] _RAND_854;
  reg [31:0] _RAND_855;
  reg [31:0] _RAND_856;
  reg [31:0] _RAND_857;
  reg [31:0] _RAND_858;
  reg [31:0] _RAND_859;
  reg [31:0] _RAND_860;
  reg [31:0] _RAND_861;
  reg [31:0] _RAND_862;
  reg [31:0] _RAND_863;
  reg [31:0] _RAND_864;
  reg [31:0] _RAND_865;
  reg [31:0] _RAND_866;
  reg [31:0] _RAND_867;
  reg [31:0] _RAND_868;
  reg [31:0] _RAND_869;
  reg [31:0] _RAND_870;
  reg [31:0] _RAND_871;
  reg [31:0] _RAND_872;
  reg [31:0] _RAND_873;
  reg [31:0] _RAND_874;
  reg [31:0] _RAND_875;
  reg [31:0] _RAND_876;
  reg [31:0] _RAND_877;
  reg [31:0] _RAND_878;
  reg [31:0] _RAND_879;
  reg [31:0] _RAND_880;
  reg [31:0] _RAND_881;
  reg [31:0] _RAND_882;
  reg [31:0] _RAND_883;
  reg [31:0] _RAND_884;
  reg [31:0] _RAND_885;
  reg [31:0] _RAND_886;
  reg [31:0] _RAND_887;
  reg [31:0] _RAND_888;
  reg [31:0] _RAND_889;
  reg [31:0] _RAND_890;
  reg [31:0] _RAND_891;
  reg [31:0] _RAND_892;
  reg [31:0] _RAND_893;
  reg [31:0] _RAND_894;
  reg [31:0] _RAND_895;
  reg [31:0] _RAND_896;
  reg [31:0] _RAND_897;
  reg [31:0] _RAND_898;
  reg [31:0] _RAND_899;
  reg [31:0] _RAND_900;
  reg [31:0] _RAND_901;
  reg [31:0] _RAND_902;
  reg [31:0] _RAND_903;
  reg [31:0] _RAND_904;
  reg [31:0] _RAND_905;
  reg [31:0] _RAND_906;
  reg [31:0] _RAND_907;
  reg [31:0] _RAND_908;
  reg [31:0] _RAND_909;
  reg [31:0] _RAND_910;
  reg [31:0] _RAND_911;
  reg [31:0] _RAND_912;
  reg [31:0] _RAND_913;
  reg [31:0] _RAND_914;
  reg [31:0] _RAND_915;
  reg [31:0] _RAND_916;
  reg [31:0] _RAND_917;
  reg [31:0] _RAND_918;
  reg [31:0] _RAND_919;
  reg [31:0] _RAND_920;
  reg [31:0] _RAND_921;
  reg [31:0] _RAND_922;
  reg [31:0] _RAND_923;
  reg [31:0] _RAND_924;
  reg [31:0] _RAND_925;
  reg [31:0] _RAND_926;
  reg [31:0] _RAND_927;
  reg [31:0] _RAND_928;
  reg [31:0] _RAND_929;
  reg [31:0] _RAND_930;
  reg [31:0] _RAND_931;
  reg [31:0] _RAND_932;
  reg [31:0] _RAND_933;
  reg [31:0] _RAND_934;
  reg [31:0] _RAND_935;
  reg [31:0] _RAND_936;
  reg [31:0] _RAND_937;
  reg [31:0] _RAND_938;
  reg [31:0] _RAND_939;
  reg [31:0] _RAND_940;
  reg [31:0] _RAND_941;
  reg [31:0] _RAND_942;
  reg [31:0] _RAND_943;
  reg [31:0] _RAND_944;
  reg [31:0] _RAND_945;
  reg [31:0] _RAND_946;
  reg [31:0] _RAND_947;
  reg [31:0] _RAND_948;
  reg [31:0] _RAND_949;
  reg [31:0] _RAND_950;
  reg [31:0] _RAND_951;
  reg [31:0] _RAND_952;
  reg [31:0] _RAND_953;
  reg [31:0] _RAND_954;
  reg [31:0] _RAND_955;
  reg [31:0] _RAND_956;
  reg [31:0] _RAND_957;
  reg [31:0] _RAND_958;
  reg [31:0] _RAND_959;
  reg [31:0] _RAND_960;
  reg [31:0] _RAND_961;
  reg [31:0] _RAND_962;
  reg [31:0] _RAND_963;
  reg [31:0] _RAND_964;
  reg [31:0] _RAND_965;
  reg [31:0] _RAND_966;
  reg [31:0] _RAND_967;
  reg [31:0] _RAND_968;
  reg [31:0] _RAND_969;
  reg [31:0] _RAND_970;
  reg [31:0] _RAND_971;
  reg [31:0] _RAND_972;
  reg [31:0] _RAND_973;
  reg [31:0] _RAND_974;
  reg [31:0] _RAND_975;
  reg [31:0] _RAND_976;
  reg [31:0] _RAND_977;
  reg [31:0] _RAND_978;
  reg [31:0] _RAND_979;
  reg [31:0] _RAND_980;
  reg [31:0] _RAND_981;
  reg [31:0] _RAND_982;
  reg [31:0] _RAND_983;
  reg [31:0] _RAND_984;
  reg [31:0] _RAND_985;
  reg [31:0] _RAND_986;
  reg [31:0] _RAND_987;
  reg [31:0] _RAND_988;
  reg [31:0] _RAND_989;
  reg [31:0] _RAND_990;
  reg [31:0] _RAND_991;
  reg [31:0] _RAND_992;
  reg [31:0] _RAND_993;
  reg [31:0] _RAND_994;
  reg [31:0] _RAND_995;
  reg [31:0] _RAND_996;
  reg [31:0] _RAND_997;
  reg [31:0] _RAND_998;
  reg [31:0] _RAND_999;
  reg [31:0] _RAND_1000;
  reg [31:0] _RAND_1001;
  reg [31:0] _RAND_1002;
  reg [31:0] _RAND_1003;
  reg [31:0] _RAND_1004;
  reg [31:0] _RAND_1005;
  reg [31:0] _RAND_1006;
  reg [31:0] _RAND_1007;
  reg [31:0] _RAND_1008;
  reg [31:0] _RAND_1009;
  reg [31:0] _RAND_1010;
  reg [31:0] _RAND_1011;
  reg [31:0] _RAND_1012;
  reg [31:0] _RAND_1013;
  reg [31:0] _RAND_1014;
  reg [31:0] _RAND_1015;
  reg [31:0] _RAND_1016;
  reg [31:0] _RAND_1017;
  reg [31:0] _RAND_1018;
  reg [31:0] _RAND_1019;
  reg [31:0] _RAND_1020;
  reg [31:0] _RAND_1021;
  reg [31:0] _RAND_1022;
  reg [31:0] _RAND_1023;
  reg [31:0] _RAND_1024;
  reg [31:0] _RAND_1025;
  reg [31:0] _RAND_1026;
  reg [31:0] _RAND_1027;
  reg [31:0] _RAND_1028;
  reg [255:0] _RAND_1029;
  reg [31:0] _RAND_1030;
  reg [31:0] _RAND_1031;
  reg [31:0] _RAND_1032;
  reg [31:0] _RAND_1033;
  reg [31:0] _RAND_1034;
  reg [31:0] _RAND_1035;
  reg [31:0] _RAND_1036;
  reg [31:0] _RAND_1037;
  reg [31:0] _RAND_1038;
`endif // RANDOMIZE_REG_INIT
  wire  rvclkhdr_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_1_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_1_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_1_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_1_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_2_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_2_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_2_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_2_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_3_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_3_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_3_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_3_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_4_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_4_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_4_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_4_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_5_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_5_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_5_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_5_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_6_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_6_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_6_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_6_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_7_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_7_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_7_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_7_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_8_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_8_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_8_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_8_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_9_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_9_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_9_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_9_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_10_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_10_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_10_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_10_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_11_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_11_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_11_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_11_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_12_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_12_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_12_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_12_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_13_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_13_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_13_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_13_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_14_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_14_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_14_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_14_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_15_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_15_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_15_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_15_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_16_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_16_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_16_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_16_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_17_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_17_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_17_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_17_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_18_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_18_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_18_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_18_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_19_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_19_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_19_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_19_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_20_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_20_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_20_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_20_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_21_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_21_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_21_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_21_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_22_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_22_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_22_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_22_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_23_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_23_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_23_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_23_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_24_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_24_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_24_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_24_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_25_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_25_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_25_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_25_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_26_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_26_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_26_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_26_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_27_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_27_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_27_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_27_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_28_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_28_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_28_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_28_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_29_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_29_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_29_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_29_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_30_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_30_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_30_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_30_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_31_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_31_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_31_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_31_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_32_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_32_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_32_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_32_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_33_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_33_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_33_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_33_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_34_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_34_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_34_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_34_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_35_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_35_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_35_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_35_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_36_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_36_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_36_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_36_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_37_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_37_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_37_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_37_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_38_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_38_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_38_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_38_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_39_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_39_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_39_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_39_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_40_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_40_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_40_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_40_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_41_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_41_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_41_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_41_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_42_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_42_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_42_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_42_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_43_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_43_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_43_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_43_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_44_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_44_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_44_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_44_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_45_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_45_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_45_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_45_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_46_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_46_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_46_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_46_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_47_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_47_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_47_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_47_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_48_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_48_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_48_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_48_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_49_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_49_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_49_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_49_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_50_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_50_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_50_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_50_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_51_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_51_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_51_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_51_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_52_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_52_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_52_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_52_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_53_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_53_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_53_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_53_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_54_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_54_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_54_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_54_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_55_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_55_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_55_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_55_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_56_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_56_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_56_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_56_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_57_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_57_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_57_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_57_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_58_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_58_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_58_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_58_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_59_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_59_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_59_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_59_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_60_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_60_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_60_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_60_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_61_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_61_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_61_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_61_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_62_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_62_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_62_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_62_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_63_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_63_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_63_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_63_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_64_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_64_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_64_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_64_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_65_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_65_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_65_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_65_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_66_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_66_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_66_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_66_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_67_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_67_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_67_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_67_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_68_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_68_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_68_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_68_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_69_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_69_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_69_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_69_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_70_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_70_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_70_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_70_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_71_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_71_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_71_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_71_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_72_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_72_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_72_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_72_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_73_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_73_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_73_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_73_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_74_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_74_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_74_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_74_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_75_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_75_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_75_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_75_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_76_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_76_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_76_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_76_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_77_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_77_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_77_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_77_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_78_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_78_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_78_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_78_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_79_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_79_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_79_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_79_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_80_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_80_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_80_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_80_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_81_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_81_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_81_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_81_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_82_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_82_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_82_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_82_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_83_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_83_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_83_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_83_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_84_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_84_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_84_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_84_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_85_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_85_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_85_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_85_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_86_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_86_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_86_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_86_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_87_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_87_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_87_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_87_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_88_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_88_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_88_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_88_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_89_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_89_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_89_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_89_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_90_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_90_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_90_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_90_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_91_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_91_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_91_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_91_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_92_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_92_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_92_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_92_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_93_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_93_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_93_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_93_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_94_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_94_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_94_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_94_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_95_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_95_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_95_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_95_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_96_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_96_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_96_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_96_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_97_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_97_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_97_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_97_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_98_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_98_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_98_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_98_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_99_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_99_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_99_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_99_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_100_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_100_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_100_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_100_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_101_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_101_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_101_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_101_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_102_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_102_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_102_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_102_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_103_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_103_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_103_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_103_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_104_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_104_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_104_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_104_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_105_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_105_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_105_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_105_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_106_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_106_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_106_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_106_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_107_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_107_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_107_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_107_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_108_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_108_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_108_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_108_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_109_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_109_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_109_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_109_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_110_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_110_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_110_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_110_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_111_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_111_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_111_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_111_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_112_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_112_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_112_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_112_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_113_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_113_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_113_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_113_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_114_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_114_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_114_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_114_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_115_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_115_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_115_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_115_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_116_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_116_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_116_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_116_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_117_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_117_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_117_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_117_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_118_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_118_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_118_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_118_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_119_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_119_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_119_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_119_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_120_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_120_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_120_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_120_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_121_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_121_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_121_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_121_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_122_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_122_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_122_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_122_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_123_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_123_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_123_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_123_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_124_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_124_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_124_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_124_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_125_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_125_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_125_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_125_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_126_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_126_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_126_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_126_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_127_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_127_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_127_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_127_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_128_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_128_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_128_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_128_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_129_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_129_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_129_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_129_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_130_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_130_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_130_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_130_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_131_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_131_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_131_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_131_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_132_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_132_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_132_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_132_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_133_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_133_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_133_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_133_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_134_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_134_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_134_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_134_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_135_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_135_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_135_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_135_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_136_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_136_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_136_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_136_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_137_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_137_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_137_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_137_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_138_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_138_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_138_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_138_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_139_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_139_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_139_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_139_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_140_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_140_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_140_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_140_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_141_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_141_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_141_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_141_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_142_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_142_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_142_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_142_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_143_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_143_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_143_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_143_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_144_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_144_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_144_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_144_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_145_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_145_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_145_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_145_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_146_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_146_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_146_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_146_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_147_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_147_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_147_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_147_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_148_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_148_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_148_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_148_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_149_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_149_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_149_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_149_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_150_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_150_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_150_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_150_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_151_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_151_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_151_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_151_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_152_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_152_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_152_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_152_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_153_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_153_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_153_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_153_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_154_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_154_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_154_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_154_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_155_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_155_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_155_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_155_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_156_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_156_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_156_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_156_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_157_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_157_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_157_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_157_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_158_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_158_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_158_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_158_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_159_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_159_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_159_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_159_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_160_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_160_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_160_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_160_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_161_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_161_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_161_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_161_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_162_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_162_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_162_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_162_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_163_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_163_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_163_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_163_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_164_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_164_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_164_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_164_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_165_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_165_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_165_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_165_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_166_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_166_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_166_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_166_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_167_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_167_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_167_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_167_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_168_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_168_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_168_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_168_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_169_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_169_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_169_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_169_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_170_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_170_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_170_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_170_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_171_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_171_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_171_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_171_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_172_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_172_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_172_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_172_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_173_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_173_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_173_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_173_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_174_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_174_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_174_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_174_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_175_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_175_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_175_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_175_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_176_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_176_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_176_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_176_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_177_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_177_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_177_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_177_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_178_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_178_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_178_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_178_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_179_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_179_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_179_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_179_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_180_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_180_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_180_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_180_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_181_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_181_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_181_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_181_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_182_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_182_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_182_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_182_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_183_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_183_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_183_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_183_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_184_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_184_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_184_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_184_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_185_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_185_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_185_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_185_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_186_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_186_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_186_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_186_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_187_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_187_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_187_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_187_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_188_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_188_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_188_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_188_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_189_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_189_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_189_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_189_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_190_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_190_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_190_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_190_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_191_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_191_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_191_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_191_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_192_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_192_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_192_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_192_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_193_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_193_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_193_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_193_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_194_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_194_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_194_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_194_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_195_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_195_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_195_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_195_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_196_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_196_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_196_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_196_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_197_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_197_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_197_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_197_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_198_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_198_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_198_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_198_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_199_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_199_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_199_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_199_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_200_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_200_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_200_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_200_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_201_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_201_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_201_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_201_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_202_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_202_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_202_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_202_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_203_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_203_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_203_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_203_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_204_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_204_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_204_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_204_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_205_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_205_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_205_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_205_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_206_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_206_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_206_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_206_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_207_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_207_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_207_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_207_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_208_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_208_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_208_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_208_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_209_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_209_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_209_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_209_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_210_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_210_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_210_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_210_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_211_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_211_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_211_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_211_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_212_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_212_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_212_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_212_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_213_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_213_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_213_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_213_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_214_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_214_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_214_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_214_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_215_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_215_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_215_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_215_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_216_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_216_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_216_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_216_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_217_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_217_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_217_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_217_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_218_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_218_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_218_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_218_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_219_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_219_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_219_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_219_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_220_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_220_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_220_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_220_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_221_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_221_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_221_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_221_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_222_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_222_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_222_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_222_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_223_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_223_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_223_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_223_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_224_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_224_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_224_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_224_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_225_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_225_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_225_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_225_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_226_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_226_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_226_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_226_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_227_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_227_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_227_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_227_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_228_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_228_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_228_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_228_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_229_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_229_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_229_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_229_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_230_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_230_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_230_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_230_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_231_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_231_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_231_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_231_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_232_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_232_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_232_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_232_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_233_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_233_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_233_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_233_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_234_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_234_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_234_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_234_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_235_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_235_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_235_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_235_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_236_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_236_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_236_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_236_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_237_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_237_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_237_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_237_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_238_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_238_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_238_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_238_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_239_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_239_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_239_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_239_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_240_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_240_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_240_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_240_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_241_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_241_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_241_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_241_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_242_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_242_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_242_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_242_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_243_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_243_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_243_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_243_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_244_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_244_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_244_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_244_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_245_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_245_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_245_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_245_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_246_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_246_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_246_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_246_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_247_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_247_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_247_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_247_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_248_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_248_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_248_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_248_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_249_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_249_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_249_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_249_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_250_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_250_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_250_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_250_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_251_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_251_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_251_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_251_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_252_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_252_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_252_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_252_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_253_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_253_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_253_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_253_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_254_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_254_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_254_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_254_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_255_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_255_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_255_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_255_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_256_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_256_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_256_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_256_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_257_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_257_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_257_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_257_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_258_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_258_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_258_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_258_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_259_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_259_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_259_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_259_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_260_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_260_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_260_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_260_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_261_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_261_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_261_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_261_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_262_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_262_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_262_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_262_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_263_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_263_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_263_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_263_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_264_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_264_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_264_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_264_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_265_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_265_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_265_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_265_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_266_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_266_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_266_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_266_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_267_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_267_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_267_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_267_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_268_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_268_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_268_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_268_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_269_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_269_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_269_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_269_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_270_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_270_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_270_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_270_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_271_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_271_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_271_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_271_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_272_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_272_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_272_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_272_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_273_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_273_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_273_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_273_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_274_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_274_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_274_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_274_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_275_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_275_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_275_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_275_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_276_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_276_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_276_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_276_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_277_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_277_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_277_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_277_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_278_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_278_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_278_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_278_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_279_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_279_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_279_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_279_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_280_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_280_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_280_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_280_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_281_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_281_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_281_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_281_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_282_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_282_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_282_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_282_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_283_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_283_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_283_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_283_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_284_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_284_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_284_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_284_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_285_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_285_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_285_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_285_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_286_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_286_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_286_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_286_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_287_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_287_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_287_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_287_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_288_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_288_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_288_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_288_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_289_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_289_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_289_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_289_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_290_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_290_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_290_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_290_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_291_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_291_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_291_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_291_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_292_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_292_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_292_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_292_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_293_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_293_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_293_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_293_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_294_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_294_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_294_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_294_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_295_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_295_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_295_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_295_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_296_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_296_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_296_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_296_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_297_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_297_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_297_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_297_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_298_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_298_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_298_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_298_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_299_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_299_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_299_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_299_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_300_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_300_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_300_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_300_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_301_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_301_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_301_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_301_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_302_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_302_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_302_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_302_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_303_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_303_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_303_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_303_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_304_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_304_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_304_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_304_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_305_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_305_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_305_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_305_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_306_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_306_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_306_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_306_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_307_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_307_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_307_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_307_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_308_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_308_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_308_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_308_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_309_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_309_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_309_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_309_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_310_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_310_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_310_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_310_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_311_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_311_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_311_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_311_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_312_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_312_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_312_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_312_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_313_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_313_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_313_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_313_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_314_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_314_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_314_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_314_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_315_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_315_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_315_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_315_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_316_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_316_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_316_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_316_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_317_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_317_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_317_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_317_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_318_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_318_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_318_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_318_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_319_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_319_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_319_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_319_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_320_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_320_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_320_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_320_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_321_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_321_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_321_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_321_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_322_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_322_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_322_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_322_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_323_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_323_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_323_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_323_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_324_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_324_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_324_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_324_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_325_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_325_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_325_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_325_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_326_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_326_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_326_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_326_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_327_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_327_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_327_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_327_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_328_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_328_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_328_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_328_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_329_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_329_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_329_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_329_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_330_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_330_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_330_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_330_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_331_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_331_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_331_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_331_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_332_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_332_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_332_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_332_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_333_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_333_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_333_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_333_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_334_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_334_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_334_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_334_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_335_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_335_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_335_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_335_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_336_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_336_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_336_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_336_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_337_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_337_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_337_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_337_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_338_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_338_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_338_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_338_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_339_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_339_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_339_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_339_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_340_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_340_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_340_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_340_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_341_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_341_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_341_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_341_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_342_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_342_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_342_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_342_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_343_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_343_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_343_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_343_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_344_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_344_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_344_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_344_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_345_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_345_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_345_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_345_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_346_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_346_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_346_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_346_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_347_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_347_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_347_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_347_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_348_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_348_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_348_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_348_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_349_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_349_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_349_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_349_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_350_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_350_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_350_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_350_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_351_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_351_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_351_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_351_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_352_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_352_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_352_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_352_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_353_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_353_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_353_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_353_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_354_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_354_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_354_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_354_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_355_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_355_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_355_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_355_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_356_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_356_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_356_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_356_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_357_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_357_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_357_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_357_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_358_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_358_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_358_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_358_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_359_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_359_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_359_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_359_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_360_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_360_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_360_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_360_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_361_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_361_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_361_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_361_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_362_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_362_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_362_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_362_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_363_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_363_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_363_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_363_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_364_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_364_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_364_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_364_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_365_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_365_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_365_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_365_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_366_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_366_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_366_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_366_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_367_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_367_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_367_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_367_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_368_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_368_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_368_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_368_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_369_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_369_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_369_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_369_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_370_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_370_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_370_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_370_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_371_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_371_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_371_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_371_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_372_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_372_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_372_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_372_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_373_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_373_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_373_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_373_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_374_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_374_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_374_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_374_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_375_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_375_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_375_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_375_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_376_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_376_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_376_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_376_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_377_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_377_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_377_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_377_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_378_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_378_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_378_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_378_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_379_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_379_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_379_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_379_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_380_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_380_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_380_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_380_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_381_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_381_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_381_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_381_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_382_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_382_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_382_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_382_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_383_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_383_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_383_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_383_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_384_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_384_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_384_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_384_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_385_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_385_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_385_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_385_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_386_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_386_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_386_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_386_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_387_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_387_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_387_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_387_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_388_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_388_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_388_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_388_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_389_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_389_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_389_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_389_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_390_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_390_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_390_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_390_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_391_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_391_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_391_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_391_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_392_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_392_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_392_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_392_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_393_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_393_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_393_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_393_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_394_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_394_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_394_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_394_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_395_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_395_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_395_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_395_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_396_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_396_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_396_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_396_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_397_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_397_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_397_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_397_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_398_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_398_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_398_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_398_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_399_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_399_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_399_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_399_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_400_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_400_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_400_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_400_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_401_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_401_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_401_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_401_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_402_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_402_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_402_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_402_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_403_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_403_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_403_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_403_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_404_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_404_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_404_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_404_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_405_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_405_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_405_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_405_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_406_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_406_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_406_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_406_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_407_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_407_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_407_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_407_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_408_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_408_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_408_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_408_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_409_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_409_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_409_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_409_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_410_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_410_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_410_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_410_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_411_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_411_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_411_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_411_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_412_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_412_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_412_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_412_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_413_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_413_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_413_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_413_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_414_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_414_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_414_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_414_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_415_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_415_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_415_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_415_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_416_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_416_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_416_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_416_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_417_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_417_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_417_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_417_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_418_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_418_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_418_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_418_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_419_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_419_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_419_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_419_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_420_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_420_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_420_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_420_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_421_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_421_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_421_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_421_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_422_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_422_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_422_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_422_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_423_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_423_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_423_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_423_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_424_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_424_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_424_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_424_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_425_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_425_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_425_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_425_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_426_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_426_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_426_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_426_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_427_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_427_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_427_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_427_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_428_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_428_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_428_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_428_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_429_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_429_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_429_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_429_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_430_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_430_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_430_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_430_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_431_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_431_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_431_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_431_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_432_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_432_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_432_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_432_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_433_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_433_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_433_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_433_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_434_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_434_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_434_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_434_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_435_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_435_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_435_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_435_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_436_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_436_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_436_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_436_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_437_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_437_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_437_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_437_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_438_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_438_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_438_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_438_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_439_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_439_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_439_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_439_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_440_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_440_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_440_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_440_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_441_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_441_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_441_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_441_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_442_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_442_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_442_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_442_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_443_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_443_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_443_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_443_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_444_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_444_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_444_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_444_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_445_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_445_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_445_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_445_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_446_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_446_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_446_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_446_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_447_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_447_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_447_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_447_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_448_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_448_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_448_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_448_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_449_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_449_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_449_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_449_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_450_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_450_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_450_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_450_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_451_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_451_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_451_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_451_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_452_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_452_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_452_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_452_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_453_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_453_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_453_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_453_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_454_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_454_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_454_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_454_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_455_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_455_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_455_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_455_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_456_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_456_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_456_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_456_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_457_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_457_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_457_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_457_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_458_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_458_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_458_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_458_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_459_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_459_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_459_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_459_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_460_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_460_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_460_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_460_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_461_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_461_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_461_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_461_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_462_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_462_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_462_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_462_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_463_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_463_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_463_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_463_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_464_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_464_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_464_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_464_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_465_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_465_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_465_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_465_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_466_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_466_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_466_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_466_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_467_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_467_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_467_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_467_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_468_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_468_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_468_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_468_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_469_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_469_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_469_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_469_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_470_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_470_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_470_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_470_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_471_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_471_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_471_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_471_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_472_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_472_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_472_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_472_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_473_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_473_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_473_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_473_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_474_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_474_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_474_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_474_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_475_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_475_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_475_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_475_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_476_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_476_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_476_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_476_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_477_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_477_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_477_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_477_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_478_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_478_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_478_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_478_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_479_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_479_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_479_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_479_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_480_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_480_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_480_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_480_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_481_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_481_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_481_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_481_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_482_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_482_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_482_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_482_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_483_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_483_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_483_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_483_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_484_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_484_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_484_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_484_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_485_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_485_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_485_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_485_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_486_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_486_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_486_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_486_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_487_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_487_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_487_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_487_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_488_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_488_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_488_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_488_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_489_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_489_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_489_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_489_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_490_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_490_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_490_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_490_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_491_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_491_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_491_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_491_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_492_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_492_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_492_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_492_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_493_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_493_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_493_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_493_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_494_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_494_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_494_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_494_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_495_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_495_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_495_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_495_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_496_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_496_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_496_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_496_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_497_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_497_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_497_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_497_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_498_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_498_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_498_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_498_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_499_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_499_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_499_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_499_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_500_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_500_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_500_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_500_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_501_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_501_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_501_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_501_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_502_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_502_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_502_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_502_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_503_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_503_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_503_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_503_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_504_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_504_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_504_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_504_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_505_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_505_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_505_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_505_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_506_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_506_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_506_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_506_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_507_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_507_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_507_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_507_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_508_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_508_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_508_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_508_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_509_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_509_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_509_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_509_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_510_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_510_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_510_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_510_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_511_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_511_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_511_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_511_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_512_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_512_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_512_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_512_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_513_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_513_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_513_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_513_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_514_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_514_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_514_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_514_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_515_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_515_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_515_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_515_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_516_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_516_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_516_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_516_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_517_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_517_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_517_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_517_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_518_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_518_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_518_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_518_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_519_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_519_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_519_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_519_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_520_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_520_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_520_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_520_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_521_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_521_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_521_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_521_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_522_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_522_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_522_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_522_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_523_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_523_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_523_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_523_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_524_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_524_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_524_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_524_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_525_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_525_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_525_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_525_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_526_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_526_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_526_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_526_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_527_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_527_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_527_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_527_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_528_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_528_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_528_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_528_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_529_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_529_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_529_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_529_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_530_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_530_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_530_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_530_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_531_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_531_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_531_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_531_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_532_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_532_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_532_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_532_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_533_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_533_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_533_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_533_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_534_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_534_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_534_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_534_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_535_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_535_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_535_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_535_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_536_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_536_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_536_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_536_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_537_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_537_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_537_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_537_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_538_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_538_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_538_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_538_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_539_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_539_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_539_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_539_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_540_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_540_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_540_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_540_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_541_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_541_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_541_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_541_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_542_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_542_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_542_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_542_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_543_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_543_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_543_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_543_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_544_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_544_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_544_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_544_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_545_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_545_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_545_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_545_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_546_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_546_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_546_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_546_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_547_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_547_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_547_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_547_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_548_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_548_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_548_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_548_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_549_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_549_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_549_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_549_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_550_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_550_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_550_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_550_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_551_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_551_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_551_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_551_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_552_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_552_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_552_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_552_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_553_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_553_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_553_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_553_io_scan_mode; // @[lib.scala 343:22]
  wire  _T_40 = io_dec_bp_dec_tlu_flush_leak_one_wb & io_dec_tlu_flush_lower_wb; // @[ifu_bp_ctl.scala 123:54]
  reg  leak_one_f_d1; // @[ifu_bp_ctl.scala 117:56]
  wire  _T_41 = ~io_dec_tlu_flush_lower_wb; // @[ifu_bp_ctl.scala 123:102]
  wire  _T_42 = leak_one_f_d1 & _T_41; // @[ifu_bp_ctl.scala 123:100]
  wire  leak_one_f = _T_40 | _T_42; // @[ifu_bp_ctl.scala 123:83]
  wire  _T = ~leak_one_f; // @[ifu_bp_ctl.scala 60:58]
  wire  exu_mp_valid = io_exu_bp_exu_mp_pkt_bits_misp & _T; // @[ifu_bp_ctl.scala 60:56]
  wire  dec_tlu_error_wb = io_dec_bp_dec_tlu_br0_r_pkt_bits_br_start_error | io_dec_bp_dec_tlu_br0_r_pkt_bits_br_error; // @[ifu_bp_ctl.scala 82:50]
  wire [7:0] _T_4 = io_ifc_fetch_addr_f[8:1] ^ io_ifc_fetch_addr_f[16:9]; // @[lib.scala 51:47]
  wire [7:0] btb_rd_addr_f = _T_4 ^ io_ifc_fetch_addr_f[24:17]; // @[lib.scala 51:85]
  wire [29:0] fetch_addr_p1_f = io_ifc_fetch_addr_f[30:1] + 30'h1; // @[ifu_bp_ctl.scala 90:51]
  wire [30:0] _T_8 = {fetch_addr_p1_f,1'h0}; // @[Cat.scala 29:58]
  wire [7:0] _T_11 = _T_8[8:1] ^ _T_8[16:9]; // @[lib.scala 51:47]
  wire [7:0] btb_rd_addr_p1_f = _T_11 ^ _T_8[24:17]; // @[lib.scala 51:85]
  wire  _T_144 = ~io_ifc_fetch_addr_f[0]; // @[ifu_bp_ctl.scala 174:40]
  wire  _T_2112 = btb_rd_addr_f == 8'h0; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_0; // @[lib.scala 374:16]
  wire [21:0] _T_2624 = _T_2112 ? btb_bank0_rd_data_way0_out_0 : 22'h0; // @[Mux.scala 27:72]
  wire  _T_2114 = btb_rd_addr_f == 8'h1; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_1; // @[lib.scala 374:16]
  wire [21:0] _T_2625 = _T_2114 ? btb_bank0_rd_data_way0_out_1 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2880 = _T_2624 | _T_2625; // @[Mux.scala 27:72]
  wire  _T_2116 = btb_rd_addr_f == 8'h2; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_2; // @[lib.scala 374:16]
  wire [21:0] _T_2626 = _T_2116 ? btb_bank0_rd_data_way0_out_2 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2881 = _T_2880 | _T_2626; // @[Mux.scala 27:72]
  wire  _T_2118 = btb_rd_addr_f == 8'h3; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_3; // @[lib.scala 374:16]
  wire [21:0] _T_2627 = _T_2118 ? btb_bank0_rd_data_way0_out_3 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2882 = _T_2881 | _T_2627; // @[Mux.scala 27:72]
  wire  _T_2120 = btb_rd_addr_f == 8'h4; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_4; // @[lib.scala 374:16]
  wire [21:0] _T_2628 = _T_2120 ? btb_bank0_rd_data_way0_out_4 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2883 = _T_2882 | _T_2628; // @[Mux.scala 27:72]
  wire  _T_2122 = btb_rd_addr_f == 8'h5; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_5; // @[lib.scala 374:16]
  wire [21:0] _T_2629 = _T_2122 ? btb_bank0_rd_data_way0_out_5 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2884 = _T_2883 | _T_2629; // @[Mux.scala 27:72]
  wire  _T_2124 = btb_rd_addr_f == 8'h6; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_6; // @[lib.scala 374:16]
  wire [21:0] _T_2630 = _T_2124 ? btb_bank0_rd_data_way0_out_6 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2885 = _T_2884 | _T_2630; // @[Mux.scala 27:72]
  wire  _T_2126 = btb_rd_addr_f == 8'h7; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_7; // @[lib.scala 374:16]
  wire [21:0] _T_2631 = _T_2126 ? btb_bank0_rd_data_way0_out_7 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2886 = _T_2885 | _T_2631; // @[Mux.scala 27:72]
  wire  _T_2128 = btb_rd_addr_f == 8'h8; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_8; // @[lib.scala 374:16]
  wire [21:0] _T_2632 = _T_2128 ? btb_bank0_rd_data_way0_out_8 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2887 = _T_2886 | _T_2632; // @[Mux.scala 27:72]
  wire  _T_2130 = btb_rd_addr_f == 8'h9; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_9; // @[lib.scala 374:16]
  wire [21:0] _T_2633 = _T_2130 ? btb_bank0_rd_data_way0_out_9 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2888 = _T_2887 | _T_2633; // @[Mux.scala 27:72]
  wire  _T_2132 = btb_rd_addr_f == 8'ha; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_10; // @[lib.scala 374:16]
  wire [21:0] _T_2634 = _T_2132 ? btb_bank0_rd_data_way0_out_10 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2889 = _T_2888 | _T_2634; // @[Mux.scala 27:72]
  wire  _T_2134 = btb_rd_addr_f == 8'hb; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_11; // @[lib.scala 374:16]
  wire [21:0] _T_2635 = _T_2134 ? btb_bank0_rd_data_way0_out_11 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2890 = _T_2889 | _T_2635; // @[Mux.scala 27:72]
  wire  _T_2136 = btb_rd_addr_f == 8'hc; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_12; // @[lib.scala 374:16]
  wire [21:0] _T_2636 = _T_2136 ? btb_bank0_rd_data_way0_out_12 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2891 = _T_2890 | _T_2636; // @[Mux.scala 27:72]
  wire  _T_2138 = btb_rd_addr_f == 8'hd; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_13; // @[lib.scala 374:16]
  wire [21:0] _T_2637 = _T_2138 ? btb_bank0_rd_data_way0_out_13 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2892 = _T_2891 | _T_2637; // @[Mux.scala 27:72]
  wire  _T_2140 = btb_rd_addr_f == 8'he; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_14; // @[lib.scala 374:16]
  wire [21:0] _T_2638 = _T_2140 ? btb_bank0_rd_data_way0_out_14 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2893 = _T_2892 | _T_2638; // @[Mux.scala 27:72]
  wire  _T_2142 = btb_rd_addr_f == 8'hf; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_15; // @[lib.scala 374:16]
  wire [21:0] _T_2639 = _T_2142 ? btb_bank0_rd_data_way0_out_15 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2894 = _T_2893 | _T_2639; // @[Mux.scala 27:72]
  wire  _T_2144 = btb_rd_addr_f == 8'h10; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_16; // @[lib.scala 374:16]
  wire [21:0] _T_2640 = _T_2144 ? btb_bank0_rd_data_way0_out_16 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2895 = _T_2894 | _T_2640; // @[Mux.scala 27:72]
  wire  _T_2146 = btb_rd_addr_f == 8'h11; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_17; // @[lib.scala 374:16]
  wire [21:0] _T_2641 = _T_2146 ? btb_bank0_rd_data_way0_out_17 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2896 = _T_2895 | _T_2641; // @[Mux.scala 27:72]
  wire  _T_2148 = btb_rd_addr_f == 8'h12; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_18; // @[lib.scala 374:16]
  wire [21:0] _T_2642 = _T_2148 ? btb_bank0_rd_data_way0_out_18 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2897 = _T_2896 | _T_2642; // @[Mux.scala 27:72]
  wire  _T_2150 = btb_rd_addr_f == 8'h13; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_19; // @[lib.scala 374:16]
  wire [21:0] _T_2643 = _T_2150 ? btb_bank0_rd_data_way0_out_19 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2898 = _T_2897 | _T_2643; // @[Mux.scala 27:72]
  wire  _T_2152 = btb_rd_addr_f == 8'h14; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_20; // @[lib.scala 374:16]
  wire [21:0] _T_2644 = _T_2152 ? btb_bank0_rd_data_way0_out_20 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2899 = _T_2898 | _T_2644; // @[Mux.scala 27:72]
  wire  _T_2154 = btb_rd_addr_f == 8'h15; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_21; // @[lib.scala 374:16]
  wire [21:0] _T_2645 = _T_2154 ? btb_bank0_rd_data_way0_out_21 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2900 = _T_2899 | _T_2645; // @[Mux.scala 27:72]
  wire  _T_2156 = btb_rd_addr_f == 8'h16; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_22; // @[lib.scala 374:16]
  wire [21:0] _T_2646 = _T_2156 ? btb_bank0_rd_data_way0_out_22 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2901 = _T_2900 | _T_2646; // @[Mux.scala 27:72]
  wire  _T_2158 = btb_rd_addr_f == 8'h17; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_23; // @[lib.scala 374:16]
  wire [21:0] _T_2647 = _T_2158 ? btb_bank0_rd_data_way0_out_23 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2902 = _T_2901 | _T_2647; // @[Mux.scala 27:72]
  wire  _T_2160 = btb_rd_addr_f == 8'h18; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_24; // @[lib.scala 374:16]
  wire [21:0] _T_2648 = _T_2160 ? btb_bank0_rd_data_way0_out_24 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2903 = _T_2902 | _T_2648; // @[Mux.scala 27:72]
  wire  _T_2162 = btb_rd_addr_f == 8'h19; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_25; // @[lib.scala 374:16]
  wire [21:0] _T_2649 = _T_2162 ? btb_bank0_rd_data_way0_out_25 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2904 = _T_2903 | _T_2649; // @[Mux.scala 27:72]
  wire  _T_2164 = btb_rd_addr_f == 8'h1a; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_26; // @[lib.scala 374:16]
  wire [21:0] _T_2650 = _T_2164 ? btb_bank0_rd_data_way0_out_26 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2905 = _T_2904 | _T_2650; // @[Mux.scala 27:72]
  wire  _T_2166 = btb_rd_addr_f == 8'h1b; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_27; // @[lib.scala 374:16]
  wire [21:0] _T_2651 = _T_2166 ? btb_bank0_rd_data_way0_out_27 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2906 = _T_2905 | _T_2651; // @[Mux.scala 27:72]
  wire  _T_2168 = btb_rd_addr_f == 8'h1c; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_28; // @[lib.scala 374:16]
  wire [21:0] _T_2652 = _T_2168 ? btb_bank0_rd_data_way0_out_28 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2907 = _T_2906 | _T_2652; // @[Mux.scala 27:72]
  wire  _T_2170 = btb_rd_addr_f == 8'h1d; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_29; // @[lib.scala 374:16]
  wire [21:0] _T_2653 = _T_2170 ? btb_bank0_rd_data_way0_out_29 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2908 = _T_2907 | _T_2653; // @[Mux.scala 27:72]
  wire  _T_2172 = btb_rd_addr_f == 8'h1e; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_30; // @[lib.scala 374:16]
  wire [21:0] _T_2654 = _T_2172 ? btb_bank0_rd_data_way0_out_30 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2909 = _T_2908 | _T_2654; // @[Mux.scala 27:72]
  wire  _T_2174 = btb_rd_addr_f == 8'h1f; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_31; // @[lib.scala 374:16]
  wire [21:0] _T_2655 = _T_2174 ? btb_bank0_rd_data_way0_out_31 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2910 = _T_2909 | _T_2655; // @[Mux.scala 27:72]
  wire  _T_2176 = btb_rd_addr_f == 8'h20; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_32; // @[lib.scala 374:16]
  wire [21:0] _T_2656 = _T_2176 ? btb_bank0_rd_data_way0_out_32 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2911 = _T_2910 | _T_2656; // @[Mux.scala 27:72]
  wire  _T_2178 = btb_rd_addr_f == 8'h21; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_33; // @[lib.scala 374:16]
  wire [21:0] _T_2657 = _T_2178 ? btb_bank0_rd_data_way0_out_33 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2912 = _T_2911 | _T_2657; // @[Mux.scala 27:72]
  wire  _T_2180 = btb_rd_addr_f == 8'h22; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_34; // @[lib.scala 374:16]
  wire [21:0] _T_2658 = _T_2180 ? btb_bank0_rd_data_way0_out_34 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2913 = _T_2912 | _T_2658; // @[Mux.scala 27:72]
  wire  _T_2182 = btb_rd_addr_f == 8'h23; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_35; // @[lib.scala 374:16]
  wire [21:0] _T_2659 = _T_2182 ? btb_bank0_rd_data_way0_out_35 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2914 = _T_2913 | _T_2659; // @[Mux.scala 27:72]
  wire  _T_2184 = btb_rd_addr_f == 8'h24; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_36; // @[lib.scala 374:16]
  wire [21:0] _T_2660 = _T_2184 ? btb_bank0_rd_data_way0_out_36 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2915 = _T_2914 | _T_2660; // @[Mux.scala 27:72]
  wire  _T_2186 = btb_rd_addr_f == 8'h25; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_37; // @[lib.scala 374:16]
  wire [21:0] _T_2661 = _T_2186 ? btb_bank0_rd_data_way0_out_37 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2916 = _T_2915 | _T_2661; // @[Mux.scala 27:72]
  wire  _T_2188 = btb_rd_addr_f == 8'h26; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_38; // @[lib.scala 374:16]
  wire [21:0] _T_2662 = _T_2188 ? btb_bank0_rd_data_way0_out_38 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2917 = _T_2916 | _T_2662; // @[Mux.scala 27:72]
  wire  _T_2190 = btb_rd_addr_f == 8'h27; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_39; // @[lib.scala 374:16]
  wire [21:0] _T_2663 = _T_2190 ? btb_bank0_rd_data_way0_out_39 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2918 = _T_2917 | _T_2663; // @[Mux.scala 27:72]
  wire  _T_2192 = btb_rd_addr_f == 8'h28; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_40; // @[lib.scala 374:16]
  wire [21:0] _T_2664 = _T_2192 ? btb_bank0_rd_data_way0_out_40 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2919 = _T_2918 | _T_2664; // @[Mux.scala 27:72]
  wire  _T_2194 = btb_rd_addr_f == 8'h29; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_41; // @[lib.scala 374:16]
  wire [21:0] _T_2665 = _T_2194 ? btb_bank0_rd_data_way0_out_41 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2920 = _T_2919 | _T_2665; // @[Mux.scala 27:72]
  wire  _T_2196 = btb_rd_addr_f == 8'h2a; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_42; // @[lib.scala 374:16]
  wire [21:0] _T_2666 = _T_2196 ? btb_bank0_rd_data_way0_out_42 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2921 = _T_2920 | _T_2666; // @[Mux.scala 27:72]
  wire  _T_2198 = btb_rd_addr_f == 8'h2b; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_43; // @[lib.scala 374:16]
  wire [21:0] _T_2667 = _T_2198 ? btb_bank0_rd_data_way0_out_43 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2922 = _T_2921 | _T_2667; // @[Mux.scala 27:72]
  wire  _T_2200 = btb_rd_addr_f == 8'h2c; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_44; // @[lib.scala 374:16]
  wire [21:0] _T_2668 = _T_2200 ? btb_bank0_rd_data_way0_out_44 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2923 = _T_2922 | _T_2668; // @[Mux.scala 27:72]
  wire  _T_2202 = btb_rd_addr_f == 8'h2d; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_45; // @[lib.scala 374:16]
  wire [21:0] _T_2669 = _T_2202 ? btb_bank0_rd_data_way0_out_45 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2924 = _T_2923 | _T_2669; // @[Mux.scala 27:72]
  wire  _T_2204 = btb_rd_addr_f == 8'h2e; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_46; // @[lib.scala 374:16]
  wire [21:0] _T_2670 = _T_2204 ? btb_bank0_rd_data_way0_out_46 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2925 = _T_2924 | _T_2670; // @[Mux.scala 27:72]
  wire  _T_2206 = btb_rd_addr_f == 8'h2f; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_47; // @[lib.scala 374:16]
  wire [21:0] _T_2671 = _T_2206 ? btb_bank0_rd_data_way0_out_47 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2926 = _T_2925 | _T_2671; // @[Mux.scala 27:72]
  wire  _T_2208 = btb_rd_addr_f == 8'h30; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_48; // @[lib.scala 374:16]
  wire [21:0] _T_2672 = _T_2208 ? btb_bank0_rd_data_way0_out_48 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2927 = _T_2926 | _T_2672; // @[Mux.scala 27:72]
  wire  _T_2210 = btb_rd_addr_f == 8'h31; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_49; // @[lib.scala 374:16]
  wire [21:0] _T_2673 = _T_2210 ? btb_bank0_rd_data_way0_out_49 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2928 = _T_2927 | _T_2673; // @[Mux.scala 27:72]
  wire  _T_2212 = btb_rd_addr_f == 8'h32; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_50; // @[lib.scala 374:16]
  wire [21:0] _T_2674 = _T_2212 ? btb_bank0_rd_data_way0_out_50 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2929 = _T_2928 | _T_2674; // @[Mux.scala 27:72]
  wire  _T_2214 = btb_rd_addr_f == 8'h33; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_51; // @[lib.scala 374:16]
  wire [21:0] _T_2675 = _T_2214 ? btb_bank0_rd_data_way0_out_51 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2930 = _T_2929 | _T_2675; // @[Mux.scala 27:72]
  wire  _T_2216 = btb_rd_addr_f == 8'h34; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_52; // @[lib.scala 374:16]
  wire [21:0] _T_2676 = _T_2216 ? btb_bank0_rd_data_way0_out_52 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2931 = _T_2930 | _T_2676; // @[Mux.scala 27:72]
  wire  _T_2218 = btb_rd_addr_f == 8'h35; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_53; // @[lib.scala 374:16]
  wire [21:0] _T_2677 = _T_2218 ? btb_bank0_rd_data_way0_out_53 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2932 = _T_2931 | _T_2677; // @[Mux.scala 27:72]
  wire  _T_2220 = btb_rd_addr_f == 8'h36; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_54; // @[lib.scala 374:16]
  wire [21:0] _T_2678 = _T_2220 ? btb_bank0_rd_data_way0_out_54 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2933 = _T_2932 | _T_2678; // @[Mux.scala 27:72]
  wire  _T_2222 = btb_rd_addr_f == 8'h37; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_55; // @[lib.scala 374:16]
  wire [21:0] _T_2679 = _T_2222 ? btb_bank0_rd_data_way0_out_55 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2934 = _T_2933 | _T_2679; // @[Mux.scala 27:72]
  wire  _T_2224 = btb_rd_addr_f == 8'h38; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_56; // @[lib.scala 374:16]
  wire [21:0] _T_2680 = _T_2224 ? btb_bank0_rd_data_way0_out_56 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2935 = _T_2934 | _T_2680; // @[Mux.scala 27:72]
  wire  _T_2226 = btb_rd_addr_f == 8'h39; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_57; // @[lib.scala 374:16]
  wire [21:0] _T_2681 = _T_2226 ? btb_bank0_rd_data_way0_out_57 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2936 = _T_2935 | _T_2681; // @[Mux.scala 27:72]
  wire  _T_2228 = btb_rd_addr_f == 8'h3a; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_58; // @[lib.scala 374:16]
  wire [21:0] _T_2682 = _T_2228 ? btb_bank0_rd_data_way0_out_58 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2937 = _T_2936 | _T_2682; // @[Mux.scala 27:72]
  wire  _T_2230 = btb_rd_addr_f == 8'h3b; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_59; // @[lib.scala 374:16]
  wire [21:0] _T_2683 = _T_2230 ? btb_bank0_rd_data_way0_out_59 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2938 = _T_2937 | _T_2683; // @[Mux.scala 27:72]
  wire  _T_2232 = btb_rd_addr_f == 8'h3c; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_60; // @[lib.scala 374:16]
  wire [21:0] _T_2684 = _T_2232 ? btb_bank0_rd_data_way0_out_60 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2939 = _T_2938 | _T_2684; // @[Mux.scala 27:72]
  wire  _T_2234 = btb_rd_addr_f == 8'h3d; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_61; // @[lib.scala 374:16]
  wire [21:0] _T_2685 = _T_2234 ? btb_bank0_rd_data_way0_out_61 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2940 = _T_2939 | _T_2685; // @[Mux.scala 27:72]
  wire  _T_2236 = btb_rd_addr_f == 8'h3e; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_62; // @[lib.scala 374:16]
  wire [21:0] _T_2686 = _T_2236 ? btb_bank0_rd_data_way0_out_62 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2941 = _T_2940 | _T_2686; // @[Mux.scala 27:72]
  wire  _T_2238 = btb_rd_addr_f == 8'h3f; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_63; // @[lib.scala 374:16]
  wire [21:0] _T_2687 = _T_2238 ? btb_bank0_rd_data_way0_out_63 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2942 = _T_2941 | _T_2687; // @[Mux.scala 27:72]
  wire  _T_2240 = btb_rd_addr_f == 8'h40; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_64; // @[lib.scala 374:16]
  wire [21:0] _T_2688 = _T_2240 ? btb_bank0_rd_data_way0_out_64 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2943 = _T_2942 | _T_2688; // @[Mux.scala 27:72]
  wire  _T_2242 = btb_rd_addr_f == 8'h41; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_65; // @[lib.scala 374:16]
  wire [21:0] _T_2689 = _T_2242 ? btb_bank0_rd_data_way0_out_65 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2944 = _T_2943 | _T_2689; // @[Mux.scala 27:72]
  wire  _T_2244 = btb_rd_addr_f == 8'h42; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_66; // @[lib.scala 374:16]
  wire [21:0] _T_2690 = _T_2244 ? btb_bank0_rd_data_way0_out_66 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2945 = _T_2944 | _T_2690; // @[Mux.scala 27:72]
  wire  _T_2246 = btb_rd_addr_f == 8'h43; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_67; // @[lib.scala 374:16]
  wire [21:0] _T_2691 = _T_2246 ? btb_bank0_rd_data_way0_out_67 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2946 = _T_2945 | _T_2691; // @[Mux.scala 27:72]
  wire  _T_2248 = btb_rd_addr_f == 8'h44; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_68; // @[lib.scala 374:16]
  wire [21:0] _T_2692 = _T_2248 ? btb_bank0_rd_data_way0_out_68 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2947 = _T_2946 | _T_2692; // @[Mux.scala 27:72]
  wire  _T_2250 = btb_rd_addr_f == 8'h45; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_69; // @[lib.scala 374:16]
  wire [21:0] _T_2693 = _T_2250 ? btb_bank0_rd_data_way0_out_69 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2948 = _T_2947 | _T_2693; // @[Mux.scala 27:72]
  wire  _T_2252 = btb_rd_addr_f == 8'h46; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_70; // @[lib.scala 374:16]
  wire [21:0] _T_2694 = _T_2252 ? btb_bank0_rd_data_way0_out_70 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2949 = _T_2948 | _T_2694; // @[Mux.scala 27:72]
  wire  _T_2254 = btb_rd_addr_f == 8'h47; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_71; // @[lib.scala 374:16]
  wire [21:0] _T_2695 = _T_2254 ? btb_bank0_rd_data_way0_out_71 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2950 = _T_2949 | _T_2695; // @[Mux.scala 27:72]
  wire  _T_2256 = btb_rd_addr_f == 8'h48; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_72; // @[lib.scala 374:16]
  wire [21:0] _T_2696 = _T_2256 ? btb_bank0_rd_data_way0_out_72 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2951 = _T_2950 | _T_2696; // @[Mux.scala 27:72]
  wire  _T_2258 = btb_rd_addr_f == 8'h49; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_73; // @[lib.scala 374:16]
  wire [21:0] _T_2697 = _T_2258 ? btb_bank0_rd_data_way0_out_73 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2952 = _T_2951 | _T_2697; // @[Mux.scala 27:72]
  wire  _T_2260 = btb_rd_addr_f == 8'h4a; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_74; // @[lib.scala 374:16]
  wire [21:0] _T_2698 = _T_2260 ? btb_bank0_rd_data_way0_out_74 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2953 = _T_2952 | _T_2698; // @[Mux.scala 27:72]
  wire  _T_2262 = btb_rd_addr_f == 8'h4b; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_75; // @[lib.scala 374:16]
  wire [21:0] _T_2699 = _T_2262 ? btb_bank0_rd_data_way0_out_75 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2954 = _T_2953 | _T_2699; // @[Mux.scala 27:72]
  wire  _T_2264 = btb_rd_addr_f == 8'h4c; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_76; // @[lib.scala 374:16]
  wire [21:0] _T_2700 = _T_2264 ? btb_bank0_rd_data_way0_out_76 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2955 = _T_2954 | _T_2700; // @[Mux.scala 27:72]
  wire  _T_2266 = btb_rd_addr_f == 8'h4d; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_77; // @[lib.scala 374:16]
  wire [21:0] _T_2701 = _T_2266 ? btb_bank0_rd_data_way0_out_77 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2956 = _T_2955 | _T_2701; // @[Mux.scala 27:72]
  wire  _T_2268 = btb_rd_addr_f == 8'h4e; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_78; // @[lib.scala 374:16]
  wire [21:0] _T_2702 = _T_2268 ? btb_bank0_rd_data_way0_out_78 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2957 = _T_2956 | _T_2702; // @[Mux.scala 27:72]
  wire  _T_2270 = btb_rd_addr_f == 8'h4f; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_79; // @[lib.scala 374:16]
  wire [21:0] _T_2703 = _T_2270 ? btb_bank0_rd_data_way0_out_79 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2958 = _T_2957 | _T_2703; // @[Mux.scala 27:72]
  wire  _T_2272 = btb_rd_addr_f == 8'h50; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_80; // @[lib.scala 374:16]
  wire [21:0] _T_2704 = _T_2272 ? btb_bank0_rd_data_way0_out_80 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2959 = _T_2958 | _T_2704; // @[Mux.scala 27:72]
  wire  _T_2274 = btb_rd_addr_f == 8'h51; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_81; // @[lib.scala 374:16]
  wire [21:0] _T_2705 = _T_2274 ? btb_bank0_rd_data_way0_out_81 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2960 = _T_2959 | _T_2705; // @[Mux.scala 27:72]
  wire  _T_2276 = btb_rd_addr_f == 8'h52; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_82; // @[lib.scala 374:16]
  wire [21:0] _T_2706 = _T_2276 ? btb_bank0_rd_data_way0_out_82 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2961 = _T_2960 | _T_2706; // @[Mux.scala 27:72]
  wire  _T_2278 = btb_rd_addr_f == 8'h53; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_83; // @[lib.scala 374:16]
  wire [21:0] _T_2707 = _T_2278 ? btb_bank0_rd_data_way0_out_83 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2962 = _T_2961 | _T_2707; // @[Mux.scala 27:72]
  wire  _T_2280 = btb_rd_addr_f == 8'h54; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_84; // @[lib.scala 374:16]
  wire [21:0] _T_2708 = _T_2280 ? btb_bank0_rd_data_way0_out_84 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2963 = _T_2962 | _T_2708; // @[Mux.scala 27:72]
  wire  _T_2282 = btb_rd_addr_f == 8'h55; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_85; // @[lib.scala 374:16]
  wire [21:0] _T_2709 = _T_2282 ? btb_bank0_rd_data_way0_out_85 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2964 = _T_2963 | _T_2709; // @[Mux.scala 27:72]
  wire  _T_2284 = btb_rd_addr_f == 8'h56; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_86; // @[lib.scala 374:16]
  wire [21:0] _T_2710 = _T_2284 ? btb_bank0_rd_data_way0_out_86 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2965 = _T_2964 | _T_2710; // @[Mux.scala 27:72]
  wire  _T_2286 = btb_rd_addr_f == 8'h57; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_87; // @[lib.scala 374:16]
  wire [21:0] _T_2711 = _T_2286 ? btb_bank0_rd_data_way0_out_87 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2966 = _T_2965 | _T_2711; // @[Mux.scala 27:72]
  wire  _T_2288 = btb_rd_addr_f == 8'h58; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_88; // @[lib.scala 374:16]
  wire [21:0] _T_2712 = _T_2288 ? btb_bank0_rd_data_way0_out_88 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2967 = _T_2966 | _T_2712; // @[Mux.scala 27:72]
  wire  _T_2290 = btb_rd_addr_f == 8'h59; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_89; // @[lib.scala 374:16]
  wire [21:0] _T_2713 = _T_2290 ? btb_bank0_rd_data_way0_out_89 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2968 = _T_2967 | _T_2713; // @[Mux.scala 27:72]
  wire  _T_2292 = btb_rd_addr_f == 8'h5a; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_90; // @[lib.scala 374:16]
  wire [21:0] _T_2714 = _T_2292 ? btb_bank0_rd_data_way0_out_90 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2969 = _T_2968 | _T_2714; // @[Mux.scala 27:72]
  wire  _T_2294 = btb_rd_addr_f == 8'h5b; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_91; // @[lib.scala 374:16]
  wire [21:0] _T_2715 = _T_2294 ? btb_bank0_rd_data_way0_out_91 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2970 = _T_2969 | _T_2715; // @[Mux.scala 27:72]
  wire  _T_2296 = btb_rd_addr_f == 8'h5c; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_92; // @[lib.scala 374:16]
  wire [21:0] _T_2716 = _T_2296 ? btb_bank0_rd_data_way0_out_92 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2971 = _T_2970 | _T_2716; // @[Mux.scala 27:72]
  wire  _T_2298 = btb_rd_addr_f == 8'h5d; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_93; // @[lib.scala 374:16]
  wire [21:0] _T_2717 = _T_2298 ? btb_bank0_rd_data_way0_out_93 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2972 = _T_2971 | _T_2717; // @[Mux.scala 27:72]
  wire  _T_2300 = btb_rd_addr_f == 8'h5e; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_94; // @[lib.scala 374:16]
  wire [21:0] _T_2718 = _T_2300 ? btb_bank0_rd_data_way0_out_94 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2973 = _T_2972 | _T_2718; // @[Mux.scala 27:72]
  wire  _T_2302 = btb_rd_addr_f == 8'h5f; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_95; // @[lib.scala 374:16]
  wire [21:0] _T_2719 = _T_2302 ? btb_bank0_rd_data_way0_out_95 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2974 = _T_2973 | _T_2719; // @[Mux.scala 27:72]
  wire  _T_2304 = btb_rd_addr_f == 8'h60; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_96; // @[lib.scala 374:16]
  wire [21:0] _T_2720 = _T_2304 ? btb_bank0_rd_data_way0_out_96 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2975 = _T_2974 | _T_2720; // @[Mux.scala 27:72]
  wire  _T_2306 = btb_rd_addr_f == 8'h61; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_97; // @[lib.scala 374:16]
  wire [21:0] _T_2721 = _T_2306 ? btb_bank0_rd_data_way0_out_97 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2976 = _T_2975 | _T_2721; // @[Mux.scala 27:72]
  wire  _T_2308 = btb_rd_addr_f == 8'h62; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_98; // @[lib.scala 374:16]
  wire [21:0] _T_2722 = _T_2308 ? btb_bank0_rd_data_way0_out_98 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2977 = _T_2976 | _T_2722; // @[Mux.scala 27:72]
  wire  _T_2310 = btb_rd_addr_f == 8'h63; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_99; // @[lib.scala 374:16]
  wire [21:0] _T_2723 = _T_2310 ? btb_bank0_rd_data_way0_out_99 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2978 = _T_2977 | _T_2723; // @[Mux.scala 27:72]
  wire  _T_2312 = btb_rd_addr_f == 8'h64; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_100; // @[lib.scala 374:16]
  wire [21:0] _T_2724 = _T_2312 ? btb_bank0_rd_data_way0_out_100 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2979 = _T_2978 | _T_2724; // @[Mux.scala 27:72]
  wire  _T_2314 = btb_rd_addr_f == 8'h65; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_101; // @[lib.scala 374:16]
  wire [21:0] _T_2725 = _T_2314 ? btb_bank0_rd_data_way0_out_101 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2980 = _T_2979 | _T_2725; // @[Mux.scala 27:72]
  wire  _T_2316 = btb_rd_addr_f == 8'h66; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_102; // @[lib.scala 374:16]
  wire [21:0] _T_2726 = _T_2316 ? btb_bank0_rd_data_way0_out_102 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2981 = _T_2980 | _T_2726; // @[Mux.scala 27:72]
  wire  _T_2318 = btb_rd_addr_f == 8'h67; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_103; // @[lib.scala 374:16]
  wire [21:0] _T_2727 = _T_2318 ? btb_bank0_rd_data_way0_out_103 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2982 = _T_2981 | _T_2727; // @[Mux.scala 27:72]
  wire  _T_2320 = btb_rd_addr_f == 8'h68; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_104; // @[lib.scala 374:16]
  wire [21:0] _T_2728 = _T_2320 ? btb_bank0_rd_data_way0_out_104 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2983 = _T_2982 | _T_2728; // @[Mux.scala 27:72]
  wire  _T_2322 = btb_rd_addr_f == 8'h69; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_105; // @[lib.scala 374:16]
  wire [21:0] _T_2729 = _T_2322 ? btb_bank0_rd_data_way0_out_105 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2984 = _T_2983 | _T_2729; // @[Mux.scala 27:72]
  wire  _T_2324 = btb_rd_addr_f == 8'h6a; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_106; // @[lib.scala 374:16]
  wire [21:0] _T_2730 = _T_2324 ? btb_bank0_rd_data_way0_out_106 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2985 = _T_2984 | _T_2730; // @[Mux.scala 27:72]
  wire  _T_2326 = btb_rd_addr_f == 8'h6b; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_107; // @[lib.scala 374:16]
  wire [21:0] _T_2731 = _T_2326 ? btb_bank0_rd_data_way0_out_107 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2986 = _T_2985 | _T_2731; // @[Mux.scala 27:72]
  wire  _T_2328 = btb_rd_addr_f == 8'h6c; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_108; // @[lib.scala 374:16]
  wire [21:0] _T_2732 = _T_2328 ? btb_bank0_rd_data_way0_out_108 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2987 = _T_2986 | _T_2732; // @[Mux.scala 27:72]
  wire  _T_2330 = btb_rd_addr_f == 8'h6d; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_109; // @[lib.scala 374:16]
  wire [21:0] _T_2733 = _T_2330 ? btb_bank0_rd_data_way0_out_109 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2988 = _T_2987 | _T_2733; // @[Mux.scala 27:72]
  wire  _T_2332 = btb_rd_addr_f == 8'h6e; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_110; // @[lib.scala 374:16]
  wire [21:0] _T_2734 = _T_2332 ? btb_bank0_rd_data_way0_out_110 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2989 = _T_2988 | _T_2734; // @[Mux.scala 27:72]
  wire  _T_2334 = btb_rd_addr_f == 8'h6f; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_111; // @[lib.scala 374:16]
  wire [21:0] _T_2735 = _T_2334 ? btb_bank0_rd_data_way0_out_111 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2990 = _T_2989 | _T_2735; // @[Mux.scala 27:72]
  wire  _T_2336 = btb_rd_addr_f == 8'h70; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_112; // @[lib.scala 374:16]
  wire [21:0] _T_2736 = _T_2336 ? btb_bank0_rd_data_way0_out_112 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2991 = _T_2990 | _T_2736; // @[Mux.scala 27:72]
  wire  _T_2338 = btb_rd_addr_f == 8'h71; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_113; // @[lib.scala 374:16]
  wire [21:0] _T_2737 = _T_2338 ? btb_bank0_rd_data_way0_out_113 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2992 = _T_2991 | _T_2737; // @[Mux.scala 27:72]
  wire  _T_2340 = btb_rd_addr_f == 8'h72; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_114; // @[lib.scala 374:16]
  wire [21:0] _T_2738 = _T_2340 ? btb_bank0_rd_data_way0_out_114 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2993 = _T_2992 | _T_2738; // @[Mux.scala 27:72]
  wire  _T_2342 = btb_rd_addr_f == 8'h73; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_115; // @[lib.scala 374:16]
  wire [21:0] _T_2739 = _T_2342 ? btb_bank0_rd_data_way0_out_115 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2994 = _T_2993 | _T_2739; // @[Mux.scala 27:72]
  wire  _T_2344 = btb_rd_addr_f == 8'h74; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_116; // @[lib.scala 374:16]
  wire [21:0] _T_2740 = _T_2344 ? btb_bank0_rd_data_way0_out_116 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2995 = _T_2994 | _T_2740; // @[Mux.scala 27:72]
  wire  _T_2346 = btb_rd_addr_f == 8'h75; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_117; // @[lib.scala 374:16]
  wire [21:0] _T_2741 = _T_2346 ? btb_bank0_rd_data_way0_out_117 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2996 = _T_2995 | _T_2741; // @[Mux.scala 27:72]
  wire  _T_2348 = btb_rd_addr_f == 8'h76; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_118; // @[lib.scala 374:16]
  wire [21:0] _T_2742 = _T_2348 ? btb_bank0_rd_data_way0_out_118 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2997 = _T_2996 | _T_2742; // @[Mux.scala 27:72]
  wire  _T_2350 = btb_rd_addr_f == 8'h77; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_119; // @[lib.scala 374:16]
  wire [21:0] _T_2743 = _T_2350 ? btb_bank0_rd_data_way0_out_119 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2998 = _T_2997 | _T_2743; // @[Mux.scala 27:72]
  wire  _T_2352 = btb_rd_addr_f == 8'h78; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_120; // @[lib.scala 374:16]
  wire [21:0] _T_2744 = _T_2352 ? btb_bank0_rd_data_way0_out_120 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2999 = _T_2998 | _T_2744; // @[Mux.scala 27:72]
  wire  _T_2354 = btb_rd_addr_f == 8'h79; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_121; // @[lib.scala 374:16]
  wire [21:0] _T_2745 = _T_2354 ? btb_bank0_rd_data_way0_out_121 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3000 = _T_2999 | _T_2745; // @[Mux.scala 27:72]
  wire  _T_2356 = btb_rd_addr_f == 8'h7a; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_122; // @[lib.scala 374:16]
  wire [21:0] _T_2746 = _T_2356 ? btb_bank0_rd_data_way0_out_122 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3001 = _T_3000 | _T_2746; // @[Mux.scala 27:72]
  wire  _T_2358 = btb_rd_addr_f == 8'h7b; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_123; // @[lib.scala 374:16]
  wire [21:0] _T_2747 = _T_2358 ? btb_bank0_rd_data_way0_out_123 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3002 = _T_3001 | _T_2747; // @[Mux.scala 27:72]
  wire  _T_2360 = btb_rd_addr_f == 8'h7c; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_124; // @[lib.scala 374:16]
  wire [21:0] _T_2748 = _T_2360 ? btb_bank0_rd_data_way0_out_124 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3003 = _T_3002 | _T_2748; // @[Mux.scala 27:72]
  wire  _T_2362 = btb_rd_addr_f == 8'h7d; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_125; // @[lib.scala 374:16]
  wire [21:0] _T_2749 = _T_2362 ? btb_bank0_rd_data_way0_out_125 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3004 = _T_3003 | _T_2749; // @[Mux.scala 27:72]
  wire  _T_2364 = btb_rd_addr_f == 8'h7e; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_126; // @[lib.scala 374:16]
  wire [21:0] _T_2750 = _T_2364 ? btb_bank0_rd_data_way0_out_126 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3005 = _T_3004 | _T_2750; // @[Mux.scala 27:72]
  wire  _T_2366 = btb_rd_addr_f == 8'h7f; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_127; // @[lib.scala 374:16]
  wire [21:0] _T_2751 = _T_2366 ? btb_bank0_rd_data_way0_out_127 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3006 = _T_3005 | _T_2751; // @[Mux.scala 27:72]
  wire  _T_2368 = btb_rd_addr_f == 8'h80; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_128; // @[lib.scala 374:16]
  wire [21:0] _T_2752 = _T_2368 ? btb_bank0_rd_data_way0_out_128 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3007 = _T_3006 | _T_2752; // @[Mux.scala 27:72]
  wire  _T_2370 = btb_rd_addr_f == 8'h81; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_129; // @[lib.scala 374:16]
  wire [21:0] _T_2753 = _T_2370 ? btb_bank0_rd_data_way0_out_129 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3008 = _T_3007 | _T_2753; // @[Mux.scala 27:72]
  wire  _T_2372 = btb_rd_addr_f == 8'h82; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_130; // @[lib.scala 374:16]
  wire [21:0] _T_2754 = _T_2372 ? btb_bank0_rd_data_way0_out_130 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3009 = _T_3008 | _T_2754; // @[Mux.scala 27:72]
  wire  _T_2374 = btb_rd_addr_f == 8'h83; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_131; // @[lib.scala 374:16]
  wire [21:0] _T_2755 = _T_2374 ? btb_bank0_rd_data_way0_out_131 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3010 = _T_3009 | _T_2755; // @[Mux.scala 27:72]
  wire  _T_2376 = btb_rd_addr_f == 8'h84; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_132; // @[lib.scala 374:16]
  wire [21:0] _T_2756 = _T_2376 ? btb_bank0_rd_data_way0_out_132 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3011 = _T_3010 | _T_2756; // @[Mux.scala 27:72]
  wire  _T_2378 = btb_rd_addr_f == 8'h85; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_133; // @[lib.scala 374:16]
  wire [21:0] _T_2757 = _T_2378 ? btb_bank0_rd_data_way0_out_133 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3012 = _T_3011 | _T_2757; // @[Mux.scala 27:72]
  wire  _T_2380 = btb_rd_addr_f == 8'h86; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_134; // @[lib.scala 374:16]
  wire [21:0] _T_2758 = _T_2380 ? btb_bank0_rd_data_way0_out_134 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3013 = _T_3012 | _T_2758; // @[Mux.scala 27:72]
  wire  _T_2382 = btb_rd_addr_f == 8'h87; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_135; // @[lib.scala 374:16]
  wire [21:0] _T_2759 = _T_2382 ? btb_bank0_rd_data_way0_out_135 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3014 = _T_3013 | _T_2759; // @[Mux.scala 27:72]
  wire  _T_2384 = btb_rd_addr_f == 8'h88; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_136; // @[lib.scala 374:16]
  wire [21:0] _T_2760 = _T_2384 ? btb_bank0_rd_data_way0_out_136 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3015 = _T_3014 | _T_2760; // @[Mux.scala 27:72]
  wire  _T_2386 = btb_rd_addr_f == 8'h89; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_137; // @[lib.scala 374:16]
  wire [21:0] _T_2761 = _T_2386 ? btb_bank0_rd_data_way0_out_137 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3016 = _T_3015 | _T_2761; // @[Mux.scala 27:72]
  wire  _T_2388 = btb_rd_addr_f == 8'h8a; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_138; // @[lib.scala 374:16]
  wire [21:0] _T_2762 = _T_2388 ? btb_bank0_rd_data_way0_out_138 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3017 = _T_3016 | _T_2762; // @[Mux.scala 27:72]
  wire  _T_2390 = btb_rd_addr_f == 8'h8b; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_139; // @[lib.scala 374:16]
  wire [21:0] _T_2763 = _T_2390 ? btb_bank0_rd_data_way0_out_139 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3018 = _T_3017 | _T_2763; // @[Mux.scala 27:72]
  wire  _T_2392 = btb_rd_addr_f == 8'h8c; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_140; // @[lib.scala 374:16]
  wire [21:0] _T_2764 = _T_2392 ? btb_bank0_rd_data_way0_out_140 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3019 = _T_3018 | _T_2764; // @[Mux.scala 27:72]
  wire  _T_2394 = btb_rd_addr_f == 8'h8d; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_141; // @[lib.scala 374:16]
  wire [21:0] _T_2765 = _T_2394 ? btb_bank0_rd_data_way0_out_141 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3020 = _T_3019 | _T_2765; // @[Mux.scala 27:72]
  wire  _T_2396 = btb_rd_addr_f == 8'h8e; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_142; // @[lib.scala 374:16]
  wire [21:0] _T_2766 = _T_2396 ? btb_bank0_rd_data_way0_out_142 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3021 = _T_3020 | _T_2766; // @[Mux.scala 27:72]
  wire  _T_2398 = btb_rd_addr_f == 8'h8f; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_143; // @[lib.scala 374:16]
  wire [21:0] _T_2767 = _T_2398 ? btb_bank0_rd_data_way0_out_143 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3022 = _T_3021 | _T_2767; // @[Mux.scala 27:72]
  wire  _T_2400 = btb_rd_addr_f == 8'h90; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_144; // @[lib.scala 374:16]
  wire [21:0] _T_2768 = _T_2400 ? btb_bank0_rd_data_way0_out_144 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3023 = _T_3022 | _T_2768; // @[Mux.scala 27:72]
  wire  _T_2402 = btb_rd_addr_f == 8'h91; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_145; // @[lib.scala 374:16]
  wire [21:0] _T_2769 = _T_2402 ? btb_bank0_rd_data_way0_out_145 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3024 = _T_3023 | _T_2769; // @[Mux.scala 27:72]
  wire  _T_2404 = btb_rd_addr_f == 8'h92; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_146; // @[lib.scala 374:16]
  wire [21:0] _T_2770 = _T_2404 ? btb_bank0_rd_data_way0_out_146 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3025 = _T_3024 | _T_2770; // @[Mux.scala 27:72]
  wire  _T_2406 = btb_rd_addr_f == 8'h93; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_147; // @[lib.scala 374:16]
  wire [21:0] _T_2771 = _T_2406 ? btb_bank0_rd_data_way0_out_147 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3026 = _T_3025 | _T_2771; // @[Mux.scala 27:72]
  wire  _T_2408 = btb_rd_addr_f == 8'h94; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_148; // @[lib.scala 374:16]
  wire [21:0] _T_2772 = _T_2408 ? btb_bank0_rd_data_way0_out_148 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3027 = _T_3026 | _T_2772; // @[Mux.scala 27:72]
  wire  _T_2410 = btb_rd_addr_f == 8'h95; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_149; // @[lib.scala 374:16]
  wire [21:0] _T_2773 = _T_2410 ? btb_bank0_rd_data_way0_out_149 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3028 = _T_3027 | _T_2773; // @[Mux.scala 27:72]
  wire  _T_2412 = btb_rd_addr_f == 8'h96; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_150; // @[lib.scala 374:16]
  wire [21:0] _T_2774 = _T_2412 ? btb_bank0_rd_data_way0_out_150 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3029 = _T_3028 | _T_2774; // @[Mux.scala 27:72]
  wire  _T_2414 = btb_rd_addr_f == 8'h97; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_151; // @[lib.scala 374:16]
  wire [21:0] _T_2775 = _T_2414 ? btb_bank0_rd_data_way0_out_151 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3030 = _T_3029 | _T_2775; // @[Mux.scala 27:72]
  wire  _T_2416 = btb_rd_addr_f == 8'h98; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_152; // @[lib.scala 374:16]
  wire [21:0] _T_2776 = _T_2416 ? btb_bank0_rd_data_way0_out_152 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3031 = _T_3030 | _T_2776; // @[Mux.scala 27:72]
  wire  _T_2418 = btb_rd_addr_f == 8'h99; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_153; // @[lib.scala 374:16]
  wire [21:0] _T_2777 = _T_2418 ? btb_bank0_rd_data_way0_out_153 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3032 = _T_3031 | _T_2777; // @[Mux.scala 27:72]
  wire  _T_2420 = btb_rd_addr_f == 8'h9a; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_154; // @[lib.scala 374:16]
  wire [21:0] _T_2778 = _T_2420 ? btb_bank0_rd_data_way0_out_154 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3033 = _T_3032 | _T_2778; // @[Mux.scala 27:72]
  wire  _T_2422 = btb_rd_addr_f == 8'h9b; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_155; // @[lib.scala 374:16]
  wire [21:0] _T_2779 = _T_2422 ? btb_bank0_rd_data_way0_out_155 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3034 = _T_3033 | _T_2779; // @[Mux.scala 27:72]
  wire  _T_2424 = btb_rd_addr_f == 8'h9c; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_156; // @[lib.scala 374:16]
  wire [21:0] _T_2780 = _T_2424 ? btb_bank0_rd_data_way0_out_156 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3035 = _T_3034 | _T_2780; // @[Mux.scala 27:72]
  wire  _T_2426 = btb_rd_addr_f == 8'h9d; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_157; // @[lib.scala 374:16]
  wire [21:0] _T_2781 = _T_2426 ? btb_bank0_rd_data_way0_out_157 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3036 = _T_3035 | _T_2781; // @[Mux.scala 27:72]
  wire  _T_2428 = btb_rd_addr_f == 8'h9e; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_158; // @[lib.scala 374:16]
  wire [21:0] _T_2782 = _T_2428 ? btb_bank0_rd_data_way0_out_158 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3037 = _T_3036 | _T_2782; // @[Mux.scala 27:72]
  wire  _T_2430 = btb_rd_addr_f == 8'h9f; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_159; // @[lib.scala 374:16]
  wire [21:0] _T_2783 = _T_2430 ? btb_bank0_rd_data_way0_out_159 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3038 = _T_3037 | _T_2783; // @[Mux.scala 27:72]
  wire  _T_2432 = btb_rd_addr_f == 8'ha0; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_160; // @[lib.scala 374:16]
  wire [21:0] _T_2784 = _T_2432 ? btb_bank0_rd_data_way0_out_160 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3039 = _T_3038 | _T_2784; // @[Mux.scala 27:72]
  wire  _T_2434 = btb_rd_addr_f == 8'ha1; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_161; // @[lib.scala 374:16]
  wire [21:0] _T_2785 = _T_2434 ? btb_bank0_rd_data_way0_out_161 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3040 = _T_3039 | _T_2785; // @[Mux.scala 27:72]
  wire  _T_2436 = btb_rd_addr_f == 8'ha2; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_162; // @[lib.scala 374:16]
  wire [21:0] _T_2786 = _T_2436 ? btb_bank0_rd_data_way0_out_162 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3041 = _T_3040 | _T_2786; // @[Mux.scala 27:72]
  wire  _T_2438 = btb_rd_addr_f == 8'ha3; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_163; // @[lib.scala 374:16]
  wire [21:0] _T_2787 = _T_2438 ? btb_bank0_rd_data_way0_out_163 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3042 = _T_3041 | _T_2787; // @[Mux.scala 27:72]
  wire  _T_2440 = btb_rd_addr_f == 8'ha4; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_164; // @[lib.scala 374:16]
  wire [21:0] _T_2788 = _T_2440 ? btb_bank0_rd_data_way0_out_164 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3043 = _T_3042 | _T_2788; // @[Mux.scala 27:72]
  wire  _T_2442 = btb_rd_addr_f == 8'ha5; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_165; // @[lib.scala 374:16]
  wire [21:0] _T_2789 = _T_2442 ? btb_bank0_rd_data_way0_out_165 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3044 = _T_3043 | _T_2789; // @[Mux.scala 27:72]
  wire  _T_2444 = btb_rd_addr_f == 8'ha6; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_166; // @[lib.scala 374:16]
  wire [21:0] _T_2790 = _T_2444 ? btb_bank0_rd_data_way0_out_166 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3045 = _T_3044 | _T_2790; // @[Mux.scala 27:72]
  wire  _T_2446 = btb_rd_addr_f == 8'ha7; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_167; // @[lib.scala 374:16]
  wire [21:0] _T_2791 = _T_2446 ? btb_bank0_rd_data_way0_out_167 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3046 = _T_3045 | _T_2791; // @[Mux.scala 27:72]
  wire  _T_2448 = btb_rd_addr_f == 8'ha8; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_168; // @[lib.scala 374:16]
  wire [21:0] _T_2792 = _T_2448 ? btb_bank0_rd_data_way0_out_168 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3047 = _T_3046 | _T_2792; // @[Mux.scala 27:72]
  wire  _T_2450 = btb_rd_addr_f == 8'ha9; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_169; // @[lib.scala 374:16]
  wire [21:0] _T_2793 = _T_2450 ? btb_bank0_rd_data_way0_out_169 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3048 = _T_3047 | _T_2793; // @[Mux.scala 27:72]
  wire  _T_2452 = btb_rd_addr_f == 8'haa; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_170; // @[lib.scala 374:16]
  wire [21:0] _T_2794 = _T_2452 ? btb_bank0_rd_data_way0_out_170 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3049 = _T_3048 | _T_2794; // @[Mux.scala 27:72]
  wire  _T_2454 = btb_rd_addr_f == 8'hab; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_171; // @[lib.scala 374:16]
  wire [21:0] _T_2795 = _T_2454 ? btb_bank0_rd_data_way0_out_171 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3050 = _T_3049 | _T_2795; // @[Mux.scala 27:72]
  wire  _T_2456 = btb_rd_addr_f == 8'hac; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_172; // @[lib.scala 374:16]
  wire [21:0] _T_2796 = _T_2456 ? btb_bank0_rd_data_way0_out_172 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3051 = _T_3050 | _T_2796; // @[Mux.scala 27:72]
  wire  _T_2458 = btb_rd_addr_f == 8'had; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_173; // @[lib.scala 374:16]
  wire [21:0] _T_2797 = _T_2458 ? btb_bank0_rd_data_way0_out_173 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3052 = _T_3051 | _T_2797; // @[Mux.scala 27:72]
  wire  _T_2460 = btb_rd_addr_f == 8'hae; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_174; // @[lib.scala 374:16]
  wire [21:0] _T_2798 = _T_2460 ? btb_bank0_rd_data_way0_out_174 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3053 = _T_3052 | _T_2798; // @[Mux.scala 27:72]
  wire  _T_2462 = btb_rd_addr_f == 8'haf; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_175; // @[lib.scala 374:16]
  wire [21:0] _T_2799 = _T_2462 ? btb_bank0_rd_data_way0_out_175 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3054 = _T_3053 | _T_2799; // @[Mux.scala 27:72]
  wire  _T_2464 = btb_rd_addr_f == 8'hb0; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_176; // @[lib.scala 374:16]
  wire [21:0] _T_2800 = _T_2464 ? btb_bank0_rd_data_way0_out_176 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3055 = _T_3054 | _T_2800; // @[Mux.scala 27:72]
  wire  _T_2466 = btb_rd_addr_f == 8'hb1; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_177; // @[lib.scala 374:16]
  wire [21:0] _T_2801 = _T_2466 ? btb_bank0_rd_data_way0_out_177 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3056 = _T_3055 | _T_2801; // @[Mux.scala 27:72]
  wire  _T_2468 = btb_rd_addr_f == 8'hb2; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_178; // @[lib.scala 374:16]
  wire [21:0] _T_2802 = _T_2468 ? btb_bank0_rd_data_way0_out_178 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3057 = _T_3056 | _T_2802; // @[Mux.scala 27:72]
  wire  _T_2470 = btb_rd_addr_f == 8'hb3; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_179; // @[lib.scala 374:16]
  wire [21:0] _T_2803 = _T_2470 ? btb_bank0_rd_data_way0_out_179 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3058 = _T_3057 | _T_2803; // @[Mux.scala 27:72]
  wire  _T_2472 = btb_rd_addr_f == 8'hb4; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_180; // @[lib.scala 374:16]
  wire [21:0] _T_2804 = _T_2472 ? btb_bank0_rd_data_way0_out_180 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3059 = _T_3058 | _T_2804; // @[Mux.scala 27:72]
  wire  _T_2474 = btb_rd_addr_f == 8'hb5; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_181; // @[lib.scala 374:16]
  wire [21:0] _T_2805 = _T_2474 ? btb_bank0_rd_data_way0_out_181 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3060 = _T_3059 | _T_2805; // @[Mux.scala 27:72]
  wire  _T_2476 = btb_rd_addr_f == 8'hb6; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_182; // @[lib.scala 374:16]
  wire [21:0] _T_2806 = _T_2476 ? btb_bank0_rd_data_way0_out_182 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3061 = _T_3060 | _T_2806; // @[Mux.scala 27:72]
  wire  _T_2478 = btb_rd_addr_f == 8'hb7; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_183; // @[lib.scala 374:16]
  wire [21:0] _T_2807 = _T_2478 ? btb_bank0_rd_data_way0_out_183 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3062 = _T_3061 | _T_2807; // @[Mux.scala 27:72]
  wire  _T_2480 = btb_rd_addr_f == 8'hb8; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_184; // @[lib.scala 374:16]
  wire [21:0] _T_2808 = _T_2480 ? btb_bank0_rd_data_way0_out_184 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3063 = _T_3062 | _T_2808; // @[Mux.scala 27:72]
  wire  _T_2482 = btb_rd_addr_f == 8'hb9; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_185; // @[lib.scala 374:16]
  wire [21:0] _T_2809 = _T_2482 ? btb_bank0_rd_data_way0_out_185 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3064 = _T_3063 | _T_2809; // @[Mux.scala 27:72]
  wire  _T_2484 = btb_rd_addr_f == 8'hba; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_186; // @[lib.scala 374:16]
  wire [21:0] _T_2810 = _T_2484 ? btb_bank0_rd_data_way0_out_186 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3065 = _T_3064 | _T_2810; // @[Mux.scala 27:72]
  wire  _T_2486 = btb_rd_addr_f == 8'hbb; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_187; // @[lib.scala 374:16]
  wire [21:0] _T_2811 = _T_2486 ? btb_bank0_rd_data_way0_out_187 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3066 = _T_3065 | _T_2811; // @[Mux.scala 27:72]
  wire  _T_2488 = btb_rd_addr_f == 8'hbc; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_188; // @[lib.scala 374:16]
  wire [21:0] _T_2812 = _T_2488 ? btb_bank0_rd_data_way0_out_188 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3067 = _T_3066 | _T_2812; // @[Mux.scala 27:72]
  wire  _T_2490 = btb_rd_addr_f == 8'hbd; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_189; // @[lib.scala 374:16]
  wire [21:0] _T_2813 = _T_2490 ? btb_bank0_rd_data_way0_out_189 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3068 = _T_3067 | _T_2813; // @[Mux.scala 27:72]
  wire  _T_2492 = btb_rd_addr_f == 8'hbe; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_190; // @[lib.scala 374:16]
  wire [21:0] _T_2814 = _T_2492 ? btb_bank0_rd_data_way0_out_190 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3069 = _T_3068 | _T_2814; // @[Mux.scala 27:72]
  wire  _T_2494 = btb_rd_addr_f == 8'hbf; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_191; // @[lib.scala 374:16]
  wire [21:0] _T_2815 = _T_2494 ? btb_bank0_rd_data_way0_out_191 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3070 = _T_3069 | _T_2815; // @[Mux.scala 27:72]
  wire  _T_2496 = btb_rd_addr_f == 8'hc0; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_192; // @[lib.scala 374:16]
  wire [21:0] _T_2816 = _T_2496 ? btb_bank0_rd_data_way0_out_192 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3071 = _T_3070 | _T_2816; // @[Mux.scala 27:72]
  wire  _T_2498 = btb_rd_addr_f == 8'hc1; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_193; // @[lib.scala 374:16]
  wire [21:0] _T_2817 = _T_2498 ? btb_bank0_rd_data_way0_out_193 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3072 = _T_3071 | _T_2817; // @[Mux.scala 27:72]
  wire  _T_2500 = btb_rd_addr_f == 8'hc2; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_194; // @[lib.scala 374:16]
  wire [21:0] _T_2818 = _T_2500 ? btb_bank0_rd_data_way0_out_194 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3073 = _T_3072 | _T_2818; // @[Mux.scala 27:72]
  wire  _T_2502 = btb_rd_addr_f == 8'hc3; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_195; // @[lib.scala 374:16]
  wire [21:0] _T_2819 = _T_2502 ? btb_bank0_rd_data_way0_out_195 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3074 = _T_3073 | _T_2819; // @[Mux.scala 27:72]
  wire  _T_2504 = btb_rd_addr_f == 8'hc4; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_196; // @[lib.scala 374:16]
  wire [21:0] _T_2820 = _T_2504 ? btb_bank0_rd_data_way0_out_196 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3075 = _T_3074 | _T_2820; // @[Mux.scala 27:72]
  wire  _T_2506 = btb_rd_addr_f == 8'hc5; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_197; // @[lib.scala 374:16]
  wire [21:0] _T_2821 = _T_2506 ? btb_bank0_rd_data_way0_out_197 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3076 = _T_3075 | _T_2821; // @[Mux.scala 27:72]
  wire  _T_2508 = btb_rd_addr_f == 8'hc6; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_198; // @[lib.scala 374:16]
  wire [21:0] _T_2822 = _T_2508 ? btb_bank0_rd_data_way0_out_198 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3077 = _T_3076 | _T_2822; // @[Mux.scala 27:72]
  wire  _T_2510 = btb_rd_addr_f == 8'hc7; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_199; // @[lib.scala 374:16]
  wire [21:0] _T_2823 = _T_2510 ? btb_bank0_rd_data_way0_out_199 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3078 = _T_3077 | _T_2823; // @[Mux.scala 27:72]
  wire  _T_2512 = btb_rd_addr_f == 8'hc8; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_200; // @[lib.scala 374:16]
  wire [21:0] _T_2824 = _T_2512 ? btb_bank0_rd_data_way0_out_200 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3079 = _T_3078 | _T_2824; // @[Mux.scala 27:72]
  wire  _T_2514 = btb_rd_addr_f == 8'hc9; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_201; // @[lib.scala 374:16]
  wire [21:0] _T_2825 = _T_2514 ? btb_bank0_rd_data_way0_out_201 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3080 = _T_3079 | _T_2825; // @[Mux.scala 27:72]
  wire  _T_2516 = btb_rd_addr_f == 8'hca; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_202; // @[lib.scala 374:16]
  wire [21:0] _T_2826 = _T_2516 ? btb_bank0_rd_data_way0_out_202 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3081 = _T_3080 | _T_2826; // @[Mux.scala 27:72]
  wire  _T_2518 = btb_rd_addr_f == 8'hcb; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_203; // @[lib.scala 374:16]
  wire [21:0] _T_2827 = _T_2518 ? btb_bank0_rd_data_way0_out_203 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3082 = _T_3081 | _T_2827; // @[Mux.scala 27:72]
  wire  _T_2520 = btb_rd_addr_f == 8'hcc; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_204; // @[lib.scala 374:16]
  wire [21:0] _T_2828 = _T_2520 ? btb_bank0_rd_data_way0_out_204 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3083 = _T_3082 | _T_2828; // @[Mux.scala 27:72]
  wire  _T_2522 = btb_rd_addr_f == 8'hcd; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_205; // @[lib.scala 374:16]
  wire [21:0] _T_2829 = _T_2522 ? btb_bank0_rd_data_way0_out_205 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3084 = _T_3083 | _T_2829; // @[Mux.scala 27:72]
  wire  _T_2524 = btb_rd_addr_f == 8'hce; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_206; // @[lib.scala 374:16]
  wire [21:0] _T_2830 = _T_2524 ? btb_bank0_rd_data_way0_out_206 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3085 = _T_3084 | _T_2830; // @[Mux.scala 27:72]
  wire  _T_2526 = btb_rd_addr_f == 8'hcf; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_207; // @[lib.scala 374:16]
  wire [21:0] _T_2831 = _T_2526 ? btb_bank0_rd_data_way0_out_207 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3086 = _T_3085 | _T_2831; // @[Mux.scala 27:72]
  wire  _T_2528 = btb_rd_addr_f == 8'hd0; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_208; // @[lib.scala 374:16]
  wire [21:0] _T_2832 = _T_2528 ? btb_bank0_rd_data_way0_out_208 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3087 = _T_3086 | _T_2832; // @[Mux.scala 27:72]
  wire  _T_2530 = btb_rd_addr_f == 8'hd1; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_209; // @[lib.scala 374:16]
  wire [21:0] _T_2833 = _T_2530 ? btb_bank0_rd_data_way0_out_209 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3088 = _T_3087 | _T_2833; // @[Mux.scala 27:72]
  wire  _T_2532 = btb_rd_addr_f == 8'hd2; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_210; // @[lib.scala 374:16]
  wire [21:0] _T_2834 = _T_2532 ? btb_bank0_rd_data_way0_out_210 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3089 = _T_3088 | _T_2834; // @[Mux.scala 27:72]
  wire  _T_2534 = btb_rd_addr_f == 8'hd3; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_211; // @[lib.scala 374:16]
  wire [21:0] _T_2835 = _T_2534 ? btb_bank0_rd_data_way0_out_211 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3090 = _T_3089 | _T_2835; // @[Mux.scala 27:72]
  wire  _T_2536 = btb_rd_addr_f == 8'hd4; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_212; // @[lib.scala 374:16]
  wire [21:0] _T_2836 = _T_2536 ? btb_bank0_rd_data_way0_out_212 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3091 = _T_3090 | _T_2836; // @[Mux.scala 27:72]
  wire  _T_2538 = btb_rd_addr_f == 8'hd5; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_213; // @[lib.scala 374:16]
  wire [21:0] _T_2837 = _T_2538 ? btb_bank0_rd_data_way0_out_213 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3092 = _T_3091 | _T_2837; // @[Mux.scala 27:72]
  wire  _T_2540 = btb_rd_addr_f == 8'hd6; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_214; // @[lib.scala 374:16]
  wire [21:0] _T_2838 = _T_2540 ? btb_bank0_rd_data_way0_out_214 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3093 = _T_3092 | _T_2838; // @[Mux.scala 27:72]
  wire  _T_2542 = btb_rd_addr_f == 8'hd7; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_215; // @[lib.scala 374:16]
  wire [21:0] _T_2839 = _T_2542 ? btb_bank0_rd_data_way0_out_215 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3094 = _T_3093 | _T_2839; // @[Mux.scala 27:72]
  wire  _T_2544 = btb_rd_addr_f == 8'hd8; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_216; // @[lib.scala 374:16]
  wire [21:0] _T_2840 = _T_2544 ? btb_bank0_rd_data_way0_out_216 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3095 = _T_3094 | _T_2840; // @[Mux.scala 27:72]
  wire  _T_2546 = btb_rd_addr_f == 8'hd9; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_217; // @[lib.scala 374:16]
  wire [21:0] _T_2841 = _T_2546 ? btb_bank0_rd_data_way0_out_217 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3096 = _T_3095 | _T_2841; // @[Mux.scala 27:72]
  wire  _T_2548 = btb_rd_addr_f == 8'hda; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_218; // @[lib.scala 374:16]
  wire [21:0] _T_2842 = _T_2548 ? btb_bank0_rd_data_way0_out_218 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3097 = _T_3096 | _T_2842; // @[Mux.scala 27:72]
  wire  _T_2550 = btb_rd_addr_f == 8'hdb; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_219; // @[lib.scala 374:16]
  wire [21:0] _T_2843 = _T_2550 ? btb_bank0_rd_data_way0_out_219 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3098 = _T_3097 | _T_2843; // @[Mux.scala 27:72]
  wire  _T_2552 = btb_rd_addr_f == 8'hdc; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_220; // @[lib.scala 374:16]
  wire [21:0] _T_2844 = _T_2552 ? btb_bank0_rd_data_way0_out_220 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3099 = _T_3098 | _T_2844; // @[Mux.scala 27:72]
  wire  _T_2554 = btb_rd_addr_f == 8'hdd; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_221; // @[lib.scala 374:16]
  wire [21:0] _T_2845 = _T_2554 ? btb_bank0_rd_data_way0_out_221 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3100 = _T_3099 | _T_2845; // @[Mux.scala 27:72]
  wire  _T_2556 = btb_rd_addr_f == 8'hde; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_222; // @[lib.scala 374:16]
  wire [21:0] _T_2846 = _T_2556 ? btb_bank0_rd_data_way0_out_222 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3101 = _T_3100 | _T_2846; // @[Mux.scala 27:72]
  wire  _T_2558 = btb_rd_addr_f == 8'hdf; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_223; // @[lib.scala 374:16]
  wire [21:0] _T_2847 = _T_2558 ? btb_bank0_rd_data_way0_out_223 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3102 = _T_3101 | _T_2847; // @[Mux.scala 27:72]
  wire  _T_2560 = btb_rd_addr_f == 8'he0; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_224; // @[lib.scala 374:16]
  wire [21:0] _T_2848 = _T_2560 ? btb_bank0_rd_data_way0_out_224 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3103 = _T_3102 | _T_2848; // @[Mux.scala 27:72]
  wire  _T_2562 = btb_rd_addr_f == 8'he1; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_225; // @[lib.scala 374:16]
  wire [21:0] _T_2849 = _T_2562 ? btb_bank0_rd_data_way0_out_225 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3104 = _T_3103 | _T_2849; // @[Mux.scala 27:72]
  wire  _T_2564 = btb_rd_addr_f == 8'he2; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_226; // @[lib.scala 374:16]
  wire [21:0] _T_2850 = _T_2564 ? btb_bank0_rd_data_way0_out_226 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3105 = _T_3104 | _T_2850; // @[Mux.scala 27:72]
  wire  _T_2566 = btb_rd_addr_f == 8'he3; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_227; // @[lib.scala 374:16]
  wire [21:0] _T_2851 = _T_2566 ? btb_bank0_rd_data_way0_out_227 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3106 = _T_3105 | _T_2851; // @[Mux.scala 27:72]
  wire  _T_2568 = btb_rd_addr_f == 8'he4; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_228; // @[lib.scala 374:16]
  wire [21:0] _T_2852 = _T_2568 ? btb_bank0_rd_data_way0_out_228 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3107 = _T_3106 | _T_2852; // @[Mux.scala 27:72]
  wire  _T_2570 = btb_rd_addr_f == 8'he5; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_229; // @[lib.scala 374:16]
  wire [21:0] _T_2853 = _T_2570 ? btb_bank0_rd_data_way0_out_229 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3108 = _T_3107 | _T_2853; // @[Mux.scala 27:72]
  wire  _T_2572 = btb_rd_addr_f == 8'he6; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_230; // @[lib.scala 374:16]
  wire [21:0] _T_2854 = _T_2572 ? btb_bank0_rd_data_way0_out_230 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3109 = _T_3108 | _T_2854; // @[Mux.scala 27:72]
  wire  _T_2574 = btb_rd_addr_f == 8'he7; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_231; // @[lib.scala 374:16]
  wire [21:0] _T_2855 = _T_2574 ? btb_bank0_rd_data_way0_out_231 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3110 = _T_3109 | _T_2855; // @[Mux.scala 27:72]
  wire  _T_2576 = btb_rd_addr_f == 8'he8; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_232; // @[lib.scala 374:16]
  wire [21:0] _T_2856 = _T_2576 ? btb_bank0_rd_data_way0_out_232 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3111 = _T_3110 | _T_2856; // @[Mux.scala 27:72]
  wire  _T_2578 = btb_rd_addr_f == 8'he9; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_233; // @[lib.scala 374:16]
  wire [21:0] _T_2857 = _T_2578 ? btb_bank0_rd_data_way0_out_233 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3112 = _T_3111 | _T_2857; // @[Mux.scala 27:72]
  wire  _T_2580 = btb_rd_addr_f == 8'hea; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_234; // @[lib.scala 374:16]
  wire [21:0] _T_2858 = _T_2580 ? btb_bank0_rd_data_way0_out_234 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3113 = _T_3112 | _T_2858; // @[Mux.scala 27:72]
  wire  _T_2582 = btb_rd_addr_f == 8'heb; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_235; // @[lib.scala 374:16]
  wire [21:0] _T_2859 = _T_2582 ? btb_bank0_rd_data_way0_out_235 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3114 = _T_3113 | _T_2859; // @[Mux.scala 27:72]
  wire  _T_2584 = btb_rd_addr_f == 8'hec; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_236; // @[lib.scala 374:16]
  wire [21:0] _T_2860 = _T_2584 ? btb_bank0_rd_data_way0_out_236 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3115 = _T_3114 | _T_2860; // @[Mux.scala 27:72]
  wire  _T_2586 = btb_rd_addr_f == 8'hed; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_237; // @[lib.scala 374:16]
  wire [21:0] _T_2861 = _T_2586 ? btb_bank0_rd_data_way0_out_237 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3116 = _T_3115 | _T_2861; // @[Mux.scala 27:72]
  wire  _T_2588 = btb_rd_addr_f == 8'hee; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_238; // @[lib.scala 374:16]
  wire [21:0] _T_2862 = _T_2588 ? btb_bank0_rd_data_way0_out_238 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3117 = _T_3116 | _T_2862; // @[Mux.scala 27:72]
  wire  _T_2590 = btb_rd_addr_f == 8'hef; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_239; // @[lib.scala 374:16]
  wire [21:0] _T_2863 = _T_2590 ? btb_bank0_rd_data_way0_out_239 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3118 = _T_3117 | _T_2863; // @[Mux.scala 27:72]
  wire  _T_2592 = btb_rd_addr_f == 8'hf0; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_240; // @[lib.scala 374:16]
  wire [21:0] _T_2864 = _T_2592 ? btb_bank0_rd_data_way0_out_240 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3119 = _T_3118 | _T_2864; // @[Mux.scala 27:72]
  wire  _T_2594 = btb_rd_addr_f == 8'hf1; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_241; // @[lib.scala 374:16]
  wire [21:0] _T_2865 = _T_2594 ? btb_bank0_rd_data_way0_out_241 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3120 = _T_3119 | _T_2865; // @[Mux.scala 27:72]
  wire  _T_2596 = btb_rd_addr_f == 8'hf2; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_242; // @[lib.scala 374:16]
  wire [21:0] _T_2866 = _T_2596 ? btb_bank0_rd_data_way0_out_242 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3121 = _T_3120 | _T_2866; // @[Mux.scala 27:72]
  wire  _T_2598 = btb_rd_addr_f == 8'hf3; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_243; // @[lib.scala 374:16]
  wire [21:0] _T_2867 = _T_2598 ? btb_bank0_rd_data_way0_out_243 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3122 = _T_3121 | _T_2867; // @[Mux.scala 27:72]
  wire  _T_2600 = btb_rd_addr_f == 8'hf4; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_244; // @[lib.scala 374:16]
  wire [21:0] _T_2868 = _T_2600 ? btb_bank0_rd_data_way0_out_244 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3123 = _T_3122 | _T_2868; // @[Mux.scala 27:72]
  wire  _T_2602 = btb_rd_addr_f == 8'hf5; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_245; // @[lib.scala 374:16]
  wire [21:0] _T_2869 = _T_2602 ? btb_bank0_rd_data_way0_out_245 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3124 = _T_3123 | _T_2869; // @[Mux.scala 27:72]
  wire  _T_2604 = btb_rd_addr_f == 8'hf6; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_246; // @[lib.scala 374:16]
  wire [21:0] _T_2870 = _T_2604 ? btb_bank0_rd_data_way0_out_246 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3125 = _T_3124 | _T_2870; // @[Mux.scala 27:72]
  wire  _T_2606 = btb_rd_addr_f == 8'hf7; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_247; // @[lib.scala 374:16]
  wire [21:0] _T_2871 = _T_2606 ? btb_bank0_rd_data_way0_out_247 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3126 = _T_3125 | _T_2871; // @[Mux.scala 27:72]
  wire  _T_2608 = btb_rd_addr_f == 8'hf8; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_248; // @[lib.scala 374:16]
  wire [21:0] _T_2872 = _T_2608 ? btb_bank0_rd_data_way0_out_248 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3127 = _T_3126 | _T_2872; // @[Mux.scala 27:72]
  wire  _T_2610 = btb_rd_addr_f == 8'hf9; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_249; // @[lib.scala 374:16]
  wire [21:0] _T_2873 = _T_2610 ? btb_bank0_rd_data_way0_out_249 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3128 = _T_3127 | _T_2873; // @[Mux.scala 27:72]
  wire  _T_2612 = btb_rd_addr_f == 8'hfa; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_250; // @[lib.scala 374:16]
  wire [21:0] _T_2874 = _T_2612 ? btb_bank0_rd_data_way0_out_250 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3129 = _T_3128 | _T_2874; // @[Mux.scala 27:72]
  wire  _T_2614 = btb_rd_addr_f == 8'hfb; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_251; // @[lib.scala 374:16]
  wire [21:0] _T_2875 = _T_2614 ? btb_bank0_rd_data_way0_out_251 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3130 = _T_3129 | _T_2875; // @[Mux.scala 27:72]
  wire  _T_2616 = btb_rd_addr_f == 8'hfc; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_252; // @[lib.scala 374:16]
  wire [21:0] _T_2876 = _T_2616 ? btb_bank0_rd_data_way0_out_252 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3131 = _T_3130 | _T_2876; // @[Mux.scala 27:72]
  wire  _T_2618 = btb_rd_addr_f == 8'hfd; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_253; // @[lib.scala 374:16]
  wire [21:0] _T_2877 = _T_2618 ? btb_bank0_rd_data_way0_out_253 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3132 = _T_3131 | _T_2877; // @[Mux.scala 27:72]
  wire  _T_2620 = btb_rd_addr_f == 8'hfe; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_254; // @[lib.scala 374:16]
  wire [21:0] _T_2878 = _T_2620 ? btb_bank0_rd_data_way0_out_254 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3133 = _T_3132 | _T_2878; // @[Mux.scala 27:72]
  wire  _T_2622 = btb_rd_addr_f == 8'hff; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_255; // @[lib.scala 374:16]
  wire [21:0] _T_2879 = _T_2622 ? btb_bank0_rd_data_way0_out_255 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] btb_bank0_rd_data_way0_f = _T_3133 | _T_2879; // @[Mux.scala 27:72]
  wire [4:0] _T_25 = io_ifc_fetch_addr_f[13:9] ^ io_ifc_fetch_addr_f[18:14]; // @[lib.scala 42:111]
  wire [4:0] fetch_rd_tag_f = _T_25 ^ io_ifc_fetch_addr_f[23:19]; // @[lib.scala 42:111]
  wire  _T_46 = btb_bank0_rd_data_way0_f[21:17] == fetch_rd_tag_f; // @[ifu_bp_ctl.scala 127:97]
  wire  _T_47 = btb_bank0_rd_data_way0_f[0] & _T_46; // @[ifu_bp_ctl.scala 127:55]
  reg  dec_tlu_way_wb_f; // @[ifu_bp_ctl.scala 118:59]
  wire  _T_19 = io_exu_bp_exu_i0_br_index_r == btb_rd_addr_f; // @[ifu_bp_ctl.scala 102:72]
  wire  branch_error_collision_f = dec_tlu_error_wb & _T_19; // @[ifu_bp_ctl.scala 102:51]
  wire  branch_error_bank_conflict_f = branch_error_collision_f & dec_tlu_error_wb; // @[ifu_bp_ctl.scala 106:63]
  wire  _T_48 = dec_tlu_way_wb_f & branch_error_bank_conflict_f; // @[ifu_bp_ctl.scala 128:44]
  wire  _T_49 = ~_T_48; // @[ifu_bp_ctl.scala 128:25]
  wire  _T_50 = _T_47 & _T_49; // @[ifu_bp_ctl.scala 127:117]
  wire  _T_51 = _T_50 & io_ifc_fetch_req_f; // @[ifu_bp_ctl.scala 128:76]
  wire  tag_match_way0_f = _T_51 & _T; // @[ifu_bp_ctl.scala 128:97]
  wire  _T_82 = btb_bank0_rd_data_way0_f[3] ^ btb_bank0_rd_data_way0_f[4]; // @[ifu_bp_ctl.scala 142:91]
  wire  _T_83 = tag_match_way0_f & _T_82; // @[ifu_bp_ctl.scala 142:56]
  wire  _T_87 = ~_T_82; // @[ifu_bp_ctl.scala 143:58]
  wire  _T_88 = tag_match_way0_f & _T_87; // @[ifu_bp_ctl.scala 143:56]
  wire [1:0] tag_match_way0_expanded_f = {_T_83,_T_88}; // @[Cat.scala 29:58]
  wire [21:0] _T_127 = tag_match_way0_expanded_f[1] ? btb_bank0_rd_data_way0_f : 22'h0; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_0; // @[lib.scala 374:16]
  wire [21:0] _T_3648 = _T_2112 ? btb_bank0_rd_data_way1_out_0 : 22'h0; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_1; // @[lib.scala 374:16]
  wire [21:0] _T_3649 = _T_2114 ? btb_bank0_rd_data_way1_out_1 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3904 = _T_3648 | _T_3649; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_2; // @[lib.scala 374:16]
  wire [21:0] _T_3650 = _T_2116 ? btb_bank0_rd_data_way1_out_2 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3905 = _T_3904 | _T_3650; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_3; // @[lib.scala 374:16]
  wire [21:0] _T_3651 = _T_2118 ? btb_bank0_rd_data_way1_out_3 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3906 = _T_3905 | _T_3651; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_4; // @[lib.scala 374:16]
  wire [21:0] _T_3652 = _T_2120 ? btb_bank0_rd_data_way1_out_4 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3907 = _T_3906 | _T_3652; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_5; // @[lib.scala 374:16]
  wire [21:0] _T_3653 = _T_2122 ? btb_bank0_rd_data_way1_out_5 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3908 = _T_3907 | _T_3653; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_6; // @[lib.scala 374:16]
  wire [21:0] _T_3654 = _T_2124 ? btb_bank0_rd_data_way1_out_6 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3909 = _T_3908 | _T_3654; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_7; // @[lib.scala 374:16]
  wire [21:0] _T_3655 = _T_2126 ? btb_bank0_rd_data_way1_out_7 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3910 = _T_3909 | _T_3655; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_8; // @[lib.scala 374:16]
  wire [21:0] _T_3656 = _T_2128 ? btb_bank0_rd_data_way1_out_8 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3911 = _T_3910 | _T_3656; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_9; // @[lib.scala 374:16]
  wire [21:0] _T_3657 = _T_2130 ? btb_bank0_rd_data_way1_out_9 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3912 = _T_3911 | _T_3657; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_10; // @[lib.scala 374:16]
  wire [21:0] _T_3658 = _T_2132 ? btb_bank0_rd_data_way1_out_10 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3913 = _T_3912 | _T_3658; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_11; // @[lib.scala 374:16]
  wire [21:0] _T_3659 = _T_2134 ? btb_bank0_rd_data_way1_out_11 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3914 = _T_3913 | _T_3659; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_12; // @[lib.scala 374:16]
  wire [21:0] _T_3660 = _T_2136 ? btb_bank0_rd_data_way1_out_12 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3915 = _T_3914 | _T_3660; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_13; // @[lib.scala 374:16]
  wire [21:0] _T_3661 = _T_2138 ? btb_bank0_rd_data_way1_out_13 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3916 = _T_3915 | _T_3661; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_14; // @[lib.scala 374:16]
  wire [21:0] _T_3662 = _T_2140 ? btb_bank0_rd_data_way1_out_14 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3917 = _T_3916 | _T_3662; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_15; // @[lib.scala 374:16]
  wire [21:0] _T_3663 = _T_2142 ? btb_bank0_rd_data_way1_out_15 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3918 = _T_3917 | _T_3663; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_16; // @[lib.scala 374:16]
  wire [21:0] _T_3664 = _T_2144 ? btb_bank0_rd_data_way1_out_16 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3919 = _T_3918 | _T_3664; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_17; // @[lib.scala 374:16]
  wire [21:0] _T_3665 = _T_2146 ? btb_bank0_rd_data_way1_out_17 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3920 = _T_3919 | _T_3665; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_18; // @[lib.scala 374:16]
  wire [21:0] _T_3666 = _T_2148 ? btb_bank0_rd_data_way1_out_18 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3921 = _T_3920 | _T_3666; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_19; // @[lib.scala 374:16]
  wire [21:0] _T_3667 = _T_2150 ? btb_bank0_rd_data_way1_out_19 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3922 = _T_3921 | _T_3667; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_20; // @[lib.scala 374:16]
  wire [21:0] _T_3668 = _T_2152 ? btb_bank0_rd_data_way1_out_20 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3923 = _T_3922 | _T_3668; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_21; // @[lib.scala 374:16]
  wire [21:0] _T_3669 = _T_2154 ? btb_bank0_rd_data_way1_out_21 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3924 = _T_3923 | _T_3669; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_22; // @[lib.scala 374:16]
  wire [21:0] _T_3670 = _T_2156 ? btb_bank0_rd_data_way1_out_22 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3925 = _T_3924 | _T_3670; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_23; // @[lib.scala 374:16]
  wire [21:0] _T_3671 = _T_2158 ? btb_bank0_rd_data_way1_out_23 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3926 = _T_3925 | _T_3671; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_24; // @[lib.scala 374:16]
  wire [21:0] _T_3672 = _T_2160 ? btb_bank0_rd_data_way1_out_24 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3927 = _T_3926 | _T_3672; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_25; // @[lib.scala 374:16]
  wire [21:0] _T_3673 = _T_2162 ? btb_bank0_rd_data_way1_out_25 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3928 = _T_3927 | _T_3673; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_26; // @[lib.scala 374:16]
  wire [21:0] _T_3674 = _T_2164 ? btb_bank0_rd_data_way1_out_26 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3929 = _T_3928 | _T_3674; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_27; // @[lib.scala 374:16]
  wire [21:0] _T_3675 = _T_2166 ? btb_bank0_rd_data_way1_out_27 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3930 = _T_3929 | _T_3675; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_28; // @[lib.scala 374:16]
  wire [21:0] _T_3676 = _T_2168 ? btb_bank0_rd_data_way1_out_28 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3931 = _T_3930 | _T_3676; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_29; // @[lib.scala 374:16]
  wire [21:0] _T_3677 = _T_2170 ? btb_bank0_rd_data_way1_out_29 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3932 = _T_3931 | _T_3677; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_30; // @[lib.scala 374:16]
  wire [21:0] _T_3678 = _T_2172 ? btb_bank0_rd_data_way1_out_30 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3933 = _T_3932 | _T_3678; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_31; // @[lib.scala 374:16]
  wire [21:0] _T_3679 = _T_2174 ? btb_bank0_rd_data_way1_out_31 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3934 = _T_3933 | _T_3679; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_32; // @[lib.scala 374:16]
  wire [21:0] _T_3680 = _T_2176 ? btb_bank0_rd_data_way1_out_32 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3935 = _T_3934 | _T_3680; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_33; // @[lib.scala 374:16]
  wire [21:0] _T_3681 = _T_2178 ? btb_bank0_rd_data_way1_out_33 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3936 = _T_3935 | _T_3681; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_34; // @[lib.scala 374:16]
  wire [21:0] _T_3682 = _T_2180 ? btb_bank0_rd_data_way1_out_34 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3937 = _T_3936 | _T_3682; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_35; // @[lib.scala 374:16]
  wire [21:0] _T_3683 = _T_2182 ? btb_bank0_rd_data_way1_out_35 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3938 = _T_3937 | _T_3683; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_36; // @[lib.scala 374:16]
  wire [21:0] _T_3684 = _T_2184 ? btb_bank0_rd_data_way1_out_36 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3939 = _T_3938 | _T_3684; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_37; // @[lib.scala 374:16]
  wire [21:0] _T_3685 = _T_2186 ? btb_bank0_rd_data_way1_out_37 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3940 = _T_3939 | _T_3685; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_38; // @[lib.scala 374:16]
  wire [21:0] _T_3686 = _T_2188 ? btb_bank0_rd_data_way1_out_38 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3941 = _T_3940 | _T_3686; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_39; // @[lib.scala 374:16]
  wire [21:0] _T_3687 = _T_2190 ? btb_bank0_rd_data_way1_out_39 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3942 = _T_3941 | _T_3687; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_40; // @[lib.scala 374:16]
  wire [21:0] _T_3688 = _T_2192 ? btb_bank0_rd_data_way1_out_40 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3943 = _T_3942 | _T_3688; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_41; // @[lib.scala 374:16]
  wire [21:0] _T_3689 = _T_2194 ? btb_bank0_rd_data_way1_out_41 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3944 = _T_3943 | _T_3689; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_42; // @[lib.scala 374:16]
  wire [21:0] _T_3690 = _T_2196 ? btb_bank0_rd_data_way1_out_42 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3945 = _T_3944 | _T_3690; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_43; // @[lib.scala 374:16]
  wire [21:0] _T_3691 = _T_2198 ? btb_bank0_rd_data_way1_out_43 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3946 = _T_3945 | _T_3691; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_44; // @[lib.scala 374:16]
  wire [21:0] _T_3692 = _T_2200 ? btb_bank0_rd_data_way1_out_44 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3947 = _T_3946 | _T_3692; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_45; // @[lib.scala 374:16]
  wire [21:0] _T_3693 = _T_2202 ? btb_bank0_rd_data_way1_out_45 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3948 = _T_3947 | _T_3693; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_46; // @[lib.scala 374:16]
  wire [21:0] _T_3694 = _T_2204 ? btb_bank0_rd_data_way1_out_46 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3949 = _T_3948 | _T_3694; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_47; // @[lib.scala 374:16]
  wire [21:0] _T_3695 = _T_2206 ? btb_bank0_rd_data_way1_out_47 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3950 = _T_3949 | _T_3695; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_48; // @[lib.scala 374:16]
  wire [21:0] _T_3696 = _T_2208 ? btb_bank0_rd_data_way1_out_48 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3951 = _T_3950 | _T_3696; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_49; // @[lib.scala 374:16]
  wire [21:0] _T_3697 = _T_2210 ? btb_bank0_rd_data_way1_out_49 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3952 = _T_3951 | _T_3697; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_50; // @[lib.scala 374:16]
  wire [21:0] _T_3698 = _T_2212 ? btb_bank0_rd_data_way1_out_50 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3953 = _T_3952 | _T_3698; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_51; // @[lib.scala 374:16]
  wire [21:0] _T_3699 = _T_2214 ? btb_bank0_rd_data_way1_out_51 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3954 = _T_3953 | _T_3699; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_52; // @[lib.scala 374:16]
  wire [21:0] _T_3700 = _T_2216 ? btb_bank0_rd_data_way1_out_52 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3955 = _T_3954 | _T_3700; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_53; // @[lib.scala 374:16]
  wire [21:0] _T_3701 = _T_2218 ? btb_bank0_rd_data_way1_out_53 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3956 = _T_3955 | _T_3701; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_54; // @[lib.scala 374:16]
  wire [21:0] _T_3702 = _T_2220 ? btb_bank0_rd_data_way1_out_54 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3957 = _T_3956 | _T_3702; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_55; // @[lib.scala 374:16]
  wire [21:0] _T_3703 = _T_2222 ? btb_bank0_rd_data_way1_out_55 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3958 = _T_3957 | _T_3703; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_56; // @[lib.scala 374:16]
  wire [21:0] _T_3704 = _T_2224 ? btb_bank0_rd_data_way1_out_56 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3959 = _T_3958 | _T_3704; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_57; // @[lib.scala 374:16]
  wire [21:0] _T_3705 = _T_2226 ? btb_bank0_rd_data_way1_out_57 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3960 = _T_3959 | _T_3705; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_58; // @[lib.scala 374:16]
  wire [21:0] _T_3706 = _T_2228 ? btb_bank0_rd_data_way1_out_58 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3961 = _T_3960 | _T_3706; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_59; // @[lib.scala 374:16]
  wire [21:0] _T_3707 = _T_2230 ? btb_bank0_rd_data_way1_out_59 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3962 = _T_3961 | _T_3707; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_60; // @[lib.scala 374:16]
  wire [21:0] _T_3708 = _T_2232 ? btb_bank0_rd_data_way1_out_60 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3963 = _T_3962 | _T_3708; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_61; // @[lib.scala 374:16]
  wire [21:0] _T_3709 = _T_2234 ? btb_bank0_rd_data_way1_out_61 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3964 = _T_3963 | _T_3709; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_62; // @[lib.scala 374:16]
  wire [21:0] _T_3710 = _T_2236 ? btb_bank0_rd_data_way1_out_62 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3965 = _T_3964 | _T_3710; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_63; // @[lib.scala 374:16]
  wire [21:0] _T_3711 = _T_2238 ? btb_bank0_rd_data_way1_out_63 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3966 = _T_3965 | _T_3711; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_64; // @[lib.scala 374:16]
  wire [21:0] _T_3712 = _T_2240 ? btb_bank0_rd_data_way1_out_64 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3967 = _T_3966 | _T_3712; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_65; // @[lib.scala 374:16]
  wire [21:0] _T_3713 = _T_2242 ? btb_bank0_rd_data_way1_out_65 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3968 = _T_3967 | _T_3713; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_66; // @[lib.scala 374:16]
  wire [21:0] _T_3714 = _T_2244 ? btb_bank0_rd_data_way1_out_66 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3969 = _T_3968 | _T_3714; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_67; // @[lib.scala 374:16]
  wire [21:0] _T_3715 = _T_2246 ? btb_bank0_rd_data_way1_out_67 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3970 = _T_3969 | _T_3715; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_68; // @[lib.scala 374:16]
  wire [21:0] _T_3716 = _T_2248 ? btb_bank0_rd_data_way1_out_68 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3971 = _T_3970 | _T_3716; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_69; // @[lib.scala 374:16]
  wire [21:0] _T_3717 = _T_2250 ? btb_bank0_rd_data_way1_out_69 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3972 = _T_3971 | _T_3717; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_70; // @[lib.scala 374:16]
  wire [21:0] _T_3718 = _T_2252 ? btb_bank0_rd_data_way1_out_70 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3973 = _T_3972 | _T_3718; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_71; // @[lib.scala 374:16]
  wire [21:0] _T_3719 = _T_2254 ? btb_bank0_rd_data_way1_out_71 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3974 = _T_3973 | _T_3719; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_72; // @[lib.scala 374:16]
  wire [21:0] _T_3720 = _T_2256 ? btb_bank0_rd_data_way1_out_72 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3975 = _T_3974 | _T_3720; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_73; // @[lib.scala 374:16]
  wire [21:0] _T_3721 = _T_2258 ? btb_bank0_rd_data_way1_out_73 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3976 = _T_3975 | _T_3721; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_74; // @[lib.scala 374:16]
  wire [21:0] _T_3722 = _T_2260 ? btb_bank0_rd_data_way1_out_74 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3977 = _T_3976 | _T_3722; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_75; // @[lib.scala 374:16]
  wire [21:0] _T_3723 = _T_2262 ? btb_bank0_rd_data_way1_out_75 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3978 = _T_3977 | _T_3723; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_76; // @[lib.scala 374:16]
  wire [21:0] _T_3724 = _T_2264 ? btb_bank0_rd_data_way1_out_76 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3979 = _T_3978 | _T_3724; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_77; // @[lib.scala 374:16]
  wire [21:0] _T_3725 = _T_2266 ? btb_bank0_rd_data_way1_out_77 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3980 = _T_3979 | _T_3725; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_78; // @[lib.scala 374:16]
  wire [21:0] _T_3726 = _T_2268 ? btb_bank0_rd_data_way1_out_78 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3981 = _T_3980 | _T_3726; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_79; // @[lib.scala 374:16]
  wire [21:0] _T_3727 = _T_2270 ? btb_bank0_rd_data_way1_out_79 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3982 = _T_3981 | _T_3727; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_80; // @[lib.scala 374:16]
  wire [21:0] _T_3728 = _T_2272 ? btb_bank0_rd_data_way1_out_80 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3983 = _T_3982 | _T_3728; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_81; // @[lib.scala 374:16]
  wire [21:0] _T_3729 = _T_2274 ? btb_bank0_rd_data_way1_out_81 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3984 = _T_3983 | _T_3729; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_82; // @[lib.scala 374:16]
  wire [21:0] _T_3730 = _T_2276 ? btb_bank0_rd_data_way1_out_82 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3985 = _T_3984 | _T_3730; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_83; // @[lib.scala 374:16]
  wire [21:0] _T_3731 = _T_2278 ? btb_bank0_rd_data_way1_out_83 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3986 = _T_3985 | _T_3731; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_84; // @[lib.scala 374:16]
  wire [21:0] _T_3732 = _T_2280 ? btb_bank0_rd_data_way1_out_84 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3987 = _T_3986 | _T_3732; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_85; // @[lib.scala 374:16]
  wire [21:0] _T_3733 = _T_2282 ? btb_bank0_rd_data_way1_out_85 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3988 = _T_3987 | _T_3733; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_86; // @[lib.scala 374:16]
  wire [21:0] _T_3734 = _T_2284 ? btb_bank0_rd_data_way1_out_86 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3989 = _T_3988 | _T_3734; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_87; // @[lib.scala 374:16]
  wire [21:0] _T_3735 = _T_2286 ? btb_bank0_rd_data_way1_out_87 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3990 = _T_3989 | _T_3735; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_88; // @[lib.scala 374:16]
  wire [21:0] _T_3736 = _T_2288 ? btb_bank0_rd_data_way1_out_88 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3991 = _T_3990 | _T_3736; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_89; // @[lib.scala 374:16]
  wire [21:0] _T_3737 = _T_2290 ? btb_bank0_rd_data_way1_out_89 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3992 = _T_3991 | _T_3737; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_90; // @[lib.scala 374:16]
  wire [21:0] _T_3738 = _T_2292 ? btb_bank0_rd_data_way1_out_90 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3993 = _T_3992 | _T_3738; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_91; // @[lib.scala 374:16]
  wire [21:0] _T_3739 = _T_2294 ? btb_bank0_rd_data_way1_out_91 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3994 = _T_3993 | _T_3739; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_92; // @[lib.scala 374:16]
  wire [21:0] _T_3740 = _T_2296 ? btb_bank0_rd_data_way1_out_92 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3995 = _T_3994 | _T_3740; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_93; // @[lib.scala 374:16]
  wire [21:0] _T_3741 = _T_2298 ? btb_bank0_rd_data_way1_out_93 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3996 = _T_3995 | _T_3741; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_94; // @[lib.scala 374:16]
  wire [21:0] _T_3742 = _T_2300 ? btb_bank0_rd_data_way1_out_94 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3997 = _T_3996 | _T_3742; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_95; // @[lib.scala 374:16]
  wire [21:0] _T_3743 = _T_2302 ? btb_bank0_rd_data_way1_out_95 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3998 = _T_3997 | _T_3743; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_96; // @[lib.scala 374:16]
  wire [21:0] _T_3744 = _T_2304 ? btb_bank0_rd_data_way1_out_96 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3999 = _T_3998 | _T_3744; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_97; // @[lib.scala 374:16]
  wire [21:0] _T_3745 = _T_2306 ? btb_bank0_rd_data_way1_out_97 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4000 = _T_3999 | _T_3745; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_98; // @[lib.scala 374:16]
  wire [21:0] _T_3746 = _T_2308 ? btb_bank0_rd_data_way1_out_98 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4001 = _T_4000 | _T_3746; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_99; // @[lib.scala 374:16]
  wire [21:0] _T_3747 = _T_2310 ? btb_bank0_rd_data_way1_out_99 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4002 = _T_4001 | _T_3747; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_100; // @[lib.scala 374:16]
  wire [21:0] _T_3748 = _T_2312 ? btb_bank0_rd_data_way1_out_100 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4003 = _T_4002 | _T_3748; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_101; // @[lib.scala 374:16]
  wire [21:0] _T_3749 = _T_2314 ? btb_bank0_rd_data_way1_out_101 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4004 = _T_4003 | _T_3749; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_102; // @[lib.scala 374:16]
  wire [21:0] _T_3750 = _T_2316 ? btb_bank0_rd_data_way1_out_102 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4005 = _T_4004 | _T_3750; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_103; // @[lib.scala 374:16]
  wire [21:0] _T_3751 = _T_2318 ? btb_bank0_rd_data_way1_out_103 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4006 = _T_4005 | _T_3751; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_104; // @[lib.scala 374:16]
  wire [21:0] _T_3752 = _T_2320 ? btb_bank0_rd_data_way1_out_104 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4007 = _T_4006 | _T_3752; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_105; // @[lib.scala 374:16]
  wire [21:0] _T_3753 = _T_2322 ? btb_bank0_rd_data_way1_out_105 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4008 = _T_4007 | _T_3753; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_106; // @[lib.scala 374:16]
  wire [21:0] _T_3754 = _T_2324 ? btb_bank0_rd_data_way1_out_106 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4009 = _T_4008 | _T_3754; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_107; // @[lib.scala 374:16]
  wire [21:0] _T_3755 = _T_2326 ? btb_bank0_rd_data_way1_out_107 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4010 = _T_4009 | _T_3755; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_108; // @[lib.scala 374:16]
  wire [21:0] _T_3756 = _T_2328 ? btb_bank0_rd_data_way1_out_108 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4011 = _T_4010 | _T_3756; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_109; // @[lib.scala 374:16]
  wire [21:0] _T_3757 = _T_2330 ? btb_bank0_rd_data_way1_out_109 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4012 = _T_4011 | _T_3757; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_110; // @[lib.scala 374:16]
  wire [21:0] _T_3758 = _T_2332 ? btb_bank0_rd_data_way1_out_110 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4013 = _T_4012 | _T_3758; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_111; // @[lib.scala 374:16]
  wire [21:0] _T_3759 = _T_2334 ? btb_bank0_rd_data_way1_out_111 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4014 = _T_4013 | _T_3759; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_112; // @[lib.scala 374:16]
  wire [21:0] _T_3760 = _T_2336 ? btb_bank0_rd_data_way1_out_112 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4015 = _T_4014 | _T_3760; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_113; // @[lib.scala 374:16]
  wire [21:0] _T_3761 = _T_2338 ? btb_bank0_rd_data_way1_out_113 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4016 = _T_4015 | _T_3761; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_114; // @[lib.scala 374:16]
  wire [21:0] _T_3762 = _T_2340 ? btb_bank0_rd_data_way1_out_114 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4017 = _T_4016 | _T_3762; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_115; // @[lib.scala 374:16]
  wire [21:0] _T_3763 = _T_2342 ? btb_bank0_rd_data_way1_out_115 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4018 = _T_4017 | _T_3763; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_116; // @[lib.scala 374:16]
  wire [21:0] _T_3764 = _T_2344 ? btb_bank0_rd_data_way1_out_116 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4019 = _T_4018 | _T_3764; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_117; // @[lib.scala 374:16]
  wire [21:0] _T_3765 = _T_2346 ? btb_bank0_rd_data_way1_out_117 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4020 = _T_4019 | _T_3765; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_118; // @[lib.scala 374:16]
  wire [21:0] _T_3766 = _T_2348 ? btb_bank0_rd_data_way1_out_118 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4021 = _T_4020 | _T_3766; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_119; // @[lib.scala 374:16]
  wire [21:0] _T_3767 = _T_2350 ? btb_bank0_rd_data_way1_out_119 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4022 = _T_4021 | _T_3767; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_120; // @[lib.scala 374:16]
  wire [21:0] _T_3768 = _T_2352 ? btb_bank0_rd_data_way1_out_120 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4023 = _T_4022 | _T_3768; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_121; // @[lib.scala 374:16]
  wire [21:0] _T_3769 = _T_2354 ? btb_bank0_rd_data_way1_out_121 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4024 = _T_4023 | _T_3769; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_122; // @[lib.scala 374:16]
  wire [21:0] _T_3770 = _T_2356 ? btb_bank0_rd_data_way1_out_122 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4025 = _T_4024 | _T_3770; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_123; // @[lib.scala 374:16]
  wire [21:0] _T_3771 = _T_2358 ? btb_bank0_rd_data_way1_out_123 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4026 = _T_4025 | _T_3771; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_124; // @[lib.scala 374:16]
  wire [21:0] _T_3772 = _T_2360 ? btb_bank0_rd_data_way1_out_124 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4027 = _T_4026 | _T_3772; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_125; // @[lib.scala 374:16]
  wire [21:0] _T_3773 = _T_2362 ? btb_bank0_rd_data_way1_out_125 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4028 = _T_4027 | _T_3773; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_126; // @[lib.scala 374:16]
  wire [21:0] _T_3774 = _T_2364 ? btb_bank0_rd_data_way1_out_126 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4029 = _T_4028 | _T_3774; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_127; // @[lib.scala 374:16]
  wire [21:0] _T_3775 = _T_2366 ? btb_bank0_rd_data_way1_out_127 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4030 = _T_4029 | _T_3775; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_128; // @[lib.scala 374:16]
  wire [21:0] _T_3776 = _T_2368 ? btb_bank0_rd_data_way1_out_128 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4031 = _T_4030 | _T_3776; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_129; // @[lib.scala 374:16]
  wire [21:0] _T_3777 = _T_2370 ? btb_bank0_rd_data_way1_out_129 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4032 = _T_4031 | _T_3777; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_130; // @[lib.scala 374:16]
  wire [21:0] _T_3778 = _T_2372 ? btb_bank0_rd_data_way1_out_130 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4033 = _T_4032 | _T_3778; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_131; // @[lib.scala 374:16]
  wire [21:0] _T_3779 = _T_2374 ? btb_bank0_rd_data_way1_out_131 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4034 = _T_4033 | _T_3779; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_132; // @[lib.scala 374:16]
  wire [21:0] _T_3780 = _T_2376 ? btb_bank0_rd_data_way1_out_132 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4035 = _T_4034 | _T_3780; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_133; // @[lib.scala 374:16]
  wire [21:0] _T_3781 = _T_2378 ? btb_bank0_rd_data_way1_out_133 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4036 = _T_4035 | _T_3781; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_134; // @[lib.scala 374:16]
  wire [21:0] _T_3782 = _T_2380 ? btb_bank0_rd_data_way1_out_134 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4037 = _T_4036 | _T_3782; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_135; // @[lib.scala 374:16]
  wire [21:0] _T_3783 = _T_2382 ? btb_bank0_rd_data_way1_out_135 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4038 = _T_4037 | _T_3783; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_136; // @[lib.scala 374:16]
  wire [21:0] _T_3784 = _T_2384 ? btb_bank0_rd_data_way1_out_136 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4039 = _T_4038 | _T_3784; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_137; // @[lib.scala 374:16]
  wire [21:0] _T_3785 = _T_2386 ? btb_bank0_rd_data_way1_out_137 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4040 = _T_4039 | _T_3785; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_138; // @[lib.scala 374:16]
  wire [21:0] _T_3786 = _T_2388 ? btb_bank0_rd_data_way1_out_138 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4041 = _T_4040 | _T_3786; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_139; // @[lib.scala 374:16]
  wire [21:0] _T_3787 = _T_2390 ? btb_bank0_rd_data_way1_out_139 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4042 = _T_4041 | _T_3787; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_140; // @[lib.scala 374:16]
  wire [21:0] _T_3788 = _T_2392 ? btb_bank0_rd_data_way1_out_140 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4043 = _T_4042 | _T_3788; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_141; // @[lib.scala 374:16]
  wire [21:0] _T_3789 = _T_2394 ? btb_bank0_rd_data_way1_out_141 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4044 = _T_4043 | _T_3789; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_142; // @[lib.scala 374:16]
  wire [21:0] _T_3790 = _T_2396 ? btb_bank0_rd_data_way1_out_142 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4045 = _T_4044 | _T_3790; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_143; // @[lib.scala 374:16]
  wire [21:0] _T_3791 = _T_2398 ? btb_bank0_rd_data_way1_out_143 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4046 = _T_4045 | _T_3791; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_144; // @[lib.scala 374:16]
  wire [21:0] _T_3792 = _T_2400 ? btb_bank0_rd_data_way1_out_144 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4047 = _T_4046 | _T_3792; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_145; // @[lib.scala 374:16]
  wire [21:0] _T_3793 = _T_2402 ? btb_bank0_rd_data_way1_out_145 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4048 = _T_4047 | _T_3793; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_146; // @[lib.scala 374:16]
  wire [21:0] _T_3794 = _T_2404 ? btb_bank0_rd_data_way1_out_146 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4049 = _T_4048 | _T_3794; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_147; // @[lib.scala 374:16]
  wire [21:0] _T_3795 = _T_2406 ? btb_bank0_rd_data_way1_out_147 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4050 = _T_4049 | _T_3795; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_148; // @[lib.scala 374:16]
  wire [21:0] _T_3796 = _T_2408 ? btb_bank0_rd_data_way1_out_148 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4051 = _T_4050 | _T_3796; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_149; // @[lib.scala 374:16]
  wire [21:0] _T_3797 = _T_2410 ? btb_bank0_rd_data_way1_out_149 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4052 = _T_4051 | _T_3797; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_150; // @[lib.scala 374:16]
  wire [21:0] _T_3798 = _T_2412 ? btb_bank0_rd_data_way1_out_150 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4053 = _T_4052 | _T_3798; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_151; // @[lib.scala 374:16]
  wire [21:0] _T_3799 = _T_2414 ? btb_bank0_rd_data_way1_out_151 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4054 = _T_4053 | _T_3799; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_152; // @[lib.scala 374:16]
  wire [21:0] _T_3800 = _T_2416 ? btb_bank0_rd_data_way1_out_152 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4055 = _T_4054 | _T_3800; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_153; // @[lib.scala 374:16]
  wire [21:0] _T_3801 = _T_2418 ? btb_bank0_rd_data_way1_out_153 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4056 = _T_4055 | _T_3801; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_154; // @[lib.scala 374:16]
  wire [21:0] _T_3802 = _T_2420 ? btb_bank0_rd_data_way1_out_154 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4057 = _T_4056 | _T_3802; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_155; // @[lib.scala 374:16]
  wire [21:0] _T_3803 = _T_2422 ? btb_bank0_rd_data_way1_out_155 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4058 = _T_4057 | _T_3803; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_156; // @[lib.scala 374:16]
  wire [21:0] _T_3804 = _T_2424 ? btb_bank0_rd_data_way1_out_156 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4059 = _T_4058 | _T_3804; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_157; // @[lib.scala 374:16]
  wire [21:0] _T_3805 = _T_2426 ? btb_bank0_rd_data_way1_out_157 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4060 = _T_4059 | _T_3805; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_158; // @[lib.scala 374:16]
  wire [21:0] _T_3806 = _T_2428 ? btb_bank0_rd_data_way1_out_158 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4061 = _T_4060 | _T_3806; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_159; // @[lib.scala 374:16]
  wire [21:0] _T_3807 = _T_2430 ? btb_bank0_rd_data_way1_out_159 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4062 = _T_4061 | _T_3807; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_160; // @[lib.scala 374:16]
  wire [21:0] _T_3808 = _T_2432 ? btb_bank0_rd_data_way1_out_160 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4063 = _T_4062 | _T_3808; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_161; // @[lib.scala 374:16]
  wire [21:0] _T_3809 = _T_2434 ? btb_bank0_rd_data_way1_out_161 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4064 = _T_4063 | _T_3809; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_162; // @[lib.scala 374:16]
  wire [21:0] _T_3810 = _T_2436 ? btb_bank0_rd_data_way1_out_162 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4065 = _T_4064 | _T_3810; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_163; // @[lib.scala 374:16]
  wire [21:0] _T_3811 = _T_2438 ? btb_bank0_rd_data_way1_out_163 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4066 = _T_4065 | _T_3811; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_164; // @[lib.scala 374:16]
  wire [21:0] _T_3812 = _T_2440 ? btb_bank0_rd_data_way1_out_164 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4067 = _T_4066 | _T_3812; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_165; // @[lib.scala 374:16]
  wire [21:0] _T_3813 = _T_2442 ? btb_bank0_rd_data_way1_out_165 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4068 = _T_4067 | _T_3813; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_166; // @[lib.scala 374:16]
  wire [21:0] _T_3814 = _T_2444 ? btb_bank0_rd_data_way1_out_166 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4069 = _T_4068 | _T_3814; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_167; // @[lib.scala 374:16]
  wire [21:0] _T_3815 = _T_2446 ? btb_bank0_rd_data_way1_out_167 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4070 = _T_4069 | _T_3815; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_168; // @[lib.scala 374:16]
  wire [21:0] _T_3816 = _T_2448 ? btb_bank0_rd_data_way1_out_168 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4071 = _T_4070 | _T_3816; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_169; // @[lib.scala 374:16]
  wire [21:0] _T_3817 = _T_2450 ? btb_bank0_rd_data_way1_out_169 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4072 = _T_4071 | _T_3817; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_170; // @[lib.scala 374:16]
  wire [21:0] _T_3818 = _T_2452 ? btb_bank0_rd_data_way1_out_170 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4073 = _T_4072 | _T_3818; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_171; // @[lib.scala 374:16]
  wire [21:0] _T_3819 = _T_2454 ? btb_bank0_rd_data_way1_out_171 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4074 = _T_4073 | _T_3819; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_172; // @[lib.scala 374:16]
  wire [21:0] _T_3820 = _T_2456 ? btb_bank0_rd_data_way1_out_172 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4075 = _T_4074 | _T_3820; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_173; // @[lib.scala 374:16]
  wire [21:0] _T_3821 = _T_2458 ? btb_bank0_rd_data_way1_out_173 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4076 = _T_4075 | _T_3821; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_174; // @[lib.scala 374:16]
  wire [21:0] _T_3822 = _T_2460 ? btb_bank0_rd_data_way1_out_174 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4077 = _T_4076 | _T_3822; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_175; // @[lib.scala 374:16]
  wire [21:0] _T_3823 = _T_2462 ? btb_bank0_rd_data_way1_out_175 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4078 = _T_4077 | _T_3823; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_176; // @[lib.scala 374:16]
  wire [21:0] _T_3824 = _T_2464 ? btb_bank0_rd_data_way1_out_176 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4079 = _T_4078 | _T_3824; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_177; // @[lib.scala 374:16]
  wire [21:0] _T_3825 = _T_2466 ? btb_bank0_rd_data_way1_out_177 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4080 = _T_4079 | _T_3825; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_178; // @[lib.scala 374:16]
  wire [21:0] _T_3826 = _T_2468 ? btb_bank0_rd_data_way1_out_178 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4081 = _T_4080 | _T_3826; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_179; // @[lib.scala 374:16]
  wire [21:0] _T_3827 = _T_2470 ? btb_bank0_rd_data_way1_out_179 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4082 = _T_4081 | _T_3827; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_180; // @[lib.scala 374:16]
  wire [21:0] _T_3828 = _T_2472 ? btb_bank0_rd_data_way1_out_180 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4083 = _T_4082 | _T_3828; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_181; // @[lib.scala 374:16]
  wire [21:0] _T_3829 = _T_2474 ? btb_bank0_rd_data_way1_out_181 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4084 = _T_4083 | _T_3829; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_182; // @[lib.scala 374:16]
  wire [21:0] _T_3830 = _T_2476 ? btb_bank0_rd_data_way1_out_182 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4085 = _T_4084 | _T_3830; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_183; // @[lib.scala 374:16]
  wire [21:0] _T_3831 = _T_2478 ? btb_bank0_rd_data_way1_out_183 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4086 = _T_4085 | _T_3831; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_184; // @[lib.scala 374:16]
  wire [21:0] _T_3832 = _T_2480 ? btb_bank0_rd_data_way1_out_184 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4087 = _T_4086 | _T_3832; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_185; // @[lib.scala 374:16]
  wire [21:0] _T_3833 = _T_2482 ? btb_bank0_rd_data_way1_out_185 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4088 = _T_4087 | _T_3833; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_186; // @[lib.scala 374:16]
  wire [21:0] _T_3834 = _T_2484 ? btb_bank0_rd_data_way1_out_186 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4089 = _T_4088 | _T_3834; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_187; // @[lib.scala 374:16]
  wire [21:0] _T_3835 = _T_2486 ? btb_bank0_rd_data_way1_out_187 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4090 = _T_4089 | _T_3835; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_188; // @[lib.scala 374:16]
  wire [21:0] _T_3836 = _T_2488 ? btb_bank0_rd_data_way1_out_188 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4091 = _T_4090 | _T_3836; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_189; // @[lib.scala 374:16]
  wire [21:0] _T_3837 = _T_2490 ? btb_bank0_rd_data_way1_out_189 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4092 = _T_4091 | _T_3837; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_190; // @[lib.scala 374:16]
  wire [21:0] _T_3838 = _T_2492 ? btb_bank0_rd_data_way1_out_190 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4093 = _T_4092 | _T_3838; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_191; // @[lib.scala 374:16]
  wire [21:0] _T_3839 = _T_2494 ? btb_bank0_rd_data_way1_out_191 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4094 = _T_4093 | _T_3839; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_192; // @[lib.scala 374:16]
  wire [21:0] _T_3840 = _T_2496 ? btb_bank0_rd_data_way1_out_192 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4095 = _T_4094 | _T_3840; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_193; // @[lib.scala 374:16]
  wire [21:0] _T_3841 = _T_2498 ? btb_bank0_rd_data_way1_out_193 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4096 = _T_4095 | _T_3841; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_194; // @[lib.scala 374:16]
  wire [21:0] _T_3842 = _T_2500 ? btb_bank0_rd_data_way1_out_194 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4097 = _T_4096 | _T_3842; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_195; // @[lib.scala 374:16]
  wire [21:0] _T_3843 = _T_2502 ? btb_bank0_rd_data_way1_out_195 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4098 = _T_4097 | _T_3843; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_196; // @[lib.scala 374:16]
  wire [21:0] _T_3844 = _T_2504 ? btb_bank0_rd_data_way1_out_196 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4099 = _T_4098 | _T_3844; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_197; // @[lib.scala 374:16]
  wire [21:0] _T_3845 = _T_2506 ? btb_bank0_rd_data_way1_out_197 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4100 = _T_4099 | _T_3845; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_198; // @[lib.scala 374:16]
  wire [21:0] _T_3846 = _T_2508 ? btb_bank0_rd_data_way1_out_198 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4101 = _T_4100 | _T_3846; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_199; // @[lib.scala 374:16]
  wire [21:0] _T_3847 = _T_2510 ? btb_bank0_rd_data_way1_out_199 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4102 = _T_4101 | _T_3847; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_200; // @[lib.scala 374:16]
  wire [21:0] _T_3848 = _T_2512 ? btb_bank0_rd_data_way1_out_200 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4103 = _T_4102 | _T_3848; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_201; // @[lib.scala 374:16]
  wire [21:0] _T_3849 = _T_2514 ? btb_bank0_rd_data_way1_out_201 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4104 = _T_4103 | _T_3849; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_202; // @[lib.scala 374:16]
  wire [21:0] _T_3850 = _T_2516 ? btb_bank0_rd_data_way1_out_202 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4105 = _T_4104 | _T_3850; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_203; // @[lib.scala 374:16]
  wire [21:0] _T_3851 = _T_2518 ? btb_bank0_rd_data_way1_out_203 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4106 = _T_4105 | _T_3851; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_204; // @[lib.scala 374:16]
  wire [21:0] _T_3852 = _T_2520 ? btb_bank0_rd_data_way1_out_204 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4107 = _T_4106 | _T_3852; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_205; // @[lib.scala 374:16]
  wire [21:0] _T_3853 = _T_2522 ? btb_bank0_rd_data_way1_out_205 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4108 = _T_4107 | _T_3853; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_206; // @[lib.scala 374:16]
  wire [21:0] _T_3854 = _T_2524 ? btb_bank0_rd_data_way1_out_206 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4109 = _T_4108 | _T_3854; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_207; // @[lib.scala 374:16]
  wire [21:0] _T_3855 = _T_2526 ? btb_bank0_rd_data_way1_out_207 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4110 = _T_4109 | _T_3855; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_208; // @[lib.scala 374:16]
  wire [21:0] _T_3856 = _T_2528 ? btb_bank0_rd_data_way1_out_208 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4111 = _T_4110 | _T_3856; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_209; // @[lib.scala 374:16]
  wire [21:0] _T_3857 = _T_2530 ? btb_bank0_rd_data_way1_out_209 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4112 = _T_4111 | _T_3857; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_210; // @[lib.scala 374:16]
  wire [21:0] _T_3858 = _T_2532 ? btb_bank0_rd_data_way1_out_210 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4113 = _T_4112 | _T_3858; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_211; // @[lib.scala 374:16]
  wire [21:0] _T_3859 = _T_2534 ? btb_bank0_rd_data_way1_out_211 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4114 = _T_4113 | _T_3859; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_212; // @[lib.scala 374:16]
  wire [21:0] _T_3860 = _T_2536 ? btb_bank0_rd_data_way1_out_212 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4115 = _T_4114 | _T_3860; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_213; // @[lib.scala 374:16]
  wire [21:0] _T_3861 = _T_2538 ? btb_bank0_rd_data_way1_out_213 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4116 = _T_4115 | _T_3861; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_214; // @[lib.scala 374:16]
  wire [21:0] _T_3862 = _T_2540 ? btb_bank0_rd_data_way1_out_214 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4117 = _T_4116 | _T_3862; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_215; // @[lib.scala 374:16]
  wire [21:0] _T_3863 = _T_2542 ? btb_bank0_rd_data_way1_out_215 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4118 = _T_4117 | _T_3863; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_216; // @[lib.scala 374:16]
  wire [21:0] _T_3864 = _T_2544 ? btb_bank0_rd_data_way1_out_216 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4119 = _T_4118 | _T_3864; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_217; // @[lib.scala 374:16]
  wire [21:0] _T_3865 = _T_2546 ? btb_bank0_rd_data_way1_out_217 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4120 = _T_4119 | _T_3865; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_218; // @[lib.scala 374:16]
  wire [21:0] _T_3866 = _T_2548 ? btb_bank0_rd_data_way1_out_218 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4121 = _T_4120 | _T_3866; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_219; // @[lib.scala 374:16]
  wire [21:0] _T_3867 = _T_2550 ? btb_bank0_rd_data_way1_out_219 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4122 = _T_4121 | _T_3867; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_220; // @[lib.scala 374:16]
  wire [21:0] _T_3868 = _T_2552 ? btb_bank0_rd_data_way1_out_220 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4123 = _T_4122 | _T_3868; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_221; // @[lib.scala 374:16]
  wire [21:0] _T_3869 = _T_2554 ? btb_bank0_rd_data_way1_out_221 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4124 = _T_4123 | _T_3869; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_222; // @[lib.scala 374:16]
  wire [21:0] _T_3870 = _T_2556 ? btb_bank0_rd_data_way1_out_222 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4125 = _T_4124 | _T_3870; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_223; // @[lib.scala 374:16]
  wire [21:0] _T_3871 = _T_2558 ? btb_bank0_rd_data_way1_out_223 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4126 = _T_4125 | _T_3871; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_224; // @[lib.scala 374:16]
  wire [21:0] _T_3872 = _T_2560 ? btb_bank0_rd_data_way1_out_224 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4127 = _T_4126 | _T_3872; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_225; // @[lib.scala 374:16]
  wire [21:0] _T_3873 = _T_2562 ? btb_bank0_rd_data_way1_out_225 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4128 = _T_4127 | _T_3873; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_226; // @[lib.scala 374:16]
  wire [21:0] _T_3874 = _T_2564 ? btb_bank0_rd_data_way1_out_226 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4129 = _T_4128 | _T_3874; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_227; // @[lib.scala 374:16]
  wire [21:0] _T_3875 = _T_2566 ? btb_bank0_rd_data_way1_out_227 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4130 = _T_4129 | _T_3875; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_228; // @[lib.scala 374:16]
  wire [21:0] _T_3876 = _T_2568 ? btb_bank0_rd_data_way1_out_228 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4131 = _T_4130 | _T_3876; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_229; // @[lib.scala 374:16]
  wire [21:0] _T_3877 = _T_2570 ? btb_bank0_rd_data_way1_out_229 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4132 = _T_4131 | _T_3877; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_230; // @[lib.scala 374:16]
  wire [21:0] _T_3878 = _T_2572 ? btb_bank0_rd_data_way1_out_230 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4133 = _T_4132 | _T_3878; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_231; // @[lib.scala 374:16]
  wire [21:0] _T_3879 = _T_2574 ? btb_bank0_rd_data_way1_out_231 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4134 = _T_4133 | _T_3879; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_232; // @[lib.scala 374:16]
  wire [21:0] _T_3880 = _T_2576 ? btb_bank0_rd_data_way1_out_232 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4135 = _T_4134 | _T_3880; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_233; // @[lib.scala 374:16]
  wire [21:0] _T_3881 = _T_2578 ? btb_bank0_rd_data_way1_out_233 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4136 = _T_4135 | _T_3881; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_234; // @[lib.scala 374:16]
  wire [21:0] _T_3882 = _T_2580 ? btb_bank0_rd_data_way1_out_234 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4137 = _T_4136 | _T_3882; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_235; // @[lib.scala 374:16]
  wire [21:0] _T_3883 = _T_2582 ? btb_bank0_rd_data_way1_out_235 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4138 = _T_4137 | _T_3883; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_236; // @[lib.scala 374:16]
  wire [21:0] _T_3884 = _T_2584 ? btb_bank0_rd_data_way1_out_236 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4139 = _T_4138 | _T_3884; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_237; // @[lib.scala 374:16]
  wire [21:0] _T_3885 = _T_2586 ? btb_bank0_rd_data_way1_out_237 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4140 = _T_4139 | _T_3885; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_238; // @[lib.scala 374:16]
  wire [21:0] _T_3886 = _T_2588 ? btb_bank0_rd_data_way1_out_238 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4141 = _T_4140 | _T_3886; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_239; // @[lib.scala 374:16]
  wire [21:0] _T_3887 = _T_2590 ? btb_bank0_rd_data_way1_out_239 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4142 = _T_4141 | _T_3887; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_240; // @[lib.scala 374:16]
  wire [21:0] _T_3888 = _T_2592 ? btb_bank0_rd_data_way1_out_240 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4143 = _T_4142 | _T_3888; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_241; // @[lib.scala 374:16]
  wire [21:0] _T_3889 = _T_2594 ? btb_bank0_rd_data_way1_out_241 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4144 = _T_4143 | _T_3889; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_242; // @[lib.scala 374:16]
  wire [21:0] _T_3890 = _T_2596 ? btb_bank0_rd_data_way1_out_242 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4145 = _T_4144 | _T_3890; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_243; // @[lib.scala 374:16]
  wire [21:0] _T_3891 = _T_2598 ? btb_bank0_rd_data_way1_out_243 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4146 = _T_4145 | _T_3891; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_244; // @[lib.scala 374:16]
  wire [21:0] _T_3892 = _T_2600 ? btb_bank0_rd_data_way1_out_244 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4147 = _T_4146 | _T_3892; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_245; // @[lib.scala 374:16]
  wire [21:0] _T_3893 = _T_2602 ? btb_bank0_rd_data_way1_out_245 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4148 = _T_4147 | _T_3893; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_246; // @[lib.scala 374:16]
  wire [21:0] _T_3894 = _T_2604 ? btb_bank0_rd_data_way1_out_246 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4149 = _T_4148 | _T_3894; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_247; // @[lib.scala 374:16]
  wire [21:0] _T_3895 = _T_2606 ? btb_bank0_rd_data_way1_out_247 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4150 = _T_4149 | _T_3895; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_248; // @[lib.scala 374:16]
  wire [21:0] _T_3896 = _T_2608 ? btb_bank0_rd_data_way1_out_248 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4151 = _T_4150 | _T_3896; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_249; // @[lib.scala 374:16]
  wire [21:0] _T_3897 = _T_2610 ? btb_bank0_rd_data_way1_out_249 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4152 = _T_4151 | _T_3897; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_250; // @[lib.scala 374:16]
  wire [21:0] _T_3898 = _T_2612 ? btb_bank0_rd_data_way1_out_250 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4153 = _T_4152 | _T_3898; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_251; // @[lib.scala 374:16]
  wire [21:0] _T_3899 = _T_2614 ? btb_bank0_rd_data_way1_out_251 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4154 = _T_4153 | _T_3899; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_252; // @[lib.scala 374:16]
  wire [21:0] _T_3900 = _T_2616 ? btb_bank0_rd_data_way1_out_252 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4155 = _T_4154 | _T_3900; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_253; // @[lib.scala 374:16]
  wire [21:0] _T_3901 = _T_2618 ? btb_bank0_rd_data_way1_out_253 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4156 = _T_4155 | _T_3901; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_254; // @[lib.scala 374:16]
  wire [21:0] _T_3902 = _T_2620 ? btb_bank0_rd_data_way1_out_254 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4157 = _T_4156 | _T_3902; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_255; // @[lib.scala 374:16]
  wire [21:0] _T_3903 = _T_2622 ? btb_bank0_rd_data_way1_out_255 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] btb_bank0_rd_data_way1_f = _T_4157 | _T_3903; // @[Mux.scala 27:72]
  wire  _T_55 = btb_bank0_rd_data_way1_f[21:17] == fetch_rd_tag_f; // @[ifu_bp_ctl.scala 131:97]
  wire  _T_56 = btb_bank0_rd_data_way1_f[0] & _T_55; // @[ifu_bp_ctl.scala 131:55]
  wire  _T_59 = _T_56 & _T_49; // @[ifu_bp_ctl.scala 131:117]
  wire  _T_60 = _T_59 & io_ifc_fetch_req_f; // @[ifu_bp_ctl.scala 132:76]
  wire  tag_match_way1_f = _T_60 & _T; // @[ifu_bp_ctl.scala 132:97]
  wire  _T_91 = btb_bank0_rd_data_way1_f[3] ^ btb_bank0_rd_data_way1_f[4]; // @[ifu_bp_ctl.scala 145:91]
  wire  _T_92 = tag_match_way1_f & _T_91; // @[ifu_bp_ctl.scala 145:56]
  wire  _T_96 = ~_T_91; // @[ifu_bp_ctl.scala 146:58]
  wire  _T_97 = tag_match_way1_f & _T_96; // @[ifu_bp_ctl.scala 146:56]
  wire [1:0] tag_match_way1_expanded_f = {_T_92,_T_97}; // @[Cat.scala 29:58]
  wire [21:0] _T_128 = tag_match_way1_expanded_f[1] ? btb_bank0_rd_data_way1_f : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] btb_bank0o_rd_data_f = _T_127 | _T_128; // @[Mux.scala 27:72]
  wire [21:0] _T_146 = _T_144 ? btb_bank0o_rd_data_f : 22'h0; // @[Mux.scala 27:72]
  wire  _T_4160 = btb_rd_addr_p1_f == 8'h0; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4672 = _T_4160 ? btb_bank0_rd_data_way0_out_0 : 22'h0; // @[Mux.scala 27:72]
  wire  _T_4162 = btb_rd_addr_p1_f == 8'h1; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4673 = _T_4162 ? btb_bank0_rd_data_way0_out_1 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4928 = _T_4672 | _T_4673; // @[Mux.scala 27:72]
  wire  _T_4164 = btb_rd_addr_p1_f == 8'h2; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4674 = _T_4164 ? btb_bank0_rd_data_way0_out_2 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4929 = _T_4928 | _T_4674; // @[Mux.scala 27:72]
  wire  _T_4166 = btb_rd_addr_p1_f == 8'h3; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4675 = _T_4166 ? btb_bank0_rd_data_way0_out_3 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4930 = _T_4929 | _T_4675; // @[Mux.scala 27:72]
  wire  _T_4168 = btb_rd_addr_p1_f == 8'h4; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4676 = _T_4168 ? btb_bank0_rd_data_way0_out_4 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4931 = _T_4930 | _T_4676; // @[Mux.scala 27:72]
  wire  _T_4170 = btb_rd_addr_p1_f == 8'h5; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4677 = _T_4170 ? btb_bank0_rd_data_way0_out_5 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4932 = _T_4931 | _T_4677; // @[Mux.scala 27:72]
  wire  _T_4172 = btb_rd_addr_p1_f == 8'h6; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4678 = _T_4172 ? btb_bank0_rd_data_way0_out_6 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4933 = _T_4932 | _T_4678; // @[Mux.scala 27:72]
  wire  _T_4174 = btb_rd_addr_p1_f == 8'h7; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4679 = _T_4174 ? btb_bank0_rd_data_way0_out_7 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4934 = _T_4933 | _T_4679; // @[Mux.scala 27:72]
  wire  _T_4176 = btb_rd_addr_p1_f == 8'h8; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4680 = _T_4176 ? btb_bank0_rd_data_way0_out_8 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4935 = _T_4934 | _T_4680; // @[Mux.scala 27:72]
  wire  _T_4178 = btb_rd_addr_p1_f == 8'h9; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4681 = _T_4178 ? btb_bank0_rd_data_way0_out_9 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4936 = _T_4935 | _T_4681; // @[Mux.scala 27:72]
  wire  _T_4180 = btb_rd_addr_p1_f == 8'ha; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4682 = _T_4180 ? btb_bank0_rd_data_way0_out_10 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4937 = _T_4936 | _T_4682; // @[Mux.scala 27:72]
  wire  _T_4182 = btb_rd_addr_p1_f == 8'hb; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4683 = _T_4182 ? btb_bank0_rd_data_way0_out_11 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4938 = _T_4937 | _T_4683; // @[Mux.scala 27:72]
  wire  _T_4184 = btb_rd_addr_p1_f == 8'hc; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4684 = _T_4184 ? btb_bank0_rd_data_way0_out_12 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4939 = _T_4938 | _T_4684; // @[Mux.scala 27:72]
  wire  _T_4186 = btb_rd_addr_p1_f == 8'hd; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4685 = _T_4186 ? btb_bank0_rd_data_way0_out_13 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4940 = _T_4939 | _T_4685; // @[Mux.scala 27:72]
  wire  _T_4188 = btb_rd_addr_p1_f == 8'he; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4686 = _T_4188 ? btb_bank0_rd_data_way0_out_14 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4941 = _T_4940 | _T_4686; // @[Mux.scala 27:72]
  wire  _T_4190 = btb_rd_addr_p1_f == 8'hf; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4687 = _T_4190 ? btb_bank0_rd_data_way0_out_15 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4942 = _T_4941 | _T_4687; // @[Mux.scala 27:72]
  wire  _T_4192 = btb_rd_addr_p1_f == 8'h10; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4688 = _T_4192 ? btb_bank0_rd_data_way0_out_16 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4943 = _T_4942 | _T_4688; // @[Mux.scala 27:72]
  wire  _T_4194 = btb_rd_addr_p1_f == 8'h11; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4689 = _T_4194 ? btb_bank0_rd_data_way0_out_17 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4944 = _T_4943 | _T_4689; // @[Mux.scala 27:72]
  wire  _T_4196 = btb_rd_addr_p1_f == 8'h12; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4690 = _T_4196 ? btb_bank0_rd_data_way0_out_18 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4945 = _T_4944 | _T_4690; // @[Mux.scala 27:72]
  wire  _T_4198 = btb_rd_addr_p1_f == 8'h13; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4691 = _T_4198 ? btb_bank0_rd_data_way0_out_19 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4946 = _T_4945 | _T_4691; // @[Mux.scala 27:72]
  wire  _T_4200 = btb_rd_addr_p1_f == 8'h14; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4692 = _T_4200 ? btb_bank0_rd_data_way0_out_20 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4947 = _T_4946 | _T_4692; // @[Mux.scala 27:72]
  wire  _T_4202 = btb_rd_addr_p1_f == 8'h15; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4693 = _T_4202 ? btb_bank0_rd_data_way0_out_21 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4948 = _T_4947 | _T_4693; // @[Mux.scala 27:72]
  wire  _T_4204 = btb_rd_addr_p1_f == 8'h16; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4694 = _T_4204 ? btb_bank0_rd_data_way0_out_22 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4949 = _T_4948 | _T_4694; // @[Mux.scala 27:72]
  wire  _T_4206 = btb_rd_addr_p1_f == 8'h17; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4695 = _T_4206 ? btb_bank0_rd_data_way0_out_23 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4950 = _T_4949 | _T_4695; // @[Mux.scala 27:72]
  wire  _T_4208 = btb_rd_addr_p1_f == 8'h18; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4696 = _T_4208 ? btb_bank0_rd_data_way0_out_24 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4951 = _T_4950 | _T_4696; // @[Mux.scala 27:72]
  wire  _T_4210 = btb_rd_addr_p1_f == 8'h19; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4697 = _T_4210 ? btb_bank0_rd_data_way0_out_25 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4952 = _T_4951 | _T_4697; // @[Mux.scala 27:72]
  wire  _T_4212 = btb_rd_addr_p1_f == 8'h1a; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4698 = _T_4212 ? btb_bank0_rd_data_way0_out_26 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4953 = _T_4952 | _T_4698; // @[Mux.scala 27:72]
  wire  _T_4214 = btb_rd_addr_p1_f == 8'h1b; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4699 = _T_4214 ? btb_bank0_rd_data_way0_out_27 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4954 = _T_4953 | _T_4699; // @[Mux.scala 27:72]
  wire  _T_4216 = btb_rd_addr_p1_f == 8'h1c; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4700 = _T_4216 ? btb_bank0_rd_data_way0_out_28 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4955 = _T_4954 | _T_4700; // @[Mux.scala 27:72]
  wire  _T_4218 = btb_rd_addr_p1_f == 8'h1d; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4701 = _T_4218 ? btb_bank0_rd_data_way0_out_29 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4956 = _T_4955 | _T_4701; // @[Mux.scala 27:72]
  wire  _T_4220 = btb_rd_addr_p1_f == 8'h1e; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4702 = _T_4220 ? btb_bank0_rd_data_way0_out_30 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4957 = _T_4956 | _T_4702; // @[Mux.scala 27:72]
  wire  _T_4222 = btb_rd_addr_p1_f == 8'h1f; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4703 = _T_4222 ? btb_bank0_rd_data_way0_out_31 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4958 = _T_4957 | _T_4703; // @[Mux.scala 27:72]
  wire  _T_4224 = btb_rd_addr_p1_f == 8'h20; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4704 = _T_4224 ? btb_bank0_rd_data_way0_out_32 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4959 = _T_4958 | _T_4704; // @[Mux.scala 27:72]
  wire  _T_4226 = btb_rd_addr_p1_f == 8'h21; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4705 = _T_4226 ? btb_bank0_rd_data_way0_out_33 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4960 = _T_4959 | _T_4705; // @[Mux.scala 27:72]
  wire  _T_4228 = btb_rd_addr_p1_f == 8'h22; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4706 = _T_4228 ? btb_bank0_rd_data_way0_out_34 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4961 = _T_4960 | _T_4706; // @[Mux.scala 27:72]
  wire  _T_4230 = btb_rd_addr_p1_f == 8'h23; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4707 = _T_4230 ? btb_bank0_rd_data_way0_out_35 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4962 = _T_4961 | _T_4707; // @[Mux.scala 27:72]
  wire  _T_4232 = btb_rd_addr_p1_f == 8'h24; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4708 = _T_4232 ? btb_bank0_rd_data_way0_out_36 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4963 = _T_4962 | _T_4708; // @[Mux.scala 27:72]
  wire  _T_4234 = btb_rd_addr_p1_f == 8'h25; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4709 = _T_4234 ? btb_bank0_rd_data_way0_out_37 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4964 = _T_4963 | _T_4709; // @[Mux.scala 27:72]
  wire  _T_4236 = btb_rd_addr_p1_f == 8'h26; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4710 = _T_4236 ? btb_bank0_rd_data_way0_out_38 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4965 = _T_4964 | _T_4710; // @[Mux.scala 27:72]
  wire  _T_4238 = btb_rd_addr_p1_f == 8'h27; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4711 = _T_4238 ? btb_bank0_rd_data_way0_out_39 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4966 = _T_4965 | _T_4711; // @[Mux.scala 27:72]
  wire  _T_4240 = btb_rd_addr_p1_f == 8'h28; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4712 = _T_4240 ? btb_bank0_rd_data_way0_out_40 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4967 = _T_4966 | _T_4712; // @[Mux.scala 27:72]
  wire  _T_4242 = btb_rd_addr_p1_f == 8'h29; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4713 = _T_4242 ? btb_bank0_rd_data_way0_out_41 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4968 = _T_4967 | _T_4713; // @[Mux.scala 27:72]
  wire  _T_4244 = btb_rd_addr_p1_f == 8'h2a; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4714 = _T_4244 ? btb_bank0_rd_data_way0_out_42 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4969 = _T_4968 | _T_4714; // @[Mux.scala 27:72]
  wire  _T_4246 = btb_rd_addr_p1_f == 8'h2b; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4715 = _T_4246 ? btb_bank0_rd_data_way0_out_43 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4970 = _T_4969 | _T_4715; // @[Mux.scala 27:72]
  wire  _T_4248 = btb_rd_addr_p1_f == 8'h2c; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4716 = _T_4248 ? btb_bank0_rd_data_way0_out_44 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4971 = _T_4970 | _T_4716; // @[Mux.scala 27:72]
  wire  _T_4250 = btb_rd_addr_p1_f == 8'h2d; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4717 = _T_4250 ? btb_bank0_rd_data_way0_out_45 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4972 = _T_4971 | _T_4717; // @[Mux.scala 27:72]
  wire  _T_4252 = btb_rd_addr_p1_f == 8'h2e; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4718 = _T_4252 ? btb_bank0_rd_data_way0_out_46 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4973 = _T_4972 | _T_4718; // @[Mux.scala 27:72]
  wire  _T_4254 = btb_rd_addr_p1_f == 8'h2f; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4719 = _T_4254 ? btb_bank0_rd_data_way0_out_47 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4974 = _T_4973 | _T_4719; // @[Mux.scala 27:72]
  wire  _T_4256 = btb_rd_addr_p1_f == 8'h30; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4720 = _T_4256 ? btb_bank0_rd_data_way0_out_48 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4975 = _T_4974 | _T_4720; // @[Mux.scala 27:72]
  wire  _T_4258 = btb_rd_addr_p1_f == 8'h31; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4721 = _T_4258 ? btb_bank0_rd_data_way0_out_49 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4976 = _T_4975 | _T_4721; // @[Mux.scala 27:72]
  wire  _T_4260 = btb_rd_addr_p1_f == 8'h32; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4722 = _T_4260 ? btb_bank0_rd_data_way0_out_50 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4977 = _T_4976 | _T_4722; // @[Mux.scala 27:72]
  wire  _T_4262 = btb_rd_addr_p1_f == 8'h33; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4723 = _T_4262 ? btb_bank0_rd_data_way0_out_51 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4978 = _T_4977 | _T_4723; // @[Mux.scala 27:72]
  wire  _T_4264 = btb_rd_addr_p1_f == 8'h34; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4724 = _T_4264 ? btb_bank0_rd_data_way0_out_52 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4979 = _T_4978 | _T_4724; // @[Mux.scala 27:72]
  wire  _T_4266 = btb_rd_addr_p1_f == 8'h35; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4725 = _T_4266 ? btb_bank0_rd_data_way0_out_53 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4980 = _T_4979 | _T_4725; // @[Mux.scala 27:72]
  wire  _T_4268 = btb_rd_addr_p1_f == 8'h36; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4726 = _T_4268 ? btb_bank0_rd_data_way0_out_54 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4981 = _T_4980 | _T_4726; // @[Mux.scala 27:72]
  wire  _T_4270 = btb_rd_addr_p1_f == 8'h37; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4727 = _T_4270 ? btb_bank0_rd_data_way0_out_55 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4982 = _T_4981 | _T_4727; // @[Mux.scala 27:72]
  wire  _T_4272 = btb_rd_addr_p1_f == 8'h38; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4728 = _T_4272 ? btb_bank0_rd_data_way0_out_56 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4983 = _T_4982 | _T_4728; // @[Mux.scala 27:72]
  wire  _T_4274 = btb_rd_addr_p1_f == 8'h39; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4729 = _T_4274 ? btb_bank0_rd_data_way0_out_57 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4984 = _T_4983 | _T_4729; // @[Mux.scala 27:72]
  wire  _T_4276 = btb_rd_addr_p1_f == 8'h3a; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4730 = _T_4276 ? btb_bank0_rd_data_way0_out_58 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4985 = _T_4984 | _T_4730; // @[Mux.scala 27:72]
  wire  _T_4278 = btb_rd_addr_p1_f == 8'h3b; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4731 = _T_4278 ? btb_bank0_rd_data_way0_out_59 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4986 = _T_4985 | _T_4731; // @[Mux.scala 27:72]
  wire  _T_4280 = btb_rd_addr_p1_f == 8'h3c; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4732 = _T_4280 ? btb_bank0_rd_data_way0_out_60 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4987 = _T_4986 | _T_4732; // @[Mux.scala 27:72]
  wire  _T_4282 = btb_rd_addr_p1_f == 8'h3d; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4733 = _T_4282 ? btb_bank0_rd_data_way0_out_61 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4988 = _T_4987 | _T_4733; // @[Mux.scala 27:72]
  wire  _T_4284 = btb_rd_addr_p1_f == 8'h3e; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4734 = _T_4284 ? btb_bank0_rd_data_way0_out_62 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4989 = _T_4988 | _T_4734; // @[Mux.scala 27:72]
  wire  _T_4286 = btb_rd_addr_p1_f == 8'h3f; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4735 = _T_4286 ? btb_bank0_rd_data_way0_out_63 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4990 = _T_4989 | _T_4735; // @[Mux.scala 27:72]
  wire  _T_4288 = btb_rd_addr_p1_f == 8'h40; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4736 = _T_4288 ? btb_bank0_rd_data_way0_out_64 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4991 = _T_4990 | _T_4736; // @[Mux.scala 27:72]
  wire  _T_4290 = btb_rd_addr_p1_f == 8'h41; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4737 = _T_4290 ? btb_bank0_rd_data_way0_out_65 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4992 = _T_4991 | _T_4737; // @[Mux.scala 27:72]
  wire  _T_4292 = btb_rd_addr_p1_f == 8'h42; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4738 = _T_4292 ? btb_bank0_rd_data_way0_out_66 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4993 = _T_4992 | _T_4738; // @[Mux.scala 27:72]
  wire  _T_4294 = btb_rd_addr_p1_f == 8'h43; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4739 = _T_4294 ? btb_bank0_rd_data_way0_out_67 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4994 = _T_4993 | _T_4739; // @[Mux.scala 27:72]
  wire  _T_4296 = btb_rd_addr_p1_f == 8'h44; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4740 = _T_4296 ? btb_bank0_rd_data_way0_out_68 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4995 = _T_4994 | _T_4740; // @[Mux.scala 27:72]
  wire  _T_4298 = btb_rd_addr_p1_f == 8'h45; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4741 = _T_4298 ? btb_bank0_rd_data_way0_out_69 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4996 = _T_4995 | _T_4741; // @[Mux.scala 27:72]
  wire  _T_4300 = btb_rd_addr_p1_f == 8'h46; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4742 = _T_4300 ? btb_bank0_rd_data_way0_out_70 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4997 = _T_4996 | _T_4742; // @[Mux.scala 27:72]
  wire  _T_4302 = btb_rd_addr_p1_f == 8'h47; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4743 = _T_4302 ? btb_bank0_rd_data_way0_out_71 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4998 = _T_4997 | _T_4743; // @[Mux.scala 27:72]
  wire  _T_4304 = btb_rd_addr_p1_f == 8'h48; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4744 = _T_4304 ? btb_bank0_rd_data_way0_out_72 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4999 = _T_4998 | _T_4744; // @[Mux.scala 27:72]
  wire  _T_4306 = btb_rd_addr_p1_f == 8'h49; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4745 = _T_4306 ? btb_bank0_rd_data_way0_out_73 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5000 = _T_4999 | _T_4745; // @[Mux.scala 27:72]
  wire  _T_4308 = btb_rd_addr_p1_f == 8'h4a; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4746 = _T_4308 ? btb_bank0_rd_data_way0_out_74 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5001 = _T_5000 | _T_4746; // @[Mux.scala 27:72]
  wire  _T_4310 = btb_rd_addr_p1_f == 8'h4b; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4747 = _T_4310 ? btb_bank0_rd_data_way0_out_75 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5002 = _T_5001 | _T_4747; // @[Mux.scala 27:72]
  wire  _T_4312 = btb_rd_addr_p1_f == 8'h4c; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4748 = _T_4312 ? btb_bank0_rd_data_way0_out_76 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5003 = _T_5002 | _T_4748; // @[Mux.scala 27:72]
  wire  _T_4314 = btb_rd_addr_p1_f == 8'h4d; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4749 = _T_4314 ? btb_bank0_rd_data_way0_out_77 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5004 = _T_5003 | _T_4749; // @[Mux.scala 27:72]
  wire  _T_4316 = btb_rd_addr_p1_f == 8'h4e; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4750 = _T_4316 ? btb_bank0_rd_data_way0_out_78 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5005 = _T_5004 | _T_4750; // @[Mux.scala 27:72]
  wire  _T_4318 = btb_rd_addr_p1_f == 8'h4f; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4751 = _T_4318 ? btb_bank0_rd_data_way0_out_79 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5006 = _T_5005 | _T_4751; // @[Mux.scala 27:72]
  wire  _T_4320 = btb_rd_addr_p1_f == 8'h50; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4752 = _T_4320 ? btb_bank0_rd_data_way0_out_80 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5007 = _T_5006 | _T_4752; // @[Mux.scala 27:72]
  wire  _T_4322 = btb_rd_addr_p1_f == 8'h51; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4753 = _T_4322 ? btb_bank0_rd_data_way0_out_81 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5008 = _T_5007 | _T_4753; // @[Mux.scala 27:72]
  wire  _T_4324 = btb_rd_addr_p1_f == 8'h52; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4754 = _T_4324 ? btb_bank0_rd_data_way0_out_82 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5009 = _T_5008 | _T_4754; // @[Mux.scala 27:72]
  wire  _T_4326 = btb_rd_addr_p1_f == 8'h53; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4755 = _T_4326 ? btb_bank0_rd_data_way0_out_83 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5010 = _T_5009 | _T_4755; // @[Mux.scala 27:72]
  wire  _T_4328 = btb_rd_addr_p1_f == 8'h54; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4756 = _T_4328 ? btb_bank0_rd_data_way0_out_84 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5011 = _T_5010 | _T_4756; // @[Mux.scala 27:72]
  wire  _T_4330 = btb_rd_addr_p1_f == 8'h55; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4757 = _T_4330 ? btb_bank0_rd_data_way0_out_85 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5012 = _T_5011 | _T_4757; // @[Mux.scala 27:72]
  wire  _T_4332 = btb_rd_addr_p1_f == 8'h56; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4758 = _T_4332 ? btb_bank0_rd_data_way0_out_86 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5013 = _T_5012 | _T_4758; // @[Mux.scala 27:72]
  wire  _T_4334 = btb_rd_addr_p1_f == 8'h57; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4759 = _T_4334 ? btb_bank0_rd_data_way0_out_87 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5014 = _T_5013 | _T_4759; // @[Mux.scala 27:72]
  wire  _T_4336 = btb_rd_addr_p1_f == 8'h58; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4760 = _T_4336 ? btb_bank0_rd_data_way0_out_88 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5015 = _T_5014 | _T_4760; // @[Mux.scala 27:72]
  wire  _T_4338 = btb_rd_addr_p1_f == 8'h59; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4761 = _T_4338 ? btb_bank0_rd_data_way0_out_89 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5016 = _T_5015 | _T_4761; // @[Mux.scala 27:72]
  wire  _T_4340 = btb_rd_addr_p1_f == 8'h5a; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4762 = _T_4340 ? btb_bank0_rd_data_way0_out_90 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5017 = _T_5016 | _T_4762; // @[Mux.scala 27:72]
  wire  _T_4342 = btb_rd_addr_p1_f == 8'h5b; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4763 = _T_4342 ? btb_bank0_rd_data_way0_out_91 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5018 = _T_5017 | _T_4763; // @[Mux.scala 27:72]
  wire  _T_4344 = btb_rd_addr_p1_f == 8'h5c; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4764 = _T_4344 ? btb_bank0_rd_data_way0_out_92 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5019 = _T_5018 | _T_4764; // @[Mux.scala 27:72]
  wire  _T_4346 = btb_rd_addr_p1_f == 8'h5d; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4765 = _T_4346 ? btb_bank0_rd_data_way0_out_93 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5020 = _T_5019 | _T_4765; // @[Mux.scala 27:72]
  wire  _T_4348 = btb_rd_addr_p1_f == 8'h5e; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4766 = _T_4348 ? btb_bank0_rd_data_way0_out_94 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5021 = _T_5020 | _T_4766; // @[Mux.scala 27:72]
  wire  _T_4350 = btb_rd_addr_p1_f == 8'h5f; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4767 = _T_4350 ? btb_bank0_rd_data_way0_out_95 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5022 = _T_5021 | _T_4767; // @[Mux.scala 27:72]
  wire  _T_4352 = btb_rd_addr_p1_f == 8'h60; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4768 = _T_4352 ? btb_bank0_rd_data_way0_out_96 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5023 = _T_5022 | _T_4768; // @[Mux.scala 27:72]
  wire  _T_4354 = btb_rd_addr_p1_f == 8'h61; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4769 = _T_4354 ? btb_bank0_rd_data_way0_out_97 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5024 = _T_5023 | _T_4769; // @[Mux.scala 27:72]
  wire  _T_4356 = btb_rd_addr_p1_f == 8'h62; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4770 = _T_4356 ? btb_bank0_rd_data_way0_out_98 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5025 = _T_5024 | _T_4770; // @[Mux.scala 27:72]
  wire  _T_4358 = btb_rd_addr_p1_f == 8'h63; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4771 = _T_4358 ? btb_bank0_rd_data_way0_out_99 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5026 = _T_5025 | _T_4771; // @[Mux.scala 27:72]
  wire  _T_4360 = btb_rd_addr_p1_f == 8'h64; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4772 = _T_4360 ? btb_bank0_rd_data_way0_out_100 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5027 = _T_5026 | _T_4772; // @[Mux.scala 27:72]
  wire  _T_4362 = btb_rd_addr_p1_f == 8'h65; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4773 = _T_4362 ? btb_bank0_rd_data_way0_out_101 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5028 = _T_5027 | _T_4773; // @[Mux.scala 27:72]
  wire  _T_4364 = btb_rd_addr_p1_f == 8'h66; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4774 = _T_4364 ? btb_bank0_rd_data_way0_out_102 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5029 = _T_5028 | _T_4774; // @[Mux.scala 27:72]
  wire  _T_4366 = btb_rd_addr_p1_f == 8'h67; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4775 = _T_4366 ? btb_bank0_rd_data_way0_out_103 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5030 = _T_5029 | _T_4775; // @[Mux.scala 27:72]
  wire  _T_4368 = btb_rd_addr_p1_f == 8'h68; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4776 = _T_4368 ? btb_bank0_rd_data_way0_out_104 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5031 = _T_5030 | _T_4776; // @[Mux.scala 27:72]
  wire  _T_4370 = btb_rd_addr_p1_f == 8'h69; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4777 = _T_4370 ? btb_bank0_rd_data_way0_out_105 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5032 = _T_5031 | _T_4777; // @[Mux.scala 27:72]
  wire  _T_4372 = btb_rd_addr_p1_f == 8'h6a; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4778 = _T_4372 ? btb_bank0_rd_data_way0_out_106 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5033 = _T_5032 | _T_4778; // @[Mux.scala 27:72]
  wire  _T_4374 = btb_rd_addr_p1_f == 8'h6b; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4779 = _T_4374 ? btb_bank0_rd_data_way0_out_107 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5034 = _T_5033 | _T_4779; // @[Mux.scala 27:72]
  wire  _T_4376 = btb_rd_addr_p1_f == 8'h6c; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4780 = _T_4376 ? btb_bank0_rd_data_way0_out_108 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5035 = _T_5034 | _T_4780; // @[Mux.scala 27:72]
  wire  _T_4378 = btb_rd_addr_p1_f == 8'h6d; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4781 = _T_4378 ? btb_bank0_rd_data_way0_out_109 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5036 = _T_5035 | _T_4781; // @[Mux.scala 27:72]
  wire  _T_4380 = btb_rd_addr_p1_f == 8'h6e; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4782 = _T_4380 ? btb_bank0_rd_data_way0_out_110 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5037 = _T_5036 | _T_4782; // @[Mux.scala 27:72]
  wire  _T_4382 = btb_rd_addr_p1_f == 8'h6f; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4783 = _T_4382 ? btb_bank0_rd_data_way0_out_111 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5038 = _T_5037 | _T_4783; // @[Mux.scala 27:72]
  wire  _T_4384 = btb_rd_addr_p1_f == 8'h70; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4784 = _T_4384 ? btb_bank0_rd_data_way0_out_112 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5039 = _T_5038 | _T_4784; // @[Mux.scala 27:72]
  wire  _T_4386 = btb_rd_addr_p1_f == 8'h71; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4785 = _T_4386 ? btb_bank0_rd_data_way0_out_113 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5040 = _T_5039 | _T_4785; // @[Mux.scala 27:72]
  wire  _T_4388 = btb_rd_addr_p1_f == 8'h72; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4786 = _T_4388 ? btb_bank0_rd_data_way0_out_114 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5041 = _T_5040 | _T_4786; // @[Mux.scala 27:72]
  wire  _T_4390 = btb_rd_addr_p1_f == 8'h73; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4787 = _T_4390 ? btb_bank0_rd_data_way0_out_115 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5042 = _T_5041 | _T_4787; // @[Mux.scala 27:72]
  wire  _T_4392 = btb_rd_addr_p1_f == 8'h74; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4788 = _T_4392 ? btb_bank0_rd_data_way0_out_116 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5043 = _T_5042 | _T_4788; // @[Mux.scala 27:72]
  wire  _T_4394 = btb_rd_addr_p1_f == 8'h75; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4789 = _T_4394 ? btb_bank0_rd_data_way0_out_117 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5044 = _T_5043 | _T_4789; // @[Mux.scala 27:72]
  wire  _T_4396 = btb_rd_addr_p1_f == 8'h76; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4790 = _T_4396 ? btb_bank0_rd_data_way0_out_118 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5045 = _T_5044 | _T_4790; // @[Mux.scala 27:72]
  wire  _T_4398 = btb_rd_addr_p1_f == 8'h77; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4791 = _T_4398 ? btb_bank0_rd_data_way0_out_119 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5046 = _T_5045 | _T_4791; // @[Mux.scala 27:72]
  wire  _T_4400 = btb_rd_addr_p1_f == 8'h78; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4792 = _T_4400 ? btb_bank0_rd_data_way0_out_120 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5047 = _T_5046 | _T_4792; // @[Mux.scala 27:72]
  wire  _T_4402 = btb_rd_addr_p1_f == 8'h79; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4793 = _T_4402 ? btb_bank0_rd_data_way0_out_121 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5048 = _T_5047 | _T_4793; // @[Mux.scala 27:72]
  wire  _T_4404 = btb_rd_addr_p1_f == 8'h7a; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4794 = _T_4404 ? btb_bank0_rd_data_way0_out_122 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5049 = _T_5048 | _T_4794; // @[Mux.scala 27:72]
  wire  _T_4406 = btb_rd_addr_p1_f == 8'h7b; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4795 = _T_4406 ? btb_bank0_rd_data_way0_out_123 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5050 = _T_5049 | _T_4795; // @[Mux.scala 27:72]
  wire  _T_4408 = btb_rd_addr_p1_f == 8'h7c; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4796 = _T_4408 ? btb_bank0_rd_data_way0_out_124 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5051 = _T_5050 | _T_4796; // @[Mux.scala 27:72]
  wire  _T_4410 = btb_rd_addr_p1_f == 8'h7d; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4797 = _T_4410 ? btb_bank0_rd_data_way0_out_125 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5052 = _T_5051 | _T_4797; // @[Mux.scala 27:72]
  wire  _T_4412 = btb_rd_addr_p1_f == 8'h7e; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4798 = _T_4412 ? btb_bank0_rd_data_way0_out_126 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5053 = _T_5052 | _T_4798; // @[Mux.scala 27:72]
  wire  _T_4414 = btb_rd_addr_p1_f == 8'h7f; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4799 = _T_4414 ? btb_bank0_rd_data_way0_out_127 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5054 = _T_5053 | _T_4799; // @[Mux.scala 27:72]
  wire  _T_4416 = btb_rd_addr_p1_f == 8'h80; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4800 = _T_4416 ? btb_bank0_rd_data_way0_out_128 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5055 = _T_5054 | _T_4800; // @[Mux.scala 27:72]
  wire  _T_4418 = btb_rd_addr_p1_f == 8'h81; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4801 = _T_4418 ? btb_bank0_rd_data_way0_out_129 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5056 = _T_5055 | _T_4801; // @[Mux.scala 27:72]
  wire  _T_4420 = btb_rd_addr_p1_f == 8'h82; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4802 = _T_4420 ? btb_bank0_rd_data_way0_out_130 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5057 = _T_5056 | _T_4802; // @[Mux.scala 27:72]
  wire  _T_4422 = btb_rd_addr_p1_f == 8'h83; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4803 = _T_4422 ? btb_bank0_rd_data_way0_out_131 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5058 = _T_5057 | _T_4803; // @[Mux.scala 27:72]
  wire  _T_4424 = btb_rd_addr_p1_f == 8'h84; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4804 = _T_4424 ? btb_bank0_rd_data_way0_out_132 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5059 = _T_5058 | _T_4804; // @[Mux.scala 27:72]
  wire  _T_4426 = btb_rd_addr_p1_f == 8'h85; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4805 = _T_4426 ? btb_bank0_rd_data_way0_out_133 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5060 = _T_5059 | _T_4805; // @[Mux.scala 27:72]
  wire  _T_4428 = btb_rd_addr_p1_f == 8'h86; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4806 = _T_4428 ? btb_bank0_rd_data_way0_out_134 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5061 = _T_5060 | _T_4806; // @[Mux.scala 27:72]
  wire  _T_4430 = btb_rd_addr_p1_f == 8'h87; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4807 = _T_4430 ? btb_bank0_rd_data_way0_out_135 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5062 = _T_5061 | _T_4807; // @[Mux.scala 27:72]
  wire  _T_4432 = btb_rd_addr_p1_f == 8'h88; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4808 = _T_4432 ? btb_bank0_rd_data_way0_out_136 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5063 = _T_5062 | _T_4808; // @[Mux.scala 27:72]
  wire  _T_4434 = btb_rd_addr_p1_f == 8'h89; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4809 = _T_4434 ? btb_bank0_rd_data_way0_out_137 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5064 = _T_5063 | _T_4809; // @[Mux.scala 27:72]
  wire  _T_4436 = btb_rd_addr_p1_f == 8'h8a; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4810 = _T_4436 ? btb_bank0_rd_data_way0_out_138 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5065 = _T_5064 | _T_4810; // @[Mux.scala 27:72]
  wire  _T_4438 = btb_rd_addr_p1_f == 8'h8b; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4811 = _T_4438 ? btb_bank0_rd_data_way0_out_139 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5066 = _T_5065 | _T_4811; // @[Mux.scala 27:72]
  wire  _T_4440 = btb_rd_addr_p1_f == 8'h8c; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4812 = _T_4440 ? btb_bank0_rd_data_way0_out_140 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5067 = _T_5066 | _T_4812; // @[Mux.scala 27:72]
  wire  _T_4442 = btb_rd_addr_p1_f == 8'h8d; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4813 = _T_4442 ? btb_bank0_rd_data_way0_out_141 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5068 = _T_5067 | _T_4813; // @[Mux.scala 27:72]
  wire  _T_4444 = btb_rd_addr_p1_f == 8'h8e; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4814 = _T_4444 ? btb_bank0_rd_data_way0_out_142 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5069 = _T_5068 | _T_4814; // @[Mux.scala 27:72]
  wire  _T_4446 = btb_rd_addr_p1_f == 8'h8f; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4815 = _T_4446 ? btb_bank0_rd_data_way0_out_143 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5070 = _T_5069 | _T_4815; // @[Mux.scala 27:72]
  wire  _T_4448 = btb_rd_addr_p1_f == 8'h90; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4816 = _T_4448 ? btb_bank0_rd_data_way0_out_144 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5071 = _T_5070 | _T_4816; // @[Mux.scala 27:72]
  wire  _T_4450 = btb_rd_addr_p1_f == 8'h91; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4817 = _T_4450 ? btb_bank0_rd_data_way0_out_145 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5072 = _T_5071 | _T_4817; // @[Mux.scala 27:72]
  wire  _T_4452 = btb_rd_addr_p1_f == 8'h92; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4818 = _T_4452 ? btb_bank0_rd_data_way0_out_146 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5073 = _T_5072 | _T_4818; // @[Mux.scala 27:72]
  wire  _T_4454 = btb_rd_addr_p1_f == 8'h93; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4819 = _T_4454 ? btb_bank0_rd_data_way0_out_147 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5074 = _T_5073 | _T_4819; // @[Mux.scala 27:72]
  wire  _T_4456 = btb_rd_addr_p1_f == 8'h94; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4820 = _T_4456 ? btb_bank0_rd_data_way0_out_148 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5075 = _T_5074 | _T_4820; // @[Mux.scala 27:72]
  wire  _T_4458 = btb_rd_addr_p1_f == 8'h95; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4821 = _T_4458 ? btb_bank0_rd_data_way0_out_149 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5076 = _T_5075 | _T_4821; // @[Mux.scala 27:72]
  wire  _T_4460 = btb_rd_addr_p1_f == 8'h96; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4822 = _T_4460 ? btb_bank0_rd_data_way0_out_150 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5077 = _T_5076 | _T_4822; // @[Mux.scala 27:72]
  wire  _T_4462 = btb_rd_addr_p1_f == 8'h97; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4823 = _T_4462 ? btb_bank0_rd_data_way0_out_151 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5078 = _T_5077 | _T_4823; // @[Mux.scala 27:72]
  wire  _T_4464 = btb_rd_addr_p1_f == 8'h98; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4824 = _T_4464 ? btb_bank0_rd_data_way0_out_152 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5079 = _T_5078 | _T_4824; // @[Mux.scala 27:72]
  wire  _T_4466 = btb_rd_addr_p1_f == 8'h99; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4825 = _T_4466 ? btb_bank0_rd_data_way0_out_153 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5080 = _T_5079 | _T_4825; // @[Mux.scala 27:72]
  wire  _T_4468 = btb_rd_addr_p1_f == 8'h9a; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4826 = _T_4468 ? btb_bank0_rd_data_way0_out_154 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5081 = _T_5080 | _T_4826; // @[Mux.scala 27:72]
  wire  _T_4470 = btb_rd_addr_p1_f == 8'h9b; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4827 = _T_4470 ? btb_bank0_rd_data_way0_out_155 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5082 = _T_5081 | _T_4827; // @[Mux.scala 27:72]
  wire  _T_4472 = btb_rd_addr_p1_f == 8'h9c; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4828 = _T_4472 ? btb_bank0_rd_data_way0_out_156 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5083 = _T_5082 | _T_4828; // @[Mux.scala 27:72]
  wire  _T_4474 = btb_rd_addr_p1_f == 8'h9d; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4829 = _T_4474 ? btb_bank0_rd_data_way0_out_157 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5084 = _T_5083 | _T_4829; // @[Mux.scala 27:72]
  wire  _T_4476 = btb_rd_addr_p1_f == 8'h9e; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4830 = _T_4476 ? btb_bank0_rd_data_way0_out_158 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5085 = _T_5084 | _T_4830; // @[Mux.scala 27:72]
  wire  _T_4478 = btb_rd_addr_p1_f == 8'h9f; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4831 = _T_4478 ? btb_bank0_rd_data_way0_out_159 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5086 = _T_5085 | _T_4831; // @[Mux.scala 27:72]
  wire  _T_4480 = btb_rd_addr_p1_f == 8'ha0; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4832 = _T_4480 ? btb_bank0_rd_data_way0_out_160 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5087 = _T_5086 | _T_4832; // @[Mux.scala 27:72]
  wire  _T_4482 = btb_rd_addr_p1_f == 8'ha1; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4833 = _T_4482 ? btb_bank0_rd_data_way0_out_161 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5088 = _T_5087 | _T_4833; // @[Mux.scala 27:72]
  wire  _T_4484 = btb_rd_addr_p1_f == 8'ha2; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4834 = _T_4484 ? btb_bank0_rd_data_way0_out_162 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5089 = _T_5088 | _T_4834; // @[Mux.scala 27:72]
  wire  _T_4486 = btb_rd_addr_p1_f == 8'ha3; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4835 = _T_4486 ? btb_bank0_rd_data_way0_out_163 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5090 = _T_5089 | _T_4835; // @[Mux.scala 27:72]
  wire  _T_4488 = btb_rd_addr_p1_f == 8'ha4; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4836 = _T_4488 ? btb_bank0_rd_data_way0_out_164 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5091 = _T_5090 | _T_4836; // @[Mux.scala 27:72]
  wire  _T_4490 = btb_rd_addr_p1_f == 8'ha5; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4837 = _T_4490 ? btb_bank0_rd_data_way0_out_165 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5092 = _T_5091 | _T_4837; // @[Mux.scala 27:72]
  wire  _T_4492 = btb_rd_addr_p1_f == 8'ha6; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4838 = _T_4492 ? btb_bank0_rd_data_way0_out_166 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5093 = _T_5092 | _T_4838; // @[Mux.scala 27:72]
  wire  _T_4494 = btb_rd_addr_p1_f == 8'ha7; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4839 = _T_4494 ? btb_bank0_rd_data_way0_out_167 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5094 = _T_5093 | _T_4839; // @[Mux.scala 27:72]
  wire  _T_4496 = btb_rd_addr_p1_f == 8'ha8; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4840 = _T_4496 ? btb_bank0_rd_data_way0_out_168 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5095 = _T_5094 | _T_4840; // @[Mux.scala 27:72]
  wire  _T_4498 = btb_rd_addr_p1_f == 8'ha9; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4841 = _T_4498 ? btb_bank0_rd_data_way0_out_169 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5096 = _T_5095 | _T_4841; // @[Mux.scala 27:72]
  wire  _T_4500 = btb_rd_addr_p1_f == 8'haa; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4842 = _T_4500 ? btb_bank0_rd_data_way0_out_170 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5097 = _T_5096 | _T_4842; // @[Mux.scala 27:72]
  wire  _T_4502 = btb_rd_addr_p1_f == 8'hab; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4843 = _T_4502 ? btb_bank0_rd_data_way0_out_171 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5098 = _T_5097 | _T_4843; // @[Mux.scala 27:72]
  wire  _T_4504 = btb_rd_addr_p1_f == 8'hac; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4844 = _T_4504 ? btb_bank0_rd_data_way0_out_172 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5099 = _T_5098 | _T_4844; // @[Mux.scala 27:72]
  wire  _T_4506 = btb_rd_addr_p1_f == 8'had; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4845 = _T_4506 ? btb_bank0_rd_data_way0_out_173 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5100 = _T_5099 | _T_4845; // @[Mux.scala 27:72]
  wire  _T_4508 = btb_rd_addr_p1_f == 8'hae; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4846 = _T_4508 ? btb_bank0_rd_data_way0_out_174 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5101 = _T_5100 | _T_4846; // @[Mux.scala 27:72]
  wire  _T_4510 = btb_rd_addr_p1_f == 8'haf; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4847 = _T_4510 ? btb_bank0_rd_data_way0_out_175 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5102 = _T_5101 | _T_4847; // @[Mux.scala 27:72]
  wire  _T_4512 = btb_rd_addr_p1_f == 8'hb0; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4848 = _T_4512 ? btb_bank0_rd_data_way0_out_176 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5103 = _T_5102 | _T_4848; // @[Mux.scala 27:72]
  wire  _T_4514 = btb_rd_addr_p1_f == 8'hb1; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4849 = _T_4514 ? btb_bank0_rd_data_way0_out_177 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5104 = _T_5103 | _T_4849; // @[Mux.scala 27:72]
  wire  _T_4516 = btb_rd_addr_p1_f == 8'hb2; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4850 = _T_4516 ? btb_bank0_rd_data_way0_out_178 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5105 = _T_5104 | _T_4850; // @[Mux.scala 27:72]
  wire  _T_4518 = btb_rd_addr_p1_f == 8'hb3; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4851 = _T_4518 ? btb_bank0_rd_data_way0_out_179 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5106 = _T_5105 | _T_4851; // @[Mux.scala 27:72]
  wire  _T_4520 = btb_rd_addr_p1_f == 8'hb4; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4852 = _T_4520 ? btb_bank0_rd_data_way0_out_180 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5107 = _T_5106 | _T_4852; // @[Mux.scala 27:72]
  wire  _T_4522 = btb_rd_addr_p1_f == 8'hb5; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4853 = _T_4522 ? btb_bank0_rd_data_way0_out_181 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5108 = _T_5107 | _T_4853; // @[Mux.scala 27:72]
  wire  _T_4524 = btb_rd_addr_p1_f == 8'hb6; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4854 = _T_4524 ? btb_bank0_rd_data_way0_out_182 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5109 = _T_5108 | _T_4854; // @[Mux.scala 27:72]
  wire  _T_4526 = btb_rd_addr_p1_f == 8'hb7; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4855 = _T_4526 ? btb_bank0_rd_data_way0_out_183 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5110 = _T_5109 | _T_4855; // @[Mux.scala 27:72]
  wire  _T_4528 = btb_rd_addr_p1_f == 8'hb8; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4856 = _T_4528 ? btb_bank0_rd_data_way0_out_184 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5111 = _T_5110 | _T_4856; // @[Mux.scala 27:72]
  wire  _T_4530 = btb_rd_addr_p1_f == 8'hb9; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4857 = _T_4530 ? btb_bank0_rd_data_way0_out_185 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5112 = _T_5111 | _T_4857; // @[Mux.scala 27:72]
  wire  _T_4532 = btb_rd_addr_p1_f == 8'hba; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4858 = _T_4532 ? btb_bank0_rd_data_way0_out_186 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5113 = _T_5112 | _T_4858; // @[Mux.scala 27:72]
  wire  _T_4534 = btb_rd_addr_p1_f == 8'hbb; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4859 = _T_4534 ? btb_bank0_rd_data_way0_out_187 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5114 = _T_5113 | _T_4859; // @[Mux.scala 27:72]
  wire  _T_4536 = btb_rd_addr_p1_f == 8'hbc; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4860 = _T_4536 ? btb_bank0_rd_data_way0_out_188 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5115 = _T_5114 | _T_4860; // @[Mux.scala 27:72]
  wire  _T_4538 = btb_rd_addr_p1_f == 8'hbd; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4861 = _T_4538 ? btb_bank0_rd_data_way0_out_189 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5116 = _T_5115 | _T_4861; // @[Mux.scala 27:72]
  wire  _T_4540 = btb_rd_addr_p1_f == 8'hbe; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4862 = _T_4540 ? btb_bank0_rd_data_way0_out_190 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5117 = _T_5116 | _T_4862; // @[Mux.scala 27:72]
  wire  _T_4542 = btb_rd_addr_p1_f == 8'hbf; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4863 = _T_4542 ? btb_bank0_rd_data_way0_out_191 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5118 = _T_5117 | _T_4863; // @[Mux.scala 27:72]
  wire  _T_4544 = btb_rd_addr_p1_f == 8'hc0; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4864 = _T_4544 ? btb_bank0_rd_data_way0_out_192 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5119 = _T_5118 | _T_4864; // @[Mux.scala 27:72]
  wire  _T_4546 = btb_rd_addr_p1_f == 8'hc1; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4865 = _T_4546 ? btb_bank0_rd_data_way0_out_193 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5120 = _T_5119 | _T_4865; // @[Mux.scala 27:72]
  wire  _T_4548 = btb_rd_addr_p1_f == 8'hc2; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4866 = _T_4548 ? btb_bank0_rd_data_way0_out_194 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5121 = _T_5120 | _T_4866; // @[Mux.scala 27:72]
  wire  _T_4550 = btb_rd_addr_p1_f == 8'hc3; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4867 = _T_4550 ? btb_bank0_rd_data_way0_out_195 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5122 = _T_5121 | _T_4867; // @[Mux.scala 27:72]
  wire  _T_4552 = btb_rd_addr_p1_f == 8'hc4; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4868 = _T_4552 ? btb_bank0_rd_data_way0_out_196 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5123 = _T_5122 | _T_4868; // @[Mux.scala 27:72]
  wire  _T_4554 = btb_rd_addr_p1_f == 8'hc5; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4869 = _T_4554 ? btb_bank0_rd_data_way0_out_197 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5124 = _T_5123 | _T_4869; // @[Mux.scala 27:72]
  wire  _T_4556 = btb_rd_addr_p1_f == 8'hc6; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4870 = _T_4556 ? btb_bank0_rd_data_way0_out_198 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5125 = _T_5124 | _T_4870; // @[Mux.scala 27:72]
  wire  _T_4558 = btb_rd_addr_p1_f == 8'hc7; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4871 = _T_4558 ? btb_bank0_rd_data_way0_out_199 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5126 = _T_5125 | _T_4871; // @[Mux.scala 27:72]
  wire  _T_4560 = btb_rd_addr_p1_f == 8'hc8; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4872 = _T_4560 ? btb_bank0_rd_data_way0_out_200 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5127 = _T_5126 | _T_4872; // @[Mux.scala 27:72]
  wire  _T_4562 = btb_rd_addr_p1_f == 8'hc9; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4873 = _T_4562 ? btb_bank0_rd_data_way0_out_201 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5128 = _T_5127 | _T_4873; // @[Mux.scala 27:72]
  wire  _T_4564 = btb_rd_addr_p1_f == 8'hca; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4874 = _T_4564 ? btb_bank0_rd_data_way0_out_202 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5129 = _T_5128 | _T_4874; // @[Mux.scala 27:72]
  wire  _T_4566 = btb_rd_addr_p1_f == 8'hcb; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4875 = _T_4566 ? btb_bank0_rd_data_way0_out_203 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5130 = _T_5129 | _T_4875; // @[Mux.scala 27:72]
  wire  _T_4568 = btb_rd_addr_p1_f == 8'hcc; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4876 = _T_4568 ? btb_bank0_rd_data_way0_out_204 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5131 = _T_5130 | _T_4876; // @[Mux.scala 27:72]
  wire  _T_4570 = btb_rd_addr_p1_f == 8'hcd; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4877 = _T_4570 ? btb_bank0_rd_data_way0_out_205 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5132 = _T_5131 | _T_4877; // @[Mux.scala 27:72]
  wire  _T_4572 = btb_rd_addr_p1_f == 8'hce; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4878 = _T_4572 ? btb_bank0_rd_data_way0_out_206 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5133 = _T_5132 | _T_4878; // @[Mux.scala 27:72]
  wire  _T_4574 = btb_rd_addr_p1_f == 8'hcf; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4879 = _T_4574 ? btb_bank0_rd_data_way0_out_207 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5134 = _T_5133 | _T_4879; // @[Mux.scala 27:72]
  wire  _T_4576 = btb_rd_addr_p1_f == 8'hd0; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4880 = _T_4576 ? btb_bank0_rd_data_way0_out_208 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5135 = _T_5134 | _T_4880; // @[Mux.scala 27:72]
  wire  _T_4578 = btb_rd_addr_p1_f == 8'hd1; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4881 = _T_4578 ? btb_bank0_rd_data_way0_out_209 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5136 = _T_5135 | _T_4881; // @[Mux.scala 27:72]
  wire  _T_4580 = btb_rd_addr_p1_f == 8'hd2; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4882 = _T_4580 ? btb_bank0_rd_data_way0_out_210 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5137 = _T_5136 | _T_4882; // @[Mux.scala 27:72]
  wire  _T_4582 = btb_rd_addr_p1_f == 8'hd3; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4883 = _T_4582 ? btb_bank0_rd_data_way0_out_211 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5138 = _T_5137 | _T_4883; // @[Mux.scala 27:72]
  wire  _T_4584 = btb_rd_addr_p1_f == 8'hd4; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4884 = _T_4584 ? btb_bank0_rd_data_way0_out_212 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5139 = _T_5138 | _T_4884; // @[Mux.scala 27:72]
  wire  _T_4586 = btb_rd_addr_p1_f == 8'hd5; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4885 = _T_4586 ? btb_bank0_rd_data_way0_out_213 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5140 = _T_5139 | _T_4885; // @[Mux.scala 27:72]
  wire  _T_4588 = btb_rd_addr_p1_f == 8'hd6; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4886 = _T_4588 ? btb_bank0_rd_data_way0_out_214 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5141 = _T_5140 | _T_4886; // @[Mux.scala 27:72]
  wire  _T_4590 = btb_rd_addr_p1_f == 8'hd7; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4887 = _T_4590 ? btb_bank0_rd_data_way0_out_215 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5142 = _T_5141 | _T_4887; // @[Mux.scala 27:72]
  wire  _T_4592 = btb_rd_addr_p1_f == 8'hd8; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4888 = _T_4592 ? btb_bank0_rd_data_way0_out_216 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5143 = _T_5142 | _T_4888; // @[Mux.scala 27:72]
  wire  _T_4594 = btb_rd_addr_p1_f == 8'hd9; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4889 = _T_4594 ? btb_bank0_rd_data_way0_out_217 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5144 = _T_5143 | _T_4889; // @[Mux.scala 27:72]
  wire  _T_4596 = btb_rd_addr_p1_f == 8'hda; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4890 = _T_4596 ? btb_bank0_rd_data_way0_out_218 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5145 = _T_5144 | _T_4890; // @[Mux.scala 27:72]
  wire  _T_4598 = btb_rd_addr_p1_f == 8'hdb; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4891 = _T_4598 ? btb_bank0_rd_data_way0_out_219 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5146 = _T_5145 | _T_4891; // @[Mux.scala 27:72]
  wire  _T_4600 = btb_rd_addr_p1_f == 8'hdc; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4892 = _T_4600 ? btb_bank0_rd_data_way0_out_220 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5147 = _T_5146 | _T_4892; // @[Mux.scala 27:72]
  wire  _T_4602 = btb_rd_addr_p1_f == 8'hdd; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4893 = _T_4602 ? btb_bank0_rd_data_way0_out_221 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5148 = _T_5147 | _T_4893; // @[Mux.scala 27:72]
  wire  _T_4604 = btb_rd_addr_p1_f == 8'hde; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4894 = _T_4604 ? btb_bank0_rd_data_way0_out_222 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5149 = _T_5148 | _T_4894; // @[Mux.scala 27:72]
  wire  _T_4606 = btb_rd_addr_p1_f == 8'hdf; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4895 = _T_4606 ? btb_bank0_rd_data_way0_out_223 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5150 = _T_5149 | _T_4895; // @[Mux.scala 27:72]
  wire  _T_4608 = btb_rd_addr_p1_f == 8'he0; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4896 = _T_4608 ? btb_bank0_rd_data_way0_out_224 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5151 = _T_5150 | _T_4896; // @[Mux.scala 27:72]
  wire  _T_4610 = btb_rd_addr_p1_f == 8'he1; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4897 = _T_4610 ? btb_bank0_rd_data_way0_out_225 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5152 = _T_5151 | _T_4897; // @[Mux.scala 27:72]
  wire  _T_4612 = btb_rd_addr_p1_f == 8'he2; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4898 = _T_4612 ? btb_bank0_rd_data_way0_out_226 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5153 = _T_5152 | _T_4898; // @[Mux.scala 27:72]
  wire  _T_4614 = btb_rd_addr_p1_f == 8'he3; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4899 = _T_4614 ? btb_bank0_rd_data_way0_out_227 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5154 = _T_5153 | _T_4899; // @[Mux.scala 27:72]
  wire  _T_4616 = btb_rd_addr_p1_f == 8'he4; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4900 = _T_4616 ? btb_bank0_rd_data_way0_out_228 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5155 = _T_5154 | _T_4900; // @[Mux.scala 27:72]
  wire  _T_4618 = btb_rd_addr_p1_f == 8'he5; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4901 = _T_4618 ? btb_bank0_rd_data_way0_out_229 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5156 = _T_5155 | _T_4901; // @[Mux.scala 27:72]
  wire  _T_4620 = btb_rd_addr_p1_f == 8'he6; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4902 = _T_4620 ? btb_bank0_rd_data_way0_out_230 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5157 = _T_5156 | _T_4902; // @[Mux.scala 27:72]
  wire  _T_4622 = btb_rd_addr_p1_f == 8'he7; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4903 = _T_4622 ? btb_bank0_rd_data_way0_out_231 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5158 = _T_5157 | _T_4903; // @[Mux.scala 27:72]
  wire  _T_4624 = btb_rd_addr_p1_f == 8'he8; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4904 = _T_4624 ? btb_bank0_rd_data_way0_out_232 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5159 = _T_5158 | _T_4904; // @[Mux.scala 27:72]
  wire  _T_4626 = btb_rd_addr_p1_f == 8'he9; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4905 = _T_4626 ? btb_bank0_rd_data_way0_out_233 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5160 = _T_5159 | _T_4905; // @[Mux.scala 27:72]
  wire  _T_4628 = btb_rd_addr_p1_f == 8'hea; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4906 = _T_4628 ? btb_bank0_rd_data_way0_out_234 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5161 = _T_5160 | _T_4906; // @[Mux.scala 27:72]
  wire  _T_4630 = btb_rd_addr_p1_f == 8'heb; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4907 = _T_4630 ? btb_bank0_rd_data_way0_out_235 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5162 = _T_5161 | _T_4907; // @[Mux.scala 27:72]
  wire  _T_4632 = btb_rd_addr_p1_f == 8'hec; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4908 = _T_4632 ? btb_bank0_rd_data_way0_out_236 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5163 = _T_5162 | _T_4908; // @[Mux.scala 27:72]
  wire  _T_4634 = btb_rd_addr_p1_f == 8'hed; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4909 = _T_4634 ? btb_bank0_rd_data_way0_out_237 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5164 = _T_5163 | _T_4909; // @[Mux.scala 27:72]
  wire  _T_4636 = btb_rd_addr_p1_f == 8'hee; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4910 = _T_4636 ? btb_bank0_rd_data_way0_out_238 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5165 = _T_5164 | _T_4910; // @[Mux.scala 27:72]
  wire  _T_4638 = btb_rd_addr_p1_f == 8'hef; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4911 = _T_4638 ? btb_bank0_rd_data_way0_out_239 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5166 = _T_5165 | _T_4911; // @[Mux.scala 27:72]
  wire  _T_4640 = btb_rd_addr_p1_f == 8'hf0; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4912 = _T_4640 ? btb_bank0_rd_data_way0_out_240 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5167 = _T_5166 | _T_4912; // @[Mux.scala 27:72]
  wire  _T_4642 = btb_rd_addr_p1_f == 8'hf1; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4913 = _T_4642 ? btb_bank0_rd_data_way0_out_241 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5168 = _T_5167 | _T_4913; // @[Mux.scala 27:72]
  wire  _T_4644 = btb_rd_addr_p1_f == 8'hf2; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4914 = _T_4644 ? btb_bank0_rd_data_way0_out_242 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5169 = _T_5168 | _T_4914; // @[Mux.scala 27:72]
  wire  _T_4646 = btb_rd_addr_p1_f == 8'hf3; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4915 = _T_4646 ? btb_bank0_rd_data_way0_out_243 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5170 = _T_5169 | _T_4915; // @[Mux.scala 27:72]
  wire  _T_4648 = btb_rd_addr_p1_f == 8'hf4; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4916 = _T_4648 ? btb_bank0_rd_data_way0_out_244 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5171 = _T_5170 | _T_4916; // @[Mux.scala 27:72]
  wire  _T_4650 = btb_rd_addr_p1_f == 8'hf5; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4917 = _T_4650 ? btb_bank0_rd_data_way0_out_245 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5172 = _T_5171 | _T_4917; // @[Mux.scala 27:72]
  wire  _T_4652 = btb_rd_addr_p1_f == 8'hf6; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4918 = _T_4652 ? btb_bank0_rd_data_way0_out_246 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5173 = _T_5172 | _T_4918; // @[Mux.scala 27:72]
  wire  _T_4654 = btb_rd_addr_p1_f == 8'hf7; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4919 = _T_4654 ? btb_bank0_rd_data_way0_out_247 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5174 = _T_5173 | _T_4919; // @[Mux.scala 27:72]
  wire  _T_4656 = btb_rd_addr_p1_f == 8'hf8; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4920 = _T_4656 ? btb_bank0_rd_data_way0_out_248 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5175 = _T_5174 | _T_4920; // @[Mux.scala 27:72]
  wire  _T_4658 = btb_rd_addr_p1_f == 8'hf9; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4921 = _T_4658 ? btb_bank0_rd_data_way0_out_249 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5176 = _T_5175 | _T_4921; // @[Mux.scala 27:72]
  wire  _T_4660 = btb_rd_addr_p1_f == 8'hfa; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4922 = _T_4660 ? btb_bank0_rd_data_way0_out_250 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5177 = _T_5176 | _T_4922; // @[Mux.scala 27:72]
  wire  _T_4662 = btb_rd_addr_p1_f == 8'hfb; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4923 = _T_4662 ? btb_bank0_rd_data_way0_out_251 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5178 = _T_5177 | _T_4923; // @[Mux.scala 27:72]
  wire  _T_4664 = btb_rd_addr_p1_f == 8'hfc; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4924 = _T_4664 ? btb_bank0_rd_data_way0_out_252 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5179 = _T_5178 | _T_4924; // @[Mux.scala 27:72]
  wire  _T_4666 = btb_rd_addr_p1_f == 8'hfd; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4925 = _T_4666 ? btb_bank0_rd_data_way0_out_253 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5180 = _T_5179 | _T_4925; // @[Mux.scala 27:72]
  wire  _T_4668 = btb_rd_addr_p1_f == 8'hfe; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4926 = _T_4668 ? btb_bank0_rd_data_way0_out_254 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5181 = _T_5180 | _T_4926; // @[Mux.scala 27:72]
  wire  _T_4670 = btb_rd_addr_p1_f == 8'hff; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4927 = _T_4670 ? btb_bank0_rd_data_way0_out_255 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] btb_bank0_rd_data_way0_p1_f = _T_5181 | _T_4927; // @[Mux.scala 27:72]
  wire [4:0] _T_31 = _T_8[13:9] ^ _T_8[18:14]; // @[lib.scala 42:111]
  wire [4:0] fetch_rd_tag_p1_f = _T_31 ^ _T_8[23:19]; // @[lib.scala 42:111]
  wire  _T_64 = btb_bank0_rd_data_way0_p1_f[21:17] == fetch_rd_tag_p1_f; // @[ifu_bp_ctl.scala 135:106]
  wire  _T_65 = btb_bank0_rd_data_way0_p1_f[0] & _T_64; // @[ifu_bp_ctl.scala 135:61]
  wire  _T_20 = io_exu_bp_exu_i0_br_index_r == btb_rd_addr_p1_f; // @[ifu_bp_ctl.scala 103:75]
  wire  branch_error_collision_p1_f = dec_tlu_error_wb & _T_20; // @[ifu_bp_ctl.scala 103:54]
  wire  branch_error_bank_conflict_p1_f = branch_error_collision_p1_f & dec_tlu_error_wb; // @[ifu_bp_ctl.scala 107:69]
  wire  _T_66 = dec_tlu_way_wb_f & branch_error_bank_conflict_p1_f; // @[ifu_bp_ctl.scala 136:24]
  wire  _T_67 = ~_T_66; // @[ifu_bp_ctl.scala 136:5]
  wire  _T_68 = _T_65 & _T_67; // @[ifu_bp_ctl.scala 135:129]
  wire  _T_69 = _T_68 & io_ifc_fetch_req_f; // @[ifu_bp_ctl.scala 136:59]
  wire  tag_match_way0_p1_f = _T_69 & _T; // @[ifu_bp_ctl.scala 136:80]
  wire  _T_100 = btb_bank0_rd_data_way0_p1_f[3] ^ btb_bank0_rd_data_way0_p1_f[4]; // @[ifu_bp_ctl.scala 148:100]
  wire  _T_101 = tag_match_way0_p1_f & _T_100; // @[ifu_bp_ctl.scala 148:62]
  wire  _T_105 = ~_T_100; // @[ifu_bp_ctl.scala 149:64]
  wire  _T_106 = tag_match_way0_p1_f & _T_105; // @[ifu_bp_ctl.scala 149:62]
  wire [1:0] tag_match_way0_expanded_p1_f = {_T_101,_T_106}; // @[Cat.scala 29:58]
  wire [21:0] _T_134 = tag_match_way0_expanded_p1_f[0] ? btb_bank0_rd_data_way0_p1_f : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5696 = _T_4160 ? btb_bank0_rd_data_way1_out_0 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5697 = _T_4162 ? btb_bank0_rd_data_way1_out_1 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5952 = _T_5696 | _T_5697; // @[Mux.scala 27:72]
  wire [21:0] _T_5698 = _T_4164 ? btb_bank0_rd_data_way1_out_2 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5953 = _T_5952 | _T_5698; // @[Mux.scala 27:72]
  wire [21:0] _T_5699 = _T_4166 ? btb_bank0_rd_data_way1_out_3 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5954 = _T_5953 | _T_5699; // @[Mux.scala 27:72]
  wire [21:0] _T_5700 = _T_4168 ? btb_bank0_rd_data_way1_out_4 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5955 = _T_5954 | _T_5700; // @[Mux.scala 27:72]
  wire [21:0] _T_5701 = _T_4170 ? btb_bank0_rd_data_way1_out_5 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5956 = _T_5955 | _T_5701; // @[Mux.scala 27:72]
  wire [21:0] _T_5702 = _T_4172 ? btb_bank0_rd_data_way1_out_6 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5957 = _T_5956 | _T_5702; // @[Mux.scala 27:72]
  wire [21:0] _T_5703 = _T_4174 ? btb_bank0_rd_data_way1_out_7 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5958 = _T_5957 | _T_5703; // @[Mux.scala 27:72]
  wire [21:0] _T_5704 = _T_4176 ? btb_bank0_rd_data_way1_out_8 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5959 = _T_5958 | _T_5704; // @[Mux.scala 27:72]
  wire [21:0] _T_5705 = _T_4178 ? btb_bank0_rd_data_way1_out_9 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5960 = _T_5959 | _T_5705; // @[Mux.scala 27:72]
  wire [21:0] _T_5706 = _T_4180 ? btb_bank0_rd_data_way1_out_10 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5961 = _T_5960 | _T_5706; // @[Mux.scala 27:72]
  wire [21:0] _T_5707 = _T_4182 ? btb_bank0_rd_data_way1_out_11 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5962 = _T_5961 | _T_5707; // @[Mux.scala 27:72]
  wire [21:0] _T_5708 = _T_4184 ? btb_bank0_rd_data_way1_out_12 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5963 = _T_5962 | _T_5708; // @[Mux.scala 27:72]
  wire [21:0] _T_5709 = _T_4186 ? btb_bank0_rd_data_way1_out_13 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5964 = _T_5963 | _T_5709; // @[Mux.scala 27:72]
  wire [21:0] _T_5710 = _T_4188 ? btb_bank0_rd_data_way1_out_14 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5965 = _T_5964 | _T_5710; // @[Mux.scala 27:72]
  wire [21:0] _T_5711 = _T_4190 ? btb_bank0_rd_data_way1_out_15 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5966 = _T_5965 | _T_5711; // @[Mux.scala 27:72]
  wire [21:0] _T_5712 = _T_4192 ? btb_bank0_rd_data_way1_out_16 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5967 = _T_5966 | _T_5712; // @[Mux.scala 27:72]
  wire [21:0] _T_5713 = _T_4194 ? btb_bank0_rd_data_way1_out_17 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5968 = _T_5967 | _T_5713; // @[Mux.scala 27:72]
  wire [21:0] _T_5714 = _T_4196 ? btb_bank0_rd_data_way1_out_18 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5969 = _T_5968 | _T_5714; // @[Mux.scala 27:72]
  wire [21:0] _T_5715 = _T_4198 ? btb_bank0_rd_data_way1_out_19 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5970 = _T_5969 | _T_5715; // @[Mux.scala 27:72]
  wire [21:0] _T_5716 = _T_4200 ? btb_bank0_rd_data_way1_out_20 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5971 = _T_5970 | _T_5716; // @[Mux.scala 27:72]
  wire [21:0] _T_5717 = _T_4202 ? btb_bank0_rd_data_way1_out_21 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5972 = _T_5971 | _T_5717; // @[Mux.scala 27:72]
  wire [21:0] _T_5718 = _T_4204 ? btb_bank0_rd_data_way1_out_22 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5973 = _T_5972 | _T_5718; // @[Mux.scala 27:72]
  wire [21:0] _T_5719 = _T_4206 ? btb_bank0_rd_data_way1_out_23 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5974 = _T_5973 | _T_5719; // @[Mux.scala 27:72]
  wire [21:0] _T_5720 = _T_4208 ? btb_bank0_rd_data_way1_out_24 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5975 = _T_5974 | _T_5720; // @[Mux.scala 27:72]
  wire [21:0] _T_5721 = _T_4210 ? btb_bank0_rd_data_way1_out_25 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5976 = _T_5975 | _T_5721; // @[Mux.scala 27:72]
  wire [21:0] _T_5722 = _T_4212 ? btb_bank0_rd_data_way1_out_26 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5977 = _T_5976 | _T_5722; // @[Mux.scala 27:72]
  wire [21:0] _T_5723 = _T_4214 ? btb_bank0_rd_data_way1_out_27 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5978 = _T_5977 | _T_5723; // @[Mux.scala 27:72]
  wire [21:0] _T_5724 = _T_4216 ? btb_bank0_rd_data_way1_out_28 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5979 = _T_5978 | _T_5724; // @[Mux.scala 27:72]
  wire [21:0] _T_5725 = _T_4218 ? btb_bank0_rd_data_way1_out_29 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5980 = _T_5979 | _T_5725; // @[Mux.scala 27:72]
  wire [21:0] _T_5726 = _T_4220 ? btb_bank0_rd_data_way1_out_30 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5981 = _T_5980 | _T_5726; // @[Mux.scala 27:72]
  wire [21:0] _T_5727 = _T_4222 ? btb_bank0_rd_data_way1_out_31 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5982 = _T_5981 | _T_5727; // @[Mux.scala 27:72]
  wire [21:0] _T_5728 = _T_4224 ? btb_bank0_rd_data_way1_out_32 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5983 = _T_5982 | _T_5728; // @[Mux.scala 27:72]
  wire [21:0] _T_5729 = _T_4226 ? btb_bank0_rd_data_way1_out_33 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5984 = _T_5983 | _T_5729; // @[Mux.scala 27:72]
  wire [21:0] _T_5730 = _T_4228 ? btb_bank0_rd_data_way1_out_34 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5985 = _T_5984 | _T_5730; // @[Mux.scala 27:72]
  wire [21:0] _T_5731 = _T_4230 ? btb_bank0_rd_data_way1_out_35 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5986 = _T_5985 | _T_5731; // @[Mux.scala 27:72]
  wire [21:0] _T_5732 = _T_4232 ? btb_bank0_rd_data_way1_out_36 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5987 = _T_5986 | _T_5732; // @[Mux.scala 27:72]
  wire [21:0] _T_5733 = _T_4234 ? btb_bank0_rd_data_way1_out_37 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5988 = _T_5987 | _T_5733; // @[Mux.scala 27:72]
  wire [21:0] _T_5734 = _T_4236 ? btb_bank0_rd_data_way1_out_38 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5989 = _T_5988 | _T_5734; // @[Mux.scala 27:72]
  wire [21:0] _T_5735 = _T_4238 ? btb_bank0_rd_data_way1_out_39 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5990 = _T_5989 | _T_5735; // @[Mux.scala 27:72]
  wire [21:0] _T_5736 = _T_4240 ? btb_bank0_rd_data_way1_out_40 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5991 = _T_5990 | _T_5736; // @[Mux.scala 27:72]
  wire [21:0] _T_5737 = _T_4242 ? btb_bank0_rd_data_way1_out_41 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5992 = _T_5991 | _T_5737; // @[Mux.scala 27:72]
  wire [21:0] _T_5738 = _T_4244 ? btb_bank0_rd_data_way1_out_42 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5993 = _T_5992 | _T_5738; // @[Mux.scala 27:72]
  wire [21:0] _T_5739 = _T_4246 ? btb_bank0_rd_data_way1_out_43 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5994 = _T_5993 | _T_5739; // @[Mux.scala 27:72]
  wire [21:0] _T_5740 = _T_4248 ? btb_bank0_rd_data_way1_out_44 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5995 = _T_5994 | _T_5740; // @[Mux.scala 27:72]
  wire [21:0] _T_5741 = _T_4250 ? btb_bank0_rd_data_way1_out_45 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5996 = _T_5995 | _T_5741; // @[Mux.scala 27:72]
  wire [21:0] _T_5742 = _T_4252 ? btb_bank0_rd_data_way1_out_46 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5997 = _T_5996 | _T_5742; // @[Mux.scala 27:72]
  wire [21:0] _T_5743 = _T_4254 ? btb_bank0_rd_data_way1_out_47 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5998 = _T_5997 | _T_5743; // @[Mux.scala 27:72]
  wire [21:0] _T_5744 = _T_4256 ? btb_bank0_rd_data_way1_out_48 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5999 = _T_5998 | _T_5744; // @[Mux.scala 27:72]
  wire [21:0] _T_5745 = _T_4258 ? btb_bank0_rd_data_way1_out_49 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6000 = _T_5999 | _T_5745; // @[Mux.scala 27:72]
  wire [21:0] _T_5746 = _T_4260 ? btb_bank0_rd_data_way1_out_50 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6001 = _T_6000 | _T_5746; // @[Mux.scala 27:72]
  wire [21:0] _T_5747 = _T_4262 ? btb_bank0_rd_data_way1_out_51 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6002 = _T_6001 | _T_5747; // @[Mux.scala 27:72]
  wire [21:0] _T_5748 = _T_4264 ? btb_bank0_rd_data_way1_out_52 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6003 = _T_6002 | _T_5748; // @[Mux.scala 27:72]
  wire [21:0] _T_5749 = _T_4266 ? btb_bank0_rd_data_way1_out_53 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6004 = _T_6003 | _T_5749; // @[Mux.scala 27:72]
  wire [21:0] _T_5750 = _T_4268 ? btb_bank0_rd_data_way1_out_54 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6005 = _T_6004 | _T_5750; // @[Mux.scala 27:72]
  wire [21:0] _T_5751 = _T_4270 ? btb_bank0_rd_data_way1_out_55 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6006 = _T_6005 | _T_5751; // @[Mux.scala 27:72]
  wire [21:0] _T_5752 = _T_4272 ? btb_bank0_rd_data_way1_out_56 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6007 = _T_6006 | _T_5752; // @[Mux.scala 27:72]
  wire [21:0] _T_5753 = _T_4274 ? btb_bank0_rd_data_way1_out_57 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6008 = _T_6007 | _T_5753; // @[Mux.scala 27:72]
  wire [21:0] _T_5754 = _T_4276 ? btb_bank0_rd_data_way1_out_58 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6009 = _T_6008 | _T_5754; // @[Mux.scala 27:72]
  wire [21:0] _T_5755 = _T_4278 ? btb_bank0_rd_data_way1_out_59 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6010 = _T_6009 | _T_5755; // @[Mux.scala 27:72]
  wire [21:0] _T_5756 = _T_4280 ? btb_bank0_rd_data_way1_out_60 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6011 = _T_6010 | _T_5756; // @[Mux.scala 27:72]
  wire [21:0] _T_5757 = _T_4282 ? btb_bank0_rd_data_way1_out_61 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6012 = _T_6011 | _T_5757; // @[Mux.scala 27:72]
  wire [21:0] _T_5758 = _T_4284 ? btb_bank0_rd_data_way1_out_62 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6013 = _T_6012 | _T_5758; // @[Mux.scala 27:72]
  wire [21:0] _T_5759 = _T_4286 ? btb_bank0_rd_data_way1_out_63 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6014 = _T_6013 | _T_5759; // @[Mux.scala 27:72]
  wire [21:0] _T_5760 = _T_4288 ? btb_bank0_rd_data_way1_out_64 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6015 = _T_6014 | _T_5760; // @[Mux.scala 27:72]
  wire [21:0] _T_5761 = _T_4290 ? btb_bank0_rd_data_way1_out_65 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6016 = _T_6015 | _T_5761; // @[Mux.scala 27:72]
  wire [21:0] _T_5762 = _T_4292 ? btb_bank0_rd_data_way1_out_66 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6017 = _T_6016 | _T_5762; // @[Mux.scala 27:72]
  wire [21:0] _T_5763 = _T_4294 ? btb_bank0_rd_data_way1_out_67 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6018 = _T_6017 | _T_5763; // @[Mux.scala 27:72]
  wire [21:0] _T_5764 = _T_4296 ? btb_bank0_rd_data_way1_out_68 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6019 = _T_6018 | _T_5764; // @[Mux.scala 27:72]
  wire [21:0] _T_5765 = _T_4298 ? btb_bank0_rd_data_way1_out_69 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6020 = _T_6019 | _T_5765; // @[Mux.scala 27:72]
  wire [21:0] _T_5766 = _T_4300 ? btb_bank0_rd_data_way1_out_70 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6021 = _T_6020 | _T_5766; // @[Mux.scala 27:72]
  wire [21:0] _T_5767 = _T_4302 ? btb_bank0_rd_data_way1_out_71 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6022 = _T_6021 | _T_5767; // @[Mux.scala 27:72]
  wire [21:0] _T_5768 = _T_4304 ? btb_bank0_rd_data_way1_out_72 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6023 = _T_6022 | _T_5768; // @[Mux.scala 27:72]
  wire [21:0] _T_5769 = _T_4306 ? btb_bank0_rd_data_way1_out_73 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6024 = _T_6023 | _T_5769; // @[Mux.scala 27:72]
  wire [21:0] _T_5770 = _T_4308 ? btb_bank0_rd_data_way1_out_74 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6025 = _T_6024 | _T_5770; // @[Mux.scala 27:72]
  wire [21:0] _T_5771 = _T_4310 ? btb_bank0_rd_data_way1_out_75 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6026 = _T_6025 | _T_5771; // @[Mux.scala 27:72]
  wire [21:0] _T_5772 = _T_4312 ? btb_bank0_rd_data_way1_out_76 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6027 = _T_6026 | _T_5772; // @[Mux.scala 27:72]
  wire [21:0] _T_5773 = _T_4314 ? btb_bank0_rd_data_way1_out_77 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6028 = _T_6027 | _T_5773; // @[Mux.scala 27:72]
  wire [21:0] _T_5774 = _T_4316 ? btb_bank0_rd_data_way1_out_78 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6029 = _T_6028 | _T_5774; // @[Mux.scala 27:72]
  wire [21:0] _T_5775 = _T_4318 ? btb_bank0_rd_data_way1_out_79 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6030 = _T_6029 | _T_5775; // @[Mux.scala 27:72]
  wire [21:0] _T_5776 = _T_4320 ? btb_bank0_rd_data_way1_out_80 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6031 = _T_6030 | _T_5776; // @[Mux.scala 27:72]
  wire [21:0] _T_5777 = _T_4322 ? btb_bank0_rd_data_way1_out_81 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6032 = _T_6031 | _T_5777; // @[Mux.scala 27:72]
  wire [21:0] _T_5778 = _T_4324 ? btb_bank0_rd_data_way1_out_82 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6033 = _T_6032 | _T_5778; // @[Mux.scala 27:72]
  wire [21:0] _T_5779 = _T_4326 ? btb_bank0_rd_data_way1_out_83 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6034 = _T_6033 | _T_5779; // @[Mux.scala 27:72]
  wire [21:0] _T_5780 = _T_4328 ? btb_bank0_rd_data_way1_out_84 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6035 = _T_6034 | _T_5780; // @[Mux.scala 27:72]
  wire [21:0] _T_5781 = _T_4330 ? btb_bank0_rd_data_way1_out_85 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6036 = _T_6035 | _T_5781; // @[Mux.scala 27:72]
  wire [21:0] _T_5782 = _T_4332 ? btb_bank0_rd_data_way1_out_86 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6037 = _T_6036 | _T_5782; // @[Mux.scala 27:72]
  wire [21:0] _T_5783 = _T_4334 ? btb_bank0_rd_data_way1_out_87 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6038 = _T_6037 | _T_5783; // @[Mux.scala 27:72]
  wire [21:0] _T_5784 = _T_4336 ? btb_bank0_rd_data_way1_out_88 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6039 = _T_6038 | _T_5784; // @[Mux.scala 27:72]
  wire [21:0] _T_5785 = _T_4338 ? btb_bank0_rd_data_way1_out_89 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6040 = _T_6039 | _T_5785; // @[Mux.scala 27:72]
  wire [21:0] _T_5786 = _T_4340 ? btb_bank0_rd_data_way1_out_90 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6041 = _T_6040 | _T_5786; // @[Mux.scala 27:72]
  wire [21:0] _T_5787 = _T_4342 ? btb_bank0_rd_data_way1_out_91 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6042 = _T_6041 | _T_5787; // @[Mux.scala 27:72]
  wire [21:0] _T_5788 = _T_4344 ? btb_bank0_rd_data_way1_out_92 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6043 = _T_6042 | _T_5788; // @[Mux.scala 27:72]
  wire [21:0] _T_5789 = _T_4346 ? btb_bank0_rd_data_way1_out_93 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6044 = _T_6043 | _T_5789; // @[Mux.scala 27:72]
  wire [21:0] _T_5790 = _T_4348 ? btb_bank0_rd_data_way1_out_94 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6045 = _T_6044 | _T_5790; // @[Mux.scala 27:72]
  wire [21:0] _T_5791 = _T_4350 ? btb_bank0_rd_data_way1_out_95 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6046 = _T_6045 | _T_5791; // @[Mux.scala 27:72]
  wire [21:0] _T_5792 = _T_4352 ? btb_bank0_rd_data_way1_out_96 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6047 = _T_6046 | _T_5792; // @[Mux.scala 27:72]
  wire [21:0] _T_5793 = _T_4354 ? btb_bank0_rd_data_way1_out_97 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6048 = _T_6047 | _T_5793; // @[Mux.scala 27:72]
  wire [21:0] _T_5794 = _T_4356 ? btb_bank0_rd_data_way1_out_98 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6049 = _T_6048 | _T_5794; // @[Mux.scala 27:72]
  wire [21:0] _T_5795 = _T_4358 ? btb_bank0_rd_data_way1_out_99 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6050 = _T_6049 | _T_5795; // @[Mux.scala 27:72]
  wire [21:0] _T_5796 = _T_4360 ? btb_bank0_rd_data_way1_out_100 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6051 = _T_6050 | _T_5796; // @[Mux.scala 27:72]
  wire [21:0] _T_5797 = _T_4362 ? btb_bank0_rd_data_way1_out_101 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6052 = _T_6051 | _T_5797; // @[Mux.scala 27:72]
  wire [21:0] _T_5798 = _T_4364 ? btb_bank0_rd_data_way1_out_102 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6053 = _T_6052 | _T_5798; // @[Mux.scala 27:72]
  wire [21:0] _T_5799 = _T_4366 ? btb_bank0_rd_data_way1_out_103 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6054 = _T_6053 | _T_5799; // @[Mux.scala 27:72]
  wire [21:0] _T_5800 = _T_4368 ? btb_bank0_rd_data_way1_out_104 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6055 = _T_6054 | _T_5800; // @[Mux.scala 27:72]
  wire [21:0] _T_5801 = _T_4370 ? btb_bank0_rd_data_way1_out_105 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6056 = _T_6055 | _T_5801; // @[Mux.scala 27:72]
  wire [21:0] _T_5802 = _T_4372 ? btb_bank0_rd_data_way1_out_106 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6057 = _T_6056 | _T_5802; // @[Mux.scala 27:72]
  wire [21:0] _T_5803 = _T_4374 ? btb_bank0_rd_data_way1_out_107 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6058 = _T_6057 | _T_5803; // @[Mux.scala 27:72]
  wire [21:0] _T_5804 = _T_4376 ? btb_bank0_rd_data_way1_out_108 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6059 = _T_6058 | _T_5804; // @[Mux.scala 27:72]
  wire [21:0] _T_5805 = _T_4378 ? btb_bank0_rd_data_way1_out_109 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6060 = _T_6059 | _T_5805; // @[Mux.scala 27:72]
  wire [21:0] _T_5806 = _T_4380 ? btb_bank0_rd_data_way1_out_110 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6061 = _T_6060 | _T_5806; // @[Mux.scala 27:72]
  wire [21:0] _T_5807 = _T_4382 ? btb_bank0_rd_data_way1_out_111 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6062 = _T_6061 | _T_5807; // @[Mux.scala 27:72]
  wire [21:0] _T_5808 = _T_4384 ? btb_bank0_rd_data_way1_out_112 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6063 = _T_6062 | _T_5808; // @[Mux.scala 27:72]
  wire [21:0] _T_5809 = _T_4386 ? btb_bank0_rd_data_way1_out_113 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6064 = _T_6063 | _T_5809; // @[Mux.scala 27:72]
  wire [21:0] _T_5810 = _T_4388 ? btb_bank0_rd_data_way1_out_114 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6065 = _T_6064 | _T_5810; // @[Mux.scala 27:72]
  wire [21:0] _T_5811 = _T_4390 ? btb_bank0_rd_data_way1_out_115 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6066 = _T_6065 | _T_5811; // @[Mux.scala 27:72]
  wire [21:0] _T_5812 = _T_4392 ? btb_bank0_rd_data_way1_out_116 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6067 = _T_6066 | _T_5812; // @[Mux.scala 27:72]
  wire [21:0] _T_5813 = _T_4394 ? btb_bank0_rd_data_way1_out_117 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6068 = _T_6067 | _T_5813; // @[Mux.scala 27:72]
  wire [21:0] _T_5814 = _T_4396 ? btb_bank0_rd_data_way1_out_118 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6069 = _T_6068 | _T_5814; // @[Mux.scala 27:72]
  wire [21:0] _T_5815 = _T_4398 ? btb_bank0_rd_data_way1_out_119 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6070 = _T_6069 | _T_5815; // @[Mux.scala 27:72]
  wire [21:0] _T_5816 = _T_4400 ? btb_bank0_rd_data_way1_out_120 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6071 = _T_6070 | _T_5816; // @[Mux.scala 27:72]
  wire [21:0] _T_5817 = _T_4402 ? btb_bank0_rd_data_way1_out_121 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6072 = _T_6071 | _T_5817; // @[Mux.scala 27:72]
  wire [21:0] _T_5818 = _T_4404 ? btb_bank0_rd_data_way1_out_122 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6073 = _T_6072 | _T_5818; // @[Mux.scala 27:72]
  wire [21:0] _T_5819 = _T_4406 ? btb_bank0_rd_data_way1_out_123 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6074 = _T_6073 | _T_5819; // @[Mux.scala 27:72]
  wire [21:0] _T_5820 = _T_4408 ? btb_bank0_rd_data_way1_out_124 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6075 = _T_6074 | _T_5820; // @[Mux.scala 27:72]
  wire [21:0] _T_5821 = _T_4410 ? btb_bank0_rd_data_way1_out_125 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6076 = _T_6075 | _T_5821; // @[Mux.scala 27:72]
  wire [21:0] _T_5822 = _T_4412 ? btb_bank0_rd_data_way1_out_126 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6077 = _T_6076 | _T_5822; // @[Mux.scala 27:72]
  wire [21:0] _T_5823 = _T_4414 ? btb_bank0_rd_data_way1_out_127 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6078 = _T_6077 | _T_5823; // @[Mux.scala 27:72]
  wire [21:0] _T_5824 = _T_4416 ? btb_bank0_rd_data_way1_out_128 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6079 = _T_6078 | _T_5824; // @[Mux.scala 27:72]
  wire [21:0] _T_5825 = _T_4418 ? btb_bank0_rd_data_way1_out_129 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6080 = _T_6079 | _T_5825; // @[Mux.scala 27:72]
  wire [21:0] _T_5826 = _T_4420 ? btb_bank0_rd_data_way1_out_130 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6081 = _T_6080 | _T_5826; // @[Mux.scala 27:72]
  wire [21:0] _T_5827 = _T_4422 ? btb_bank0_rd_data_way1_out_131 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6082 = _T_6081 | _T_5827; // @[Mux.scala 27:72]
  wire [21:0] _T_5828 = _T_4424 ? btb_bank0_rd_data_way1_out_132 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6083 = _T_6082 | _T_5828; // @[Mux.scala 27:72]
  wire [21:0] _T_5829 = _T_4426 ? btb_bank0_rd_data_way1_out_133 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6084 = _T_6083 | _T_5829; // @[Mux.scala 27:72]
  wire [21:0] _T_5830 = _T_4428 ? btb_bank0_rd_data_way1_out_134 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6085 = _T_6084 | _T_5830; // @[Mux.scala 27:72]
  wire [21:0] _T_5831 = _T_4430 ? btb_bank0_rd_data_way1_out_135 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6086 = _T_6085 | _T_5831; // @[Mux.scala 27:72]
  wire [21:0] _T_5832 = _T_4432 ? btb_bank0_rd_data_way1_out_136 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6087 = _T_6086 | _T_5832; // @[Mux.scala 27:72]
  wire [21:0] _T_5833 = _T_4434 ? btb_bank0_rd_data_way1_out_137 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6088 = _T_6087 | _T_5833; // @[Mux.scala 27:72]
  wire [21:0] _T_5834 = _T_4436 ? btb_bank0_rd_data_way1_out_138 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6089 = _T_6088 | _T_5834; // @[Mux.scala 27:72]
  wire [21:0] _T_5835 = _T_4438 ? btb_bank0_rd_data_way1_out_139 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6090 = _T_6089 | _T_5835; // @[Mux.scala 27:72]
  wire [21:0] _T_5836 = _T_4440 ? btb_bank0_rd_data_way1_out_140 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6091 = _T_6090 | _T_5836; // @[Mux.scala 27:72]
  wire [21:0] _T_5837 = _T_4442 ? btb_bank0_rd_data_way1_out_141 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6092 = _T_6091 | _T_5837; // @[Mux.scala 27:72]
  wire [21:0] _T_5838 = _T_4444 ? btb_bank0_rd_data_way1_out_142 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6093 = _T_6092 | _T_5838; // @[Mux.scala 27:72]
  wire [21:0] _T_5839 = _T_4446 ? btb_bank0_rd_data_way1_out_143 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6094 = _T_6093 | _T_5839; // @[Mux.scala 27:72]
  wire [21:0] _T_5840 = _T_4448 ? btb_bank0_rd_data_way1_out_144 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6095 = _T_6094 | _T_5840; // @[Mux.scala 27:72]
  wire [21:0] _T_5841 = _T_4450 ? btb_bank0_rd_data_way1_out_145 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6096 = _T_6095 | _T_5841; // @[Mux.scala 27:72]
  wire [21:0] _T_5842 = _T_4452 ? btb_bank0_rd_data_way1_out_146 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6097 = _T_6096 | _T_5842; // @[Mux.scala 27:72]
  wire [21:0] _T_5843 = _T_4454 ? btb_bank0_rd_data_way1_out_147 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6098 = _T_6097 | _T_5843; // @[Mux.scala 27:72]
  wire [21:0] _T_5844 = _T_4456 ? btb_bank0_rd_data_way1_out_148 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6099 = _T_6098 | _T_5844; // @[Mux.scala 27:72]
  wire [21:0] _T_5845 = _T_4458 ? btb_bank0_rd_data_way1_out_149 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6100 = _T_6099 | _T_5845; // @[Mux.scala 27:72]
  wire [21:0] _T_5846 = _T_4460 ? btb_bank0_rd_data_way1_out_150 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6101 = _T_6100 | _T_5846; // @[Mux.scala 27:72]
  wire [21:0] _T_5847 = _T_4462 ? btb_bank0_rd_data_way1_out_151 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6102 = _T_6101 | _T_5847; // @[Mux.scala 27:72]
  wire [21:0] _T_5848 = _T_4464 ? btb_bank0_rd_data_way1_out_152 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6103 = _T_6102 | _T_5848; // @[Mux.scala 27:72]
  wire [21:0] _T_5849 = _T_4466 ? btb_bank0_rd_data_way1_out_153 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6104 = _T_6103 | _T_5849; // @[Mux.scala 27:72]
  wire [21:0] _T_5850 = _T_4468 ? btb_bank0_rd_data_way1_out_154 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6105 = _T_6104 | _T_5850; // @[Mux.scala 27:72]
  wire [21:0] _T_5851 = _T_4470 ? btb_bank0_rd_data_way1_out_155 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6106 = _T_6105 | _T_5851; // @[Mux.scala 27:72]
  wire [21:0] _T_5852 = _T_4472 ? btb_bank0_rd_data_way1_out_156 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6107 = _T_6106 | _T_5852; // @[Mux.scala 27:72]
  wire [21:0] _T_5853 = _T_4474 ? btb_bank0_rd_data_way1_out_157 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6108 = _T_6107 | _T_5853; // @[Mux.scala 27:72]
  wire [21:0] _T_5854 = _T_4476 ? btb_bank0_rd_data_way1_out_158 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6109 = _T_6108 | _T_5854; // @[Mux.scala 27:72]
  wire [21:0] _T_5855 = _T_4478 ? btb_bank0_rd_data_way1_out_159 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6110 = _T_6109 | _T_5855; // @[Mux.scala 27:72]
  wire [21:0] _T_5856 = _T_4480 ? btb_bank0_rd_data_way1_out_160 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6111 = _T_6110 | _T_5856; // @[Mux.scala 27:72]
  wire [21:0] _T_5857 = _T_4482 ? btb_bank0_rd_data_way1_out_161 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6112 = _T_6111 | _T_5857; // @[Mux.scala 27:72]
  wire [21:0] _T_5858 = _T_4484 ? btb_bank0_rd_data_way1_out_162 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6113 = _T_6112 | _T_5858; // @[Mux.scala 27:72]
  wire [21:0] _T_5859 = _T_4486 ? btb_bank0_rd_data_way1_out_163 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6114 = _T_6113 | _T_5859; // @[Mux.scala 27:72]
  wire [21:0] _T_5860 = _T_4488 ? btb_bank0_rd_data_way1_out_164 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6115 = _T_6114 | _T_5860; // @[Mux.scala 27:72]
  wire [21:0] _T_5861 = _T_4490 ? btb_bank0_rd_data_way1_out_165 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6116 = _T_6115 | _T_5861; // @[Mux.scala 27:72]
  wire [21:0] _T_5862 = _T_4492 ? btb_bank0_rd_data_way1_out_166 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6117 = _T_6116 | _T_5862; // @[Mux.scala 27:72]
  wire [21:0] _T_5863 = _T_4494 ? btb_bank0_rd_data_way1_out_167 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6118 = _T_6117 | _T_5863; // @[Mux.scala 27:72]
  wire [21:0] _T_5864 = _T_4496 ? btb_bank0_rd_data_way1_out_168 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6119 = _T_6118 | _T_5864; // @[Mux.scala 27:72]
  wire [21:0] _T_5865 = _T_4498 ? btb_bank0_rd_data_way1_out_169 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6120 = _T_6119 | _T_5865; // @[Mux.scala 27:72]
  wire [21:0] _T_5866 = _T_4500 ? btb_bank0_rd_data_way1_out_170 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6121 = _T_6120 | _T_5866; // @[Mux.scala 27:72]
  wire [21:0] _T_5867 = _T_4502 ? btb_bank0_rd_data_way1_out_171 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6122 = _T_6121 | _T_5867; // @[Mux.scala 27:72]
  wire [21:0] _T_5868 = _T_4504 ? btb_bank0_rd_data_way1_out_172 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6123 = _T_6122 | _T_5868; // @[Mux.scala 27:72]
  wire [21:0] _T_5869 = _T_4506 ? btb_bank0_rd_data_way1_out_173 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6124 = _T_6123 | _T_5869; // @[Mux.scala 27:72]
  wire [21:0] _T_5870 = _T_4508 ? btb_bank0_rd_data_way1_out_174 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6125 = _T_6124 | _T_5870; // @[Mux.scala 27:72]
  wire [21:0] _T_5871 = _T_4510 ? btb_bank0_rd_data_way1_out_175 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6126 = _T_6125 | _T_5871; // @[Mux.scala 27:72]
  wire [21:0] _T_5872 = _T_4512 ? btb_bank0_rd_data_way1_out_176 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6127 = _T_6126 | _T_5872; // @[Mux.scala 27:72]
  wire [21:0] _T_5873 = _T_4514 ? btb_bank0_rd_data_way1_out_177 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6128 = _T_6127 | _T_5873; // @[Mux.scala 27:72]
  wire [21:0] _T_5874 = _T_4516 ? btb_bank0_rd_data_way1_out_178 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6129 = _T_6128 | _T_5874; // @[Mux.scala 27:72]
  wire [21:0] _T_5875 = _T_4518 ? btb_bank0_rd_data_way1_out_179 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6130 = _T_6129 | _T_5875; // @[Mux.scala 27:72]
  wire [21:0] _T_5876 = _T_4520 ? btb_bank0_rd_data_way1_out_180 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6131 = _T_6130 | _T_5876; // @[Mux.scala 27:72]
  wire [21:0] _T_5877 = _T_4522 ? btb_bank0_rd_data_way1_out_181 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6132 = _T_6131 | _T_5877; // @[Mux.scala 27:72]
  wire [21:0] _T_5878 = _T_4524 ? btb_bank0_rd_data_way1_out_182 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6133 = _T_6132 | _T_5878; // @[Mux.scala 27:72]
  wire [21:0] _T_5879 = _T_4526 ? btb_bank0_rd_data_way1_out_183 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6134 = _T_6133 | _T_5879; // @[Mux.scala 27:72]
  wire [21:0] _T_5880 = _T_4528 ? btb_bank0_rd_data_way1_out_184 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6135 = _T_6134 | _T_5880; // @[Mux.scala 27:72]
  wire [21:0] _T_5881 = _T_4530 ? btb_bank0_rd_data_way1_out_185 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6136 = _T_6135 | _T_5881; // @[Mux.scala 27:72]
  wire [21:0] _T_5882 = _T_4532 ? btb_bank0_rd_data_way1_out_186 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6137 = _T_6136 | _T_5882; // @[Mux.scala 27:72]
  wire [21:0] _T_5883 = _T_4534 ? btb_bank0_rd_data_way1_out_187 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6138 = _T_6137 | _T_5883; // @[Mux.scala 27:72]
  wire [21:0] _T_5884 = _T_4536 ? btb_bank0_rd_data_way1_out_188 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6139 = _T_6138 | _T_5884; // @[Mux.scala 27:72]
  wire [21:0] _T_5885 = _T_4538 ? btb_bank0_rd_data_way1_out_189 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6140 = _T_6139 | _T_5885; // @[Mux.scala 27:72]
  wire [21:0] _T_5886 = _T_4540 ? btb_bank0_rd_data_way1_out_190 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6141 = _T_6140 | _T_5886; // @[Mux.scala 27:72]
  wire [21:0] _T_5887 = _T_4542 ? btb_bank0_rd_data_way1_out_191 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6142 = _T_6141 | _T_5887; // @[Mux.scala 27:72]
  wire [21:0] _T_5888 = _T_4544 ? btb_bank0_rd_data_way1_out_192 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6143 = _T_6142 | _T_5888; // @[Mux.scala 27:72]
  wire [21:0] _T_5889 = _T_4546 ? btb_bank0_rd_data_way1_out_193 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6144 = _T_6143 | _T_5889; // @[Mux.scala 27:72]
  wire [21:0] _T_5890 = _T_4548 ? btb_bank0_rd_data_way1_out_194 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6145 = _T_6144 | _T_5890; // @[Mux.scala 27:72]
  wire [21:0] _T_5891 = _T_4550 ? btb_bank0_rd_data_way1_out_195 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6146 = _T_6145 | _T_5891; // @[Mux.scala 27:72]
  wire [21:0] _T_5892 = _T_4552 ? btb_bank0_rd_data_way1_out_196 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6147 = _T_6146 | _T_5892; // @[Mux.scala 27:72]
  wire [21:0] _T_5893 = _T_4554 ? btb_bank0_rd_data_way1_out_197 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6148 = _T_6147 | _T_5893; // @[Mux.scala 27:72]
  wire [21:0] _T_5894 = _T_4556 ? btb_bank0_rd_data_way1_out_198 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6149 = _T_6148 | _T_5894; // @[Mux.scala 27:72]
  wire [21:0] _T_5895 = _T_4558 ? btb_bank0_rd_data_way1_out_199 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6150 = _T_6149 | _T_5895; // @[Mux.scala 27:72]
  wire [21:0] _T_5896 = _T_4560 ? btb_bank0_rd_data_way1_out_200 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6151 = _T_6150 | _T_5896; // @[Mux.scala 27:72]
  wire [21:0] _T_5897 = _T_4562 ? btb_bank0_rd_data_way1_out_201 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6152 = _T_6151 | _T_5897; // @[Mux.scala 27:72]
  wire [21:0] _T_5898 = _T_4564 ? btb_bank0_rd_data_way1_out_202 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6153 = _T_6152 | _T_5898; // @[Mux.scala 27:72]
  wire [21:0] _T_5899 = _T_4566 ? btb_bank0_rd_data_way1_out_203 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6154 = _T_6153 | _T_5899; // @[Mux.scala 27:72]
  wire [21:0] _T_5900 = _T_4568 ? btb_bank0_rd_data_way1_out_204 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6155 = _T_6154 | _T_5900; // @[Mux.scala 27:72]
  wire [21:0] _T_5901 = _T_4570 ? btb_bank0_rd_data_way1_out_205 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6156 = _T_6155 | _T_5901; // @[Mux.scala 27:72]
  wire [21:0] _T_5902 = _T_4572 ? btb_bank0_rd_data_way1_out_206 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6157 = _T_6156 | _T_5902; // @[Mux.scala 27:72]
  wire [21:0] _T_5903 = _T_4574 ? btb_bank0_rd_data_way1_out_207 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6158 = _T_6157 | _T_5903; // @[Mux.scala 27:72]
  wire [21:0] _T_5904 = _T_4576 ? btb_bank0_rd_data_way1_out_208 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6159 = _T_6158 | _T_5904; // @[Mux.scala 27:72]
  wire [21:0] _T_5905 = _T_4578 ? btb_bank0_rd_data_way1_out_209 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6160 = _T_6159 | _T_5905; // @[Mux.scala 27:72]
  wire [21:0] _T_5906 = _T_4580 ? btb_bank0_rd_data_way1_out_210 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6161 = _T_6160 | _T_5906; // @[Mux.scala 27:72]
  wire [21:0] _T_5907 = _T_4582 ? btb_bank0_rd_data_way1_out_211 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6162 = _T_6161 | _T_5907; // @[Mux.scala 27:72]
  wire [21:0] _T_5908 = _T_4584 ? btb_bank0_rd_data_way1_out_212 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6163 = _T_6162 | _T_5908; // @[Mux.scala 27:72]
  wire [21:0] _T_5909 = _T_4586 ? btb_bank0_rd_data_way1_out_213 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6164 = _T_6163 | _T_5909; // @[Mux.scala 27:72]
  wire [21:0] _T_5910 = _T_4588 ? btb_bank0_rd_data_way1_out_214 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6165 = _T_6164 | _T_5910; // @[Mux.scala 27:72]
  wire [21:0] _T_5911 = _T_4590 ? btb_bank0_rd_data_way1_out_215 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6166 = _T_6165 | _T_5911; // @[Mux.scala 27:72]
  wire [21:0] _T_5912 = _T_4592 ? btb_bank0_rd_data_way1_out_216 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6167 = _T_6166 | _T_5912; // @[Mux.scala 27:72]
  wire [21:0] _T_5913 = _T_4594 ? btb_bank0_rd_data_way1_out_217 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6168 = _T_6167 | _T_5913; // @[Mux.scala 27:72]
  wire [21:0] _T_5914 = _T_4596 ? btb_bank0_rd_data_way1_out_218 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6169 = _T_6168 | _T_5914; // @[Mux.scala 27:72]
  wire [21:0] _T_5915 = _T_4598 ? btb_bank0_rd_data_way1_out_219 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6170 = _T_6169 | _T_5915; // @[Mux.scala 27:72]
  wire [21:0] _T_5916 = _T_4600 ? btb_bank0_rd_data_way1_out_220 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6171 = _T_6170 | _T_5916; // @[Mux.scala 27:72]
  wire [21:0] _T_5917 = _T_4602 ? btb_bank0_rd_data_way1_out_221 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6172 = _T_6171 | _T_5917; // @[Mux.scala 27:72]
  wire [21:0] _T_5918 = _T_4604 ? btb_bank0_rd_data_way1_out_222 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6173 = _T_6172 | _T_5918; // @[Mux.scala 27:72]
  wire [21:0] _T_5919 = _T_4606 ? btb_bank0_rd_data_way1_out_223 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6174 = _T_6173 | _T_5919; // @[Mux.scala 27:72]
  wire [21:0] _T_5920 = _T_4608 ? btb_bank0_rd_data_way1_out_224 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6175 = _T_6174 | _T_5920; // @[Mux.scala 27:72]
  wire [21:0] _T_5921 = _T_4610 ? btb_bank0_rd_data_way1_out_225 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6176 = _T_6175 | _T_5921; // @[Mux.scala 27:72]
  wire [21:0] _T_5922 = _T_4612 ? btb_bank0_rd_data_way1_out_226 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6177 = _T_6176 | _T_5922; // @[Mux.scala 27:72]
  wire [21:0] _T_5923 = _T_4614 ? btb_bank0_rd_data_way1_out_227 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6178 = _T_6177 | _T_5923; // @[Mux.scala 27:72]
  wire [21:0] _T_5924 = _T_4616 ? btb_bank0_rd_data_way1_out_228 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6179 = _T_6178 | _T_5924; // @[Mux.scala 27:72]
  wire [21:0] _T_5925 = _T_4618 ? btb_bank0_rd_data_way1_out_229 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6180 = _T_6179 | _T_5925; // @[Mux.scala 27:72]
  wire [21:0] _T_5926 = _T_4620 ? btb_bank0_rd_data_way1_out_230 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6181 = _T_6180 | _T_5926; // @[Mux.scala 27:72]
  wire [21:0] _T_5927 = _T_4622 ? btb_bank0_rd_data_way1_out_231 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6182 = _T_6181 | _T_5927; // @[Mux.scala 27:72]
  wire [21:0] _T_5928 = _T_4624 ? btb_bank0_rd_data_way1_out_232 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6183 = _T_6182 | _T_5928; // @[Mux.scala 27:72]
  wire [21:0] _T_5929 = _T_4626 ? btb_bank0_rd_data_way1_out_233 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6184 = _T_6183 | _T_5929; // @[Mux.scala 27:72]
  wire [21:0] _T_5930 = _T_4628 ? btb_bank0_rd_data_way1_out_234 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6185 = _T_6184 | _T_5930; // @[Mux.scala 27:72]
  wire [21:0] _T_5931 = _T_4630 ? btb_bank0_rd_data_way1_out_235 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6186 = _T_6185 | _T_5931; // @[Mux.scala 27:72]
  wire [21:0] _T_5932 = _T_4632 ? btb_bank0_rd_data_way1_out_236 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6187 = _T_6186 | _T_5932; // @[Mux.scala 27:72]
  wire [21:0] _T_5933 = _T_4634 ? btb_bank0_rd_data_way1_out_237 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6188 = _T_6187 | _T_5933; // @[Mux.scala 27:72]
  wire [21:0] _T_5934 = _T_4636 ? btb_bank0_rd_data_way1_out_238 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6189 = _T_6188 | _T_5934; // @[Mux.scala 27:72]
  wire [21:0] _T_5935 = _T_4638 ? btb_bank0_rd_data_way1_out_239 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6190 = _T_6189 | _T_5935; // @[Mux.scala 27:72]
  wire [21:0] _T_5936 = _T_4640 ? btb_bank0_rd_data_way1_out_240 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6191 = _T_6190 | _T_5936; // @[Mux.scala 27:72]
  wire [21:0] _T_5937 = _T_4642 ? btb_bank0_rd_data_way1_out_241 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6192 = _T_6191 | _T_5937; // @[Mux.scala 27:72]
  wire [21:0] _T_5938 = _T_4644 ? btb_bank0_rd_data_way1_out_242 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6193 = _T_6192 | _T_5938; // @[Mux.scala 27:72]
  wire [21:0] _T_5939 = _T_4646 ? btb_bank0_rd_data_way1_out_243 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6194 = _T_6193 | _T_5939; // @[Mux.scala 27:72]
  wire [21:0] _T_5940 = _T_4648 ? btb_bank0_rd_data_way1_out_244 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6195 = _T_6194 | _T_5940; // @[Mux.scala 27:72]
  wire [21:0] _T_5941 = _T_4650 ? btb_bank0_rd_data_way1_out_245 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6196 = _T_6195 | _T_5941; // @[Mux.scala 27:72]
  wire [21:0] _T_5942 = _T_4652 ? btb_bank0_rd_data_way1_out_246 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6197 = _T_6196 | _T_5942; // @[Mux.scala 27:72]
  wire [21:0] _T_5943 = _T_4654 ? btb_bank0_rd_data_way1_out_247 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6198 = _T_6197 | _T_5943; // @[Mux.scala 27:72]
  wire [21:0] _T_5944 = _T_4656 ? btb_bank0_rd_data_way1_out_248 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6199 = _T_6198 | _T_5944; // @[Mux.scala 27:72]
  wire [21:0] _T_5945 = _T_4658 ? btb_bank0_rd_data_way1_out_249 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6200 = _T_6199 | _T_5945; // @[Mux.scala 27:72]
  wire [21:0] _T_5946 = _T_4660 ? btb_bank0_rd_data_way1_out_250 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6201 = _T_6200 | _T_5946; // @[Mux.scala 27:72]
  wire [21:0] _T_5947 = _T_4662 ? btb_bank0_rd_data_way1_out_251 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6202 = _T_6201 | _T_5947; // @[Mux.scala 27:72]
  wire [21:0] _T_5948 = _T_4664 ? btb_bank0_rd_data_way1_out_252 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6203 = _T_6202 | _T_5948; // @[Mux.scala 27:72]
  wire [21:0] _T_5949 = _T_4666 ? btb_bank0_rd_data_way1_out_253 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6204 = _T_6203 | _T_5949; // @[Mux.scala 27:72]
  wire [21:0] _T_5950 = _T_4668 ? btb_bank0_rd_data_way1_out_254 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6205 = _T_6204 | _T_5950; // @[Mux.scala 27:72]
  wire [21:0] _T_5951 = _T_4670 ? btb_bank0_rd_data_way1_out_255 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] btb_bank0_rd_data_way1_p1_f = _T_6205 | _T_5951; // @[Mux.scala 27:72]
  wire  _T_73 = btb_bank0_rd_data_way1_p1_f[21:17] == fetch_rd_tag_p1_f; // @[ifu_bp_ctl.scala 138:106]
  wire  _T_74 = btb_bank0_rd_data_way1_p1_f[0] & _T_73; // @[ifu_bp_ctl.scala 138:61]
  wire  _T_77 = _T_74 & _T_67; // @[ifu_bp_ctl.scala 138:129]
  wire  _T_78 = _T_77 & io_ifc_fetch_req_f; // @[ifu_bp_ctl.scala 139:59]
  wire  tag_match_way1_p1_f = _T_78 & _T; // @[ifu_bp_ctl.scala 139:80]
  wire  _T_109 = btb_bank0_rd_data_way1_p1_f[3] ^ btb_bank0_rd_data_way1_p1_f[4]; // @[ifu_bp_ctl.scala 151:100]
  wire  _T_110 = tag_match_way1_p1_f & _T_109; // @[ifu_bp_ctl.scala 151:62]
  wire  _T_114 = ~_T_109; // @[ifu_bp_ctl.scala 152:64]
  wire  _T_115 = tag_match_way1_p1_f & _T_114; // @[ifu_bp_ctl.scala 152:62]
  wire [1:0] tag_match_way1_expanded_p1_f = {_T_110,_T_115}; // @[Cat.scala 29:58]
  wire [21:0] _T_135 = tag_match_way1_expanded_p1_f[0] ? btb_bank0_rd_data_way1_p1_f : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] btb_bank0e_rd_data_p1_f = _T_134 | _T_135; // @[Mux.scala 27:72]
  wire [21:0] _T_147 = io_ifc_fetch_addr_f[0] ? btb_bank0e_rd_data_p1_f : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] btb_vbank1_rd_data_f = _T_146 | _T_147; // @[Mux.scala 27:72]
  wire  _T_243 = btb_vbank1_rd_data_f[2] | btb_vbank1_rd_data_f[1]; // @[ifu_bp_ctl.scala 264:59]
  wire [21:0] _T_120 = tag_match_way0_expanded_f[0] ? btb_bank0_rd_data_way0_f : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_121 = tag_match_way1_expanded_f[0] ? btb_bank0_rd_data_way1_f : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] btb_bank0e_rd_data_f = _T_120 | _T_121; // @[Mux.scala 27:72]
  wire [21:0] _T_140 = _T_144 ? btb_bank0e_rd_data_f : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_141 = io_ifc_fetch_addr_f[0] ? btb_bank0o_rd_data_f : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] btb_vbank0_rd_data_f = _T_140 | _T_141; // @[Mux.scala 27:72]
  wire  _T_246 = btb_vbank0_rd_data_f[2] | btb_vbank0_rd_data_f[1]; // @[ifu_bp_ctl.scala 265:59]
  wire [1:0] bht_force_taken_f = {_T_243,_T_246}; // @[Cat.scala 29:58]
  wire [9:0] _T_570 = {btb_rd_addr_f,2'h0}; // @[Cat.scala 29:58]
  reg [7:0] fghr; // @[ifu_bp_ctl.scala 323:44]
  wire [7:0] bht_rd_addr_f = _T_570[9:2] ^ fghr; // @[lib.scala 56:35]
  wire  _T_21408 = bht_rd_addr_f == 8'h0; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_0; // @[Reg.scala 27:20]
  wire [1:0] _T_21920 = _T_21408 ? bht_bank_rd_data_out_1_0 : 2'h0; // @[Mux.scala 27:72]
  wire  _T_21410 = bht_rd_addr_f == 8'h1; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_1; // @[Reg.scala 27:20]
  wire [1:0] _T_21921 = _T_21410 ? bht_bank_rd_data_out_1_1 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22176 = _T_21920 | _T_21921; // @[Mux.scala 27:72]
  wire  _T_21412 = bht_rd_addr_f == 8'h2; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_2; // @[Reg.scala 27:20]
  wire [1:0] _T_21922 = _T_21412 ? bht_bank_rd_data_out_1_2 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22177 = _T_22176 | _T_21922; // @[Mux.scala 27:72]
  wire  _T_21414 = bht_rd_addr_f == 8'h3; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_3; // @[Reg.scala 27:20]
  wire [1:0] _T_21923 = _T_21414 ? bht_bank_rd_data_out_1_3 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22178 = _T_22177 | _T_21923; // @[Mux.scala 27:72]
  wire  _T_21416 = bht_rd_addr_f == 8'h4; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_4; // @[Reg.scala 27:20]
  wire [1:0] _T_21924 = _T_21416 ? bht_bank_rd_data_out_1_4 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22179 = _T_22178 | _T_21924; // @[Mux.scala 27:72]
  wire  _T_21418 = bht_rd_addr_f == 8'h5; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_5; // @[Reg.scala 27:20]
  wire [1:0] _T_21925 = _T_21418 ? bht_bank_rd_data_out_1_5 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22180 = _T_22179 | _T_21925; // @[Mux.scala 27:72]
  wire  _T_21420 = bht_rd_addr_f == 8'h6; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_6; // @[Reg.scala 27:20]
  wire [1:0] _T_21926 = _T_21420 ? bht_bank_rd_data_out_1_6 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22181 = _T_22180 | _T_21926; // @[Mux.scala 27:72]
  wire  _T_21422 = bht_rd_addr_f == 8'h7; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_7; // @[Reg.scala 27:20]
  wire [1:0] _T_21927 = _T_21422 ? bht_bank_rd_data_out_1_7 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22182 = _T_22181 | _T_21927; // @[Mux.scala 27:72]
  wire  _T_21424 = bht_rd_addr_f == 8'h8; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_8; // @[Reg.scala 27:20]
  wire [1:0] _T_21928 = _T_21424 ? bht_bank_rd_data_out_1_8 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22183 = _T_22182 | _T_21928; // @[Mux.scala 27:72]
  wire  _T_21426 = bht_rd_addr_f == 8'h9; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_9; // @[Reg.scala 27:20]
  wire [1:0] _T_21929 = _T_21426 ? bht_bank_rd_data_out_1_9 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22184 = _T_22183 | _T_21929; // @[Mux.scala 27:72]
  wire  _T_21428 = bht_rd_addr_f == 8'ha; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_10; // @[Reg.scala 27:20]
  wire [1:0] _T_21930 = _T_21428 ? bht_bank_rd_data_out_1_10 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22185 = _T_22184 | _T_21930; // @[Mux.scala 27:72]
  wire  _T_21430 = bht_rd_addr_f == 8'hb; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_11; // @[Reg.scala 27:20]
  wire [1:0] _T_21931 = _T_21430 ? bht_bank_rd_data_out_1_11 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22186 = _T_22185 | _T_21931; // @[Mux.scala 27:72]
  wire  _T_21432 = bht_rd_addr_f == 8'hc; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_12; // @[Reg.scala 27:20]
  wire [1:0] _T_21932 = _T_21432 ? bht_bank_rd_data_out_1_12 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22187 = _T_22186 | _T_21932; // @[Mux.scala 27:72]
  wire  _T_21434 = bht_rd_addr_f == 8'hd; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_13; // @[Reg.scala 27:20]
  wire [1:0] _T_21933 = _T_21434 ? bht_bank_rd_data_out_1_13 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22188 = _T_22187 | _T_21933; // @[Mux.scala 27:72]
  wire  _T_21436 = bht_rd_addr_f == 8'he; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_14; // @[Reg.scala 27:20]
  wire [1:0] _T_21934 = _T_21436 ? bht_bank_rd_data_out_1_14 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22189 = _T_22188 | _T_21934; // @[Mux.scala 27:72]
  wire  _T_21438 = bht_rd_addr_f == 8'hf; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_15; // @[Reg.scala 27:20]
  wire [1:0] _T_21935 = _T_21438 ? bht_bank_rd_data_out_1_15 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22190 = _T_22189 | _T_21935; // @[Mux.scala 27:72]
  wire  _T_21440 = bht_rd_addr_f == 8'h10; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_16; // @[Reg.scala 27:20]
  wire [1:0] _T_21936 = _T_21440 ? bht_bank_rd_data_out_1_16 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22191 = _T_22190 | _T_21936; // @[Mux.scala 27:72]
  wire  _T_21442 = bht_rd_addr_f == 8'h11; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_17; // @[Reg.scala 27:20]
  wire [1:0] _T_21937 = _T_21442 ? bht_bank_rd_data_out_1_17 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22192 = _T_22191 | _T_21937; // @[Mux.scala 27:72]
  wire  _T_21444 = bht_rd_addr_f == 8'h12; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_18; // @[Reg.scala 27:20]
  wire [1:0] _T_21938 = _T_21444 ? bht_bank_rd_data_out_1_18 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22193 = _T_22192 | _T_21938; // @[Mux.scala 27:72]
  wire  _T_21446 = bht_rd_addr_f == 8'h13; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_19; // @[Reg.scala 27:20]
  wire [1:0] _T_21939 = _T_21446 ? bht_bank_rd_data_out_1_19 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22194 = _T_22193 | _T_21939; // @[Mux.scala 27:72]
  wire  _T_21448 = bht_rd_addr_f == 8'h14; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_20; // @[Reg.scala 27:20]
  wire [1:0] _T_21940 = _T_21448 ? bht_bank_rd_data_out_1_20 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22195 = _T_22194 | _T_21940; // @[Mux.scala 27:72]
  wire  _T_21450 = bht_rd_addr_f == 8'h15; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_21; // @[Reg.scala 27:20]
  wire [1:0] _T_21941 = _T_21450 ? bht_bank_rd_data_out_1_21 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22196 = _T_22195 | _T_21941; // @[Mux.scala 27:72]
  wire  _T_21452 = bht_rd_addr_f == 8'h16; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_22; // @[Reg.scala 27:20]
  wire [1:0] _T_21942 = _T_21452 ? bht_bank_rd_data_out_1_22 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22197 = _T_22196 | _T_21942; // @[Mux.scala 27:72]
  wire  _T_21454 = bht_rd_addr_f == 8'h17; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_23; // @[Reg.scala 27:20]
  wire [1:0] _T_21943 = _T_21454 ? bht_bank_rd_data_out_1_23 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22198 = _T_22197 | _T_21943; // @[Mux.scala 27:72]
  wire  _T_21456 = bht_rd_addr_f == 8'h18; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_24; // @[Reg.scala 27:20]
  wire [1:0] _T_21944 = _T_21456 ? bht_bank_rd_data_out_1_24 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22199 = _T_22198 | _T_21944; // @[Mux.scala 27:72]
  wire  _T_21458 = bht_rd_addr_f == 8'h19; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_25; // @[Reg.scala 27:20]
  wire [1:0] _T_21945 = _T_21458 ? bht_bank_rd_data_out_1_25 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22200 = _T_22199 | _T_21945; // @[Mux.scala 27:72]
  wire  _T_21460 = bht_rd_addr_f == 8'h1a; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_26; // @[Reg.scala 27:20]
  wire [1:0] _T_21946 = _T_21460 ? bht_bank_rd_data_out_1_26 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22201 = _T_22200 | _T_21946; // @[Mux.scala 27:72]
  wire  _T_21462 = bht_rd_addr_f == 8'h1b; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_27; // @[Reg.scala 27:20]
  wire [1:0] _T_21947 = _T_21462 ? bht_bank_rd_data_out_1_27 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22202 = _T_22201 | _T_21947; // @[Mux.scala 27:72]
  wire  _T_21464 = bht_rd_addr_f == 8'h1c; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_28; // @[Reg.scala 27:20]
  wire [1:0] _T_21948 = _T_21464 ? bht_bank_rd_data_out_1_28 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22203 = _T_22202 | _T_21948; // @[Mux.scala 27:72]
  wire  _T_21466 = bht_rd_addr_f == 8'h1d; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_29; // @[Reg.scala 27:20]
  wire [1:0] _T_21949 = _T_21466 ? bht_bank_rd_data_out_1_29 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22204 = _T_22203 | _T_21949; // @[Mux.scala 27:72]
  wire  _T_21468 = bht_rd_addr_f == 8'h1e; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_30; // @[Reg.scala 27:20]
  wire [1:0] _T_21950 = _T_21468 ? bht_bank_rd_data_out_1_30 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22205 = _T_22204 | _T_21950; // @[Mux.scala 27:72]
  wire  _T_21470 = bht_rd_addr_f == 8'h1f; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_31; // @[Reg.scala 27:20]
  wire [1:0] _T_21951 = _T_21470 ? bht_bank_rd_data_out_1_31 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22206 = _T_22205 | _T_21951; // @[Mux.scala 27:72]
  wire  _T_21472 = bht_rd_addr_f == 8'h20; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_32; // @[Reg.scala 27:20]
  wire [1:0] _T_21952 = _T_21472 ? bht_bank_rd_data_out_1_32 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22207 = _T_22206 | _T_21952; // @[Mux.scala 27:72]
  wire  _T_21474 = bht_rd_addr_f == 8'h21; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_33; // @[Reg.scala 27:20]
  wire [1:0] _T_21953 = _T_21474 ? bht_bank_rd_data_out_1_33 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22208 = _T_22207 | _T_21953; // @[Mux.scala 27:72]
  wire  _T_21476 = bht_rd_addr_f == 8'h22; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_34; // @[Reg.scala 27:20]
  wire [1:0] _T_21954 = _T_21476 ? bht_bank_rd_data_out_1_34 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22209 = _T_22208 | _T_21954; // @[Mux.scala 27:72]
  wire  _T_21478 = bht_rd_addr_f == 8'h23; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_35; // @[Reg.scala 27:20]
  wire [1:0] _T_21955 = _T_21478 ? bht_bank_rd_data_out_1_35 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22210 = _T_22209 | _T_21955; // @[Mux.scala 27:72]
  wire  _T_21480 = bht_rd_addr_f == 8'h24; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_36; // @[Reg.scala 27:20]
  wire [1:0] _T_21956 = _T_21480 ? bht_bank_rd_data_out_1_36 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22211 = _T_22210 | _T_21956; // @[Mux.scala 27:72]
  wire  _T_21482 = bht_rd_addr_f == 8'h25; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_37; // @[Reg.scala 27:20]
  wire [1:0] _T_21957 = _T_21482 ? bht_bank_rd_data_out_1_37 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22212 = _T_22211 | _T_21957; // @[Mux.scala 27:72]
  wire  _T_21484 = bht_rd_addr_f == 8'h26; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_38; // @[Reg.scala 27:20]
  wire [1:0] _T_21958 = _T_21484 ? bht_bank_rd_data_out_1_38 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22213 = _T_22212 | _T_21958; // @[Mux.scala 27:72]
  wire  _T_21486 = bht_rd_addr_f == 8'h27; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_39; // @[Reg.scala 27:20]
  wire [1:0] _T_21959 = _T_21486 ? bht_bank_rd_data_out_1_39 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22214 = _T_22213 | _T_21959; // @[Mux.scala 27:72]
  wire  _T_21488 = bht_rd_addr_f == 8'h28; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_40; // @[Reg.scala 27:20]
  wire [1:0] _T_21960 = _T_21488 ? bht_bank_rd_data_out_1_40 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22215 = _T_22214 | _T_21960; // @[Mux.scala 27:72]
  wire  _T_21490 = bht_rd_addr_f == 8'h29; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_41; // @[Reg.scala 27:20]
  wire [1:0] _T_21961 = _T_21490 ? bht_bank_rd_data_out_1_41 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22216 = _T_22215 | _T_21961; // @[Mux.scala 27:72]
  wire  _T_21492 = bht_rd_addr_f == 8'h2a; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_42; // @[Reg.scala 27:20]
  wire [1:0] _T_21962 = _T_21492 ? bht_bank_rd_data_out_1_42 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22217 = _T_22216 | _T_21962; // @[Mux.scala 27:72]
  wire  _T_21494 = bht_rd_addr_f == 8'h2b; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_43; // @[Reg.scala 27:20]
  wire [1:0] _T_21963 = _T_21494 ? bht_bank_rd_data_out_1_43 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22218 = _T_22217 | _T_21963; // @[Mux.scala 27:72]
  wire  _T_21496 = bht_rd_addr_f == 8'h2c; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_44; // @[Reg.scala 27:20]
  wire [1:0] _T_21964 = _T_21496 ? bht_bank_rd_data_out_1_44 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22219 = _T_22218 | _T_21964; // @[Mux.scala 27:72]
  wire  _T_21498 = bht_rd_addr_f == 8'h2d; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_45; // @[Reg.scala 27:20]
  wire [1:0] _T_21965 = _T_21498 ? bht_bank_rd_data_out_1_45 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22220 = _T_22219 | _T_21965; // @[Mux.scala 27:72]
  wire  _T_21500 = bht_rd_addr_f == 8'h2e; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_46; // @[Reg.scala 27:20]
  wire [1:0] _T_21966 = _T_21500 ? bht_bank_rd_data_out_1_46 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22221 = _T_22220 | _T_21966; // @[Mux.scala 27:72]
  wire  _T_21502 = bht_rd_addr_f == 8'h2f; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_47; // @[Reg.scala 27:20]
  wire [1:0] _T_21967 = _T_21502 ? bht_bank_rd_data_out_1_47 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22222 = _T_22221 | _T_21967; // @[Mux.scala 27:72]
  wire  _T_21504 = bht_rd_addr_f == 8'h30; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_48; // @[Reg.scala 27:20]
  wire [1:0] _T_21968 = _T_21504 ? bht_bank_rd_data_out_1_48 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22223 = _T_22222 | _T_21968; // @[Mux.scala 27:72]
  wire  _T_21506 = bht_rd_addr_f == 8'h31; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_49; // @[Reg.scala 27:20]
  wire [1:0] _T_21969 = _T_21506 ? bht_bank_rd_data_out_1_49 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22224 = _T_22223 | _T_21969; // @[Mux.scala 27:72]
  wire  _T_21508 = bht_rd_addr_f == 8'h32; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_50; // @[Reg.scala 27:20]
  wire [1:0] _T_21970 = _T_21508 ? bht_bank_rd_data_out_1_50 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22225 = _T_22224 | _T_21970; // @[Mux.scala 27:72]
  wire  _T_21510 = bht_rd_addr_f == 8'h33; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_51; // @[Reg.scala 27:20]
  wire [1:0] _T_21971 = _T_21510 ? bht_bank_rd_data_out_1_51 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22226 = _T_22225 | _T_21971; // @[Mux.scala 27:72]
  wire  _T_21512 = bht_rd_addr_f == 8'h34; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_52; // @[Reg.scala 27:20]
  wire [1:0] _T_21972 = _T_21512 ? bht_bank_rd_data_out_1_52 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22227 = _T_22226 | _T_21972; // @[Mux.scala 27:72]
  wire  _T_21514 = bht_rd_addr_f == 8'h35; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_53; // @[Reg.scala 27:20]
  wire [1:0] _T_21973 = _T_21514 ? bht_bank_rd_data_out_1_53 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22228 = _T_22227 | _T_21973; // @[Mux.scala 27:72]
  wire  _T_21516 = bht_rd_addr_f == 8'h36; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_54; // @[Reg.scala 27:20]
  wire [1:0] _T_21974 = _T_21516 ? bht_bank_rd_data_out_1_54 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22229 = _T_22228 | _T_21974; // @[Mux.scala 27:72]
  wire  _T_21518 = bht_rd_addr_f == 8'h37; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_55; // @[Reg.scala 27:20]
  wire [1:0] _T_21975 = _T_21518 ? bht_bank_rd_data_out_1_55 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22230 = _T_22229 | _T_21975; // @[Mux.scala 27:72]
  wire  _T_21520 = bht_rd_addr_f == 8'h38; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_56; // @[Reg.scala 27:20]
  wire [1:0] _T_21976 = _T_21520 ? bht_bank_rd_data_out_1_56 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22231 = _T_22230 | _T_21976; // @[Mux.scala 27:72]
  wire  _T_21522 = bht_rd_addr_f == 8'h39; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_57; // @[Reg.scala 27:20]
  wire [1:0] _T_21977 = _T_21522 ? bht_bank_rd_data_out_1_57 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22232 = _T_22231 | _T_21977; // @[Mux.scala 27:72]
  wire  _T_21524 = bht_rd_addr_f == 8'h3a; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_58; // @[Reg.scala 27:20]
  wire [1:0] _T_21978 = _T_21524 ? bht_bank_rd_data_out_1_58 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22233 = _T_22232 | _T_21978; // @[Mux.scala 27:72]
  wire  _T_21526 = bht_rd_addr_f == 8'h3b; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_59; // @[Reg.scala 27:20]
  wire [1:0] _T_21979 = _T_21526 ? bht_bank_rd_data_out_1_59 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22234 = _T_22233 | _T_21979; // @[Mux.scala 27:72]
  wire  _T_21528 = bht_rd_addr_f == 8'h3c; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_60; // @[Reg.scala 27:20]
  wire [1:0] _T_21980 = _T_21528 ? bht_bank_rd_data_out_1_60 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22235 = _T_22234 | _T_21980; // @[Mux.scala 27:72]
  wire  _T_21530 = bht_rd_addr_f == 8'h3d; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_61; // @[Reg.scala 27:20]
  wire [1:0] _T_21981 = _T_21530 ? bht_bank_rd_data_out_1_61 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22236 = _T_22235 | _T_21981; // @[Mux.scala 27:72]
  wire  _T_21532 = bht_rd_addr_f == 8'h3e; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_62; // @[Reg.scala 27:20]
  wire [1:0] _T_21982 = _T_21532 ? bht_bank_rd_data_out_1_62 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22237 = _T_22236 | _T_21982; // @[Mux.scala 27:72]
  wire  _T_21534 = bht_rd_addr_f == 8'h3f; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_63; // @[Reg.scala 27:20]
  wire [1:0] _T_21983 = _T_21534 ? bht_bank_rd_data_out_1_63 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22238 = _T_22237 | _T_21983; // @[Mux.scala 27:72]
  wire  _T_21536 = bht_rd_addr_f == 8'h40; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_64; // @[Reg.scala 27:20]
  wire [1:0] _T_21984 = _T_21536 ? bht_bank_rd_data_out_1_64 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22239 = _T_22238 | _T_21984; // @[Mux.scala 27:72]
  wire  _T_21538 = bht_rd_addr_f == 8'h41; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_65; // @[Reg.scala 27:20]
  wire [1:0] _T_21985 = _T_21538 ? bht_bank_rd_data_out_1_65 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22240 = _T_22239 | _T_21985; // @[Mux.scala 27:72]
  wire  _T_21540 = bht_rd_addr_f == 8'h42; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_66; // @[Reg.scala 27:20]
  wire [1:0] _T_21986 = _T_21540 ? bht_bank_rd_data_out_1_66 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22241 = _T_22240 | _T_21986; // @[Mux.scala 27:72]
  wire  _T_21542 = bht_rd_addr_f == 8'h43; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_67; // @[Reg.scala 27:20]
  wire [1:0] _T_21987 = _T_21542 ? bht_bank_rd_data_out_1_67 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22242 = _T_22241 | _T_21987; // @[Mux.scala 27:72]
  wire  _T_21544 = bht_rd_addr_f == 8'h44; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_68; // @[Reg.scala 27:20]
  wire [1:0] _T_21988 = _T_21544 ? bht_bank_rd_data_out_1_68 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22243 = _T_22242 | _T_21988; // @[Mux.scala 27:72]
  wire  _T_21546 = bht_rd_addr_f == 8'h45; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_69; // @[Reg.scala 27:20]
  wire [1:0] _T_21989 = _T_21546 ? bht_bank_rd_data_out_1_69 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22244 = _T_22243 | _T_21989; // @[Mux.scala 27:72]
  wire  _T_21548 = bht_rd_addr_f == 8'h46; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_70; // @[Reg.scala 27:20]
  wire [1:0] _T_21990 = _T_21548 ? bht_bank_rd_data_out_1_70 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22245 = _T_22244 | _T_21990; // @[Mux.scala 27:72]
  wire  _T_21550 = bht_rd_addr_f == 8'h47; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_71; // @[Reg.scala 27:20]
  wire [1:0] _T_21991 = _T_21550 ? bht_bank_rd_data_out_1_71 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22246 = _T_22245 | _T_21991; // @[Mux.scala 27:72]
  wire  _T_21552 = bht_rd_addr_f == 8'h48; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_72; // @[Reg.scala 27:20]
  wire [1:0] _T_21992 = _T_21552 ? bht_bank_rd_data_out_1_72 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22247 = _T_22246 | _T_21992; // @[Mux.scala 27:72]
  wire  _T_21554 = bht_rd_addr_f == 8'h49; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_73; // @[Reg.scala 27:20]
  wire [1:0] _T_21993 = _T_21554 ? bht_bank_rd_data_out_1_73 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22248 = _T_22247 | _T_21993; // @[Mux.scala 27:72]
  wire  _T_21556 = bht_rd_addr_f == 8'h4a; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_74; // @[Reg.scala 27:20]
  wire [1:0] _T_21994 = _T_21556 ? bht_bank_rd_data_out_1_74 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22249 = _T_22248 | _T_21994; // @[Mux.scala 27:72]
  wire  _T_21558 = bht_rd_addr_f == 8'h4b; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_75; // @[Reg.scala 27:20]
  wire [1:0] _T_21995 = _T_21558 ? bht_bank_rd_data_out_1_75 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22250 = _T_22249 | _T_21995; // @[Mux.scala 27:72]
  wire  _T_21560 = bht_rd_addr_f == 8'h4c; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_76; // @[Reg.scala 27:20]
  wire [1:0] _T_21996 = _T_21560 ? bht_bank_rd_data_out_1_76 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22251 = _T_22250 | _T_21996; // @[Mux.scala 27:72]
  wire  _T_21562 = bht_rd_addr_f == 8'h4d; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_77; // @[Reg.scala 27:20]
  wire [1:0] _T_21997 = _T_21562 ? bht_bank_rd_data_out_1_77 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22252 = _T_22251 | _T_21997; // @[Mux.scala 27:72]
  wire  _T_21564 = bht_rd_addr_f == 8'h4e; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_78; // @[Reg.scala 27:20]
  wire [1:0] _T_21998 = _T_21564 ? bht_bank_rd_data_out_1_78 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22253 = _T_22252 | _T_21998; // @[Mux.scala 27:72]
  wire  _T_21566 = bht_rd_addr_f == 8'h4f; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_79; // @[Reg.scala 27:20]
  wire [1:0] _T_21999 = _T_21566 ? bht_bank_rd_data_out_1_79 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22254 = _T_22253 | _T_21999; // @[Mux.scala 27:72]
  wire  _T_21568 = bht_rd_addr_f == 8'h50; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_80; // @[Reg.scala 27:20]
  wire [1:0] _T_22000 = _T_21568 ? bht_bank_rd_data_out_1_80 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22255 = _T_22254 | _T_22000; // @[Mux.scala 27:72]
  wire  _T_21570 = bht_rd_addr_f == 8'h51; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_81; // @[Reg.scala 27:20]
  wire [1:0] _T_22001 = _T_21570 ? bht_bank_rd_data_out_1_81 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22256 = _T_22255 | _T_22001; // @[Mux.scala 27:72]
  wire  _T_21572 = bht_rd_addr_f == 8'h52; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_82; // @[Reg.scala 27:20]
  wire [1:0] _T_22002 = _T_21572 ? bht_bank_rd_data_out_1_82 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22257 = _T_22256 | _T_22002; // @[Mux.scala 27:72]
  wire  _T_21574 = bht_rd_addr_f == 8'h53; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_83; // @[Reg.scala 27:20]
  wire [1:0] _T_22003 = _T_21574 ? bht_bank_rd_data_out_1_83 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22258 = _T_22257 | _T_22003; // @[Mux.scala 27:72]
  wire  _T_21576 = bht_rd_addr_f == 8'h54; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_84; // @[Reg.scala 27:20]
  wire [1:0] _T_22004 = _T_21576 ? bht_bank_rd_data_out_1_84 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22259 = _T_22258 | _T_22004; // @[Mux.scala 27:72]
  wire  _T_21578 = bht_rd_addr_f == 8'h55; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_85; // @[Reg.scala 27:20]
  wire [1:0] _T_22005 = _T_21578 ? bht_bank_rd_data_out_1_85 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22260 = _T_22259 | _T_22005; // @[Mux.scala 27:72]
  wire  _T_21580 = bht_rd_addr_f == 8'h56; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_86; // @[Reg.scala 27:20]
  wire [1:0] _T_22006 = _T_21580 ? bht_bank_rd_data_out_1_86 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22261 = _T_22260 | _T_22006; // @[Mux.scala 27:72]
  wire  _T_21582 = bht_rd_addr_f == 8'h57; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_87; // @[Reg.scala 27:20]
  wire [1:0] _T_22007 = _T_21582 ? bht_bank_rd_data_out_1_87 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22262 = _T_22261 | _T_22007; // @[Mux.scala 27:72]
  wire  _T_21584 = bht_rd_addr_f == 8'h58; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_88; // @[Reg.scala 27:20]
  wire [1:0] _T_22008 = _T_21584 ? bht_bank_rd_data_out_1_88 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22263 = _T_22262 | _T_22008; // @[Mux.scala 27:72]
  wire  _T_21586 = bht_rd_addr_f == 8'h59; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_89; // @[Reg.scala 27:20]
  wire [1:0] _T_22009 = _T_21586 ? bht_bank_rd_data_out_1_89 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22264 = _T_22263 | _T_22009; // @[Mux.scala 27:72]
  wire  _T_21588 = bht_rd_addr_f == 8'h5a; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_90; // @[Reg.scala 27:20]
  wire [1:0] _T_22010 = _T_21588 ? bht_bank_rd_data_out_1_90 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22265 = _T_22264 | _T_22010; // @[Mux.scala 27:72]
  wire  _T_21590 = bht_rd_addr_f == 8'h5b; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_91; // @[Reg.scala 27:20]
  wire [1:0] _T_22011 = _T_21590 ? bht_bank_rd_data_out_1_91 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22266 = _T_22265 | _T_22011; // @[Mux.scala 27:72]
  wire  _T_21592 = bht_rd_addr_f == 8'h5c; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_92; // @[Reg.scala 27:20]
  wire [1:0] _T_22012 = _T_21592 ? bht_bank_rd_data_out_1_92 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22267 = _T_22266 | _T_22012; // @[Mux.scala 27:72]
  wire  _T_21594 = bht_rd_addr_f == 8'h5d; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_93; // @[Reg.scala 27:20]
  wire [1:0] _T_22013 = _T_21594 ? bht_bank_rd_data_out_1_93 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22268 = _T_22267 | _T_22013; // @[Mux.scala 27:72]
  wire  _T_21596 = bht_rd_addr_f == 8'h5e; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_94; // @[Reg.scala 27:20]
  wire [1:0] _T_22014 = _T_21596 ? bht_bank_rd_data_out_1_94 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22269 = _T_22268 | _T_22014; // @[Mux.scala 27:72]
  wire  _T_21598 = bht_rd_addr_f == 8'h5f; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_95; // @[Reg.scala 27:20]
  wire [1:0] _T_22015 = _T_21598 ? bht_bank_rd_data_out_1_95 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22270 = _T_22269 | _T_22015; // @[Mux.scala 27:72]
  wire  _T_21600 = bht_rd_addr_f == 8'h60; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_96; // @[Reg.scala 27:20]
  wire [1:0] _T_22016 = _T_21600 ? bht_bank_rd_data_out_1_96 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22271 = _T_22270 | _T_22016; // @[Mux.scala 27:72]
  wire  _T_21602 = bht_rd_addr_f == 8'h61; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_97; // @[Reg.scala 27:20]
  wire [1:0] _T_22017 = _T_21602 ? bht_bank_rd_data_out_1_97 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22272 = _T_22271 | _T_22017; // @[Mux.scala 27:72]
  wire  _T_21604 = bht_rd_addr_f == 8'h62; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_98; // @[Reg.scala 27:20]
  wire [1:0] _T_22018 = _T_21604 ? bht_bank_rd_data_out_1_98 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22273 = _T_22272 | _T_22018; // @[Mux.scala 27:72]
  wire  _T_21606 = bht_rd_addr_f == 8'h63; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_99; // @[Reg.scala 27:20]
  wire [1:0] _T_22019 = _T_21606 ? bht_bank_rd_data_out_1_99 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22274 = _T_22273 | _T_22019; // @[Mux.scala 27:72]
  wire  _T_21608 = bht_rd_addr_f == 8'h64; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_100; // @[Reg.scala 27:20]
  wire [1:0] _T_22020 = _T_21608 ? bht_bank_rd_data_out_1_100 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22275 = _T_22274 | _T_22020; // @[Mux.scala 27:72]
  wire  _T_21610 = bht_rd_addr_f == 8'h65; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_101; // @[Reg.scala 27:20]
  wire [1:0] _T_22021 = _T_21610 ? bht_bank_rd_data_out_1_101 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22276 = _T_22275 | _T_22021; // @[Mux.scala 27:72]
  wire  _T_21612 = bht_rd_addr_f == 8'h66; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_102; // @[Reg.scala 27:20]
  wire [1:0] _T_22022 = _T_21612 ? bht_bank_rd_data_out_1_102 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22277 = _T_22276 | _T_22022; // @[Mux.scala 27:72]
  wire  _T_21614 = bht_rd_addr_f == 8'h67; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_103; // @[Reg.scala 27:20]
  wire [1:0] _T_22023 = _T_21614 ? bht_bank_rd_data_out_1_103 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22278 = _T_22277 | _T_22023; // @[Mux.scala 27:72]
  wire  _T_21616 = bht_rd_addr_f == 8'h68; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_104; // @[Reg.scala 27:20]
  wire [1:0] _T_22024 = _T_21616 ? bht_bank_rd_data_out_1_104 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22279 = _T_22278 | _T_22024; // @[Mux.scala 27:72]
  wire  _T_21618 = bht_rd_addr_f == 8'h69; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_105; // @[Reg.scala 27:20]
  wire [1:0] _T_22025 = _T_21618 ? bht_bank_rd_data_out_1_105 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22280 = _T_22279 | _T_22025; // @[Mux.scala 27:72]
  wire  _T_21620 = bht_rd_addr_f == 8'h6a; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_106; // @[Reg.scala 27:20]
  wire [1:0] _T_22026 = _T_21620 ? bht_bank_rd_data_out_1_106 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22281 = _T_22280 | _T_22026; // @[Mux.scala 27:72]
  wire  _T_21622 = bht_rd_addr_f == 8'h6b; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_107; // @[Reg.scala 27:20]
  wire [1:0] _T_22027 = _T_21622 ? bht_bank_rd_data_out_1_107 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22282 = _T_22281 | _T_22027; // @[Mux.scala 27:72]
  wire  _T_21624 = bht_rd_addr_f == 8'h6c; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_108; // @[Reg.scala 27:20]
  wire [1:0] _T_22028 = _T_21624 ? bht_bank_rd_data_out_1_108 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22283 = _T_22282 | _T_22028; // @[Mux.scala 27:72]
  wire  _T_21626 = bht_rd_addr_f == 8'h6d; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_109; // @[Reg.scala 27:20]
  wire [1:0] _T_22029 = _T_21626 ? bht_bank_rd_data_out_1_109 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22284 = _T_22283 | _T_22029; // @[Mux.scala 27:72]
  wire  _T_21628 = bht_rd_addr_f == 8'h6e; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_110; // @[Reg.scala 27:20]
  wire [1:0] _T_22030 = _T_21628 ? bht_bank_rd_data_out_1_110 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22285 = _T_22284 | _T_22030; // @[Mux.scala 27:72]
  wire  _T_21630 = bht_rd_addr_f == 8'h6f; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_111; // @[Reg.scala 27:20]
  wire [1:0] _T_22031 = _T_21630 ? bht_bank_rd_data_out_1_111 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22286 = _T_22285 | _T_22031; // @[Mux.scala 27:72]
  wire  _T_21632 = bht_rd_addr_f == 8'h70; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_112; // @[Reg.scala 27:20]
  wire [1:0] _T_22032 = _T_21632 ? bht_bank_rd_data_out_1_112 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22287 = _T_22286 | _T_22032; // @[Mux.scala 27:72]
  wire  _T_21634 = bht_rd_addr_f == 8'h71; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_113; // @[Reg.scala 27:20]
  wire [1:0] _T_22033 = _T_21634 ? bht_bank_rd_data_out_1_113 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22288 = _T_22287 | _T_22033; // @[Mux.scala 27:72]
  wire  _T_21636 = bht_rd_addr_f == 8'h72; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_114; // @[Reg.scala 27:20]
  wire [1:0] _T_22034 = _T_21636 ? bht_bank_rd_data_out_1_114 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22289 = _T_22288 | _T_22034; // @[Mux.scala 27:72]
  wire  _T_21638 = bht_rd_addr_f == 8'h73; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_115; // @[Reg.scala 27:20]
  wire [1:0] _T_22035 = _T_21638 ? bht_bank_rd_data_out_1_115 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22290 = _T_22289 | _T_22035; // @[Mux.scala 27:72]
  wire  _T_21640 = bht_rd_addr_f == 8'h74; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_116; // @[Reg.scala 27:20]
  wire [1:0] _T_22036 = _T_21640 ? bht_bank_rd_data_out_1_116 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22291 = _T_22290 | _T_22036; // @[Mux.scala 27:72]
  wire  _T_21642 = bht_rd_addr_f == 8'h75; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_117; // @[Reg.scala 27:20]
  wire [1:0] _T_22037 = _T_21642 ? bht_bank_rd_data_out_1_117 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22292 = _T_22291 | _T_22037; // @[Mux.scala 27:72]
  wire  _T_21644 = bht_rd_addr_f == 8'h76; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_118; // @[Reg.scala 27:20]
  wire [1:0] _T_22038 = _T_21644 ? bht_bank_rd_data_out_1_118 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22293 = _T_22292 | _T_22038; // @[Mux.scala 27:72]
  wire  _T_21646 = bht_rd_addr_f == 8'h77; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_119; // @[Reg.scala 27:20]
  wire [1:0] _T_22039 = _T_21646 ? bht_bank_rd_data_out_1_119 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22294 = _T_22293 | _T_22039; // @[Mux.scala 27:72]
  wire  _T_21648 = bht_rd_addr_f == 8'h78; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_120; // @[Reg.scala 27:20]
  wire [1:0] _T_22040 = _T_21648 ? bht_bank_rd_data_out_1_120 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22295 = _T_22294 | _T_22040; // @[Mux.scala 27:72]
  wire  _T_21650 = bht_rd_addr_f == 8'h79; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_121; // @[Reg.scala 27:20]
  wire [1:0] _T_22041 = _T_21650 ? bht_bank_rd_data_out_1_121 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22296 = _T_22295 | _T_22041; // @[Mux.scala 27:72]
  wire  _T_21652 = bht_rd_addr_f == 8'h7a; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_122; // @[Reg.scala 27:20]
  wire [1:0] _T_22042 = _T_21652 ? bht_bank_rd_data_out_1_122 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22297 = _T_22296 | _T_22042; // @[Mux.scala 27:72]
  wire  _T_21654 = bht_rd_addr_f == 8'h7b; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_123; // @[Reg.scala 27:20]
  wire [1:0] _T_22043 = _T_21654 ? bht_bank_rd_data_out_1_123 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22298 = _T_22297 | _T_22043; // @[Mux.scala 27:72]
  wire  _T_21656 = bht_rd_addr_f == 8'h7c; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_124; // @[Reg.scala 27:20]
  wire [1:0] _T_22044 = _T_21656 ? bht_bank_rd_data_out_1_124 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22299 = _T_22298 | _T_22044; // @[Mux.scala 27:72]
  wire  _T_21658 = bht_rd_addr_f == 8'h7d; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_125; // @[Reg.scala 27:20]
  wire [1:0] _T_22045 = _T_21658 ? bht_bank_rd_data_out_1_125 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22300 = _T_22299 | _T_22045; // @[Mux.scala 27:72]
  wire  _T_21660 = bht_rd_addr_f == 8'h7e; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_126; // @[Reg.scala 27:20]
  wire [1:0] _T_22046 = _T_21660 ? bht_bank_rd_data_out_1_126 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22301 = _T_22300 | _T_22046; // @[Mux.scala 27:72]
  wire  _T_21662 = bht_rd_addr_f == 8'h7f; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_127; // @[Reg.scala 27:20]
  wire [1:0] _T_22047 = _T_21662 ? bht_bank_rd_data_out_1_127 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22302 = _T_22301 | _T_22047; // @[Mux.scala 27:72]
  wire  _T_21664 = bht_rd_addr_f == 8'h80; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_128; // @[Reg.scala 27:20]
  wire [1:0] _T_22048 = _T_21664 ? bht_bank_rd_data_out_1_128 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22303 = _T_22302 | _T_22048; // @[Mux.scala 27:72]
  wire  _T_21666 = bht_rd_addr_f == 8'h81; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_129; // @[Reg.scala 27:20]
  wire [1:0] _T_22049 = _T_21666 ? bht_bank_rd_data_out_1_129 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22304 = _T_22303 | _T_22049; // @[Mux.scala 27:72]
  wire  _T_21668 = bht_rd_addr_f == 8'h82; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_130; // @[Reg.scala 27:20]
  wire [1:0] _T_22050 = _T_21668 ? bht_bank_rd_data_out_1_130 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22305 = _T_22304 | _T_22050; // @[Mux.scala 27:72]
  wire  _T_21670 = bht_rd_addr_f == 8'h83; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_131; // @[Reg.scala 27:20]
  wire [1:0] _T_22051 = _T_21670 ? bht_bank_rd_data_out_1_131 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22306 = _T_22305 | _T_22051; // @[Mux.scala 27:72]
  wire  _T_21672 = bht_rd_addr_f == 8'h84; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_132; // @[Reg.scala 27:20]
  wire [1:0] _T_22052 = _T_21672 ? bht_bank_rd_data_out_1_132 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22307 = _T_22306 | _T_22052; // @[Mux.scala 27:72]
  wire  _T_21674 = bht_rd_addr_f == 8'h85; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_133; // @[Reg.scala 27:20]
  wire [1:0] _T_22053 = _T_21674 ? bht_bank_rd_data_out_1_133 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22308 = _T_22307 | _T_22053; // @[Mux.scala 27:72]
  wire  _T_21676 = bht_rd_addr_f == 8'h86; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_134; // @[Reg.scala 27:20]
  wire [1:0] _T_22054 = _T_21676 ? bht_bank_rd_data_out_1_134 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22309 = _T_22308 | _T_22054; // @[Mux.scala 27:72]
  wire  _T_21678 = bht_rd_addr_f == 8'h87; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_135; // @[Reg.scala 27:20]
  wire [1:0] _T_22055 = _T_21678 ? bht_bank_rd_data_out_1_135 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22310 = _T_22309 | _T_22055; // @[Mux.scala 27:72]
  wire  _T_21680 = bht_rd_addr_f == 8'h88; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_136; // @[Reg.scala 27:20]
  wire [1:0] _T_22056 = _T_21680 ? bht_bank_rd_data_out_1_136 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22311 = _T_22310 | _T_22056; // @[Mux.scala 27:72]
  wire  _T_21682 = bht_rd_addr_f == 8'h89; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_137; // @[Reg.scala 27:20]
  wire [1:0] _T_22057 = _T_21682 ? bht_bank_rd_data_out_1_137 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22312 = _T_22311 | _T_22057; // @[Mux.scala 27:72]
  wire  _T_21684 = bht_rd_addr_f == 8'h8a; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_138; // @[Reg.scala 27:20]
  wire [1:0] _T_22058 = _T_21684 ? bht_bank_rd_data_out_1_138 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22313 = _T_22312 | _T_22058; // @[Mux.scala 27:72]
  wire  _T_21686 = bht_rd_addr_f == 8'h8b; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_139; // @[Reg.scala 27:20]
  wire [1:0] _T_22059 = _T_21686 ? bht_bank_rd_data_out_1_139 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22314 = _T_22313 | _T_22059; // @[Mux.scala 27:72]
  wire  _T_21688 = bht_rd_addr_f == 8'h8c; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_140; // @[Reg.scala 27:20]
  wire [1:0] _T_22060 = _T_21688 ? bht_bank_rd_data_out_1_140 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22315 = _T_22314 | _T_22060; // @[Mux.scala 27:72]
  wire  _T_21690 = bht_rd_addr_f == 8'h8d; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_141; // @[Reg.scala 27:20]
  wire [1:0] _T_22061 = _T_21690 ? bht_bank_rd_data_out_1_141 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22316 = _T_22315 | _T_22061; // @[Mux.scala 27:72]
  wire  _T_21692 = bht_rd_addr_f == 8'h8e; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_142; // @[Reg.scala 27:20]
  wire [1:0] _T_22062 = _T_21692 ? bht_bank_rd_data_out_1_142 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22317 = _T_22316 | _T_22062; // @[Mux.scala 27:72]
  wire  _T_21694 = bht_rd_addr_f == 8'h8f; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_143; // @[Reg.scala 27:20]
  wire [1:0] _T_22063 = _T_21694 ? bht_bank_rd_data_out_1_143 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22318 = _T_22317 | _T_22063; // @[Mux.scala 27:72]
  wire  _T_21696 = bht_rd_addr_f == 8'h90; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_144; // @[Reg.scala 27:20]
  wire [1:0] _T_22064 = _T_21696 ? bht_bank_rd_data_out_1_144 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22319 = _T_22318 | _T_22064; // @[Mux.scala 27:72]
  wire  _T_21698 = bht_rd_addr_f == 8'h91; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_145; // @[Reg.scala 27:20]
  wire [1:0] _T_22065 = _T_21698 ? bht_bank_rd_data_out_1_145 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22320 = _T_22319 | _T_22065; // @[Mux.scala 27:72]
  wire  _T_21700 = bht_rd_addr_f == 8'h92; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_146; // @[Reg.scala 27:20]
  wire [1:0] _T_22066 = _T_21700 ? bht_bank_rd_data_out_1_146 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22321 = _T_22320 | _T_22066; // @[Mux.scala 27:72]
  wire  _T_21702 = bht_rd_addr_f == 8'h93; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_147; // @[Reg.scala 27:20]
  wire [1:0] _T_22067 = _T_21702 ? bht_bank_rd_data_out_1_147 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22322 = _T_22321 | _T_22067; // @[Mux.scala 27:72]
  wire  _T_21704 = bht_rd_addr_f == 8'h94; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_148; // @[Reg.scala 27:20]
  wire [1:0] _T_22068 = _T_21704 ? bht_bank_rd_data_out_1_148 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22323 = _T_22322 | _T_22068; // @[Mux.scala 27:72]
  wire  _T_21706 = bht_rd_addr_f == 8'h95; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_149; // @[Reg.scala 27:20]
  wire [1:0] _T_22069 = _T_21706 ? bht_bank_rd_data_out_1_149 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22324 = _T_22323 | _T_22069; // @[Mux.scala 27:72]
  wire  _T_21708 = bht_rd_addr_f == 8'h96; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_150; // @[Reg.scala 27:20]
  wire [1:0] _T_22070 = _T_21708 ? bht_bank_rd_data_out_1_150 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22325 = _T_22324 | _T_22070; // @[Mux.scala 27:72]
  wire  _T_21710 = bht_rd_addr_f == 8'h97; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_151; // @[Reg.scala 27:20]
  wire [1:0] _T_22071 = _T_21710 ? bht_bank_rd_data_out_1_151 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22326 = _T_22325 | _T_22071; // @[Mux.scala 27:72]
  wire  _T_21712 = bht_rd_addr_f == 8'h98; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_152; // @[Reg.scala 27:20]
  wire [1:0] _T_22072 = _T_21712 ? bht_bank_rd_data_out_1_152 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22327 = _T_22326 | _T_22072; // @[Mux.scala 27:72]
  wire  _T_21714 = bht_rd_addr_f == 8'h99; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_153; // @[Reg.scala 27:20]
  wire [1:0] _T_22073 = _T_21714 ? bht_bank_rd_data_out_1_153 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22328 = _T_22327 | _T_22073; // @[Mux.scala 27:72]
  wire  _T_21716 = bht_rd_addr_f == 8'h9a; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_154; // @[Reg.scala 27:20]
  wire [1:0] _T_22074 = _T_21716 ? bht_bank_rd_data_out_1_154 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22329 = _T_22328 | _T_22074; // @[Mux.scala 27:72]
  wire  _T_21718 = bht_rd_addr_f == 8'h9b; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_155; // @[Reg.scala 27:20]
  wire [1:0] _T_22075 = _T_21718 ? bht_bank_rd_data_out_1_155 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22330 = _T_22329 | _T_22075; // @[Mux.scala 27:72]
  wire  _T_21720 = bht_rd_addr_f == 8'h9c; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_156; // @[Reg.scala 27:20]
  wire [1:0] _T_22076 = _T_21720 ? bht_bank_rd_data_out_1_156 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22331 = _T_22330 | _T_22076; // @[Mux.scala 27:72]
  wire  _T_21722 = bht_rd_addr_f == 8'h9d; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_157; // @[Reg.scala 27:20]
  wire [1:0] _T_22077 = _T_21722 ? bht_bank_rd_data_out_1_157 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22332 = _T_22331 | _T_22077; // @[Mux.scala 27:72]
  wire  _T_21724 = bht_rd_addr_f == 8'h9e; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_158; // @[Reg.scala 27:20]
  wire [1:0] _T_22078 = _T_21724 ? bht_bank_rd_data_out_1_158 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22333 = _T_22332 | _T_22078; // @[Mux.scala 27:72]
  wire  _T_21726 = bht_rd_addr_f == 8'h9f; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_159; // @[Reg.scala 27:20]
  wire [1:0] _T_22079 = _T_21726 ? bht_bank_rd_data_out_1_159 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22334 = _T_22333 | _T_22079; // @[Mux.scala 27:72]
  wire  _T_21728 = bht_rd_addr_f == 8'ha0; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_160; // @[Reg.scala 27:20]
  wire [1:0] _T_22080 = _T_21728 ? bht_bank_rd_data_out_1_160 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22335 = _T_22334 | _T_22080; // @[Mux.scala 27:72]
  wire  _T_21730 = bht_rd_addr_f == 8'ha1; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_161; // @[Reg.scala 27:20]
  wire [1:0] _T_22081 = _T_21730 ? bht_bank_rd_data_out_1_161 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22336 = _T_22335 | _T_22081; // @[Mux.scala 27:72]
  wire  _T_21732 = bht_rd_addr_f == 8'ha2; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_162; // @[Reg.scala 27:20]
  wire [1:0] _T_22082 = _T_21732 ? bht_bank_rd_data_out_1_162 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22337 = _T_22336 | _T_22082; // @[Mux.scala 27:72]
  wire  _T_21734 = bht_rd_addr_f == 8'ha3; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_163; // @[Reg.scala 27:20]
  wire [1:0] _T_22083 = _T_21734 ? bht_bank_rd_data_out_1_163 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22338 = _T_22337 | _T_22083; // @[Mux.scala 27:72]
  wire  _T_21736 = bht_rd_addr_f == 8'ha4; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_164; // @[Reg.scala 27:20]
  wire [1:0] _T_22084 = _T_21736 ? bht_bank_rd_data_out_1_164 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22339 = _T_22338 | _T_22084; // @[Mux.scala 27:72]
  wire  _T_21738 = bht_rd_addr_f == 8'ha5; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_165; // @[Reg.scala 27:20]
  wire [1:0] _T_22085 = _T_21738 ? bht_bank_rd_data_out_1_165 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22340 = _T_22339 | _T_22085; // @[Mux.scala 27:72]
  wire  _T_21740 = bht_rd_addr_f == 8'ha6; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_166; // @[Reg.scala 27:20]
  wire [1:0] _T_22086 = _T_21740 ? bht_bank_rd_data_out_1_166 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22341 = _T_22340 | _T_22086; // @[Mux.scala 27:72]
  wire  _T_21742 = bht_rd_addr_f == 8'ha7; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_167; // @[Reg.scala 27:20]
  wire [1:0] _T_22087 = _T_21742 ? bht_bank_rd_data_out_1_167 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22342 = _T_22341 | _T_22087; // @[Mux.scala 27:72]
  wire  _T_21744 = bht_rd_addr_f == 8'ha8; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_168; // @[Reg.scala 27:20]
  wire [1:0] _T_22088 = _T_21744 ? bht_bank_rd_data_out_1_168 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22343 = _T_22342 | _T_22088; // @[Mux.scala 27:72]
  wire  _T_21746 = bht_rd_addr_f == 8'ha9; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_169; // @[Reg.scala 27:20]
  wire [1:0] _T_22089 = _T_21746 ? bht_bank_rd_data_out_1_169 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22344 = _T_22343 | _T_22089; // @[Mux.scala 27:72]
  wire  _T_21748 = bht_rd_addr_f == 8'haa; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_170; // @[Reg.scala 27:20]
  wire [1:0] _T_22090 = _T_21748 ? bht_bank_rd_data_out_1_170 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22345 = _T_22344 | _T_22090; // @[Mux.scala 27:72]
  wire  _T_21750 = bht_rd_addr_f == 8'hab; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_171; // @[Reg.scala 27:20]
  wire [1:0] _T_22091 = _T_21750 ? bht_bank_rd_data_out_1_171 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22346 = _T_22345 | _T_22091; // @[Mux.scala 27:72]
  wire  _T_21752 = bht_rd_addr_f == 8'hac; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_172; // @[Reg.scala 27:20]
  wire [1:0] _T_22092 = _T_21752 ? bht_bank_rd_data_out_1_172 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22347 = _T_22346 | _T_22092; // @[Mux.scala 27:72]
  wire  _T_21754 = bht_rd_addr_f == 8'had; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_173; // @[Reg.scala 27:20]
  wire [1:0] _T_22093 = _T_21754 ? bht_bank_rd_data_out_1_173 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22348 = _T_22347 | _T_22093; // @[Mux.scala 27:72]
  wire  _T_21756 = bht_rd_addr_f == 8'hae; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_174; // @[Reg.scala 27:20]
  wire [1:0] _T_22094 = _T_21756 ? bht_bank_rd_data_out_1_174 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22349 = _T_22348 | _T_22094; // @[Mux.scala 27:72]
  wire  _T_21758 = bht_rd_addr_f == 8'haf; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_175; // @[Reg.scala 27:20]
  wire [1:0] _T_22095 = _T_21758 ? bht_bank_rd_data_out_1_175 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22350 = _T_22349 | _T_22095; // @[Mux.scala 27:72]
  wire  _T_21760 = bht_rd_addr_f == 8'hb0; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_176; // @[Reg.scala 27:20]
  wire [1:0] _T_22096 = _T_21760 ? bht_bank_rd_data_out_1_176 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22351 = _T_22350 | _T_22096; // @[Mux.scala 27:72]
  wire  _T_21762 = bht_rd_addr_f == 8'hb1; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_177; // @[Reg.scala 27:20]
  wire [1:0] _T_22097 = _T_21762 ? bht_bank_rd_data_out_1_177 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22352 = _T_22351 | _T_22097; // @[Mux.scala 27:72]
  wire  _T_21764 = bht_rd_addr_f == 8'hb2; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_178; // @[Reg.scala 27:20]
  wire [1:0] _T_22098 = _T_21764 ? bht_bank_rd_data_out_1_178 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22353 = _T_22352 | _T_22098; // @[Mux.scala 27:72]
  wire  _T_21766 = bht_rd_addr_f == 8'hb3; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_179; // @[Reg.scala 27:20]
  wire [1:0] _T_22099 = _T_21766 ? bht_bank_rd_data_out_1_179 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22354 = _T_22353 | _T_22099; // @[Mux.scala 27:72]
  wire  _T_21768 = bht_rd_addr_f == 8'hb4; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_180; // @[Reg.scala 27:20]
  wire [1:0] _T_22100 = _T_21768 ? bht_bank_rd_data_out_1_180 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22355 = _T_22354 | _T_22100; // @[Mux.scala 27:72]
  wire  _T_21770 = bht_rd_addr_f == 8'hb5; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_181; // @[Reg.scala 27:20]
  wire [1:0] _T_22101 = _T_21770 ? bht_bank_rd_data_out_1_181 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22356 = _T_22355 | _T_22101; // @[Mux.scala 27:72]
  wire  _T_21772 = bht_rd_addr_f == 8'hb6; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_182; // @[Reg.scala 27:20]
  wire [1:0] _T_22102 = _T_21772 ? bht_bank_rd_data_out_1_182 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22357 = _T_22356 | _T_22102; // @[Mux.scala 27:72]
  wire  _T_21774 = bht_rd_addr_f == 8'hb7; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_183; // @[Reg.scala 27:20]
  wire [1:0] _T_22103 = _T_21774 ? bht_bank_rd_data_out_1_183 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22358 = _T_22357 | _T_22103; // @[Mux.scala 27:72]
  wire  _T_21776 = bht_rd_addr_f == 8'hb8; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_184; // @[Reg.scala 27:20]
  wire [1:0] _T_22104 = _T_21776 ? bht_bank_rd_data_out_1_184 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22359 = _T_22358 | _T_22104; // @[Mux.scala 27:72]
  wire  _T_21778 = bht_rd_addr_f == 8'hb9; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_185; // @[Reg.scala 27:20]
  wire [1:0] _T_22105 = _T_21778 ? bht_bank_rd_data_out_1_185 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22360 = _T_22359 | _T_22105; // @[Mux.scala 27:72]
  wire  _T_21780 = bht_rd_addr_f == 8'hba; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_186; // @[Reg.scala 27:20]
  wire [1:0] _T_22106 = _T_21780 ? bht_bank_rd_data_out_1_186 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22361 = _T_22360 | _T_22106; // @[Mux.scala 27:72]
  wire  _T_21782 = bht_rd_addr_f == 8'hbb; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_187; // @[Reg.scala 27:20]
  wire [1:0] _T_22107 = _T_21782 ? bht_bank_rd_data_out_1_187 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22362 = _T_22361 | _T_22107; // @[Mux.scala 27:72]
  wire  _T_21784 = bht_rd_addr_f == 8'hbc; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_188; // @[Reg.scala 27:20]
  wire [1:0] _T_22108 = _T_21784 ? bht_bank_rd_data_out_1_188 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22363 = _T_22362 | _T_22108; // @[Mux.scala 27:72]
  wire  _T_21786 = bht_rd_addr_f == 8'hbd; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_189; // @[Reg.scala 27:20]
  wire [1:0] _T_22109 = _T_21786 ? bht_bank_rd_data_out_1_189 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22364 = _T_22363 | _T_22109; // @[Mux.scala 27:72]
  wire  _T_21788 = bht_rd_addr_f == 8'hbe; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_190; // @[Reg.scala 27:20]
  wire [1:0] _T_22110 = _T_21788 ? bht_bank_rd_data_out_1_190 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22365 = _T_22364 | _T_22110; // @[Mux.scala 27:72]
  wire  _T_21790 = bht_rd_addr_f == 8'hbf; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_191; // @[Reg.scala 27:20]
  wire [1:0] _T_22111 = _T_21790 ? bht_bank_rd_data_out_1_191 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22366 = _T_22365 | _T_22111; // @[Mux.scala 27:72]
  wire  _T_21792 = bht_rd_addr_f == 8'hc0; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_192; // @[Reg.scala 27:20]
  wire [1:0] _T_22112 = _T_21792 ? bht_bank_rd_data_out_1_192 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22367 = _T_22366 | _T_22112; // @[Mux.scala 27:72]
  wire  _T_21794 = bht_rd_addr_f == 8'hc1; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_193; // @[Reg.scala 27:20]
  wire [1:0] _T_22113 = _T_21794 ? bht_bank_rd_data_out_1_193 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22368 = _T_22367 | _T_22113; // @[Mux.scala 27:72]
  wire  _T_21796 = bht_rd_addr_f == 8'hc2; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_194; // @[Reg.scala 27:20]
  wire [1:0] _T_22114 = _T_21796 ? bht_bank_rd_data_out_1_194 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22369 = _T_22368 | _T_22114; // @[Mux.scala 27:72]
  wire  _T_21798 = bht_rd_addr_f == 8'hc3; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_195; // @[Reg.scala 27:20]
  wire [1:0] _T_22115 = _T_21798 ? bht_bank_rd_data_out_1_195 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22370 = _T_22369 | _T_22115; // @[Mux.scala 27:72]
  wire  _T_21800 = bht_rd_addr_f == 8'hc4; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_196; // @[Reg.scala 27:20]
  wire [1:0] _T_22116 = _T_21800 ? bht_bank_rd_data_out_1_196 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22371 = _T_22370 | _T_22116; // @[Mux.scala 27:72]
  wire  _T_21802 = bht_rd_addr_f == 8'hc5; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_197; // @[Reg.scala 27:20]
  wire [1:0] _T_22117 = _T_21802 ? bht_bank_rd_data_out_1_197 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22372 = _T_22371 | _T_22117; // @[Mux.scala 27:72]
  wire  _T_21804 = bht_rd_addr_f == 8'hc6; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_198; // @[Reg.scala 27:20]
  wire [1:0] _T_22118 = _T_21804 ? bht_bank_rd_data_out_1_198 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22373 = _T_22372 | _T_22118; // @[Mux.scala 27:72]
  wire  _T_21806 = bht_rd_addr_f == 8'hc7; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_199; // @[Reg.scala 27:20]
  wire [1:0] _T_22119 = _T_21806 ? bht_bank_rd_data_out_1_199 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22374 = _T_22373 | _T_22119; // @[Mux.scala 27:72]
  wire  _T_21808 = bht_rd_addr_f == 8'hc8; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_200; // @[Reg.scala 27:20]
  wire [1:0] _T_22120 = _T_21808 ? bht_bank_rd_data_out_1_200 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22375 = _T_22374 | _T_22120; // @[Mux.scala 27:72]
  wire  _T_21810 = bht_rd_addr_f == 8'hc9; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_201; // @[Reg.scala 27:20]
  wire [1:0] _T_22121 = _T_21810 ? bht_bank_rd_data_out_1_201 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22376 = _T_22375 | _T_22121; // @[Mux.scala 27:72]
  wire  _T_21812 = bht_rd_addr_f == 8'hca; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_202; // @[Reg.scala 27:20]
  wire [1:0] _T_22122 = _T_21812 ? bht_bank_rd_data_out_1_202 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22377 = _T_22376 | _T_22122; // @[Mux.scala 27:72]
  wire  _T_21814 = bht_rd_addr_f == 8'hcb; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_203; // @[Reg.scala 27:20]
  wire [1:0] _T_22123 = _T_21814 ? bht_bank_rd_data_out_1_203 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22378 = _T_22377 | _T_22123; // @[Mux.scala 27:72]
  wire  _T_21816 = bht_rd_addr_f == 8'hcc; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_204; // @[Reg.scala 27:20]
  wire [1:0] _T_22124 = _T_21816 ? bht_bank_rd_data_out_1_204 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22379 = _T_22378 | _T_22124; // @[Mux.scala 27:72]
  wire  _T_21818 = bht_rd_addr_f == 8'hcd; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_205; // @[Reg.scala 27:20]
  wire [1:0] _T_22125 = _T_21818 ? bht_bank_rd_data_out_1_205 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22380 = _T_22379 | _T_22125; // @[Mux.scala 27:72]
  wire  _T_21820 = bht_rd_addr_f == 8'hce; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_206; // @[Reg.scala 27:20]
  wire [1:0] _T_22126 = _T_21820 ? bht_bank_rd_data_out_1_206 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22381 = _T_22380 | _T_22126; // @[Mux.scala 27:72]
  wire  _T_21822 = bht_rd_addr_f == 8'hcf; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_207; // @[Reg.scala 27:20]
  wire [1:0] _T_22127 = _T_21822 ? bht_bank_rd_data_out_1_207 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22382 = _T_22381 | _T_22127; // @[Mux.scala 27:72]
  wire  _T_21824 = bht_rd_addr_f == 8'hd0; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_208; // @[Reg.scala 27:20]
  wire [1:0] _T_22128 = _T_21824 ? bht_bank_rd_data_out_1_208 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22383 = _T_22382 | _T_22128; // @[Mux.scala 27:72]
  wire  _T_21826 = bht_rd_addr_f == 8'hd1; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_209; // @[Reg.scala 27:20]
  wire [1:0] _T_22129 = _T_21826 ? bht_bank_rd_data_out_1_209 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22384 = _T_22383 | _T_22129; // @[Mux.scala 27:72]
  wire  _T_21828 = bht_rd_addr_f == 8'hd2; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_210; // @[Reg.scala 27:20]
  wire [1:0] _T_22130 = _T_21828 ? bht_bank_rd_data_out_1_210 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22385 = _T_22384 | _T_22130; // @[Mux.scala 27:72]
  wire  _T_21830 = bht_rd_addr_f == 8'hd3; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_211; // @[Reg.scala 27:20]
  wire [1:0] _T_22131 = _T_21830 ? bht_bank_rd_data_out_1_211 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22386 = _T_22385 | _T_22131; // @[Mux.scala 27:72]
  wire  _T_21832 = bht_rd_addr_f == 8'hd4; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_212; // @[Reg.scala 27:20]
  wire [1:0] _T_22132 = _T_21832 ? bht_bank_rd_data_out_1_212 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22387 = _T_22386 | _T_22132; // @[Mux.scala 27:72]
  wire  _T_21834 = bht_rd_addr_f == 8'hd5; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_213; // @[Reg.scala 27:20]
  wire [1:0] _T_22133 = _T_21834 ? bht_bank_rd_data_out_1_213 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22388 = _T_22387 | _T_22133; // @[Mux.scala 27:72]
  wire  _T_21836 = bht_rd_addr_f == 8'hd6; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_214; // @[Reg.scala 27:20]
  wire [1:0] _T_22134 = _T_21836 ? bht_bank_rd_data_out_1_214 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22389 = _T_22388 | _T_22134; // @[Mux.scala 27:72]
  wire  _T_21838 = bht_rd_addr_f == 8'hd7; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_215; // @[Reg.scala 27:20]
  wire [1:0] _T_22135 = _T_21838 ? bht_bank_rd_data_out_1_215 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22390 = _T_22389 | _T_22135; // @[Mux.scala 27:72]
  wire  _T_21840 = bht_rd_addr_f == 8'hd8; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_216; // @[Reg.scala 27:20]
  wire [1:0] _T_22136 = _T_21840 ? bht_bank_rd_data_out_1_216 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22391 = _T_22390 | _T_22136; // @[Mux.scala 27:72]
  wire  _T_21842 = bht_rd_addr_f == 8'hd9; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_217; // @[Reg.scala 27:20]
  wire [1:0] _T_22137 = _T_21842 ? bht_bank_rd_data_out_1_217 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22392 = _T_22391 | _T_22137; // @[Mux.scala 27:72]
  wire  _T_21844 = bht_rd_addr_f == 8'hda; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_218; // @[Reg.scala 27:20]
  wire [1:0] _T_22138 = _T_21844 ? bht_bank_rd_data_out_1_218 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22393 = _T_22392 | _T_22138; // @[Mux.scala 27:72]
  wire  _T_21846 = bht_rd_addr_f == 8'hdb; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_219; // @[Reg.scala 27:20]
  wire [1:0] _T_22139 = _T_21846 ? bht_bank_rd_data_out_1_219 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22394 = _T_22393 | _T_22139; // @[Mux.scala 27:72]
  wire  _T_21848 = bht_rd_addr_f == 8'hdc; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_220; // @[Reg.scala 27:20]
  wire [1:0] _T_22140 = _T_21848 ? bht_bank_rd_data_out_1_220 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22395 = _T_22394 | _T_22140; // @[Mux.scala 27:72]
  wire  _T_21850 = bht_rd_addr_f == 8'hdd; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_221; // @[Reg.scala 27:20]
  wire [1:0] _T_22141 = _T_21850 ? bht_bank_rd_data_out_1_221 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22396 = _T_22395 | _T_22141; // @[Mux.scala 27:72]
  wire  _T_21852 = bht_rd_addr_f == 8'hde; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_222; // @[Reg.scala 27:20]
  wire [1:0] _T_22142 = _T_21852 ? bht_bank_rd_data_out_1_222 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22397 = _T_22396 | _T_22142; // @[Mux.scala 27:72]
  wire  _T_21854 = bht_rd_addr_f == 8'hdf; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_223; // @[Reg.scala 27:20]
  wire [1:0] _T_22143 = _T_21854 ? bht_bank_rd_data_out_1_223 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22398 = _T_22397 | _T_22143; // @[Mux.scala 27:72]
  wire  _T_21856 = bht_rd_addr_f == 8'he0; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_224; // @[Reg.scala 27:20]
  wire [1:0] _T_22144 = _T_21856 ? bht_bank_rd_data_out_1_224 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22399 = _T_22398 | _T_22144; // @[Mux.scala 27:72]
  wire  _T_21858 = bht_rd_addr_f == 8'he1; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_225; // @[Reg.scala 27:20]
  wire [1:0] _T_22145 = _T_21858 ? bht_bank_rd_data_out_1_225 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22400 = _T_22399 | _T_22145; // @[Mux.scala 27:72]
  wire  _T_21860 = bht_rd_addr_f == 8'he2; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_226; // @[Reg.scala 27:20]
  wire [1:0] _T_22146 = _T_21860 ? bht_bank_rd_data_out_1_226 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22401 = _T_22400 | _T_22146; // @[Mux.scala 27:72]
  wire  _T_21862 = bht_rd_addr_f == 8'he3; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_227; // @[Reg.scala 27:20]
  wire [1:0] _T_22147 = _T_21862 ? bht_bank_rd_data_out_1_227 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22402 = _T_22401 | _T_22147; // @[Mux.scala 27:72]
  wire  _T_21864 = bht_rd_addr_f == 8'he4; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_228; // @[Reg.scala 27:20]
  wire [1:0] _T_22148 = _T_21864 ? bht_bank_rd_data_out_1_228 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22403 = _T_22402 | _T_22148; // @[Mux.scala 27:72]
  wire  _T_21866 = bht_rd_addr_f == 8'he5; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_229; // @[Reg.scala 27:20]
  wire [1:0] _T_22149 = _T_21866 ? bht_bank_rd_data_out_1_229 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22404 = _T_22403 | _T_22149; // @[Mux.scala 27:72]
  wire  _T_21868 = bht_rd_addr_f == 8'he6; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_230; // @[Reg.scala 27:20]
  wire [1:0] _T_22150 = _T_21868 ? bht_bank_rd_data_out_1_230 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22405 = _T_22404 | _T_22150; // @[Mux.scala 27:72]
  wire  _T_21870 = bht_rd_addr_f == 8'he7; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_231; // @[Reg.scala 27:20]
  wire [1:0] _T_22151 = _T_21870 ? bht_bank_rd_data_out_1_231 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22406 = _T_22405 | _T_22151; // @[Mux.scala 27:72]
  wire  _T_21872 = bht_rd_addr_f == 8'he8; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_232; // @[Reg.scala 27:20]
  wire [1:0] _T_22152 = _T_21872 ? bht_bank_rd_data_out_1_232 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22407 = _T_22406 | _T_22152; // @[Mux.scala 27:72]
  wire  _T_21874 = bht_rd_addr_f == 8'he9; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_233; // @[Reg.scala 27:20]
  wire [1:0] _T_22153 = _T_21874 ? bht_bank_rd_data_out_1_233 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22408 = _T_22407 | _T_22153; // @[Mux.scala 27:72]
  wire  _T_21876 = bht_rd_addr_f == 8'hea; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_234; // @[Reg.scala 27:20]
  wire [1:0] _T_22154 = _T_21876 ? bht_bank_rd_data_out_1_234 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22409 = _T_22408 | _T_22154; // @[Mux.scala 27:72]
  wire  _T_21878 = bht_rd_addr_f == 8'heb; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_235; // @[Reg.scala 27:20]
  wire [1:0] _T_22155 = _T_21878 ? bht_bank_rd_data_out_1_235 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22410 = _T_22409 | _T_22155; // @[Mux.scala 27:72]
  wire  _T_21880 = bht_rd_addr_f == 8'hec; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_236; // @[Reg.scala 27:20]
  wire [1:0] _T_22156 = _T_21880 ? bht_bank_rd_data_out_1_236 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22411 = _T_22410 | _T_22156; // @[Mux.scala 27:72]
  wire  _T_21882 = bht_rd_addr_f == 8'hed; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_237; // @[Reg.scala 27:20]
  wire [1:0] _T_22157 = _T_21882 ? bht_bank_rd_data_out_1_237 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22412 = _T_22411 | _T_22157; // @[Mux.scala 27:72]
  wire  _T_21884 = bht_rd_addr_f == 8'hee; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_238; // @[Reg.scala 27:20]
  wire [1:0] _T_22158 = _T_21884 ? bht_bank_rd_data_out_1_238 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22413 = _T_22412 | _T_22158; // @[Mux.scala 27:72]
  wire  _T_21886 = bht_rd_addr_f == 8'hef; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_239; // @[Reg.scala 27:20]
  wire [1:0] _T_22159 = _T_21886 ? bht_bank_rd_data_out_1_239 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22414 = _T_22413 | _T_22159; // @[Mux.scala 27:72]
  wire  _T_21888 = bht_rd_addr_f == 8'hf0; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_240; // @[Reg.scala 27:20]
  wire [1:0] _T_22160 = _T_21888 ? bht_bank_rd_data_out_1_240 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22415 = _T_22414 | _T_22160; // @[Mux.scala 27:72]
  wire  _T_21890 = bht_rd_addr_f == 8'hf1; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_241; // @[Reg.scala 27:20]
  wire [1:0] _T_22161 = _T_21890 ? bht_bank_rd_data_out_1_241 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22416 = _T_22415 | _T_22161; // @[Mux.scala 27:72]
  wire  _T_21892 = bht_rd_addr_f == 8'hf2; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_242; // @[Reg.scala 27:20]
  wire [1:0] _T_22162 = _T_21892 ? bht_bank_rd_data_out_1_242 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22417 = _T_22416 | _T_22162; // @[Mux.scala 27:72]
  wire  _T_21894 = bht_rd_addr_f == 8'hf3; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_243; // @[Reg.scala 27:20]
  wire [1:0] _T_22163 = _T_21894 ? bht_bank_rd_data_out_1_243 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22418 = _T_22417 | _T_22163; // @[Mux.scala 27:72]
  wire  _T_21896 = bht_rd_addr_f == 8'hf4; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_244; // @[Reg.scala 27:20]
  wire [1:0] _T_22164 = _T_21896 ? bht_bank_rd_data_out_1_244 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22419 = _T_22418 | _T_22164; // @[Mux.scala 27:72]
  wire  _T_21898 = bht_rd_addr_f == 8'hf5; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_245; // @[Reg.scala 27:20]
  wire [1:0] _T_22165 = _T_21898 ? bht_bank_rd_data_out_1_245 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22420 = _T_22419 | _T_22165; // @[Mux.scala 27:72]
  wire  _T_21900 = bht_rd_addr_f == 8'hf6; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_246; // @[Reg.scala 27:20]
  wire [1:0] _T_22166 = _T_21900 ? bht_bank_rd_data_out_1_246 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22421 = _T_22420 | _T_22166; // @[Mux.scala 27:72]
  wire  _T_21902 = bht_rd_addr_f == 8'hf7; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_247; // @[Reg.scala 27:20]
  wire [1:0] _T_22167 = _T_21902 ? bht_bank_rd_data_out_1_247 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22422 = _T_22421 | _T_22167; // @[Mux.scala 27:72]
  wire  _T_21904 = bht_rd_addr_f == 8'hf8; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_248; // @[Reg.scala 27:20]
  wire [1:0] _T_22168 = _T_21904 ? bht_bank_rd_data_out_1_248 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22423 = _T_22422 | _T_22168; // @[Mux.scala 27:72]
  wire  _T_21906 = bht_rd_addr_f == 8'hf9; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_249; // @[Reg.scala 27:20]
  wire [1:0] _T_22169 = _T_21906 ? bht_bank_rd_data_out_1_249 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22424 = _T_22423 | _T_22169; // @[Mux.scala 27:72]
  wire  _T_21908 = bht_rd_addr_f == 8'hfa; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_250; // @[Reg.scala 27:20]
  wire [1:0] _T_22170 = _T_21908 ? bht_bank_rd_data_out_1_250 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22425 = _T_22424 | _T_22170; // @[Mux.scala 27:72]
  wire  _T_21910 = bht_rd_addr_f == 8'hfb; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_251; // @[Reg.scala 27:20]
  wire [1:0] _T_22171 = _T_21910 ? bht_bank_rd_data_out_1_251 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22426 = _T_22425 | _T_22171; // @[Mux.scala 27:72]
  wire  _T_21912 = bht_rd_addr_f == 8'hfc; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_252; // @[Reg.scala 27:20]
  wire [1:0] _T_22172 = _T_21912 ? bht_bank_rd_data_out_1_252 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22427 = _T_22426 | _T_22172; // @[Mux.scala 27:72]
  wire  _T_21914 = bht_rd_addr_f == 8'hfd; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_253; // @[Reg.scala 27:20]
  wire [1:0] _T_22173 = _T_21914 ? bht_bank_rd_data_out_1_253 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22428 = _T_22427 | _T_22173; // @[Mux.scala 27:72]
  wire  _T_21916 = bht_rd_addr_f == 8'hfe; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_254; // @[Reg.scala 27:20]
  wire [1:0] _T_22174 = _T_21916 ? bht_bank_rd_data_out_1_254 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22429 = _T_22428 | _T_22174; // @[Mux.scala 27:72]
  wire  _T_21918 = bht_rd_addr_f == 8'hff; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_255; // @[Reg.scala 27:20]
  wire [1:0] _T_22175 = _T_21918 ? bht_bank_rd_data_out_1_255 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] bht_bank1_rd_data_f = _T_22429 | _T_22175; // @[Mux.scala 27:72]
  wire [1:0] _T_260 = _T_144 ? bht_bank1_rd_data_f : 2'h0; // @[Mux.scala 27:72]
  wire [9:0] _T_573 = {btb_rd_addr_p1_f,2'h0}; // @[Cat.scala 29:58]
  wire [7:0] bht_rd_addr_hashed_p1_f = _T_573[9:2] ^ fghr; // @[lib.scala 56:35]
  wire  _T_22432 = bht_rd_addr_hashed_p1_f == 8'h0; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_0; // @[Reg.scala 27:20]
  wire [1:0] _T_22944 = _T_22432 ? bht_bank_rd_data_out_0_0 : 2'h0; // @[Mux.scala 27:72]
  wire  _T_22434 = bht_rd_addr_hashed_p1_f == 8'h1; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_1; // @[Reg.scala 27:20]
  wire [1:0] _T_22945 = _T_22434 ? bht_bank_rd_data_out_0_1 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23200 = _T_22944 | _T_22945; // @[Mux.scala 27:72]
  wire  _T_22436 = bht_rd_addr_hashed_p1_f == 8'h2; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_2; // @[Reg.scala 27:20]
  wire [1:0] _T_22946 = _T_22436 ? bht_bank_rd_data_out_0_2 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23201 = _T_23200 | _T_22946; // @[Mux.scala 27:72]
  wire  _T_22438 = bht_rd_addr_hashed_p1_f == 8'h3; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_3; // @[Reg.scala 27:20]
  wire [1:0] _T_22947 = _T_22438 ? bht_bank_rd_data_out_0_3 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23202 = _T_23201 | _T_22947; // @[Mux.scala 27:72]
  wire  _T_22440 = bht_rd_addr_hashed_p1_f == 8'h4; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_4; // @[Reg.scala 27:20]
  wire [1:0] _T_22948 = _T_22440 ? bht_bank_rd_data_out_0_4 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23203 = _T_23202 | _T_22948; // @[Mux.scala 27:72]
  wire  _T_22442 = bht_rd_addr_hashed_p1_f == 8'h5; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_5; // @[Reg.scala 27:20]
  wire [1:0] _T_22949 = _T_22442 ? bht_bank_rd_data_out_0_5 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23204 = _T_23203 | _T_22949; // @[Mux.scala 27:72]
  wire  _T_22444 = bht_rd_addr_hashed_p1_f == 8'h6; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_6; // @[Reg.scala 27:20]
  wire [1:0] _T_22950 = _T_22444 ? bht_bank_rd_data_out_0_6 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23205 = _T_23204 | _T_22950; // @[Mux.scala 27:72]
  wire  _T_22446 = bht_rd_addr_hashed_p1_f == 8'h7; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_7; // @[Reg.scala 27:20]
  wire [1:0] _T_22951 = _T_22446 ? bht_bank_rd_data_out_0_7 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23206 = _T_23205 | _T_22951; // @[Mux.scala 27:72]
  wire  _T_22448 = bht_rd_addr_hashed_p1_f == 8'h8; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_8; // @[Reg.scala 27:20]
  wire [1:0] _T_22952 = _T_22448 ? bht_bank_rd_data_out_0_8 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23207 = _T_23206 | _T_22952; // @[Mux.scala 27:72]
  wire  _T_22450 = bht_rd_addr_hashed_p1_f == 8'h9; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_9; // @[Reg.scala 27:20]
  wire [1:0] _T_22953 = _T_22450 ? bht_bank_rd_data_out_0_9 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23208 = _T_23207 | _T_22953; // @[Mux.scala 27:72]
  wire  _T_22452 = bht_rd_addr_hashed_p1_f == 8'ha; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_10; // @[Reg.scala 27:20]
  wire [1:0] _T_22954 = _T_22452 ? bht_bank_rd_data_out_0_10 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23209 = _T_23208 | _T_22954; // @[Mux.scala 27:72]
  wire  _T_22454 = bht_rd_addr_hashed_p1_f == 8'hb; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_11; // @[Reg.scala 27:20]
  wire [1:0] _T_22955 = _T_22454 ? bht_bank_rd_data_out_0_11 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23210 = _T_23209 | _T_22955; // @[Mux.scala 27:72]
  wire  _T_22456 = bht_rd_addr_hashed_p1_f == 8'hc; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_12; // @[Reg.scala 27:20]
  wire [1:0] _T_22956 = _T_22456 ? bht_bank_rd_data_out_0_12 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23211 = _T_23210 | _T_22956; // @[Mux.scala 27:72]
  wire  _T_22458 = bht_rd_addr_hashed_p1_f == 8'hd; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_13; // @[Reg.scala 27:20]
  wire [1:0] _T_22957 = _T_22458 ? bht_bank_rd_data_out_0_13 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23212 = _T_23211 | _T_22957; // @[Mux.scala 27:72]
  wire  _T_22460 = bht_rd_addr_hashed_p1_f == 8'he; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_14; // @[Reg.scala 27:20]
  wire [1:0] _T_22958 = _T_22460 ? bht_bank_rd_data_out_0_14 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23213 = _T_23212 | _T_22958; // @[Mux.scala 27:72]
  wire  _T_22462 = bht_rd_addr_hashed_p1_f == 8'hf; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_15; // @[Reg.scala 27:20]
  wire [1:0] _T_22959 = _T_22462 ? bht_bank_rd_data_out_0_15 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23214 = _T_23213 | _T_22959; // @[Mux.scala 27:72]
  wire  _T_22464 = bht_rd_addr_hashed_p1_f == 8'h10; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_16; // @[Reg.scala 27:20]
  wire [1:0] _T_22960 = _T_22464 ? bht_bank_rd_data_out_0_16 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23215 = _T_23214 | _T_22960; // @[Mux.scala 27:72]
  wire  _T_22466 = bht_rd_addr_hashed_p1_f == 8'h11; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_17; // @[Reg.scala 27:20]
  wire [1:0] _T_22961 = _T_22466 ? bht_bank_rd_data_out_0_17 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23216 = _T_23215 | _T_22961; // @[Mux.scala 27:72]
  wire  _T_22468 = bht_rd_addr_hashed_p1_f == 8'h12; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_18; // @[Reg.scala 27:20]
  wire [1:0] _T_22962 = _T_22468 ? bht_bank_rd_data_out_0_18 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23217 = _T_23216 | _T_22962; // @[Mux.scala 27:72]
  wire  _T_22470 = bht_rd_addr_hashed_p1_f == 8'h13; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_19; // @[Reg.scala 27:20]
  wire [1:0] _T_22963 = _T_22470 ? bht_bank_rd_data_out_0_19 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23218 = _T_23217 | _T_22963; // @[Mux.scala 27:72]
  wire  _T_22472 = bht_rd_addr_hashed_p1_f == 8'h14; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_20; // @[Reg.scala 27:20]
  wire [1:0] _T_22964 = _T_22472 ? bht_bank_rd_data_out_0_20 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23219 = _T_23218 | _T_22964; // @[Mux.scala 27:72]
  wire  _T_22474 = bht_rd_addr_hashed_p1_f == 8'h15; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_21; // @[Reg.scala 27:20]
  wire [1:0] _T_22965 = _T_22474 ? bht_bank_rd_data_out_0_21 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23220 = _T_23219 | _T_22965; // @[Mux.scala 27:72]
  wire  _T_22476 = bht_rd_addr_hashed_p1_f == 8'h16; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_22; // @[Reg.scala 27:20]
  wire [1:0] _T_22966 = _T_22476 ? bht_bank_rd_data_out_0_22 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23221 = _T_23220 | _T_22966; // @[Mux.scala 27:72]
  wire  _T_22478 = bht_rd_addr_hashed_p1_f == 8'h17; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_23; // @[Reg.scala 27:20]
  wire [1:0] _T_22967 = _T_22478 ? bht_bank_rd_data_out_0_23 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23222 = _T_23221 | _T_22967; // @[Mux.scala 27:72]
  wire  _T_22480 = bht_rd_addr_hashed_p1_f == 8'h18; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_24; // @[Reg.scala 27:20]
  wire [1:0] _T_22968 = _T_22480 ? bht_bank_rd_data_out_0_24 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23223 = _T_23222 | _T_22968; // @[Mux.scala 27:72]
  wire  _T_22482 = bht_rd_addr_hashed_p1_f == 8'h19; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_25; // @[Reg.scala 27:20]
  wire [1:0] _T_22969 = _T_22482 ? bht_bank_rd_data_out_0_25 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23224 = _T_23223 | _T_22969; // @[Mux.scala 27:72]
  wire  _T_22484 = bht_rd_addr_hashed_p1_f == 8'h1a; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_26; // @[Reg.scala 27:20]
  wire [1:0] _T_22970 = _T_22484 ? bht_bank_rd_data_out_0_26 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23225 = _T_23224 | _T_22970; // @[Mux.scala 27:72]
  wire  _T_22486 = bht_rd_addr_hashed_p1_f == 8'h1b; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_27; // @[Reg.scala 27:20]
  wire [1:0] _T_22971 = _T_22486 ? bht_bank_rd_data_out_0_27 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23226 = _T_23225 | _T_22971; // @[Mux.scala 27:72]
  wire  _T_22488 = bht_rd_addr_hashed_p1_f == 8'h1c; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_28; // @[Reg.scala 27:20]
  wire [1:0] _T_22972 = _T_22488 ? bht_bank_rd_data_out_0_28 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23227 = _T_23226 | _T_22972; // @[Mux.scala 27:72]
  wire  _T_22490 = bht_rd_addr_hashed_p1_f == 8'h1d; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_29; // @[Reg.scala 27:20]
  wire [1:0] _T_22973 = _T_22490 ? bht_bank_rd_data_out_0_29 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23228 = _T_23227 | _T_22973; // @[Mux.scala 27:72]
  wire  _T_22492 = bht_rd_addr_hashed_p1_f == 8'h1e; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_30; // @[Reg.scala 27:20]
  wire [1:0] _T_22974 = _T_22492 ? bht_bank_rd_data_out_0_30 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23229 = _T_23228 | _T_22974; // @[Mux.scala 27:72]
  wire  _T_22494 = bht_rd_addr_hashed_p1_f == 8'h1f; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_31; // @[Reg.scala 27:20]
  wire [1:0] _T_22975 = _T_22494 ? bht_bank_rd_data_out_0_31 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23230 = _T_23229 | _T_22975; // @[Mux.scala 27:72]
  wire  _T_22496 = bht_rd_addr_hashed_p1_f == 8'h20; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_32; // @[Reg.scala 27:20]
  wire [1:0] _T_22976 = _T_22496 ? bht_bank_rd_data_out_0_32 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23231 = _T_23230 | _T_22976; // @[Mux.scala 27:72]
  wire  _T_22498 = bht_rd_addr_hashed_p1_f == 8'h21; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_33; // @[Reg.scala 27:20]
  wire [1:0] _T_22977 = _T_22498 ? bht_bank_rd_data_out_0_33 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23232 = _T_23231 | _T_22977; // @[Mux.scala 27:72]
  wire  _T_22500 = bht_rd_addr_hashed_p1_f == 8'h22; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_34; // @[Reg.scala 27:20]
  wire [1:0] _T_22978 = _T_22500 ? bht_bank_rd_data_out_0_34 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23233 = _T_23232 | _T_22978; // @[Mux.scala 27:72]
  wire  _T_22502 = bht_rd_addr_hashed_p1_f == 8'h23; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_35; // @[Reg.scala 27:20]
  wire [1:0] _T_22979 = _T_22502 ? bht_bank_rd_data_out_0_35 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23234 = _T_23233 | _T_22979; // @[Mux.scala 27:72]
  wire  _T_22504 = bht_rd_addr_hashed_p1_f == 8'h24; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_36; // @[Reg.scala 27:20]
  wire [1:0] _T_22980 = _T_22504 ? bht_bank_rd_data_out_0_36 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23235 = _T_23234 | _T_22980; // @[Mux.scala 27:72]
  wire  _T_22506 = bht_rd_addr_hashed_p1_f == 8'h25; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_37; // @[Reg.scala 27:20]
  wire [1:0] _T_22981 = _T_22506 ? bht_bank_rd_data_out_0_37 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23236 = _T_23235 | _T_22981; // @[Mux.scala 27:72]
  wire  _T_22508 = bht_rd_addr_hashed_p1_f == 8'h26; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_38; // @[Reg.scala 27:20]
  wire [1:0] _T_22982 = _T_22508 ? bht_bank_rd_data_out_0_38 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23237 = _T_23236 | _T_22982; // @[Mux.scala 27:72]
  wire  _T_22510 = bht_rd_addr_hashed_p1_f == 8'h27; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_39; // @[Reg.scala 27:20]
  wire [1:0] _T_22983 = _T_22510 ? bht_bank_rd_data_out_0_39 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23238 = _T_23237 | _T_22983; // @[Mux.scala 27:72]
  wire  _T_22512 = bht_rd_addr_hashed_p1_f == 8'h28; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_40; // @[Reg.scala 27:20]
  wire [1:0] _T_22984 = _T_22512 ? bht_bank_rd_data_out_0_40 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23239 = _T_23238 | _T_22984; // @[Mux.scala 27:72]
  wire  _T_22514 = bht_rd_addr_hashed_p1_f == 8'h29; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_41; // @[Reg.scala 27:20]
  wire [1:0] _T_22985 = _T_22514 ? bht_bank_rd_data_out_0_41 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23240 = _T_23239 | _T_22985; // @[Mux.scala 27:72]
  wire  _T_22516 = bht_rd_addr_hashed_p1_f == 8'h2a; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_42; // @[Reg.scala 27:20]
  wire [1:0] _T_22986 = _T_22516 ? bht_bank_rd_data_out_0_42 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23241 = _T_23240 | _T_22986; // @[Mux.scala 27:72]
  wire  _T_22518 = bht_rd_addr_hashed_p1_f == 8'h2b; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_43; // @[Reg.scala 27:20]
  wire [1:0] _T_22987 = _T_22518 ? bht_bank_rd_data_out_0_43 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23242 = _T_23241 | _T_22987; // @[Mux.scala 27:72]
  wire  _T_22520 = bht_rd_addr_hashed_p1_f == 8'h2c; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_44; // @[Reg.scala 27:20]
  wire [1:0] _T_22988 = _T_22520 ? bht_bank_rd_data_out_0_44 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23243 = _T_23242 | _T_22988; // @[Mux.scala 27:72]
  wire  _T_22522 = bht_rd_addr_hashed_p1_f == 8'h2d; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_45; // @[Reg.scala 27:20]
  wire [1:0] _T_22989 = _T_22522 ? bht_bank_rd_data_out_0_45 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23244 = _T_23243 | _T_22989; // @[Mux.scala 27:72]
  wire  _T_22524 = bht_rd_addr_hashed_p1_f == 8'h2e; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_46; // @[Reg.scala 27:20]
  wire [1:0] _T_22990 = _T_22524 ? bht_bank_rd_data_out_0_46 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23245 = _T_23244 | _T_22990; // @[Mux.scala 27:72]
  wire  _T_22526 = bht_rd_addr_hashed_p1_f == 8'h2f; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_47; // @[Reg.scala 27:20]
  wire [1:0] _T_22991 = _T_22526 ? bht_bank_rd_data_out_0_47 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23246 = _T_23245 | _T_22991; // @[Mux.scala 27:72]
  wire  _T_22528 = bht_rd_addr_hashed_p1_f == 8'h30; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_48; // @[Reg.scala 27:20]
  wire [1:0] _T_22992 = _T_22528 ? bht_bank_rd_data_out_0_48 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23247 = _T_23246 | _T_22992; // @[Mux.scala 27:72]
  wire  _T_22530 = bht_rd_addr_hashed_p1_f == 8'h31; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_49; // @[Reg.scala 27:20]
  wire [1:0] _T_22993 = _T_22530 ? bht_bank_rd_data_out_0_49 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23248 = _T_23247 | _T_22993; // @[Mux.scala 27:72]
  wire  _T_22532 = bht_rd_addr_hashed_p1_f == 8'h32; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_50; // @[Reg.scala 27:20]
  wire [1:0] _T_22994 = _T_22532 ? bht_bank_rd_data_out_0_50 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23249 = _T_23248 | _T_22994; // @[Mux.scala 27:72]
  wire  _T_22534 = bht_rd_addr_hashed_p1_f == 8'h33; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_51; // @[Reg.scala 27:20]
  wire [1:0] _T_22995 = _T_22534 ? bht_bank_rd_data_out_0_51 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23250 = _T_23249 | _T_22995; // @[Mux.scala 27:72]
  wire  _T_22536 = bht_rd_addr_hashed_p1_f == 8'h34; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_52; // @[Reg.scala 27:20]
  wire [1:0] _T_22996 = _T_22536 ? bht_bank_rd_data_out_0_52 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23251 = _T_23250 | _T_22996; // @[Mux.scala 27:72]
  wire  _T_22538 = bht_rd_addr_hashed_p1_f == 8'h35; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_53; // @[Reg.scala 27:20]
  wire [1:0] _T_22997 = _T_22538 ? bht_bank_rd_data_out_0_53 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23252 = _T_23251 | _T_22997; // @[Mux.scala 27:72]
  wire  _T_22540 = bht_rd_addr_hashed_p1_f == 8'h36; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_54; // @[Reg.scala 27:20]
  wire [1:0] _T_22998 = _T_22540 ? bht_bank_rd_data_out_0_54 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23253 = _T_23252 | _T_22998; // @[Mux.scala 27:72]
  wire  _T_22542 = bht_rd_addr_hashed_p1_f == 8'h37; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_55; // @[Reg.scala 27:20]
  wire [1:0] _T_22999 = _T_22542 ? bht_bank_rd_data_out_0_55 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23254 = _T_23253 | _T_22999; // @[Mux.scala 27:72]
  wire  _T_22544 = bht_rd_addr_hashed_p1_f == 8'h38; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_56; // @[Reg.scala 27:20]
  wire [1:0] _T_23000 = _T_22544 ? bht_bank_rd_data_out_0_56 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23255 = _T_23254 | _T_23000; // @[Mux.scala 27:72]
  wire  _T_22546 = bht_rd_addr_hashed_p1_f == 8'h39; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_57; // @[Reg.scala 27:20]
  wire [1:0] _T_23001 = _T_22546 ? bht_bank_rd_data_out_0_57 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23256 = _T_23255 | _T_23001; // @[Mux.scala 27:72]
  wire  _T_22548 = bht_rd_addr_hashed_p1_f == 8'h3a; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_58; // @[Reg.scala 27:20]
  wire [1:0] _T_23002 = _T_22548 ? bht_bank_rd_data_out_0_58 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23257 = _T_23256 | _T_23002; // @[Mux.scala 27:72]
  wire  _T_22550 = bht_rd_addr_hashed_p1_f == 8'h3b; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_59; // @[Reg.scala 27:20]
  wire [1:0] _T_23003 = _T_22550 ? bht_bank_rd_data_out_0_59 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23258 = _T_23257 | _T_23003; // @[Mux.scala 27:72]
  wire  _T_22552 = bht_rd_addr_hashed_p1_f == 8'h3c; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_60; // @[Reg.scala 27:20]
  wire [1:0] _T_23004 = _T_22552 ? bht_bank_rd_data_out_0_60 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23259 = _T_23258 | _T_23004; // @[Mux.scala 27:72]
  wire  _T_22554 = bht_rd_addr_hashed_p1_f == 8'h3d; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_61; // @[Reg.scala 27:20]
  wire [1:0] _T_23005 = _T_22554 ? bht_bank_rd_data_out_0_61 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23260 = _T_23259 | _T_23005; // @[Mux.scala 27:72]
  wire  _T_22556 = bht_rd_addr_hashed_p1_f == 8'h3e; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_62; // @[Reg.scala 27:20]
  wire [1:0] _T_23006 = _T_22556 ? bht_bank_rd_data_out_0_62 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23261 = _T_23260 | _T_23006; // @[Mux.scala 27:72]
  wire  _T_22558 = bht_rd_addr_hashed_p1_f == 8'h3f; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_63; // @[Reg.scala 27:20]
  wire [1:0] _T_23007 = _T_22558 ? bht_bank_rd_data_out_0_63 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23262 = _T_23261 | _T_23007; // @[Mux.scala 27:72]
  wire  _T_22560 = bht_rd_addr_hashed_p1_f == 8'h40; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_64; // @[Reg.scala 27:20]
  wire [1:0] _T_23008 = _T_22560 ? bht_bank_rd_data_out_0_64 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23263 = _T_23262 | _T_23008; // @[Mux.scala 27:72]
  wire  _T_22562 = bht_rd_addr_hashed_p1_f == 8'h41; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_65; // @[Reg.scala 27:20]
  wire [1:0] _T_23009 = _T_22562 ? bht_bank_rd_data_out_0_65 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23264 = _T_23263 | _T_23009; // @[Mux.scala 27:72]
  wire  _T_22564 = bht_rd_addr_hashed_p1_f == 8'h42; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_66; // @[Reg.scala 27:20]
  wire [1:0] _T_23010 = _T_22564 ? bht_bank_rd_data_out_0_66 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23265 = _T_23264 | _T_23010; // @[Mux.scala 27:72]
  wire  _T_22566 = bht_rd_addr_hashed_p1_f == 8'h43; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_67; // @[Reg.scala 27:20]
  wire [1:0] _T_23011 = _T_22566 ? bht_bank_rd_data_out_0_67 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23266 = _T_23265 | _T_23011; // @[Mux.scala 27:72]
  wire  _T_22568 = bht_rd_addr_hashed_p1_f == 8'h44; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_68; // @[Reg.scala 27:20]
  wire [1:0] _T_23012 = _T_22568 ? bht_bank_rd_data_out_0_68 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23267 = _T_23266 | _T_23012; // @[Mux.scala 27:72]
  wire  _T_22570 = bht_rd_addr_hashed_p1_f == 8'h45; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_69; // @[Reg.scala 27:20]
  wire [1:0] _T_23013 = _T_22570 ? bht_bank_rd_data_out_0_69 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23268 = _T_23267 | _T_23013; // @[Mux.scala 27:72]
  wire  _T_22572 = bht_rd_addr_hashed_p1_f == 8'h46; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_70; // @[Reg.scala 27:20]
  wire [1:0] _T_23014 = _T_22572 ? bht_bank_rd_data_out_0_70 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23269 = _T_23268 | _T_23014; // @[Mux.scala 27:72]
  wire  _T_22574 = bht_rd_addr_hashed_p1_f == 8'h47; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_71; // @[Reg.scala 27:20]
  wire [1:0] _T_23015 = _T_22574 ? bht_bank_rd_data_out_0_71 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23270 = _T_23269 | _T_23015; // @[Mux.scala 27:72]
  wire  _T_22576 = bht_rd_addr_hashed_p1_f == 8'h48; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_72; // @[Reg.scala 27:20]
  wire [1:0] _T_23016 = _T_22576 ? bht_bank_rd_data_out_0_72 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23271 = _T_23270 | _T_23016; // @[Mux.scala 27:72]
  wire  _T_22578 = bht_rd_addr_hashed_p1_f == 8'h49; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_73; // @[Reg.scala 27:20]
  wire [1:0] _T_23017 = _T_22578 ? bht_bank_rd_data_out_0_73 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23272 = _T_23271 | _T_23017; // @[Mux.scala 27:72]
  wire  _T_22580 = bht_rd_addr_hashed_p1_f == 8'h4a; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_74; // @[Reg.scala 27:20]
  wire [1:0] _T_23018 = _T_22580 ? bht_bank_rd_data_out_0_74 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23273 = _T_23272 | _T_23018; // @[Mux.scala 27:72]
  wire  _T_22582 = bht_rd_addr_hashed_p1_f == 8'h4b; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_75; // @[Reg.scala 27:20]
  wire [1:0] _T_23019 = _T_22582 ? bht_bank_rd_data_out_0_75 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23274 = _T_23273 | _T_23019; // @[Mux.scala 27:72]
  wire  _T_22584 = bht_rd_addr_hashed_p1_f == 8'h4c; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_76; // @[Reg.scala 27:20]
  wire [1:0] _T_23020 = _T_22584 ? bht_bank_rd_data_out_0_76 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23275 = _T_23274 | _T_23020; // @[Mux.scala 27:72]
  wire  _T_22586 = bht_rd_addr_hashed_p1_f == 8'h4d; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_77; // @[Reg.scala 27:20]
  wire [1:0] _T_23021 = _T_22586 ? bht_bank_rd_data_out_0_77 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23276 = _T_23275 | _T_23021; // @[Mux.scala 27:72]
  wire  _T_22588 = bht_rd_addr_hashed_p1_f == 8'h4e; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_78; // @[Reg.scala 27:20]
  wire [1:0] _T_23022 = _T_22588 ? bht_bank_rd_data_out_0_78 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23277 = _T_23276 | _T_23022; // @[Mux.scala 27:72]
  wire  _T_22590 = bht_rd_addr_hashed_p1_f == 8'h4f; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_79; // @[Reg.scala 27:20]
  wire [1:0] _T_23023 = _T_22590 ? bht_bank_rd_data_out_0_79 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23278 = _T_23277 | _T_23023; // @[Mux.scala 27:72]
  wire  _T_22592 = bht_rd_addr_hashed_p1_f == 8'h50; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_80; // @[Reg.scala 27:20]
  wire [1:0] _T_23024 = _T_22592 ? bht_bank_rd_data_out_0_80 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23279 = _T_23278 | _T_23024; // @[Mux.scala 27:72]
  wire  _T_22594 = bht_rd_addr_hashed_p1_f == 8'h51; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_81; // @[Reg.scala 27:20]
  wire [1:0] _T_23025 = _T_22594 ? bht_bank_rd_data_out_0_81 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23280 = _T_23279 | _T_23025; // @[Mux.scala 27:72]
  wire  _T_22596 = bht_rd_addr_hashed_p1_f == 8'h52; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_82; // @[Reg.scala 27:20]
  wire [1:0] _T_23026 = _T_22596 ? bht_bank_rd_data_out_0_82 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23281 = _T_23280 | _T_23026; // @[Mux.scala 27:72]
  wire  _T_22598 = bht_rd_addr_hashed_p1_f == 8'h53; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_83; // @[Reg.scala 27:20]
  wire [1:0] _T_23027 = _T_22598 ? bht_bank_rd_data_out_0_83 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23282 = _T_23281 | _T_23027; // @[Mux.scala 27:72]
  wire  _T_22600 = bht_rd_addr_hashed_p1_f == 8'h54; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_84; // @[Reg.scala 27:20]
  wire [1:0] _T_23028 = _T_22600 ? bht_bank_rd_data_out_0_84 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23283 = _T_23282 | _T_23028; // @[Mux.scala 27:72]
  wire  _T_22602 = bht_rd_addr_hashed_p1_f == 8'h55; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_85; // @[Reg.scala 27:20]
  wire [1:0] _T_23029 = _T_22602 ? bht_bank_rd_data_out_0_85 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23284 = _T_23283 | _T_23029; // @[Mux.scala 27:72]
  wire  _T_22604 = bht_rd_addr_hashed_p1_f == 8'h56; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_86; // @[Reg.scala 27:20]
  wire [1:0] _T_23030 = _T_22604 ? bht_bank_rd_data_out_0_86 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23285 = _T_23284 | _T_23030; // @[Mux.scala 27:72]
  wire  _T_22606 = bht_rd_addr_hashed_p1_f == 8'h57; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_87; // @[Reg.scala 27:20]
  wire [1:0] _T_23031 = _T_22606 ? bht_bank_rd_data_out_0_87 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23286 = _T_23285 | _T_23031; // @[Mux.scala 27:72]
  wire  _T_22608 = bht_rd_addr_hashed_p1_f == 8'h58; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_88; // @[Reg.scala 27:20]
  wire [1:0] _T_23032 = _T_22608 ? bht_bank_rd_data_out_0_88 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23287 = _T_23286 | _T_23032; // @[Mux.scala 27:72]
  wire  _T_22610 = bht_rd_addr_hashed_p1_f == 8'h59; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_89; // @[Reg.scala 27:20]
  wire [1:0] _T_23033 = _T_22610 ? bht_bank_rd_data_out_0_89 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23288 = _T_23287 | _T_23033; // @[Mux.scala 27:72]
  wire  _T_22612 = bht_rd_addr_hashed_p1_f == 8'h5a; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_90; // @[Reg.scala 27:20]
  wire [1:0] _T_23034 = _T_22612 ? bht_bank_rd_data_out_0_90 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23289 = _T_23288 | _T_23034; // @[Mux.scala 27:72]
  wire  _T_22614 = bht_rd_addr_hashed_p1_f == 8'h5b; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_91; // @[Reg.scala 27:20]
  wire [1:0] _T_23035 = _T_22614 ? bht_bank_rd_data_out_0_91 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23290 = _T_23289 | _T_23035; // @[Mux.scala 27:72]
  wire  _T_22616 = bht_rd_addr_hashed_p1_f == 8'h5c; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_92; // @[Reg.scala 27:20]
  wire [1:0] _T_23036 = _T_22616 ? bht_bank_rd_data_out_0_92 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23291 = _T_23290 | _T_23036; // @[Mux.scala 27:72]
  wire  _T_22618 = bht_rd_addr_hashed_p1_f == 8'h5d; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_93; // @[Reg.scala 27:20]
  wire [1:0] _T_23037 = _T_22618 ? bht_bank_rd_data_out_0_93 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23292 = _T_23291 | _T_23037; // @[Mux.scala 27:72]
  wire  _T_22620 = bht_rd_addr_hashed_p1_f == 8'h5e; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_94; // @[Reg.scala 27:20]
  wire [1:0] _T_23038 = _T_22620 ? bht_bank_rd_data_out_0_94 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23293 = _T_23292 | _T_23038; // @[Mux.scala 27:72]
  wire  _T_22622 = bht_rd_addr_hashed_p1_f == 8'h5f; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_95; // @[Reg.scala 27:20]
  wire [1:0] _T_23039 = _T_22622 ? bht_bank_rd_data_out_0_95 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23294 = _T_23293 | _T_23039; // @[Mux.scala 27:72]
  wire  _T_22624 = bht_rd_addr_hashed_p1_f == 8'h60; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_96; // @[Reg.scala 27:20]
  wire [1:0] _T_23040 = _T_22624 ? bht_bank_rd_data_out_0_96 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23295 = _T_23294 | _T_23040; // @[Mux.scala 27:72]
  wire  _T_22626 = bht_rd_addr_hashed_p1_f == 8'h61; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_97; // @[Reg.scala 27:20]
  wire [1:0] _T_23041 = _T_22626 ? bht_bank_rd_data_out_0_97 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23296 = _T_23295 | _T_23041; // @[Mux.scala 27:72]
  wire  _T_22628 = bht_rd_addr_hashed_p1_f == 8'h62; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_98; // @[Reg.scala 27:20]
  wire [1:0] _T_23042 = _T_22628 ? bht_bank_rd_data_out_0_98 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23297 = _T_23296 | _T_23042; // @[Mux.scala 27:72]
  wire  _T_22630 = bht_rd_addr_hashed_p1_f == 8'h63; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_99; // @[Reg.scala 27:20]
  wire [1:0] _T_23043 = _T_22630 ? bht_bank_rd_data_out_0_99 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23298 = _T_23297 | _T_23043; // @[Mux.scala 27:72]
  wire  _T_22632 = bht_rd_addr_hashed_p1_f == 8'h64; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_100; // @[Reg.scala 27:20]
  wire [1:0] _T_23044 = _T_22632 ? bht_bank_rd_data_out_0_100 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23299 = _T_23298 | _T_23044; // @[Mux.scala 27:72]
  wire  _T_22634 = bht_rd_addr_hashed_p1_f == 8'h65; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_101; // @[Reg.scala 27:20]
  wire [1:0] _T_23045 = _T_22634 ? bht_bank_rd_data_out_0_101 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23300 = _T_23299 | _T_23045; // @[Mux.scala 27:72]
  wire  _T_22636 = bht_rd_addr_hashed_p1_f == 8'h66; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_102; // @[Reg.scala 27:20]
  wire [1:0] _T_23046 = _T_22636 ? bht_bank_rd_data_out_0_102 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23301 = _T_23300 | _T_23046; // @[Mux.scala 27:72]
  wire  _T_22638 = bht_rd_addr_hashed_p1_f == 8'h67; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_103; // @[Reg.scala 27:20]
  wire [1:0] _T_23047 = _T_22638 ? bht_bank_rd_data_out_0_103 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23302 = _T_23301 | _T_23047; // @[Mux.scala 27:72]
  wire  _T_22640 = bht_rd_addr_hashed_p1_f == 8'h68; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_104; // @[Reg.scala 27:20]
  wire [1:0] _T_23048 = _T_22640 ? bht_bank_rd_data_out_0_104 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23303 = _T_23302 | _T_23048; // @[Mux.scala 27:72]
  wire  _T_22642 = bht_rd_addr_hashed_p1_f == 8'h69; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_105; // @[Reg.scala 27:20]
  wire [1:0] _T_23049 = _T_22642 ? bht_bank_rd_data_out_0_105 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23304 = _T_23303 | _T_23049; // @[Mux.scala 27:72]
  wire  _T_22644 = bht_rd_addr_hashed_p1_f == 8'h6a; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_106; // @[Reg.scala 27:20]
  wire [1:0] _T_23050 = _T_22644 ? bht_bank_rd_data_out_0_106 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23305 = _T_23304 | _T_23050; // @[Mux.scala 27:72]
  wire  _T_22646 = bht_rd_addr_hashed_p1_f == 8'h6b; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_107; // @[Reg.scala 27:20]
  wire [1:0] _T_23051 = _T_22646 ? bht_bank_rd_data_out_0_107 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23306 = _T_23305 | _T_23051; // @[Mux.scala 27:72]
  wire  _T_22648 = bht_rd_addr_hashed_p1_f == 8'h6c; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_108; // @[Reg.scala 27:20]
  wire [1:0] _T_23052 = _T_22648 ? bht_bank_rd_data_out_0_108 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23307 = _T_23306 | _T_23052; // @[Mux.scala 27:72]
  wire  _T_22650 = bht_rd_addr_hashed_p1_f == 8'h6d; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_109; // @[Reg.scala 27:20]
  wire [1:0] _T_23053 = _T_22650 ? bht_bank_rd_data_out_0_109 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23308 = _T_23307 | _T_23053; // @[Mux.scala 27:72]
  wire  _T_22652 = bht_rd_addr_hashed_p1_f == 8'h6e; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_110; // @[Reg.scala 27:20]
  wire [1:0] _T_23054 = _T_22652 ? bht_bank_rd_data_out_0_110 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23309 = _T_23308 | _T_23054; // @[Mux.scala 27:72]
  wire  _T_22654 = bht_rd_addr_hashed_p1_f == 8'h6f; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_111; // @[Reg.scala 27:20]
  wire [1:0] _T_23055 = _T_22654 ? bht_bank_rd_data_out_0_111 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23310 = _T_23309 | _T_23055; // @[Mux.scala 27:72]
  wire  _T_22656 = bht_rd_addr_hashed_p1_f == 8'h70; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_112; // @[Reg.scala 27:20]
  wire [1:0] _T_23056 = _T_22656 ? bht_bank_rd_data_out_0_112 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23311 = _T_23310 | _T_23056; // @[Mux.scala 27:72]
  wire  _T_22658 = bht_rd_addr_hashed_p1_f == 8'h71; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_113; // @[Reg.scala 27:20]
  wire [1:0] _T_23057 = _T_22658 ? bht_bank_rd_data_out_0_113 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23312 = _T_23311 | _T_23057; // @[Mux.scala 27:72]
  wire  _T_22660 = bht_rd_addr_hashed_p1_f == 8'h72; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_114; // @[Reg.scala 27:20]
  wire [1:0] _T_23058 = _T_22660 ? bht_bank_rd_data_out_0_114 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23313 = _T_23312 | _T_23058; // @[Mux.scala 27:72]
  wire  _T_22662 = bht_rd_addr_hashed_p1_f == 8'h73; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_115; // @[Reg.scala 27:20]
  wire [1:0] _T_23059 = _T_22662 ? bht_bank_rd_data_out_0_115 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23314 = _T_23313 | _T_23059; // @[Mux.scala 27:72]
  wire  _T_22664 = bht_rd_addr_hashed_p1_f == 8'h74; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_116; // @[Reg.scala 27:20]
  wire [1:0] _T_23060 = _T_22664 ? bht_bank_rd_data_out_0_116 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23315 = _T_23314 | _T_23060; // @[Mux.scala 27:72]
  wire  _T_22666 = bht_rd_addr_hashed_p1_f == 8'h75; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_117; // @[Reg.scala 27:20]
  wire [1:0] _T_23061 = _T_22666 ? bht_bank_rd_data_out_0_117 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23316 = _T_23315 | _T_23061; // @[Mux.scala 27:72]
  wire  _T_22668 = bht_rd_addr_hashed_p1_f == 8'h76; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_118; // @[Reg.scala 27:20]
  wire [1:0] _T_23062 = _T_22668 ? bht_bank_rd_data_out_0_118 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23317 = _T_23316 | _T_23062; // @[Mux.scala 27:72]
  wire  _T_22670 = bht_rd_addr_hashed_p1_f == 8'h77; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_119; // @[Reg.scala 27:20]
  wire [1:0] _T_23063 = _T_22670 ? bht_bank_rd_data_out_0_119 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23318 = _T_23317 | _T_23063; // @[Mux.scala 27:72]
  wire  _T_22672 = bht_rd_addr_hashed_p1_f == 8'h78; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_120; // @[Reg.scala 27:20]
  wire [1:0] _T_23064 = _T_22672 ? bht_bank_rd_data_out_0_120 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23319 = _T_23318 | _T_23064; // @[Mux.scala 27:72]
  wire  _T_22674 = bht_rd_addr_hashed_p1_f == 8'h79; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_121; // @[Reg.scala 27:20]
  wire [1:0] _T_23065 = _T_22674 ? bht_bank_rd_data_out_0_121 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23320 = _T_23319 | _T_23065; // @[Mux.scala 27:72]
  wire  _T_22676 = bht_rd_addr_hashed_p1_f == 8'h7a; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_122; // @[Reg.scala 27:20]
  wire [1:0] _T_23066 = _T_22676 ? bht_bank_rd_data_out_0_122 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23321 = _T_23320 | _T_23066; // @[Mux.scala 27:72]
  wire  _T_22678 = bht_rd_addr_hashed_p1_f == 8'h7b; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_123; // @[Reg.scala 27:20]
  wire [1:0] _T_23067 = _T_22678 ? bht_bank_rd_data_out_0_123 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23322 = _T_23321 | _T_23067; // @[Mux.scala 27:72]
  wire  _T_22680 = bht_rd_addr_hashed_p1_f == 8'h7c; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_124; // @[Reg.scala 27:20]
  wire [1:0] _T_23068 = _T_22680 ? bht_bank_rd_data_out_0_124 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23323 = _T_23322 | _T_23068; // @[Mux.scala 27:72]
  wire  _T_22682 = bht_rd_addr_hashed_p1_f == 8'h7d; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_125; // @[Reg.scala 27:20]
  wire [1:0] _T_23069 = _T_22682 ? bht_bank_rd_data_out_0_125 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23324 = _T_23323 | _T_23069; // @[Mux.scala 27:72]
  wire  _T_22684 = bht_rd_addr_hashed_p1_f == 8'h7e; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_126; // @[Reg.scala 27:20]
  wire [1:0] _T_23070 = _T_22684 ? bht_bank_rd_data_out_0_126 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23325 = _T_23324 | _T_23070; // @[Mux.scala 27:72]
  wire  _T_22686 = bht_rd_addr_hashed_p1_f == 8'h7f; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_127; // @[Reg.scala 27:20]
  wire [1:0] _T_23071 = _T_22686 ? bht_bank_rd_data_out_0_127 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23326 = _T_23325 | _T_23071; // @[Mux.scala 27:72]
  wire  _T_22688 = bht_rd_addr_hashed_p1_f == 8'h80; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_128; // @[Reg.scala 27:20]
  wire [1:0] _T_23072 = _T_22688 ? bht_bank_rd_data_out_0_128 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23327 = _T_23326 | _T_23072; // @[Mux.scala 27:72]
  wire  _T_22690 = bht_rd_addr_hashed_p1_f == 8'h81; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_129; // @[Reg.scala 27:20]
  wire [1:0] _T_23073 = _T_22690 ? bht_bank_rd_data_out_0_129 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23328 = _T_23327 | _T_23073; // @[Mux.scala 27:72]
  wire  _T_22692 = bht_rd_addr_hashed_p1_f == 8'h82; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_130; // @[Reg.scala 27:20]
  wire [1:0] _T_23074 = _T_22692 ? bht_bank_rd_data_out_0_130 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23329 = _T_23328 | _T_23074; // @[Mux.scala 27:72]
  wire  _T_22694 = bht_rd_addr_hashed_p1_f == 8'h83; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_131; // @[Reg.scala 27:20]
  wire [1:0] _T_23075 = _T_22694 ? bht_bank_rd_data_out_0_131 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23330 = _T_23329 | _T_23075; // @[Mux.scala 27:72]
  wire  _T_22696 = bht_rd_addr_hashed_p1_f == 8'h84; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_132; // @[Reg.scala 27:20]
  wire [1:0] _T_23076 = _T_22696 ? bht_bank_rd_data_out_0_132 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23331 = _T_23330 | _T_23076; // @[Mux.scala 27:72]
  wire  _T_22698 = bht_rd_addr_hashed_p1_f == 8'h85; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_133; // @[Reg.scala 27:20]
  wire [1:0] _T_23077 = _T_22698 ? bht_bank_rd_data_out_0_133 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23332 = _T_23331 | _T_23077; // @[Mux.scala 27:72]
  wire  _T_22700 = bht_rd_addr_hashed_p1_f == 8'h86; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_134; // @[Reg.scala 27:20]
  wire [1:0] _T_23078 = _T_22700 ? bht_bank_rd_data_out_0_134 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23333 = _T_23332 | _T_23078; // @[Mux.scala 27:72]
  wire  _T_22702 = bht_rd_addr_hashed_p1_f == 8'h87; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_135; // @[Reg.scala 27:20]
  wire [1:0] _T_23079 = _T_22702 ? bht_bank_rd_data_out_0_135 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23334 = _T_23333 | _T_23079; // @[Mux.scala 27:72]
  wire  _T_22704 = bht_rd_addr_hashed_p1_f == 8'h88; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_136; // @[Reg.scala 27:20]
  wire [1:0] _T_23080 = _T_22704 ? bht_bank_rd_data_out_0_136 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23335 = _T_23334 | _T_23080; // @[Mux.scala 27:72]
  wire  _T_22706 = bht_rd_addr_hashed_p1_f == 8'h89; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_137; // @[Reg.scala 27:20]
  wire [1:0] _T_23081 = _T_22706 ? bht_bank_rd_data_out_0_137 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23336 = _T_23335 | _T_23081; // @[Mux.scala 27:72]
  wire  _T_22708 = bht_rd_addr_hashed_p1_f == 8'h8a; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_138; // @[Reg.scala 27:20]
  wire [1:0] _T_23082 = _T_22708 ? bht_bank_rd_data_out_0_138 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23337 = _T_23336 | _T_23082; // @[Mux.scala 27:72]
  wire  _T_22710 = bht_rd_addr_hashed_p1_f == 8'h8b; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_139; // @[Reg.scala 27:20]
  wire [1:0] _T_23083 = _T_22710 ? bht_bank_rd_data_out_0_139 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23338 = _T_23337 | _T_23083; // @[Mux.scala 27:72]
  wire  _T_22712 = bht_rd_addr_hashed_p1_f == 8'h8c; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_140; // @[Reg.scala 27:20]
  wire [1:0] _T_23084 = _T_22712 ? bht_bank_rd_data_out_0_140 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23339 = _T_23338 | _T_23084; // @[Mux.scala 27:72]
  wire  _T_22714 = bht_rd_addr_hashed_p1_f == 8'h8d; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_141; // @[Reg.scala 27:20]
  wire [1:0] _T_23085 = _T_22714 ? bht_bank_rd_data_out_0_141 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23340 = _T_23339 | _T_23085; // @[Mux.scala 27:72]
  wire  _T_22716 = bht_rd_addr_hashed_p1_f == 8'h8e; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_142; // @[Reg.scala 27:20]
  wire [1:0] _T_23086 = _T_22716 ? bht_bank_rd_data_out_0_142 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23341 = _T_23340 | _T_23086; // @[Mux.scala 27:72]
  wire  _T_22718 = bht_rd_addr_hashed_p1_f == 8'h8f; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_143; // @[Reg.scala 27:20]
  wire [1:0] _T_23087 = _T_22718 ? bht_bank_rd_data_out_0_143 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23342 = _T_23341 | _T_23087; // @[Mux.scala 27:72]
  wire  _T_22720 = bht_rd_addr_hashed_p1_f == 8'h90; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_144; // @[Reg.scala 27:20]
  wire [1:0] _T_23088 = _T_22720 ? bht_bank_rd_data_out_0_144 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23343 = _T_23342 | _T_23088; // @[Mux.scala 27:72]
  wire  _T_22722 = bht_rd_addr_hashed_p1_f == 8'h91; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_145; // @[Reg.scala 27:20]
  wire [1:0] _T_23089 = _T_22722 ? bht_bank_rd_data_out_0_145 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23344 = _T_23343 | _T_23089; // @[Mux.scala 27:72]
  wire  _T_22724 = bht_rd_addr_hashed_p1_f == 8'h92; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_146; // @[Reg.scala 27:20]
  wire [1:0] _T_23090 = _T_22724 ? bht_bank_rd_data_out_0_146 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23345 = _T_23344 | _T_23090; // @[Mux.scala 27:72]
  wire  _T_22726 = bht_rd_addr_hashed_p1_f == 8'h93; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_147; // @[Reg.scala 27:20]
  wire [1:0] _T_23091 = _T_22726 ? bht_bank_rd_data_out_0_147 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23346 = _T_23345 | _T_23091; // @[Mux.scala 27:72]
  wire  _T_22728 = bht_rd_addr_hashed_p1_f == 8'h94; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_148; // @[Reg.scala 27:20]
  wire [1:0] _T_23092 = _T_22728 ? bht_bank_rd_data_out_0_148 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23347 = _T_23346 | _T_23092; // @[Mux.scala 27:72]
  wire  _T_22730 = bht_rd_addr_hashed_p1_f == 8'h95; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_149; // @[Reg.scala 27:20]
  wire [1:0] _T_23093 = _T_22730 ? bht_bank_rd_data_out_0_149 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23348 = _T_23347 | _T_23093; // @[Mux.scala 27:72]
  wire  _T_22732 = bht_rd_addr_hashed_p1_f == 8'h96; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_150; // @[Reg.scala 27:20]
  wire [1:0] _T_23094 = _T_22732 ? bht_bank_rd_data_out_0_150 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23349 = _T_23348 | _T_23094; // @[Mux.scala 27:72]
  wire  _T_22734 = bht_rd_addr_hashed_p1_f == 8'h97; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_151; // @[Reg.scala 27:20]
  wire [1:0] _T_23095 = _T_22734 ? bht_bank_rd_data_out_0_151 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23350 = _T_23349 | _T_23095; // @[Mux.scala 27:72]
  wire  _T_22736 = bht_rd_addr_hashed_p1_f == 8'h98; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_152; // @[Reg.scala 27:20]
  wire [1:0] _T_23096 = _T_22736 ? bht_bank_rd_data_out_0_152 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23351 = _T_23350 | _T_23096; // @[Mux.scala 27:72]
  wire  _T_22738 = bht_rd_addr_hashed_p1_f == 8'h99; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_153; // @[Reg.scala 27:20]
  wire [1:0] _T_23097 = _T_22738 ? bht_bank_rd_data_out_0_153 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23352 = _T_23351 | _T_23097; // @[Mux.scala 27:72]
  wire  _T_22740 = bht_rd_addr_hashed_p1_f == 8'h9a; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_154; // @[Reg.scala 27:20]
  wire [1:0] _T_23098 = _T_22740 ? bht_bank_rd_data_out_0_154 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23353 = _T_23352 | _T_23098; // @[Mux.scala 27:72]
  wire  _T_22742 = bht_rd_addr_hashed_p1_f == 8'h9b; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_155; // @[Reg.scala 27:20]
  wire [1:0] _T_23099 = _T_22742 ? bht_bank_rd_data_out_0_155 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23354 = _T_23353 | _T_23099; // @[Mux.scala 27:72]
  wire  _T_22744 = bht_rd_addr_hashed_p1_f == 8'h9c; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_156; // @[Reg.scala 27:20]
  wire [1:0] _T_23100 = _T_22744 ? bht_bank_rd_data_out_0_156 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23355 = _T_23354 | _T_23100; // @[Mux.scala 27:72]
  wire  _T_22746 = bht_rd_addr_hashed_p1_f == 8'h9d; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_157; // @[Reg.scala 27:20]
  wire [1:0] _T_23101 = _T_22746 ? bht_bank_rd_data_out_0_157 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23356 = _T_23355 | _T_23101; // @[Mux.scala 27:72]
  wire  _T_22748 = bht_rd_addr_hashed_p1_f == 8'h9e; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_158; // @[Reg.scala 27:20]
  wire [1:0] _T_23102 = _T_22748 ? bht_bank_rd_data_out_0_158 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23357 = _T_23356 | _T_23102; // @[Mux.scala 27:72]
  wire  _T_22750 = bht_rd_addr_hashed_p1_f == 8'h9f; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_159; // @[Reg.scala 27:20]
  wire [1:0] _T_23103 = _T_22750 ? bht_bank_rd_data_out_0_159 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23358 = _T_23357 | _T_23103; // @[Mux.scala 27:72]
  wire  _T_22752 = bht_rd_addr_hashed_p1_f == 8'ha0; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_160; // @[Reg.scala 27:20]
  wire [1:0] _T_23104 = _T_22752 ? bht_bank_rd_data_out_0_160 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23359 = _T_23358 | _T_23104; // @[Mux.scala 27:72]
  wire  _T_22754 = bht_rd_addr_hashed_p1_f == 8'ha1; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_161; // @[Reg.scala 27:20]
  wire [1:0] _T_23105 = _T_22754 ? bht_bank_rd_data_out_0_161 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23360 = _T_23359 | _T_23105; // @[Mux.scala 27:72]
  wire  _T_22756 = bht_rd_addr_hashed_p1_f == 8'ha2; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_162; // @[Reg.scala 27:20]
  wire [1:0] _T_23106 = _T_22756 ? bht_bank_rd_data_out_0_162 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23361 = _T_23360 | _T_23106; // @[Mux.scala 27:72]
  wire  _T_22758 = bht_rd_addr_hashed_p1_f == 8'ha3; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_163; // @[Reg.scala 27:20]
  wire [1:0] _T_23107 = _T_22758 ? bht_bank_rd_data_out_0_163 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23362 = _T_23361 | _T_23107; // @[Mux.scala 27:72]
  wire  _T_22760 = bht_rd_addr_hashed_p1_f == 8'ha4; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_164; // @[Reg.scala 27:20]
  wire [1:0] _T_23108 = _T_22760 ? bht_bank_rd_data_out_0_164 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23363 = _T_23362 | _T_23108; // @[Mux.scala 27:72]
  wire  _T_22762 = bht_rd_addr_hashed_p1_f == 8'ha5; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_165; // @[Reg.scala 27:20]
  wire [1:0] _T_23109 = _T_22762 ? bht_bank_rd_data_out_0_165 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23364 = _T_23363 | _T_23109; // @[Mux.scala 27:72]
  wire  _T_22764 = bht_rd_addr_hashed_p1_f == 8'ha6; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_166; // @[Reg.scala 27:20]
  wire [1:0] _T_23110 = _T_22764 ? bht_bank_rd_data_out_0_166 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23365 = _T_23364 | _T_23110; // @[Mux.scala 27:72]
  wire  _T_22766 = bht_rd_addr_hashed_p1_f == 8'ha7; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_167; // @[Reg.scala 27:20]
  wire [1:0] _T_23111 = _T_22766 ? bht_bank_rd_data_out_0_167 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23366 = _T_23365 | _T_23111; // @[Mux.scala 27:72]
  wire  _T_22768 = bht_rd_addr_hashed_p1_f == 8'ha8; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_168; // @[Reg.scala 27:20]
  wire [1:0] _T_23112 = _T_22768 ? bht_bank_rd_data_out_0_168 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23367 = _T_23366 | _T_23112; // @[Mux.scala 27:72]
  wire  _T_22770 = bht_rd_addr_hashed_p1_f == 8'ha9; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_169; // @[Reg.scala 27:20]
  wire [1:0] _T_23113 = _T_22770 ? bht_bank_rd_data_out_0_169 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23368 = _T_23367 | _T_23113; // @[Mux.scala 27:72]
  wire  _T_22772 = bht_rd_addr_hashed_p1_f == 8'haa; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_170; // @[Reg.scala 27:20]
  wire [1:0] _T_23114 = _T_22772 ? bht_bank_rd_data_out_0_170 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23369 = _T_23368 | _T_23114; // @[Mux.scala 27:72]
  wire  _T_22774 = bht_rd_addr_hashed_p1_f == 8'hab; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_171; // @[Reg.scala 27:20]
  wire [1:0] _T_23115 = _T_22774 ? bht_bank_rd_data_out_0_171 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23370 = _T_23369 | _T_23115; // @[Mux.scala 27:72]
  wire  _T_22776 = bht_rd_addr_hashed_p1_f == 8'hac; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_172; // @[Reg.scala 27:20]
  wire [1:0] _T_23116 = _T_22776 ? bht_bank_rd_data_out_0_172 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23371 = _T_23370 | _T_23116; // @[Mux.scala 27:72]
  wire  _T_22778 = bht_rd_addr_hashed_p1_f == 8'had; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_173; // @[Reg.scala 27:20]
  wire [1:0] _T_23117 = _T_22778 ? bht_bank_rd_data_out_0_173 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23372 = _T_23371 | _T_23117; // @[Mux.scala 27:72]
  wire  _T_22780 = bht_rd_addr_hashed_p1_f == 8'hae; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_174; // @[Reg.scala 27:20]
  wire [1:0] _T_23118 = _T_22780 ? bht_bank_rd_data_out_0_174 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23373 = _T_23372 | _T_23118; // @[Mux.scala 27:72]
  wire  _T_22782 = bht_rd_addr_hashed_p1_f == 8'haf; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_175; // @[Reg.scala 27:20]
  wire [1:0] _T_23119 = _T_22782 ? bht_bank_rd_data_out_0_175 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23374 = _T_23373 | _T_23119; // @[Mux.scala 27:72]
  wire  _T_22784 = bht_rd_addr_hashed_p1_f == 8'hb0; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_176; // @[Reg.scala 27:20]
  wire [1:0] _T_23120 = _T_22784 ? bht_bank_rd_data_out_0_176 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23375 = _T_23374 | _T_23120; // @[Mux.scala 27:72]
  wire  _T_22786 = bht_rd_addr_hashed_p1_f == 8'hb1; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_177; // @[Reg.scala 27:20]
  wire [1:0] _T_23121 = _T_22786 ? bht_bank_rd_data_out_0_177 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23376 = _T_23375 | _T_23121; // @[Mux.scala 27:72]
  wire  _T_22788 = bht_rd_addr_hashed_p1_f == 8'hb2; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_178; // @[Reg.scala 27:20]
  wire [1:0] _T_23122 = _T_22788 ? bht_bank_rd_data_out_0_178 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23377 = _T_23376 | _T_23122; // @[Mux.scala 27:72]
  wire  _T_22790 = bht_rd_addr_hashed_p1_f == 8'hb3; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_179; // @[Reg.scala 27:20]
  wire [1:0] _T_23123 = _T_22790 ? bht_bank_rd_data_out_0_179 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23378 = _T_23377 | _T_23123; // @[Mux.scala 27:72]
  wire  _T_22792 = bht_rd_addr_hashed_p1_f == 8'hb4; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_180; // @[Reg.scala 27:20]
  wire [1:0] _T_23124 = _T_22792 ? bht_bank_rd_data_out_0_180 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23379 = _T_23378 | _T_23124; // @[Mux.scala 27:72]
  wire  _T_22794 = bht_rd_addr_hashed_p1_f == 8'hb5; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_181; // @[Reg.scala 27:20]
  wire [1:0] _T_23125 = _T_22794 ? bht_bank_rd_data_out_0_181 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23380 = _T_23379 | _T_23125; // @[Mux.scala 27:72]
  wire  _T_22796 = bht_rd_addr_hashed_p1_f == 8'hb6; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_182; // @[Reg.scala 27:20]
  wire [1:0] _T_23126 = _T_22796 ? bht_bank_rd_data_out_0_182 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23381 = _T_23380 | _T_23126; // @[Mux.scala 27:72]
  wire  _T_22798 = bht_rd_addr_hashed_p1_f == 8'hb7; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_183; // @[Reg.scala 27:20]
  wire [1:0] _T_23127 = _T_22798 ? bht_bank_rd_data_out_0_183 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23382 = _T_23381 | _T_23127; // @[Mux.scala 27:72]
  wire  _T_22800 = bht_rd_addr_hashed_p1_f == 8'hb8; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_184; // @[Reg.scala 27:20]
  wire [1:0] _T_23128 = _T_22800 ? bht_bank_rd_data_out_0_184 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23383 = _T_23382 | _T_23128; // @[Mux.scala 27:72]
  wire  _T_22802 = bht_rd_addr_hashed_p1_f == 8'hb9; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_185; // @[Reg.scala 27:20]
  wire [1:0] _T_23129 = _T_22802 ? bht_bank_rd_data_out_0_185 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23384 = _T_23383 | _T_23129; // @[Mux.scala 27:72]
  wire  _T_22804 = bht_rd_addr_hashed_p1_f == 8'hba; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_186; // @[Reg.scala 27:20]
  wire [1:0] _T_23130 = _T_22804 ? bht_bank_rd_data_out_0_186 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23385 = _T_23384 | _T_23130; // @[Mux.scala 27:72]
  wire  _T_22806 = bht_rd_addr_hashed_p1_f == 8'hbb; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_187; // @[Reg.scala 27:20]
  wire [1:0] _T_23131 = _T_22806 ? bht_bank_rd_data_out_0_187 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23386 = _T_23385 | _T_23131; // @[Mux.scala 27:72]
  wire  _T_22808 = bht_rd_addr_hashed_p1_f == 8'hbc; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_188; // @[Reg.scala 27:20]
  wire [1:0] _T_23132 = _T_22808 ? bht_bank_rd_data_out_0_188 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23387 = _T_23386 | _T_23132; // @[Mux.scala 27:72]
  wire  _T_22810 = bht_rd_addr_hashed_p1_f == 8'hbd; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_189; // @[Reg.scala 27:20]
  wire [1:0] _T_23133 = _T_22810 ? bht_bank_rd_data_out_0_189 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23388 = _T_23387 | _T_23133; // @[Mux.scala 27:72]
  wire  _T_22812 = bht_rd_addr_hashed_p1_f == 8'hbe; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_190; // @[Reg.scala 27:20]
  wire [1:0] _T_23134 = _T_22812 ? bht_bank_rd_data_out_0_190 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23389 = _T_23388 | _T_23134; // @[Mux.scala 27:72]
  wire  _T_22814 = bht_rd_addr_hashed_p1_f == 8'hbf; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_191; // @[Reg.scala 27:20]
  wire [1:0] _T_23135 = _T_22814 ? bht_bank_rd_data_out_0_191 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23390 = _T_23389 | _T_23135; // @[Mux.scala 27:72]
  wire  _T_22816 = bht_rd_addr_hashed_p1_f == 8'hc0; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_192; // @[Reg.scala 27:20]
  wire [1:0] _T_23136 = _T_22816 ? bht_bank_rd_data_out_0_192 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23391 = _T_23390 | _T_23136; // @[Mux.scala 27:72]
  wire  _T_22818 = bht_rd_addr_hashed_p1_f == 8'hc1; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_193; // @[Reg.scala 27:20]
  wire [1:0] _T_23137 = _T_22818 ? bht_bank_rd_data_out_0_193 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23392 = _T_23391 | _T_23137; // @[Mux.scala 27:72]
  wire  _T_22820 = bht_rd_addr_hashed_p1_f == 8'hc2; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_194; // @[Reg.scala 27:20]
  wire [1:0] _T_23138 = _T_22820 ? bht_bank_rd_data_out_0_194 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23393 = _T_23392 | _T_23138; // @[Mux.scala 27:72]
  wire  _T_22822 = bht_rd_addr_hashed_p1_f == 8'hc3; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_195; // @[Reg.scala 27:20]
  wire [1:0] _T_23139 = _T_22822 ? bht_bank_rd_data_out_0_195 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23394 = _T_23393 | _T_23139; // @[Mux.scala 27:72]
  wire  _T_22824 = bht_rd_addr_hashed_p1_f == 8'hc4; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_196; // @[Reg.scala 27:20]
  wire [1:0] _T_23140 = _T_22824 ? bht_bank_rd_data_out_0_196 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23395 = _T_23394 | _T_23140; // @[Mux.scala 27:72]
  wire  _T_22826 = bht_rd_addr_hashed_p1_f == 8'hc5; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_197; // @[Reg.scala 27:20]
  wire [1:0] _T_23141 = _T_22826 ? bht_bank_rd_data_out_0_197 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23396 = _T_23395 | _T_23141; // @[Mux.scala 27:72]
  wire  _T_22828 = bht_rd_addr_hashed_p1_f == 8'hc6; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_198; // @[Reg.scala 27:20]
  wire [1:0] _T_23142 = _T_22828 ? bht_bank_rd_data_out_0_198 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23397 = _T_23396 | _T_23142; // @[Mux.scala 27:72]
  wire  _T_22830 = bht_rd_addr_hashed_p1_f == 8'hc7; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_199; // @[Reg.scala 27:20]
  wire [1:0] _T_23143 = _T_22830 ? bht_bank_rd_data_out_0_199 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23398 = _T_23397 | _T_23143; // @[Mux.scala 27:72]
  wire  _T_22832 = bht_rd_addr_hashed_p1_f == 8'hc8; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_200; // @[Reg.scala 27:20]
  wire [1:0] _T_23144 = _T_22832 ? bht_bank_rd_data_out_0_200 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23399 = _T_23398 | _T_23144; // @[Mux.scala 27:72]
  wire  _T_22834 = bht_rd_addr_hashed_p1_f == 8'hc9; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_201; // @[Reg.scala 27:20]
  wire [1:0] _T_23145 = _T_22834 ? bht_bank_rd_data_out_0_201 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23400 = _T_23399 | _T_23145; // @[Mux.scala 27:72]
  wire  _T_22836 = bht_rd_addr_hashed_p1_f == 8'hca; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_202; // @[Reg.scala 27:20]
  wire [1:0] _T_23146 = _T_22836 ? bht_bank_rd_data_out_0_202 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23401 = _T_23400 | _T_23146; // @[Mux.scala 27:72]
  wire  _T_22838 = bht_rd_addr_hashed_p1_f == 8'hcb; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_203; // @[Reg.scala 27:20]
  wire [1:0] _T_23147 = _T_22838 ? bht_bank_rd_data_out_0_203 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23402 = _T_23401 | _T_23147; // @[Mux.scala 27:72]
  wire  _T_22840 = bht_rd_addr_hashed_p1_f == 8'hcc; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_204; // @[Reg.scala 27:20]
  wire [1:0] _T_23148 = _T_22840 ? bht_bank_rd_data_out_0_204 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23403 = _T_23402 | _T_23148; // @[Mux.scala 27:72]
  wire  _T_22842 = bht_rd_addr_hashed_p1_f == 8'hcd; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_205; // @[Reg.scala 27:20]
  wire [1:0] _T_23149 = _T_22842 ? bht_bank_rd_data_out_0_205 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23404 = _T_23403 | _T_23149; // @[Mux.scala 27:72]
  wire  _T_22844 = bht_rd_addr_hashed_p1_f == 8'hce; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_206; // @[Reg.scala 27:20]
  wire [1:0] _T_23150 = _T_22844 ? bht_bank_rd_data_out_0_206 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23405 = _T_23404 | _T_23150; // @[Mux.scala 27:72]
  wire  _T_22846 = bht_rd_addr_hashed_p1_f == 8'hcf; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_207; // @[Reg.scala 27:20]
  wire [1:0] _T_23151 = _T_22846 ? bht_bank_rd_data_out_0_207 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23406 = _T_23405 | _T_23151; // @[Mux.scala 27:72]
  wire  _T_22848 = bht_rd_addr_hashed_p1_f == 8'hd0; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_208; // @[Reg.scala 27:20]
  wire [1:0] _T_23152 = _T_22848 ? bht_bank_rd_data_out_0_208 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23407 = _T_23406 | _T_23152; // @[Mux.scala 27:72]
  wire  _T_22850 = bht_rd_addr_hashed_p1_f == 8'hd1; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_209; // @[Reg.scala 27:20]
  wire [1:0] _T_23153 = _T_22850 ? bht_bank_rd_data_out_0_209 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23408 = _T_23407 | _T_23153; // @[Mux.scala 27:72]
  wire  _T_22852 = bht_rd_addr_hashed_p1_f == 8'hd2; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_210; // @[Reg.scala 27:20]
  wire [1:0] _T_23154 = _T_22852 ? bht_bank_rd_data_out_0_210 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23409 = _T_23408 | _T_23154; // @[Mux.scala 27:72]
  wire  _T_22854 = bht_rd_addr_hashed_p1_f == 8'hd3; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_211; // @[Reg.scala 27:20]
  wire [1:0] _T_23155 = _T_22854 ? bht_bank_rd_data_out_0_211 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23410 = _T_23409 | _T_23155; // @[Mux.scala 27:72]
  wire  _T_22856 = bht_rd_addr_hashed_p1_f == 8'hd4; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_212; // @[Reg.scala 27:20]
  wire [1:0] _T_23156 = _T_22856 ? bht_bank_rd_data_out_0_212 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23411 = _T_23410 | _T_23156; // @[Mux.scala 27:72]
  wire  _T_22858 = bht_rd_addr_hashed_p1_f == 8'hd5; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_213; // @[Reg.scala 27:20]
  wire [1:0] _T_23157 = _T_22858 ? bht_bank_rd_data_out_0_213 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23412 = _T_23411 | _T_23157; // @[Mux.scala 27:72]
  wire  _T_22860 = bht_rd_addr_hashed_p1_f == 8'hd6; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_214; // @[Reg.scala 27:20]
  wire [1:0] _T_23158 = _T_22860 ? bht_bank_rd_data_out_0_214 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23413 = _T_23412 | _T_23158; // @[Mux.scala 27:72]
  wire  _T_22862 = bht_rd_addr_hashed_p1_f == 8'hd7; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_215; // @[Reg.scala 27:20]
  wire [1:0] _T_23159 = _T_22862 ? bht_bank_rd_data_out_0_215 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23414 = _T_23413 | _T_23159; // @[Mux.scala 27:72]
  wire  _T_22864 = bht_rd_addr_hashed_p1_f == 8'hd8; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_216; // @[Reg.scala 27:20]
  wire [1:0] _T_23160 = _T_22864 ? bht_bank_rd_data_out_0_216 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23415 = _T_23414 | _T_23160; // @[Mux.scala 27:72]
  wire  _T_22866 = bht_rd_addr_hashed_p1_f == 8'hd9; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_217; // @[Reg.scala 27:20]
  wire [1:0] _T_23161 = _T_22866 ? bht_bank_rd_data_out_0_217 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23416 = _T_23415 | _T_23161; // @[Mux.scala 27:72]
  wire  _T_22868 = bht_rd_addr_hashed_p1_f == 8'hda; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_218; // @[Reg.scala 27:20]
  wire [1:0] _T_23162 = _T_22868 ? bht_bank_rd_data_out_0_218 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23417 = _T_23416 | _T_23162; // @[Mux.scala 27:72]
  wire  _T_22870 = bht_rd_addr_hashed_p1_f == 8'hdb; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_219; // @[Reg.scala 27:20]
  wire [1:0] _T_23163 = _T_22870 ? bht_bank_rd_data_out_0_219 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23418 = _T_23417 | _T_23163; // @[Mux.scala 27:72]
  wire  _T_22872 = bht_rd_addr_hashed_p1_f == 8'hdc; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_220; // @[Reg.scala 27:20]
  wire [1:0] _T_23164 = _T_22872 ? bht_bank_rd_data_out_0_220 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23419 = _T_23418 | _T_23164; // @[Mux.scala 27:72]
  wire  _T_22874 = bht_rd_addr_hashed_p1_f == 8'hdd; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_221; // @[Reg.scala 27:20]
  wire [1:0] _T_23165 = _T_22874 ? bht_bank_rd_data_out_0_221 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23420 = _T_23419 | _T_23165; // @[Mux.scala 27:72]
  wire  _T_22876 = bht_rd_addr_hashed_p1_f == 8'hde; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_222; // @[Reg.scala 27:20]
  wire [1:0] _T_23166 = _T_22876 ? bht_bank_rd_data_out_0_222 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23421 = _T_23420 | _T_23166; // @[Mux.scala 27:72]
  wire  _T_22878 = bht_rd_addr_hashed_p1_f == 8'hdf; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_223; // @[Reg.scala 27:20]
  wire [1:0] _T_23167 = _T_22878 ? bht_bank_rd_data_out_0_223 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23422 = _T_23421 | _T_23167; // @[Mux.scala 27:72]
  wire  _T_22880 = bht_rd_addr_hashed_p1_f == 8'he0; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_224; // @[Reg.scala 27:20]
  wire [1:0] _T_23168 = _T_22880 ? bht_bank_rd_data_out_0_224 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23423 = _T_23422 | _T_23168; // @[Mux.scala 27:72]
  wire  _T_22882 = bht_rd_addr_hashed_p1_f == 8'he1; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_225; // @[Reg.scala 27:20]
  wire [1:0] _T_23169 = _T_22882 ? bht_bank_rd_data_out_0_225 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23424 = _T_23423 | _T_23169; // @[Mux.scala 27:72]
  wire  _T_22884 = bht_rd_addr_hashed_p1_f == 8'he2; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_226; // @[Reg.scala 27:20]
  wire [1:0] _T_23170 = _T_22884 ? bht_bank_rd_data_out_0_226 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23425 = _T_23424 | _T_23170; // @[Mux.scala 27:72]
  wire  _T_22886 = bht_rd_addr_hashed_p1_f == 8'he3; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_227; // @[Reg.scala 27:20]
  wire [1:0] _T_23171 = _T_22886 ? bht_bank_rd_data_out_0_227 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23426 = _T_23425 | _T_23171; // @[Mux.scala 27:72]
  wire  _T_22888 = bht_rd_addr_hashed_p1_f == 8'he4; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_228; // @[Reg.scala 27:20]
  wire [1:0] _T_23172 = _T_22888 ? bht_bank_rd_data_out_0_228 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23427 = _T_23426 | _T_23172; // @[Mux.scala 27:72]
  wire  _T_22890 = bht_rd_addr_hashed_p1_f == 8'he5; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_229; // @[Reg.scala 27:20]
  wire [1:0] _T_23173 = _T_22890 ? bht_bank_rd_data_out_0_229 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23428 = _T_23427 | _T_23173; // @[Mux.scala 27:72]
  wire  _T_22892 = bht_rd_addr_hashed_p1_f == 8'he6; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_230; // @[Reg.scala 27:20]
  wire [1:0] _T_23174 = _T_22892 ? bht_bank_rd_data_out_0_230 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23429 = _T_23428 | _T_23174; // @[Mux.scala 27:72]
  wire  _T_22894 = bht_rd_addr_hashed_p1_f == 8'he7; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_231; // @[Reg.scala 27:20]
  wire [1:0] _T_23175 = _T_22894 ? bht_bank_rd_data_out_0_231 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23430 = _T_23429 | _T_23175; // @[Mux.scala 27:72]
  wire  _T_22896 = bht_rd_addr_hashed_p1_f == 8'he8; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_232; // @[Reg.scala 27:20]
  wire [1:0] _T_23176 = _T_22896 ? bht_bank_rd_data_out_0_232 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23431 = _T_23430 | _T_23176; // @[Mux.scala 27:72]
  wire  _T_22898 = bht_rd_addr_hashed_p1_f == 8'he9; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_233; // @[Reg.scala 27:20]
  wire [1:0] _T_23177 = _T_22898 ? bht_bank_rd_data_out_0_233 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23432 = _T_23431 | _T_23177; // @[Mux.scala 27:72]
  wire  _T_22900 = bht_rd_addr_hashed_p1_f == 8'hea; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_234; // @[Reg.scala 27:20]
  wire [1:0] _T_23178 = _T_22900 ? bht_bank_rd_data_out_0_234 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23433 = _T_23432 | _T_23178; // @[Mux.scala 27:72]
  wire  _T_22902 = bht_rd_addr_hashed_p1_f == 8'heb; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_235; // @[Reg.scala 27:20]
  wire [1:0] _T_23179 = _T_22902 ? bht_bank_rd_data_out_0_235 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23434 = _T_23433 | _T_23179; // @[Mux.scala 27:72]
  wire  _T_22904 = bht_rd_addr_hashed_p1_f == 8'hec; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_236; // @[Reg.scala 27:20]
  wire [1:0] _T_23180 = _T_22904 ? bht_bank_rd_data_out_0_236 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23435 = _T_23434 | _T_23180; // @[Mux.scala 27:72]
  wire  _T_22906 = bht_rd_addr_hashed_p1_f == 8'hed; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_237; // @[Reg.scala 27:20]
  wire [1:0] _T_23181 = _T_22906 ? bht_bank_rd_data_out_0_237 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23436 = _T_23435 | _T_23181; // @[Mux.scala 27:72]
  wire  _T_22908 = bht_rd_addr_hashed_p1_f == 8'hee; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_238; // @[Reg.scala 27:20]
  wire [1:0] _T_23182 = _T_22908 ? bht_bank_rd_data_out_0_238 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23437 = _T_23436 | _T_23182; // @[Mux.scala 27:72]
  wire  _T_22910 = bht_rd_addr_hashed_p1_f == 8'hef; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_239; // @[Reg.scala 27:20]
  wire [1:0] _T_23183 = _T_22910 ? bht_bank_rd_data_out_0_239 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23438 = _T_23437 | _T_23183; // @[Mux.scala 27:72]
  wire  _T_22912 = bht_rd_addr_hashed_p1_f == 8'hf0; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_240; // @[Reg.scala 27:20]
  wire [1:0] _T_23184 = _T_22912 ? bht_bank_rd_data_out_0_240 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23439 = _T_23438 | _T_23184; // @[Mux.scala 27:72]
  wire  _T_22914 = bht_rd_addr_hashed_p1_f == 8'hf1; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_241; // @[Reg.scala 27:20]
  wire [1:0] _T_23185 = _T_22914 ? bht_bank_rd_data_out_0_241 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23440 = _T_23439 | _T_23185; // @[Mux.scala 27:72]
  wire  _T_22916 = bht_rd_addr_hashed_p1_f == 8'hf2; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_242; // @[Reg.scala 27:20]
  wire [1:0] _T_23186 = _T_22916 ? bht_bank_rd_data_out_0_242 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23441 = _T_23440 | _T_23186; // @[Mux.scala 27:72]
  wire  _T_22918 = bht_rd_addr_hashed_p1_f == 8'hf3; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_243; // @[Reg.scala 27:20]
  wire [1:0] _T_23187 = _T_22918 ? bht_bank_rd_data_out_0_243 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23442 = _T_23441 | _T_23187; // @[Mux.scala 27:72]
  wire  _T_22920 = bht_rd_addr_hashed_p1_f == 8'hf4; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_244; // @[Reg.scala 27:20]
  wire [1:0] _T_23188 = _T_22920 ? bht_bank_rd_data_out_0_244 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23443 = _T_23442 | _T_23188; // @[Mux.scala 27:72]
  wire  _T_22922 = bht_rd_addr_hashed_p1_f == 8'hf5; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_245; // @[Reg.scala 27:20]
  wire [1:0] _T_23189 = _T_22922 ? bht_bank_rd_data_out_0_245 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23444 = _T_23443 | _T_23189; // @[Mux.scala 27:72]
  wire  _T_22924 = bht_rd_addr_hashed_p1_f == 8'hf6; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_246; // @[Reg.scala 27:20]
  wire [1:0] _T_23190 = _T_22924 ? bht_bank_rd_data_out_0_246 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23445 = _T_23444 | _T_23190; // @[Mux.scala 27:72]
  wire  _T_22926 = bht_rd_addr_hashed_p1_f == 8'hf7; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_247; // @[Reg.scala 27:20]
  wire [1:0] _T_23191 = _T_22926 ? bht_bank_rd_data_out_0_247 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23446 = _T_23445 | _T_23191; // @[Mux.scala 27:72]
  wire  _T_22928 = bht_rd_addr_hashed_p1_f == 8'hf8; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_248; // @[Reg.scala 27:20]
  wire [1:0] _T_23192 = _T_22928 ? bht_bank_rd_data_out_0_248 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23447 = _T_23446 | _T_23192; // @[Mux.scala 27:72]
  wire  _T_22930 = bht_rd_addr_hashed_p1_f == 8'hf9; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_249; // @[Reg.scala 27:20]
  wire [1:0] _T_23193 = _T_22930 ? bht_bank_rd_data_out_0_249 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23448 = _T_23447 | _T_23193; // @[Mux.scala 27:72]
  wire  _T_22932 = bht_rd_addr_hashed_p1_f == 8'hfa; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_250; // @[Reg.scala 27:20]
  wire [1:0] _T_23194 = _T_22932 ? bht_bank_rd_data_out_0_250 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23449 = _T_23448 | _T_23194; // @[Mux.scala 27:72]
  wire  _T_22934 = bht_rd_addr_hashed_p1_f == 8'hfb; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_251; // @[Reg.scala 27:20]
  wire [1:0] _T_23195 = _T_22934 ? bht_bank_rd_data_out_0_251 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23450 = _T_23449 | _T_23195; // @[Mux.scala 27:72]
  wire  _T_22936 = bht_rd_addr_hashed_p1_f == 8'hfc; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_252; // @[Reg.scala 27:20]
  wire [1:0] _T_23196 = _T_22936 ? bht_bank_rd_data_out_0_252 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23451 = _T_23450 | _T_23196; // @[Mux.scala 27:72]
  wire  _T_22938 = bht_rd_addr_hashed_p1_f == 8'hfd; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_253; // @[Reg.scala 27:20]
  wire [1:0] _T_23197 = _T_22938 ? bht_bank_rd_data_out_0_253 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23452 = _T_23451 | _T_23197; // @[Mux.scala 27:72]
  wire  _T_22940 = bht_rd_addr_hashed_p1_f == 8'hfe; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_254; // @[Reg.scala 27:20]
  wire [1:0] _T_23198 = _T_22940 ? bht_bank_rd_data_out_0_254 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23453 = _T_23452 | _T_23198; // @[Mux.scala 27:72]
  wire  _T_22942 = bht_rd_addr_hashed_p1_f == 8'hff; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_255; // @[Reg.scala 27:20]
  wire [1:0] _T_23199 = _T_22942 ? bht_bank_rd_data_out_0_255 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] bht_bank0_rd_data_p1_f = _T_23453 | _T_23199; // @[Mux.scala 27:72]
  wire [1:0] _T_261 = io_ifc_fetch_addr_f[0] ? bht_bank0_rd_data_p1_f : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] bht_vbank1_rd_data_f = _T_260 | _T_261; // @[Mux.scala 27:72]
  wire  _T_265 = bht_force_taken_f[1] | bht_vbank1_rd_data_f[1]; // @[ifu_bp_ctl.scala 281:42]
  wire [1:0] wayhit_f = tag_match_way0_expanded_f | tag_match_way1_expanded_f; // @[ifu_bp_ctl.scala 155:44]
  wire [1:0] _T_159 = _T_144 ? wayhit_f : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] wayhit_p1_f = tag_match_way0_expanded_p1_f | tag_match_way1_expanded_p1_f; // @[ifu_bp_ctl.scala 157:50]
  wire [1:0] _T_158 = {wayhit_p1_f[0],wayhit_f[1]}; // @[Cat.scala 29:58]
  wire [1:0] _T_160 = io_ifc_fetch_addr_f[0] ? _T_158 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_161 = _T_159 | _T_160; // @[Mux.scala 27:72]
  wire  eoc_near = &io_ifc_fetch_addr_f[4:2]; // @[ifu_bp_ctl.scala 241:64]
  wire  _T_219 = ~eoc_near; // @[ifu_bp_ctl.scala 244:15]
  wire [1:0] _T_221 = ~io_ifc_fetch_addr_f[1:0]; // @[ifu_bp_ctl.scala 244:28]
  wire  _T_222 = |_T_221; // @[ifu_bp_ctl.scala 244:58]
  wire  eoc_mask = _T_219 | _T_222; // @[ifu_bp_ctl.scala 244:25]
  wire [1:0] _T_163 = {eoc_mask,1'h1}; // @[Cat.scala 29:58]
  wire [1:0] bht_valid_f = _T_161 & _T_163; // @[ifu_bp_ctl.scala 203:71]
  wire  _T_267 = _T_265 & bht_valid_f[1]; // @[ifu_bp_ctl.scala 281:69]
  wire [1:0] _T_20896 = _T_21408 ? bht_bank_rd_data_out_0_0 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20897 = _T_21410 ? bht_bank_rd_data_out_0_1 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21152 = _T_20896 | _T_20897; // @[Mux.scala 27:72]
  wire [1:0] _T_20898 = _T_21412 ? bht_bank_rd_data_out_0_2 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21153 = _T_21152 | _T_20898; // @[Mux.scala 27:72]
  wire [1:0] _T_20899 = _T_21414 ? bht_bank_rd_data_out_0_3 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21154 = _T_21153 | _T_20899; // @[Mux.scala 27:72]
  wire [1:0] _T_20900 = _T_21416 ? bht_bank_rd_data_out_0_4 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21155 = _T_21154 | _T_20900; // @[Mux.scala 27:72]
  wire [1:0] _T_20901 = _T_21418 ? bht_bank_rd_data_out_0_5 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21156 = _T_21155 | _T_20901; // @[Mux.scala 27:72]
  wire [1:0] _T_20902 = _T_21420 ? bht_bank_rd_data_out_0_6 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21157 = _T_21156 | _T_20902; // @[Mux.scala 27:72]
  wire [1:0] _T_20903 = _T_21422 ? bht_bank_rd_data_out_0_7 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21158 = _T_21157 | _T_20903; // @[Mux.scala 27:72]
  wire [1:0] _T_20904 = _T_21424 ? bht_bank_rd_data_out_0_8 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21159 = _T_21158 | _T_20904; // @[Mux.scala 27:72]
  wire [1:0] _T_20905 = _T_21426 ? bht_bank_rd_data_out_0_9 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21160 = _T_21159 | _T_20905; // @[Mux.scala 27:72]
  wire [1:0] _T_20906 = _T_21428 ? bht_bank_rd_data_out_0_10 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21161 = _T_21160 | _T_20906; // @[Mux.scala 27:72]
  wire [1:0] _T_20907 = _T_21430 ? bht_bank_rd_data_out_0_11 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21162 = _T_21161 | _T_20907; // @[Mux.scala 27:72]
  wire [1:0] _T_20908 = _T_21432 ? bht_bank_rd_data_out_0_12 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21163 = _T_21162 | _T_20908; // @[Mux.scala 27:72]
  wire [1:0] _T_20909 = _T_21434 ? bht_bank_rd_data_out_0_13 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21164 = _T_21163 | _T_20909; // @[Mux.scala 27:72]
  wire [1:0] _T_20910 = _T_21436 ? bht_bank_rd_data_out_0_14 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21165 = _T_21164 | _T_20910; // @[Mux.scala 27:72]
  wire [1:0] _T_20911 = _T_21438 ? bht_bank_rd_data_out_0_15 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21166 = _T_21165 | _T_20911; // @[Mux.scala 27:72]
  wire [1:0] _T_20912 = _T_21440 ? bht_bank_rd_data_out_0_16 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21167 = _T_21166 | _T_20912; // @[Mux.scala 27:72]
  wire [1:0] _T_20913 = _T_21442 ? bht_bank_rd_data_out_0_17 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21168 = _T_21167 | _T_20913; // @[Mux.scala 27:72]
  wire [1:0] _T_20914 = _T_21444 ? bht_bank_rd_data_out_0_18 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21169 = _T_21168 | _T_20914; // @[Mux.scala 27:72]
  wire [1:0] _T_20915 = _T_21446 ? bht_bank_rd_data_out_0_19 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21170 = _T_21169 | _T_20915; // @[Mux.scala 27:72]
  wire [1:0] _T_20916 = _T_21448 ? bht_bank_rd_data_out_0_20 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21171 = _T_21170 | _T_20916; // @[Mux.scala 27:72]
  wire [1:0] _T_20917 = _T_21450 ? bht_bank_rd_data_out_0_21 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21172 = _T_21171 | _T_20917; // @[Mux.scala 27:72]
  wire [1:0] _T_20918 = _T_21452 ? bht_bank_rd_data_out_0_22 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21173 = _T_21172 | _T_20918; // @[Mux.scala 27:72]
  wire [1:0] _T_20919 = _T_21454 ? bht_bank_rd_data_out_0_23 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21174 = _T_21173 | _T_20919; // @[Mux.scala 27:72]
  wire [1:0] _T_20920 = _T_21456 ? bht_bank_rd_data_out_0_24 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21175 = _T_21174 | _T_20920; // @[Mux.scala 27:72]
  wire [1:0] _T_20921 = _T_21458 ? bht_bank_rd_data_out_0_25 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21176 = _T_21175 | _T_20921; // @[Mux.scala 27:72]
  wire [1:0] _T_20922 = _T_21460 ? bht_bank_rd_data_out_0_26 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21177 = _T_21176 | _T_20922; // @[Mux.scala 27:72]
  wire [1:0] _T_20923 = _T_21462 ? bht_bank_rd_data_out_0_27 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21178 = _T_21177 | _T_20923; // @[Mux.scala 27:72]
  wire [1:0] _T_20924 = _T_21464 ? bht_bank_rd_data_out_0_28 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21179 = _T_21178 | _T_20924; // @[Mux.scala 27:72]
  wire [1:0] _T_20925 = _T_21466 ? bht_bank_rd_data_out_0_29 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21180 = _T_21179 | _T_20925; // @[Mux.scala 27:72]
  wire [1:0] _T_20926 = _T_21468 ? bht_bank_rd_data_out_0_30 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21181 = _T_21180 | _T_20926; // @[Mux.scala 27:72]
  wire [1:0] _T_20927 = _T_21470 ? bht_bank_rd_data_out_0_31 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21182 = _T_21181 | _T_20927; // @[Mux.scala 27:72]
  wire [1:0] _T_20928 = _T_21472 ? bht_bank_rd_data_out_0_32 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21183 = _T_21182 | _T_20928; // @[Mux.scala 27:72]
  wire [1:0] _T_20929 = _T_21474 ? bht_bank_rd_data_out_0_33 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21184 = _T_21183 | _T_20929; // @[Mux.scala 27:72]
  wire [1:0] _T_20930 = _T_21476 ? bht_bank_rd_data_out_0_34 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21185 = _T_21184 | _T_20930; // @[Mux.scala 27:72]
  wire [1:0] _T_20931 = _T_21478 ? bht_bank_rd_data_out_0_35 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21186 = _T_21185 | _T_20931; // @[Mux.scala 27:72]
  wire [1:0] _T_20932 = _T_21480 ? bht_bank_rd_data_out_0_36 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21187 = _T_21186 | _T_20932; // @[Mux.scala 27:72]
  wire [1:0] _T_20933 = _T_21482 ? bht_bank_rd_data_out_0_37 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21188 = _T_21187 | _T_20933; // @[Mux.scala 27:72]
  wire [1:0] _T_20934 = _T_21484 ? bht_bank_rd_data_out_0_38 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21189 = _T_21188 | _T_20934; // @[Mux.scala 27:72]
  wire [1:0] _T_20935 = _T_21486 ? bht_bank_rd_data_out_0_39 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21190 = _T_21189 | _T_20935; // @[Mux.scala 27:72]
  wire [1:0] _T_20936 = _T_21488 ? bht_bank_rd_data_out_0_40 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21191 = _T_21190 | _T_20936; // @[Mux.scala 27:72]
  wire [1:0] _T_20937 = _T_21490 ? bht_bank_rd_data_out_0_41 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21192 = _T_21191 | _T_20937; // @[Mux.scala 27:72]
  wire [1:0] _T_20938 = _T_21492 ? bht_bank_rd_data_out_0_42 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21193 = _T_21192 | _T_20938; // @[Mux.scala 27:72]
  wire [1:0] _T_20939 = _T_21494 ? bht_bank_rd_data_out_0_43 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21194 = _T_21193 | _T_20939; // @[Mux.scala 27:72]
  wire [1:0] _T_20940 = _T_21496 ? bht_bank_rd_data_out_0_44 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21195 = _T_21194 | _T_20940; // @[Mux.scala 27:72]
  wire [1:0] _T_20941 = _T_21498 ? bht_bank_rd_data_out_0_45 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21196 = _T_21195 | _T_20941; // @[Mux.scala 27:72]
  wire [1:0] _T_20942 = _T_21500 ? bht_bank_rd_data_out_0_46 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21197 = _T_21196 | _T_20942; // @[Mux.scala 27:72]
  wire [1:0] _T_20943 = _T_21502 ? bht_bank_rd_data_out_0_47 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21198 = _T_21197 | _T_20943; // @[Mux.scala 27:72]
  wire [1:0] _T_20944 = _T_21504 ? bht_bank_rd_data_out_0_48 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21199 = _T_21198 | _T_20944; // @[Mux.scala 27:72]
  wire [1:0] _T_20945 = _T_21506 ? bht_bank_rd_data_out_0_49 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21200 = _T_21199 | _T_20945; // @[Mux.scala 27:72]
  wire [1:0] _T_20946 = _T_21508 ? bht_bank_rd_data_out_0_50 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21201 = _T_21200 | _T_20946; // @[Mux.scala 27:72]
  wire [1:0] _T_20947 = _T_21510 ? bht_bank_rd_data_out_0_51 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21202 = _T_21201 | _T_20947; // @[Mux.scala 27:72]
  wire [1:0] _T_20948 = _T_21512 ? bht_bank_rd_data_out_0_52 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21203 = _T_21202 | _T_20948; // @[Mux.scala 27:72]
  wire [1:0] _T_20949 = _T_21514 ? bht_bank_rd_data_out_0_53 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21204 = _T_21203 | _T_20949; // @[Mux.scala 27:72]
  wire [1:0] _T_20950 = _T_21516 ? bht_bank_rd_data_out_0_54 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21205 = _T_21204 | _T_20950; // @[Mux.scala 27:72]
  wire [1:0] _T_20951 = _T_21518 ? bht_bank_rd_data_out_0_55 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21206 = _T_21205 | _T_20951; // @[Mux.scala 27:72]
  wire [1:0] _T_20952 = _T_21520 ? bht_bank_rd_data_out_0_56 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21207 = _T_21206 | _T_20952; // @[Mux.scala 27:72]
  wire [1:0] _T_20953 = _T_21522 ? bht_bank_rd_data_out_0_57 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21208 = _T_21207 | _T_20953; // @[Mux.scala 27:72]
  wire [1:0] _T_20954 = _T_21524 ? bht_bank_rd_data_out_0_58 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21209 = _T_21208 | _T_20954; // @[Mux.scala 27:72]
  wire [1:0] _T_20955 = _T_21526 ? bht_bank_rd_data_out_0_59 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21210 = _T_21209 | _T_20955; // @[Mux.scala 27:72]
  wire [1:0] _T_20956 = _T_21528 ? bht_bank_rd_data_out_0_60 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21211 = _T_21210 | _T_20956; // @[Mux.scala 27:72]
  wire [1:0] _T_20957 = _T_21530 ? bht_bank_rd_data_out_0_61 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21212 = _T_21211 | _T_20957; // @[Mux.scala 27:72]
  wire [1:0] _T_20958 = _T_21532 ? bht_bank_rd_data_out_0_62 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21213 = _T_21212 | _T_20958; // @[Mux.scala 27:72]
  wire [1:0] _T_20959 = _T_21534 ? bht_bank_rd_data_out_0_63 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21214 = _T_21213 | _T_20959; // @[Mux.scala 27:72]
  wire [1:0] _T_20960 = _T_21536 ? bht_bank_rd_data_out_0_64 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21215 = _T_21214 | _T_20960; // @[Mux.scala 27:72]
  wire [1:0] _T_20961 = _T_21538 ? bht_bank_rd_data_out_0_65 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21216 = _T_21215 | _T_20961; // @[Mux.scala 27:72]
  wire [1:0] _T_20962 = _T_21540 ? bht_bank_rd_data_out_0_66 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21217 = _T_21216 | _T_20962; // @[Mux.scala 27:72]
  wire [1:0] _T_20963 = _T_21542 ? bht_bank_rd_data_out_0_67 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21218 = _T_21217 | _T_20963; // @[Mux.scala 27:72]
  wire [1:0] _T_20964 = _T_21544 ? bht_bank_rd_data_out_0_68 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21219 = _T_21218 | _T_20964; // @[Mux.scala 27:72]
  wire [1:0] _T_20965 = _T_21546 ? bht_bank_rd_data_out_0_69 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21220 = _T_21219 | _T_20965; // @[Mux.scala 27:72]
  wire [1:0] _T_20966 = _T_21548 ? bht_bank_rd_data_out_0_70 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21221 = _T_21220 | _T_20966; // @[Mux.scala 27:72]
  wire [1:0] _T_20967 = _T_21550 ? bht_bank_rd_data_out_0_71 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21222 = _T_21221 | _T_20967; // @[Mux.scala 27:72]
  wire [1:0] _T_20968 = _T_21552 ? bht_bank_rd_data_out_0_72 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21223 = _T_21222 | _T_20968; // @[Mux.scala 27:72]
  wire [1:0] _T_20969 = _T_21554 ? bht_bank_rd_data_out_0_73 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21224 = _T_21223 | _T_20969; // @[Mux.scala 27:72]
  wire [1:0] _T_20970 = _T_21556 ? bht_bank_rd_data_out_0_74 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21225 = _T_21224 | _T_20970; // @[Mux.scala 27:72]
  wire [1:0] _T_20971 = _T_21558 ? bht_bank_rd_data_out_0_75 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21226 = _T_21225 | _T_20971; // @[Mux.scala 27:72]
  wire [1:0] _T_20972 = _T_21560 ? bht_bank_rd_data_out_0_76 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21227 = _T_21226 | _T_20972; // @[Mux.scala 27:72]
  wire [1:0] _T_20973 = _T_21562 ? bht_bank_rd_data_out_0_77 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21228 = _T_21227 | _T_20973; // @[Mux.scala 27:72]
  wire [1:0] _T_20974 = _T_21564 ? bht_bank_rd_data_out_0_78 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21229 = _T_21228 | _T_20974; // @[Mux.scala 27:72]
  wire [1:0] _T_20975 = _T_21566 ? bht_bank_rd_data_out_0_79 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21230 = _T_21229 | _T_20975; // @[Mux.scala 27:72]
  wire [1:0] _T_20976 = _T_21568 ? bht_bank_rd_data_out_0_80 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21231 = _T_21230 | _T_20976; // @[Mux.scala 27:72]
  wire [1:0] _T_20977 = _T_21570 ? bht_bank_rd_data_out_0_81 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21232 = _T_21231 | _T_20977; // @[Mux.scala 27:72]
  wire [1:0] _T_20978 = _T_21572 ? bht_bank_rd_data_out_0_82 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21233 = _T_21232 | _T_20978; // @[Mux.scala 27:72]
  wire [1:0] _T_20979 = _T_21574 ? bht_bank_rd_data_out_0_83 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21234 = _T_21233 | _T_20979; // @[Mux.scala 27:72]
  wire [1:0] _T_20980 = _T_21576 ? bht_bank_rd_data_out_0_84 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21235 = _T_21234 | _T_20980; // @[Mux.scala 27:72]
  wire [1:0] _T_20981 = _T_21578 ? bht_bank_rd_data_out_0_85 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21236 = _T_21235 | _T_20981; // @[Mux.scala 27:72]
  wire [1:0] _T_20982 = _T_21580 ? bht_bank_rd_data_out_0_86 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21237 = _T_21236 | _T_20982; // @[Mux.scala 27:72]
  wire [1:0] _T_20983 = _T_21582 ? bht_bank_rd_data_out_0_87 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21238 = _T_21237 | _T_20983; // @[Mux.scala 27:72]
  wire [1:0] _T_20984 = _T_21584 ? bht_bank_rd_data_out_0_88 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21239 = _T_21238 | _T_20984; // @[Mux.scala 27:72]
  wire [1:0] _T_20985 = _T_21586 ? bht_bank_rd_data_out_0_89 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21240 = _T_21239 | _T_20985; // @[Mux.scala 27:72]
  wire [1:0] _T_20986 = _T_21588 ? bht_bank_rd_data_out_0_90 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21241 = _T_21240 | _T_20986; // @[Mux.scala 27:72]
  wire [1:0] _T_20987 = _T_21590 ? bht_bank_rd_data_out_0_91 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21242 = _T_21241 | _T_20987; // @[Mux.scala 27:72]
  wire [1:0] _T_20988 = _T_21592 ? bht_bank_rd_data_out_0_92 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21243 = _T_21242 | _T_20988; // @[Mux.scala 27:72]
  wire [1:0] _T_20989 = _T_21594 ? bht_bank_rd_data_out_0_93 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21244 = _T_21243 | _T_20989; // @[Mux.scala 27:72]
  wire [1:0] _T_20990 = _T_21596 ? bht_bank_rd_data_out_0_94 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21245 = _T_21244 | _T_20990; // @[Mux.scala 27:72]
  wire [1:0] _T_20991 = _T_21598 ? bht_bank_rd_data_out_0_95 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21246 = _T_21245 | _T_20991; // @[Mux.scala 27:72]
  wire [1:0] _T_20992 = _T_21600 ? bht_bank_rd_data_out_0_96 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21247 = _T_21246 | _T_20992; // @[Mux.scala 27:72]
  wire [1:0] _T_20993 = _T_21602 ? bht_bank_rd_data_out_0_97 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21248 = _T_21247 | _T_20993; // @[Mux.scala 27:72]
  wire [1:0] _T_20994 = _T_21604 ? bht_bank_rd_data_out_0_98 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21249 = _T_21248 | _T_20994; // @[Mux.scala 27:72]
  wire [1:0] _T_20995 = _T_21606 ? bht_bank_rd_data_out_0_99 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21250 = _T_21249 | _T_20995; // @[Mux.scala 27:72]
  wire [1:0] _T_20996 = _T_21608 ? bht_bank_rd_data_out_0_100 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21251 = _T_21250 | _T_20996; // @[Mux.scala 27:72]
  wire [1:0] _T_20997 = _T_21610 ? bht_bank_rd_data_out_0_101 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21252 = _T_21251 | _T_20997; // @[Mux.scala 27:72]
  wire [1:0] _T_20998 = _T_21612 ? bht_bank_rd_data_out_0_102 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21253 = _T_21252 | _T_20998; // @[Mux.scala 27:72]
  wire [1:0] _T_20999 = _T_21614 ? bht_bank_rd_data_out_0_103 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21254 = _T_21253 | _T_20999; // @[Mux.scala 27:72]
  wire [1:0] _T_21000 = _T_21616 ? bht_bank_rd_data_out_0_104 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21255 = _T_21254 | _T_21000; // @[Mux.scala 27:72]
  wire [1:0] _T_21001 = _T_21618 ? bht_bank_rd_data_out_0_105 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21256 = _T_21255 | _T_21001; // @[Mux.scala 27:72]
  wire [1:0] _T_21002 = _T_21620 ? bht_bank_rd_data_out_0_106 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21257 = _T_21256 | _T_21002; // @[Mux.scala 27:72]
  wire [1:0] _T_21003 = _T_21622 ? bht_bank_rd_data_out_0_107 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21258 = _T_21257 | _T_21003; // @[Mux.scala 27:72]
  wire [1:0] _T_21004 = _T_21624 ? bht_bank_rd_data_out_0_108 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21259 = _T_21258 | _T_21004; // @[Mux.scala 27:72]
  wire [1:0] _T_21005 = _T_21626 ? bht_bank_rd_data_out_0_109 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21260 = _T_21259 | _T_21005; // @[Mux.scala 27:72]
  wire [1:0] _T_21006 = _T_21628 ? bht_bank_rd_data_out_0_110 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21261 = _T_21260 | _T_21006; // @[Mux.scala 27:72]
  wire [1:0] _T_21007 = _T_21630 ? bht_bank_rd_data_out_0_111 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21262 = _T_21261 | _T_21007; // @[Mux.scala 27:72]
  wire [1:0] _T_21008 = _T_21632 ? bht_bank_rd_data_out_0_112 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21263 = _T_21262 | _T_21008; // @[Mux.scala 27:72]
  wire [1:0] _T_21009 = _T_21634 ? bht_bank_rd_data_out_0_113 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21264 = _T_21263 | _T_21009; // @[Mux.scala 27:72]
  wire [1:0] _T_21010 = _T_21636 ? bht_bank_rd_data_out_0_114 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21265 = _T_21264 | _T_21010; // @[Mux.scala 27:72]
  wire [1:0] _T_21011 = _T_21638 ? bht_bank_rd_data_out_0_115 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21266 = _T_21265 | _T_21011; // @[Mux.scala 27:72]
  wire [1:0] _T_21012 = _T_21640 ? bht_bank_rd_data_out_0_116 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21267 = _T_21266 | _T_21012; // @[Mux.scala 27:72]
  wire [1:0] _T_21013 = _T_21642 ? bht_bank_rd_data_out_0_117 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21268 = _T_21267 | _T_21013; // @[Mux.scala 27:72]
  wire [1:0] _T_21014 = _T_21644 ? bht_bank_rd_data_out_0_118 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21269 = _T_21268 | _T_21014; // @[Mux.scala 27:72]
  wire [1:0] _T_21015 = _T_21646 ? bht_bank_rd_data_out_0_119 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21270 = _T_21269 | _T_21015; // @[Mux.scala 27:72]
  wire [1:0] _T_21016 = _T_21648 ? bht_bank_rd_data_out_0_120 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21271 = _T_21270 | _T_21016; // @[Mux.scala 27:72]
  wire [1:0] _T_21017 = _T_21650 ? bht_bank_rd_data_out_0_121 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21272 = _T_21271 | _T_21017; // @[Mux.scala 27:72]
  wire [1:0] _T_21018 = _T_21652 ? bht_bank_rd_data_out_0_122 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21273 = _T_21272 | _T_21018; // @[Mux.scala 27:72]
  wire [1:0] _T_21019 = _T_21654 ? bht_bank_rd_data_out_0_123 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21274 = _T_21273 | _T_21019; // @[Mux.scala 27:72]
  wire [1:0] _T_21020 = _T_21656 ? bht_bank_rd_data_out_0_124 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21275 = _T_21274 | _T_21020; // @[Mux.scala 27:72]
  wire [1:0] _T_21021 = _T_21658 ? bht_bank_rd_data_out_0_125 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21276 = _T_21275 | _T_21021; // @[Mux.scala 27:72]
  wire [1:0] _T_21022 = _T_21660 ? bht_bank_rd_data_out_0_126 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21277 = _T_21276 | _T_21022; // @[Mux.scala 27:72]
  wire [1:0] _T_21023 = _T_21662 ? bht_bank_rd_data_out_0_127 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21278 = _T_21277 | _T_21023; // @[Mux.scala 27:72]
  wire [1:0] _T_21024 = _T_21664 ? bht_bank_rd_data_out_0_128 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21279 = _T_21278 | _T_21024; // @[Mux.scala 27:72]
  wire [1:0] _T_21025 = _T_21666 ? bht_bank_rd_data_out_0_129 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21280 = _T_21279 | _T_21025; // @[Mux.scala 27:72]
  wire [1:0] _T_21026 = _T_21668 ? bht_bank_rd_data_out_0_130 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21281 = _T_21280 | _T_21026; // @[Mux.scala 27:72]
  wire [1:0] _T_21027 = _T_21670 ? bht_bank_rd_data_out_0_131 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21282 = _T_21281 | _T_21027; // @[Mux.scala 27:72]
  wire [1:0] _T_21028 = _T_21672 ? bht_bank_rd_data_out_0_132 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21283 = _T_21282 | _T_21028; // @[Mux.scala 27:72]
  wire [1:0] _T_21029 = _T_21674 ? bht_bank_rd_data_out_0_133 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21284 = _T_21283 | _T_21029; // @[Mux.scala 27:72]
  wire [1:0] _T_21030 = _T_21676 ? bht_bank_rd_data_out_0_134 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21285 = _T_21284 | _T_21030; // @[Mux.scala 27:72]
  wire [1:0] _T_21031 = _T_21678 ? bht_bank_rd_data_out_0_135 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21286 = _T_21285 | _T_21031; // @[Mux.scala 27:72]
  wire [1:0] _T_21032 = _T_21680 ? bht_bank_rd_data_out_0_136 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21287 = _T_21286 | _T_21032; // @[Mux.scala 27:72]
  wire [1:0] _T_21033 = _T_21682 ? bht_bank_rd_data_out_0_137 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21288 = _T_21287 | _T_21033; // @[Mux.scala 27:72]
  wire [1:0] _T_21034 = _T_21684 ? bht_bank_rd_data_out_0_138 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21289 = _T_21288 | _T_21034; // @[Mux.scala 27:72]
  wire [1:0] _T_21035 = _T_21686 ? bht_bank_rd_data_out_0_139 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21290 = _T_21289 | _T_21035; // @[Mux.scala 27:72]
  wire [1:0] _T_21036 = _T_21688 ? bht_bank_rd_data_out_0_140 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21291 = _T_21290 | _T_21036; // @[Mux.scala 27:72]
  wire [1:0] _T_21037 = _T_21690 ? bht_bank_rd_data_out_0_141 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21292 = _T_21291 | _T_21037; // @[Mux.scala 27:72]
  wire [1:0] _T_21038 = _T_21692 ? bht_bank_rd_data_out_0_142 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21293 = _T_21292 | _T_21038; // @[Mux.scala 27:72]
  wire [1:0] _T_21039 = _T_21694 ? bht_bank_rd_data_out_0_143 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21294 = _T_21293 | _T_21039; // @[Mux.scala 27:72]
  wire [1:0] _T_21040 = _T_21696 ? bht_bank_rd_data_out_0_144 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21295 = _T_21294 | _T_21040; // @[Mux.scala 27:72]
  wire [1:0] _T_21041 = _T_21698 ? bht_bank_rd_data_out_0_145 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21296 = _T_21295 | _T_21041; // @[Mux.scala 27:72]
  wire [1:0] _T_21042 = _T_21700 ? bht_bank_rd_data_out_0_146 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21297 = _T_21296 | _T_21042; // @[Mux.scala 27:72]
  wire [1:0] _T_21043 = _T_21702 ? bht_bank_rd_data_out_0_147 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21298 = _T_21297 | _T_21043; // @[Mux.scala 27:72]
  wire [1:0] _T_21044 = _T_21704 ? bht_bank_rd_data_out_0_148 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21299 = _T_21298 | _T_21044; // @[Mux.scala 27:72]
  wire [1:0] _T_21045 = _T_21706 ? bht_bank_rd_data_out_0_149 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21300 = _T_21299 | _T_21045; // @[Mux.scala 27:72]
  wire [1:0] _T_21046 = _T_21708 ? bht_bank_rd_data_out_0_150 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21301 = _T_21300 | _T_21046; // @[Mux.scala 27:72]
  wire [1:0] _T_21047 = _T_21710 ? bht_bank_rd_data_out_0_151 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21302 = _T_21301 | _T_21047; // @[Mux.scala 27:72]
  wire [1:0] _T_21048 = _T_21712 ? bht_bank_rd_data_out_0_152 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21303 = _T_21302 | _T_21048; // @[Mux.scala 27:72]
  wire [1:0] _T_21049 = _T_21714 ? bht_bank_rd_data_out_0_153 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21304 = _T_21303 | _T_21049; // @[Mux.scala 27:72]
  wire [1:0] _T_21050 = _T_21716 ? bht_bank_rd_data_out_0_154 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21305 = _T_21304 | _T_21050; // @[Mux.scala 27:72]
  wire [1:0] _T_21051 = _T_21718 ? bht_bank_rd_data_out_0_155 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21306 = _T_21305 | _T_21051; // @[Mux.scala 27:72]
  wire [1:0] _T_21052 = _T_21720 ? bht_bank_rd_data_out_0_156 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21307 = _T_21306 | _T_21052; // @[Mux.scala 27:72]
  wire [1:0] _T_21053 = _T_21722 ? bht_bank_rd_data_out_0_157 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21308 = _T_21307 | _T_21053; // @[Mux.scala 27:72]
  wire [1:0] _T_21054 = _T_21724 ? bht_bank_rd_data_out_0_158 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21309 = _T_21308 | _T_21054; // @[Mux.scala 27:72]
  wire [1:0] _T_21055 = _T_21726 ? bht_bank_rd_data_out_0_159 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21310 = _T_21309 | _T_21055; // @[Mux.scala 27:72]
  wire [1:0] _T_21056 = _T_21728 ? bht_bank_rd_data_out_0_160 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21311 = _T_21310 | _T_21056; // @[Mux.scala 27:72]
  wire [1:0] _T_21057 = _T_21730 ? bht_bank_rd_data_out_0_161 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21312 = _T_21311 | _T_21057; // @[Mux.scala 27:72]
  wire [1:0] _T_21058 = _T_21732 ? bht_bank_rd_data_out_0_162 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21313 = _T_21312 | _T_21058; // @[Mux.scala 27:72]
  wire [1:0] _T_21059 = _T_21734 ? bht_bank_rd_data_out_0_163 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21314 = _T_21313 | _T_21059; // @[Mux.scala 27:72]
  wire [1:0] _T_21060 = _T_21736 ? bht_bank_rd_data_out_0_164 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21315 = _T_21314 | _T_21060; // @[Mux.scala 27:72]
  wire [1:0] _T_21061 = _T_21738 ? bht_bank_rd_data_out_0_165 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21316 = _T_21315 | _T_21061; // @[Mux.scala 27:72]
  wire [1:0] _T_21062 = _T_21740 ? bht_bank_rd_data_out_0_166 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21317 = _T_21316 | _T_21062; // @[Mux.scala 27:72]
  wire [1:0] _T_21063 = _T_21742 ? bht_bank_rd_data_out_0_167 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21318 = _T_21317 | _T_21063; // @[Mux.scala 27:72]
  wire [1:0] _T_21064 = _T_21744 ? bht_bank_rd_data_out_0_168 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21319 = _T_21318 | _T_21064; // @[Mux.scala 27:72]
  wire [1:0] _T_21065 = _T_21746 ? bht_bank_rd_data_out_0_169 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21320 = _T_21319 | _T_21065; // @[Mux.scala 27:72]
  wire [1:0] _T_21066 = _T_21748 ? bht_bank_rd_data_out_0_170 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21321 = _T_21320 | _T_21066; // @[Mux.scala 27:72]
  wire [1:0] _T_21067 = _T_21750 ? bht_bank_rd_data_out_0_171 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21322 = _T_21321 | _T_21067; // @[Mux.scala 27:72]
  wire [1:0] _T_21068 = _T_21752 ? bht_bank_rd_data_out_0_172 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21323 = _T_21322 | _T_21068; // @[Mux.scala 27:72]
  wire [1:0] _T_21069 = _T_21754 ? bht_bank_rd_data_out_0_173 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21324 = _T_21323 | _T_21069; // @[Mux.scala 27:72]
  wire [1:0] _T_21070 = _T_21756 ? bht_bank_rd_data_out_0_174 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21325 = _T_21324 | _T_21070; // @[Mux.scala 27:72]
  wire [1:0] _T_21071 = _T_21758 ? bht_bank_rd_data_out_0_175 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21326 = _T_21325 | _T_21071; // @[Mux.scala 27:72]
  wire [1:0] _T_21072 = _T_21760 ? bht_bank_rd_data_out_0_176 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21327 = _T_21326 | _T_21072; // @[Mux.scala 27:72]
  wire [1:0] _T_21073 = _T_21762 ? bht_bank_rd_data_out_0_177 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21328 = _T_21327 | _T_21073; // @[Mux.scala 27:72]
  wire [1:0] _T_21074 = _T_21764 ? bht_bank_rd_data_out_0_178 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21329 = _T_21328 | _T_21074; // @[Mux.scala 27:72]
  wire [1:0] _T_21075 = _T_21766 ? bht_bank_rd_data_out_0_179 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21330 = _T_21329 | _T_21075; // @[Mux.scala 27:72]
  wire [1:0] _T_21076 = _T_21768 ? bht_bank_rd_data_out_0_180 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21331 = _T_21330 | _T_21076; // @[Mux.scala 27:72]
  wire [1:0] _T_21077 = _T_21770 ? bht_bank_rd_data_out_0_181 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21332 = _T_21331 | _T_21077; // @[Mux.scala 27:72]
  wire [1:0] _T_21078 = _T_21772 ? bht_bank_rd_data_out_0_182 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21333 = _T_21332 | _T_21078; // @[Mux.scala 27:72]
  wire [1:0] _T_21079 = _T_21774 ? bht_bank_rd_data_out_0_183 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21334 = _T_21333 | _T_21079; // @[Mux.scala 27:72]
  wire [1:0] _T_21080 = _T_21776 ? bht_bank_rd_data_out_0_184 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21335 = _T_21334 | _T_21080; // @[Mux.scala 27:72]
  wire [1:0] _T_21081 = _T_21778 ? bht_bank_rd_data_out_0_185 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21336 = _T_21335 | _T_21081; // @[Mux.scala 27:72]
  wire [1:0] _T_21082 = _T_21780 ? bht_bank_rd_data_out_0_186 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21337 = _T_21336 | _T_21082; // @[Mux.scala 27:72]
  wire [1:0] _T_21083 = _T_21782 ? bht_bank_rd_data_out_0_187 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21338 = _T_21337 | _T_21083; // @[Mux.scala 27:72]
  wire [1:0] _T_21084 = _T_21784 ? bht_bank_rd_data_out_0_188 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21339 = _T_21338 | _T_21084; // @[Mux.scala 27:72]
  wire [1:0] _T_21085 = _T_21786 ? bht_bank_rd_data_out_0_189 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21340 = _T_21339 | _T_21085; // @[Mux.scala 27:72]
  wire [1:0] _T_21086 = _T_21788 ? bht_bank_rd_data_out_0_190 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21341 = _T_21340 | _T_21086; // @[Mux.scala 27:72]
  wire [1:0] _T_21087 = _T_21790 ? bht_bank_rd_data_out_0_191 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21342 = _T_21341 | _T_21087; // @[Mux.scala 27:72]
  wire [1:0] _T_21088 = _T_21792 ? bht_bank_rd_data_out_0_192 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21343 = _T_21342 | _T_21088; // @[Mux.scala 27:72]
  wire [1:0] _T_21089 = _T_21794 ? bht_bank_rd_data_out_0_193 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21344 = _T_21343 | _T_21089; // @[Mux.scala 27:72]
  wire [1:0] _T_21090 = _T_21796 ? bht_bank_rd_data_out_0_194 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21345 = _T_21344 | _T_21090; // @[Mux.scala 27:72]
  wire [1:0] _T_21091 = _T_21798 ? bht_bank_rd_data_out_0_195 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21346 = _T_21345 | _T_21091; // @[Mux.scala 27:72]
  wire [1:0] _T_21092 = _T_21800 ? bht_bank_rd_data_out_0_196 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21347 = _T_21346 | _T_21092; // @[Mux.scala 27:72]
  wire [1:0] _T_21093 = _T_21802 ? bht_bank_rd_data_out_0_197 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21348 = _T_21347 | _T_21093; // @[Mux.scala 27:72]
  wire [1:0] _T_21094 = _T_21804 ? bht_bank_rd_data_out_0_198 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21349 = _T_21348 | _T_21094; // @[Mux.scala 27:72]
  wire [1:0] _T_21095 = _T_21806 ? bht_bank_rd_data_out_0_199 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21350 = _T_21349 | _T_21095; // @[Mux.scala 27:72]
  wire [1:0] _T_21096 = _T_21808 ? bht_bank_rd_data_out_0_200 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21351 = _T_21350 | _T_21096; // @[Mux.scala 27:72]
  wire [1:0] _T_21097 = _T_21810 ? bht_bank_rd_data_out_0_201 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21352 = _T_21351 | _T_21097; // @[Mux.scala 27:72]
  wire [1:0] _T_21098 = _T_21812 ? bht_bank_rd_data_out_0_202 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21353 = _T_21352 | _T_21098; // @[Mux.scala 27:72]
  wire [1:0] _T_21099 = _T_21814 ? bht_bank_rd_data_out_0_203 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21354 = _T_21353 | _T_21099; // @[Mux.scala 27:72]
  wire [1:0] _T_21100 = _T_21816 ? bht_bank_rd_data_out_0_204 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21355 = _T_21354 | _T_21100; // @[Mux.scala 27:72]
  wire [1:0] _T_21101 = _T_21818 ? bht_bank_rd_data_out_0_205 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21356 = _T_21355 | _T_21101; // @[Mux.scala 27:72]
  wire [1:0] _T_21102 = _T_21820 ? bht_bank_rd_data_out_0_206 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21357 = _T_21356 | _T_21102; // @[Mux.scala 27:72]
  wire [1:0] _T_21103 = _T_21822 ? bht_bank_rd_data_out_0_207 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21358 = _T_21357 | _T_21103; // @[Mux.scala 27:72]
  wire [1:0] _T_21104 = _T_21824 ? bht_bank_rd_data_out_0_208 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21359 = _T_21358 | _T_21104; // @[Mux.scala 27:72]
  wire [1:0] _T_21105 = _T_21826 ? bht_bank_rd_data_out_0_209 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21360 = _T_21359 | _T_21105; // @[Mux.scala 27:72]
  wire [1:0] _T_21106 = _T_21828 ? bht_bank_rd_data_out_0_210 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21361 = _T_21360 | _T_21106; // @[Mux.scala 27:72]
  wire [1:0] _T_21107 = _T_21830 ? bht_bank_rd_data_out_0_211 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21362 = _T_21361 | _T_21107; // @[Mux.scala 27:72]
  wire [1:0] _T_21108 = _T_21832 ? bht_bank_rd_data_out_0_212 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21363 = _T_21362 | _T_21108; // @[Mux.scala 27:72]
  wire [1:0] _T_21109 = _T_21834 ? bht_bank_rd_data_out_0_213 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21364 = _T_21363 | _T_21109; // @[Mux.scala 27:72]
  wire [1:0] _T_21110 = _T_21836 ? bht_bank_rd_data_out_0_214 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21365 = _T_21364 | _T_21110; // @[Mux.scala 27:72]
  wire [1:0] _T_21111 = _T_21838 ? bht_bank_rd_data_out_0_215 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21366 = _T_21365 | _T_21111; // @[Mux.scala 27:72]
  wire [1:0] _T_21112 = _T_21840 ? bht_bank_rd_data_out_0_216 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21367 = _T_21366 | _T_21112; // @[Mux.scala 27:72]
  wire [1:0] _T_21113 = _T_21842 ? bht_bank_rd_data_out_0_217 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21368 = _T_21367 | _T_21113; // @[Mux.scala 27:72]
  wire [1:0] _T_21114 = _T_21844 ? bht_bank_rd_data_out_0_218 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21369 = _T_21368 | _T_21114; // @[Mux.scala 27:72]
  wire [1:0] _T_21115 = _T_21846 ? bht_bank_rd_data_out_0_219 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21370 = _T_21369 | _T_21115; // @[Mux.scala 27:72]
  wire [1:0] _T_21116 = _T_21848 ? bht_bank_rd_data_out_0_220 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21371 = _T_21370 | _T_21116; // @[Mux.scala 27:72]
  wire [1:0] _T_21117 = _T_21850 ? bht_bank_rd_data_out_0_221 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21372 = _T_21371 | _T_21117; // @[Mux.scala 27:72]
  wire [1:0] _T_21118 = _T_21852 ? bht_bank_rd_data_out_0_222 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21373 = _T_21372 | _T_21118; // @[Mux.scala 27:72]
  wire [1:0] _T_21119 = _T_21854 ? bht_bank_rd_data_out_0_223 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21374 = _T_21373 | _T_21119; // @[Mux.scala 27:72]
  wire [1:0] _T_21120 = _T_21856 ? bht_bank_rd_data_out_0_224 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21375 = _T_21374 | _T_21120; // @[Mux.scala 27:72]
  wire [1:0] _T_21121 = _T_21858 ? bht_bank_rd_data_out_0_225 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21376 = _T_21375 | _T_21121; // @[Mux.scala 27:72]
  wire [1:0] _T_21122 = _T_21860 ? bht_bank_rd_data_out_0_226 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21377 = _T_21376 | _T_21122; // @[Mux.scala 27:72]
  wire [1:0] _T_21123 = _T_21862 ? bht_bank_rd_data_out_0_227 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21378 = _T_21377 | _T_21123; // @[Mux.scala 27:72]
  wire [1:0] _T_21124 = _T_21864 ? bht_bank_rd_data_out_0_228 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21379 = _T_21378 | _T_21124; // @[Mux.scala 27:72]
  wire [1:0] _T_21125 = _T_21866 ? bht_bank_rd_data_out_0_229 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21380 = _T_21379 | _T_21125; // @[Mux.scala 27:72]
  wire [1:0] _T_21126 = _T_21868 ? bht_bank_rd_data_out_0_230 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21381 = _T_21380 | _T_21126; // @[Mux.scala 27:72]
  wire [1:0] _T_21127 = _T_21870 ? bht_bank_rd_data_out_0_231 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21382 = _T_21381 | _T_21127; // @[Mux.scala 27:72]
  wire [1:0] _T_21128 = _T_21872 ? bht_bank_rd_data_out_0_232 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21383 = _T_21382 | _T_21128; // @[Mux.scala 27:72]
  wire [1:0] _T_21129 = _T_21874 ? bht_bank_rd_data_out_0_233 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21384 = _T_21383 | _T_21129; // @[Mux.scala 27:72]
  wire [1:0] _T_21130 = _T_21876 ? bht_bank_rd_data_out_0_234 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21385 = _T_21384 | _T_21130; // @[Mux.scala 27:72]
  wire [1:0] _T_21131 = _T_21878 ? bht_bank_rd_data_out_0_235 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21386 = _T_21385 | _T_21131; // @[Mux.scala 27:72]
  wire [1:0] _T_21132 = _T_21880 ? bht_bank_rd_data_out_0_236 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21387 = _T_21386 | _T_21132; // @[Mux.scala 27:72]
  wire [1:0] _T_21133 = _T_21882 ? bht_bank_rd_data_out_0_237 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21388 = _T_21387 | _T_21133; // @[Mux.scala 27:72]
  wire [1:0] _T_21134 = _T_21884 ? bht_bank_rd_data_out_0_238 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21389 = _T_21388 | _T_21134; // @[Mux.scala 27:72]
  wire [1:0] _T_21135 = _T_21886 ? bht_bank_rd_data_out_0_239 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21390 = _T_21389 | _T_21135; // @[Mux.scala 27:72]
  wire [1:0] _T_21136 = _T_21888 ? bht_bank_rd_data_out_0_240 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21391 = _T_21390 | _T_21136; // @[Mux.scala 27:72]
  wire [1:0] _T_21137 = _T_21890 ? bht_bank_rd_data_out_0_241 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21392 = _T_21391 | _T_21137; // @[Mux.scala 27:72]
  wire [1:0] _T_21138 = _T_21892 ? bht_bank_rd_data_out_0_242 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21393 = _T_21392 | _T_21138; // @[Mux.scala 27:72]
  wire [1:0] _T_21139 = _T_21894 ? bht_bank_rd_data_out_0_243 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21394 = _T_21393 | _T_21139; // @[Mux.scala 27:72]
  wire [1:0] _T_21140 = _T_21896 ? bht_bank_rd_data_out_0_244 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21395 = _T_21394 | _T_21140; // @[Mux.scala 27:72]
  wire [1:0] _T_21141 = _T_21898 ? bht_bank_rd_data_out_0_245 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21396 = _T_21395 | _T_21141; // @[Mux.scala 27:72]
  wire [1:0] _T_21142 = _T_21900 ? bht_bank_rd_data_out_0_246 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21397 = _T_21396 | _T_21142; // @[Mux.scala 27:72]
  wire [1:0] _T_21143 = _T_21902 ? bht_bank_rd_data_out_0_247 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21398 = _T_21397 | _T_21143; // @[Mux.scala 27:72]
  wire [1:0] _T_21144 = _T_21904 ? bht_bank_rd_data_out_0_248 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21399 = _T_21398 | _T_21144; // @[Mux.scala 27:72]
  wire [1:0] _T_21145 = _T_21906 ? bht_bank_rd_data_out_0_249 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21400 = _T_21399 | _T_21145; // @[Mux.scala 27:72]
  wire [1:0] _T_21146 = _T_21908 ? bht_bank_rd_data_out_0_250 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21401 = _T_21400 | _T_21146; // @[Mux.scala 27:72]
  wire [1:0] _T_21147 = _T_21910 ? bht_bank_rd_data_out_0_251 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21402 = _T_21401 | _T_21147; // @[Mux.scala 27:72]
  wire [1:0] _T_21148 = _T_21912 ? bht_bank_rd_data_out_0_252 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21403 = _T_21402 | _T_21148; // @[Mux.scala 27:72]
  wire [1:0] _T_21149 = _T_21914 ? bht_bank_rd_data_out_0_253 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21404 = _T_21403 | _T_21149; // @[Mux.scala 27:72]
  wire [1:0] _T_21150 = _T_21916 ? bht_bank_rd_data_out_0_254 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21405 = _T_21404 | _T_21150; // @[Mux.scala 27:72]
  wire [1:0] _T_21151 = _T_21918 ? bht_bank_rd_data_out_0_255 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] bht_bank0_rd_data_f = _T_21405 | _T_21151; // @[Mux.scala 27:72]
  wire [1:0] _T_252 = _T_144 ? bht_bank0_rd_data_f : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_253 = io_ifc_fetch_addr_f[0] ? bht_bank1_rd_data_f : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] bht_vbank0_rd_data_f = _T_252 | _T_253; // @[Mux.scala 27:72]
  wire  _T_270 = bht_force_taken_f[0] | bht_vbank0_rd_data_f[1]; // @[ifu_bp_ctl.scala 282:45]
  wire  _T_272 = _T_270 & bht_valid_f[0]; // @[ifu_bp_ctl.scala 282:72]
  wire [1:0] bht_dir_f = {_T_267,_T_272}; // @[Cat.scala 29:58]
  wire  _T_14 = ~bht_dir_f[0]; // @[ifu_bp_ctl.scala 96:23]
  wire [1:0] btb_sel_f = {_T_14,bht_dir_f[0]}; // @[Cat.scala 29:58]
  wire [1:0] fetch_start_f = {io_ifc_fetch_addr_f[0],_T_144}; // @[Cat.scala 29:58]
  wire  _T_32 = io_exu_bp_exu_mp_btag == fetch_rd_tag_f; // @[ifu_bp_ctl.scala 114:53]
  wire  _T_33 = _T_32 & exu_mp_valid; // @[ifu_bp_ctl.scala 114:73]
  wire  _T_34 = _T_33 & io_ifc_fetch_req_f; // @[ifu_bp_ctl.scala 114:88]
  wire  _T_35 = io_exu_bp_exu_mp_index == btb_rd_addr_f; // @[ifu_bp_ctl.scala 114:124]
  wire  fetch_mp_collision_f = _T_34 & _T_35; // @[ifu_bp_ctl.scala 114:109]
  wire  _T_36 = io_exu_bp_exu_mp_btag == fetch_rd_tag_p1_f; // @[ifu_bp_ctl.scala 115:56]
  wire  _T_37 = _T_36 & exu_mp_valid; // @[ifu_bp_ctl.scala 115:79]
  wire  _T_38 = _T_37 & io_ifc_fetch_req_f; // @[ifu_bp_ctl.scala 115:94]
  wire  _T_39 = io_exu_bp_exu_mp_index == btb_rd_addr_p1_f; // @[ifu_bp_ctl.scala 115:130]
  wire  fetch_mp_collision_p1_f = _T_38 & _T_39; // @[ifu_bp_ctl.scala 115:115]
  reg  exu_mp_way_f; // @[ifu_bp_ctl.scala 119:55]
  reg  exu_flush_final_d1; // @[ifu_bp_ctl.scala 120:61]
  wire [255:0] mp_wrindex_dec = 256'h1 << io_exu_bp_exu_mp_index; // @[ifu_bp_ctl.scala 191:28]
  wire [255:0] fetch_wrindex_dec = 256'h1 << btb_rd_addr_f; // @[ifu_bp_ctl.scala 194:31]
  wire [255:0] fetch_wrindex_p1_dec = 256'h1 << btb_rd_addr_p1_f; // @[ifu_bp_ctl.scala 197:34]
  wire [255:0] _T_150 = exu_mp_valid ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12]
  wire [255:0] mp_wrlru_b0 = mp_wrindex_dec & _T_150; // @[ifu_bp_ctl.scala 200:36]
  wire  _T_166 = bht_valid_f[0] | bht_valid_f[1]; // @[ifu_bp_ctl.scala 206:42]
  wire  _T_167 = _T_166 & io_ifc_fetch_req_f; // @[ifu_bp_ctl.scala 206:58]
  wire  lru_update_valid_f = _T_167 & _T; // @[ifu_bp_ctl.scala 206:79]
  wire [255:0] _T_170 = lru_update_valid_f ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12]
  wire [255:0] fetch_wrlru_b0 = fetch_wrindex_dec & _T_170; // @[ifu_bp_ctl.scala 208:42]
  wire [255:0] fetch_wrlru_p1_b0 = fetch_wrindex_p1_dec & _T_170; // @[ifu_bp_ctl.scala 209:48]
  wire [255:0] _T_173 = ~mp_wrlru_b0; // @[ifu_bp_ctl.scala 211:25]
  wire [255:0] _T_174 = ~fetch_wrlru_b0; // @[ifu_bp_ctl.scala 211:40]
  wire [255:0] btb_lru_b0_hold = _T_173 & _T_174; // @[ifu_bp_ctl.scala 211:38]
  wire  _T_176 = ~io_exu_bp_exu_mp_pkt_bits_way; // @[ifu_bp_ctl.scala 218:40]
  wire [255:0] _T_179 = _T_176 ? mp_wrlru_b0 : 256'h0; // @[Mux.scala 27:72]
  wire [255:0] _T_180 = tag_match_way0_f ? fetch_wrlru_b0 : 256'h0; // @[Mux.scala 27:72]
  wire [255:0] _T_181 = tag_match_way0_p1_f ? fetch_wrlru_p1_b0 : 256'h0; // @[Mux.scala 27:72]
  wire [255:0] _T_182 = _T_179 | _T_180; // @[Mux.scala 27:72]
  wire [255:0] _T_183 = _T_182 | _T_181; // @[Mux.scala 27:72]
  reg [255:0] btb_lru_b0_f; // @[lib.scala 374:16]
  wire [255:0] _T_185 = btb_lru_b0_hold & btb_lru_b0_f; // @[ifu_bp_ctl.scala 220:102]
  wire [255:0] _T_187 = fetch_wrindex_dec & btb_lru_b0_f; // @[ifu_bp_ctl.scala 223:78]
  wire  _T_188 = |_T_187; // @[ifu_bp_ctl.scala 223:94]
  wire  btb_lru_rd_f = fetch_mp_collision_f ? exu_mp_way_f : _T_188; // @[ifu_bp_ctl.scala 223:25]
  wire [255:0] _T_190 = fetch_wrindex_p1_dec & btb_lru_b0_f; // @[ifu_bp_ctl.scala 225:87]
  wire  _T_191 = |_T_190; // @[ifu_bp_ctl.scala 225:103]
  wire  btb_lru_rd_p1_f = fetch_mp_collision_p1_f ? exu_mp_way_f : _T_191; // @[ifu_bp_ctl.scala 225:28]
  wire [1:0] _T_194 = {btb_lru_rd_f,btb_lru_rd_f}; // @[Cat.scala 29:58]
  wire [1:0] _T_197 = {btb_lru_rd_p1_f,btb_lru_rd_f}; // @[Cat.scala 29:58]
  wire [1:0] _T_198 = _T_144 ? _T_194 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_199 = io_ifc_fetch_addr_f[0] ? _T_197 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] btb_vlru_rd_f = _T_198 | _T_199; // @[Mux.scala 27:72]
  wire [1:0] _T_208 = {tag_match_way1_expanded_p1_f[0],tag_match_way1_expanded_f[1]}; // @[Cat.scala 29:58]
  wire [1:0] _T_209 = _T_144 ? tag_match_way1_expanded_f : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_210 = io_ifc_fetch_addr_f[0] ? _T_208 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] tag_match_vway1_expanded_f = _T_209 | _T_210; // @[Mux.scala 27:72]
  wire [1:0] _T_212 = ~bht_valid_f; // @[ifu_bp_ctl.scala 235:52]
  wire [1:0] _T_213 = _T_212 & btb_vlru_rd_f; // @[ifu_bp_ctl.scala 235:63]
  wire [15:0] _T_230 = btb_sel_f[1] ? btb_vbank1_rd_data_f[16:1] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_231 = btb_sel_f[0] ? btb_vbank0_rd_data_f[16:1] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] btb_sel_data_f = _T_230 | _T_231; // @[Mux.scala 27:72]
  wire [11:0] btb_rd_tgt_f = btb_sel_data_f[15:4]; // @[ifu_bp_ctl.scala 251:36]
  wire  btb_rd_pc4_f = btb_sel_data_f[3]; // @[ifu_bp_ctl.scala 252:36]
  wire  btb_rd_call_f = btb_sel_data_f[1]; // @[ifu_bp_ctl.scala 253:37]
  wire  btb_rd_ret_f = btb_sel_data_f[0]; // @[ifu_bp_ctl.scala 254:36]
  wire [1:0] _T_280 = {bht_vbank1_rd_data_f[1],bht_vbank0_rd_data_f[1]}; // @[Cat.scala 29:58]
  wire [1:0] hist1_raw = bht_force_taken_f | _T_280; // @[ifu_bp_ctl.scala 288:34]
  wire [1:0] _T_234 = bht_valid_f & hist1_raw; // @[ifu_bp_ctl.scala 261:39]
  wire  _T_235 = |_T_234; // @[ifu_bp_ctl.scala 261:52]
  wire  _T_236 = _T_235 & io_ifc_fetch_req_f; // @[ifu_bp_ctl.scala 261:56]
  wire  _T_237 = ~leak_one_f_d1; // @[ifu_bp_ctl.scala 261:79]
  wire  _T_238 = _T_236 & _T_237; // @[ifu_bp_ctl.scala 261:77]
  wire  _T_239 = ~io_dec_bp_dec_tlu_bpred_disable; // @[ifu_bp_ctl.scala 261:96]
  wire  _T_275 = io_ifu_bp_hit_taken_f & btb_sel_f[1]; // @[ifu_bp_ctl.scala 285:51]
  wire  _T_276 = ~io_ifu_bp_hit_taken_f; // @[ifu_bp_ctl.scala 285:69]
  wire  _T_286 = bht_valid_f[1] & btb_vbank1_rd_data_f[4]; // @[ifu_bp_ctl.scala 294:34]
  wire  _T_289 = bht_valid_f[0] & btb_vbank0_rd_data_f[4]; // @[ifu_bp_ctl.scala 295:34]
  wire  _T_292 = ~btb_vbank1_rd_data_f[2]; // @[ifu_bp_ctl.scala 298:37]
  wire  _T_293 = bht_valid_f[1] & _T_292; // @[ifu_bp_ctl.scala 298:35]
  wire  _T_295 = _T_293 & btb_vbank1_rd_data_f[1]; // @[ifu_bp_ctl.scala 298:65]
  wire  _T_298 = ~btb_vbank0_rd_data_f[2]; // @[ifu_bp_ctl.scala 299:37]
  wire  _T_299 = bht_valid_f[0] & _T_298; // @[ifu_bp_ctl.scala 299:35]
  wire  _T_301 = _T_299 & btb_vbank0_rd_data_f[1]; // @[ifu_bp_ctl.scala 299:65]
  wire [1:0] num_valids = bht_valid_f[1] + bht_valid_f[0]; // @[ifu_bp_ctl.scala 302:35]
  wire [1:0] _T_304 = btb_sel_f & bht_dir_f; // @[ifu_bp_ctl.scala 305:28]
  wire  final_h = |_T_304; // @[ifu_bp_ctl.scala 305:41]
  wire  _T_305 = num_valids == 2'h2; // @[ifu_bp_ctl.scala 309:41]
  wire [7:0] _T_309 = {fghr[5:0],1'h0,final_h}; // @[Cat.scala 29:58]
  wire  _T_310 = num_valids == 2'h1; // @[ifu_bp_ctl.scala 310:41]
  wire [7:0] _T_313 = {fghr[6:0],final_h}; // @[Cat.scala 29:58]
  wire  _T_314 = num_valids == 2'h0; // @[ifu_bp_ctl.scala 311:41]
  wire [7:0] _T_317 = _T_305 ? _T_309 : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_318 = _T_310 ? _T_313 : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_319 = _T_314 ? fghr : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_320 = _T_317 | _T_318; // @[Mux.scala 27:72]
  wire [7:0] merged_ghr = _T_320 | _T_319; // @[Mux.scala 27:72]
  wire  _T_323 = ~exu_flush_final_d1; // @[ifu_bp_ctl.scala 320:27]
  wire  _T_324 = _T_323 & io_ifc_fetch_req_f; // @[ifu_bp_ctl.scala 320:47]
  wire  _T_325 = _T_324 & io_ic_hit_f; // @[ifu_bp_ctl.scala 320:70]
  wire  _T_327 = _T_325 & _T_237; // @[ifu_bp_ctl.scala 320:84]
  wire  _T_330 = io_ifc_fetch_req_f & io_ic_hit_f; // @[ifu_bp_ctl.scala 321:70]
  wire  _T_332 = _T_330 & _T_237; // @[ifu_bp_ctl.scala 321:84]
  wire  _T_333 = ~_T_332; // @[ifu_bp_ctl.scala 321:49]
  wire  _T_334 = _T_323 & _T_333; // @[ifu_bp_ctl.scala 321:47]
  wire [7:0] _T_336 = exu_flush_final_d1 ? io_exu_bp_exu_mp_fghr : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_337 = _T_327 ? merged_ghr : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_338 = _T_334 ? fghr : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_339 = _T_336 | _T_337; // @[Mux.scala 27:72]
  wire [1:0] _T_344 = io_dec_bp_dec_tlu_bpred_disable ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [1:0] _T_345 = ~_T_344; // @[ifu_bp_ctl.scala 330:36]
  wire  _T_349 = ~fetch_start_f[0]; // @[ifu_bp_ctl.scala 334:36]
  wire  _T_350 = bht_dir_f[0] & _T_349; // @[ifu_bp_ctl.scala 334:34]
  wire  _T_354 = _T_14 & fetch_start_f[0]; // @[ifu_bp_ctl.scala 334:72]
  wire  _T_355 = _T_350 | _T_354; // @[ifu_bp_ctl.scala 334:55]
  wire  _T_358 = bht_dir_f[0] & fetch_start_f[0]; // @[ifu_bp_ctl.scala 335:34]
  wire  _T_363 = _T_14 & _T_349; // @[ifu_bp_ctl.scala 335:71]
  wire  _T_364 = _T_358 | _T_363; // @[ifu_bp_ctl.scala 335:54]
  wire [1:0] bloc_f = {_T_355,_T_364}; // @[Cat.scala 29:58]
  wire  _T_368 = _T_14 & io_ifc_fetch_addr_f[0]; // @[ifu_bp_ctl.scala 337:35]
  wire  _T_369 = ~btb_rd_pc4_f; // @[ifu_bp_ctl.scala 337:62]
  wire  use_fa_plus = _T_368 & _T_369; // @[ifu_bp_ctl.scala 337:60]
  wire  _T_372 = fetch_start_f[0] & btb_sel_f[0]; // @[ifu_bp_ctl.scala 339:44]
  wire  btb_fg_crossing_f = _T_372 & btb_rd_pc4_f; // @[ifu_bp_ctl.scala 339:59]
  wire  bp_total_branch_offset_f = bloc_f[1] ^ btb_rd_pc4_f; // @[ifu_bp_ctl.scala 340:43]
  wire  _T_376 = io_ifc_fetch_req_f & _T_276; // @[ifu_bp_ctl.scala 342:85]
  reg [29:0] ifc_fetch_adder_prior; // @[lib.scala 374:16]
  wire  _T_381 = ~btb_fg_crossing_f; // @[ifu_bp_ctl.scala 348:32]
  wire  _T_382 = ~use_fa_plus; // @[ifu_bp_ctl.scala 348:53]
  wire  _T_383 = _T_381 & _T_382; // @[ifu_bp_ctl.scala 348:51]
  wire [29:0] _T_386 = use_fa_plus ? fetch_addr_p1_f : 30'h0; // @[Mux.scala 27:72]
  wire [29:0] _T_387 = btb_fg_crossing_f ? ifc_fetch_adder_prior : 30'h0; // @[Mux.scala 27:72]
  wire [29:0] _T_388 = _T_383 ? io_ifc_fetch_addr_f[30:1] : 30'h0; // @[Mux.scala 27:72]
  wire [29:0] _T_389 = _T_386 | _T_387; // @[Mux.scala 27:72]
  wire [29:0] adder_pc_in_f = _T_389 | _T_388; // @[Mux.scala 27:72]
  wire [31:0] _T_393 = {adder_pc_in_f,bp_total_branch_offset_f,1'h0}; // @[Cat.scala 29:58]
  wire [12:0] _T_394 = {btb_rd_tgt_f,1'h0}; // @[Cat.scala 29:58]
  wire [12:0] _T_397 = _T_393[12:1] + _T_394[12:1]; // @[lib.scala 68:31]
  wire [18:0] _T_400 = _T_393[31:13] + 19'h1; // @[lib.scala 69:27]
  wire [18:0] _T_403 = _T_393[31:13] - 19'h1; // @[lib.scala 70:27]
  wire  _T_406 = ~_T_397[12]; // @[lib.scala 72:28]
  wire  _T_407 = _T_394[12] ^ _T_406; // @[lib.scala 72:26]
  wire  _T_410 = ~_T_394[12]; // @[lib.scala 73:20]
  wire  _T_412 = _T_410 & _T_397[12]; // @[lib.scala 73:26]
  wire  _T_416 = _T_394[12] & _T_406; // @[lib.scala 74:26]
  wire [18:0] _T_418 = _T_407 ? _T_393[31:13] : 19'h0; // @[Mux.scala 27:72]
  wire [18:0] _T_419 = _T_412 ? _T_400 : 19'h0; // @[Mux.scala 27:72]
  wire [18:0] _T_420 = _T_416 ? _T_403 : 19'h0; // @[Mux.scala 27:72]
  wire [18:0] _T_421 = _T_418 | _T_419; // @[Mux.scala 27:72]
  wire [18:0] _T_422 = _T_421 | _T_420; // @[Mux.scala 27:72]
  wire [31:0] bp_btb_target_adder_f = {_T_422,_T_397[11:0],1'h0}; // @[Cat.scala 29:58]
  wire  _T_426 = ~btb_rd_call_f; // @[ifu_bp_ctl.scala 357:49]
  wire  _T_427 = btb_rd_ret_f & _T_426; // @[ifu_bp_ctl.scala 357:47]
  reg [31:0] rets_out_0; // @[lib.scala 374:16]
  wire  _T_429 = _T_427 & rets_out_0[0]; // @[ifu_bp_ctl.scala 357:64]
  wire [12:0] _T_440 = {11'h0,_T_369,1'h0}; // @[Cat.scala 29:58]
  wire [12:0] _T_443 = _T_393[12:1] + _T_440[12:1]; // @[lib.scala 68:31]
  wire  _T_452 = ~_T_443[12]; // @[lib.scala 72:28]
  wire  _T_453 = _T_440[12] ^ _T_452; // @[lib.scala 72:26]
  wire  _T_456 = ~_T_440[12]; // @[lib.scala 73:20]
  wire  _T_458 = _T_456 & _T_443[12]; // @[lib.scala 73:26]
  wire  _T_462 = _T_440[12] & _T_452; // @[lib.scala 74:26]
  wire [18:0] _T_464 = _T_453 ? _T_393[31:13] : 19'h0; // @[Mux.scala 27:72]
  wire [18:0] _T_465 = _T_458 ? _T_400 : 19'h0; // @[Mux.scala 27:72]
  wire [18:0] _T_466 = _T_462 ? _T_403 : 19'h0; // @[Mux.scala 27:72]
  wire [18:0] _T_467 = _T_464 | _T_465; // @[Mux.scala 27:72]
  wire [18:0] _T_468 = _T_467 | _T_466; // @[Mux.scala 27:72]
  wire [31:0] bp_rs_call_target_f = {_T_468,_T_443[11:0],1'h0}; // @[Cat.scala 29:58]
  wire  _T_472 = ~btb_rd_ret_f; // @[ifu_bp_ctl.scala 363:33]
  wire  _T_473 = btb_rd_call_f & _T_472; // @[ifu_bp_ctl.scala 363:31]
  wire  rs_push = _T_473 & io_ifu_bp_hit_taken_f; // @[ifu_bp_ctl.scala 363:47]
  wire  rs_pop = _T_427 & io_ifu_bp_hit_taken_f; // @[ifu_bp_ctl.scala 364:46]
  wire  _T_476 = ~rs_push; // @[ifu_bp_ctl.scala 365:17]
  wire  _T_477 = ~rs_pop; // @[ifu_bp_ctl.scala 365:28]
  wire  rs_hold = _T_476 & _T_477; // @[ifu_bp_ctl.scala 365:26]
  wire [31:0] _T_480 = {bp_rs_call_target_f[31:1],1'h1}; // @[Cat.scala 29:58]
  wire [31:0] _T_482 = rs_push ? _T_480 : 32'h0; // @[Mux.scala 27:72]
  reg [31:0] rets_out_1; // @[lib.scala 374:16]
  wire [31:0] _T_483 = rs_pop ? rets_out_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_487 = rs_push ? rets_out_0 : 32'h0; // @[Mux.scala 27:72]
  reg [31:0] rets_out_2; // @[lib.scala 374:16]
  wire [31:0] _T_488 = rs_pop ? rets_out_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_492 = rs_push ? rets_out_1 : 32'h0; // @[Mux.scala 27:72]
  reg [31:0] rets_out_3; // @[lib.scala 374:16]
  wire [31:0] _T_493 = rs_pop ? rets_out_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_497 = rs_push ? rets_out_2 : 32'h0; // @[Mux.scala 27:72]
  reg [31:0] rets_out_4; // @[lib.scala 374:16]
  wire [31:0] _T_498 = rs_pop ? rets_out_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_502 = rs_push ? rets_out_3 : 32'h0; // @[Mux.scala 27:72]
  reg [31:0] rets_out_5; // @[lib.scala 374:16]
  wire [31:0] _T_503 = rs_pop ? rets_out_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_507 = rs_push ? rets_out_4 : 32'h0; // @[Mux.scala 27:72]
  reg [31:0] rets_out_6; // @[lib.scala 374:16]
  wire [31:0] _T_508 = rs_pop ? rets_out_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_512 = rs_push ? rets_out_5 : 32'h0; // @[Mux.scala 27:72]
  reg [31:0] rets_out_7; // @[lib.scala 374:16]
  wire [31:0] _T_513 = rs_pop ? rets_out_7 : 32'h0; // @[Mux.scala 27:72]
  wire  _T_531 = ~dec_tlu_error_wb; // @[ifu_bp_ctl.scala 380:35]
  wire  btb_valid = exu_mp_valid & _T_531; // @[ifu_bp_ctl.scala 380:32]
  wire  _T_532 = io_exu_bp_exu_mp_pkt_bits_pcall | io_exu_bp_exu_mp_pkt_bits_pja; // @[ifu_bp_ctl.scala 384:89]
  wire  _T_533 = io_exu_bp_exu_mp_pkt_bits_pret | io_exu_bp_exu_mp_pkt_bits_pja; // @[ifu_bp_ctl.scala 384:113]
  wire [2:0] _T_535 = {_T_532,_T_533,btb_valid}; // @[Cat.scala 29:58]
  wire [18:0] _T_538 = {io_exu_bp_exu_mp_btag,io_exu_bp_exu_mp_pkt_bits_toffset,io_exu_bp_exu_mp_pkt_bits_pc4,io_exu_bp_exu_mp_pkt_bits_boffset}; // @[Cat.scala 29:58]
  wire  exu_mp_valid_write = exu_mp_valid & io_exu_bp_exu_mp_pkt_bits_ataken; // @[ifu_bp_ctl.scala 385:41]
  wire  _T_540 = _T_176 & exu_mp_valid_write; // @[ifu_bp_ctl.scala 388:39]
  wire  _T_542 = _T_540 & _T_531; // @[ifu_bp_ctl.scala 388:60]
  wire  _T_543 = ~io_dec_bp_dec_tlu_br0_r_pkt_bits_way; // @[ifu_bp_ctl.scala 388:87]
  wire  _T_544 = _T_543 & dec_tlu_error_wb; // @[ifu_bp_ctl.scala 388:104]
  wire  btb_wr_en_way0 = _T_542 | _T_544; // @[ifu_bp_ctl.scala 388:83]
  wire  _T_545 = io_exu_bp_exu_mp_pkt_bits_way & exu_mp_valid_write; // @[ifu_bp_ctl.scala 389:36]
  wire  _T_547 = _T_545 & _T_531; // @[ifu_bp_ctl.scala 389:57]
  wire  _T_548 = io_dec_bp_dec_tlu_br0_r_pkt_bits_way & dec_tlu_error_wb; // @[ifu_bp_ctl.scala 389:98]
  wire  btb_wr_en_way1 = _T_547 | _T_548; // @[ifu_bp_ctl.scala 389:80]
  wire [7:0] btb_wr_addr = dec_tlu_error_wb ? io_exu_bp_exu_i0_br_index_r : io_exu_bp_exu_mp_index; // @[ifu_bp_ctl.scala 392:24]
  wire  middle_of_bank = io_exu_bp_exu_mp_pkt_bits_pc4 ^ io_exu_bp_exu_mp_pkt_bits_boffset; // @[ifu_bp_ctl.scala 393:35]
  wire  _T_550 = ~io_exu_bp_exu_mp_pkt_bits_pcall; // @[ifu_bp_ctl.scala 396:43]
  wire  _T_551 = exu_mp_valid & _T_550; // @[ifu_bp_ctl.scala 396:41]
  wire  _T_552 = ~io_exu_bp_exu_mp_pkt_bits_pret; // @[ifu_bp_ctl.scala 396:58]
  wire  _T_553 = _T_551 & _T_552; // @[ifu_bp_ctl.scala 396:56]
  wire  _T_554 = ~io_exu_bp_exu_mp_pkt_bits_pja; // @[ifu_bp_ctl.scala 396:72]
  wire  _T_555 = _T_553 & _T_554; // @[ifu_bp_ctl.scala 396:70]
  wire [1:0] _T_557 = _T_555 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire  _T_558 = ~middle_of_bank; // @[ifu_bp_ctl.scala 396:106]
  wire [1:0] _T_559 = {middle_of_bank,_T_558}; // @[Cat.scala 29:58]
  wire [1:0] bht_wr_en0 = _T_557 & _T_559; // @[ifu_bp_ctl.scala 396:84]
  wire [1:0] _T_561 = io_dec_bp_dec_tlu_br0_r_pkt_valid ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire  _T_562 = ~io_dec_bp_dec_tlu_br0_r_pkt_bits_middle; // @[ifu_bp_ctl.scala 397:75]
  wire [1:0] _T_563 = {io_dec_bp_dec_tlu_br0_r_pkt_bits_middle,_T_562}; // @[Cat.scala 29:58]
  wire [1:0] bht_wr_en2 = _T_561 & _T_563; // @[ifu_bp_ctl.scala 397:46]
  wire [9:0] _T_564 = {io_exu_bp_exu_mp_index,2'h0}; // @[Cat.scala 29:58]
  wire [7:0] bht_wr_addr0 = _T_564[9:2] ^ io_exu_bp_exu_mp_eghr; // @[lib.scala 56:35]
  wire [9:0] _T_567 = {io_exu_bp_exu_i0_br_index_r,2'h0}; // @[Cat.scala 29:58]
  wire [7:0] bht_wr_addr2 = _T_567[9:2] ^ io_exu_bp_exu_i0_br_fghr_r; // @[lib.scala 56:35]
  wire  _T_576 = btb_wr_addr == 8'h0; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_579 = btb_wr_addr == 8'h1; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_582 = btb_wr_addr == 8'h2; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_585 = btb_wr_addr == 8'h3; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_588 = btb_wr_addr == 8'h4; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_591 = btb_wr_addr == 8'h5; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_594 = btb_wr_addr == 8'h6; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_597 = btb_wr_addr == 8'h7; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_600 = btb_wr_addr == 8'h8; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_603 = btb_wr_addr == 8'h9; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_606 = btb_wr_addr == 8'ha; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_609 = btb_wr_addr == 8'hb; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_612 = btb_wr_addr == 8'hc; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_615 = btb_wr_addr == 8'hd; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_618 = btb_wr_addr == 8'he; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_621 = btb_wr_addr == 8'hf; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_624 = btb_wr_addr == 8'h10; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_627 = btb_wr_addr == 8'h11; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_630 = btb_wr_addr == 8'h12; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_633 = btb_wr_addr == 8'h13; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_636 = btb_wr_addr == 8'h14; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_639 = btb_wr_addr == 8'h15; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_642 = btb_wr_addr == 8'h16; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_645 = btb_wr_addr == 8'h17; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_648 = btb_wr_addr == 8'h18; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_651 = btb_wr_addr == 8'h19; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_654 = btb_wr_addr == 8'h1a; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_657 = btb_wr_addr == 8'h1b; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_660 = btb_wr_addr == 8'h1c; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_663 = btb_wr_addr == 8'h1d; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_666 = btb_wr_addr == 8'h1e; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_669 = btb_wr_addr == 8'h1f; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_672 = btb_wr_addr == 8'h20; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_675 = btb_wr_addr == 8'h21; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_678 = btb_wr_addr == 8'h22; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_681 = btb_wr_addr == 8'h23; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_684 = btb_wr_addr == 8'h24; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_687 = btb_wr_addr == 8'h25; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_690 = btb_wr_addr == 8'h26; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_693 = btb_wr_addr == 8'h27; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_696 = btb_wr_addr == 8'h28; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_699 = btb_wr_addr == 8'h29; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_702 = btb_wr_addr == 8'h2a; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_705 = btb_wr_addr == 8'h2b; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_708 = btb_wr_addr == 8'h2c; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_711 = btb_wr_addr == 8'h2d; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_714 = btb_wr_addr == 8'h2e; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_717 = btb_wr_addr == 8'h2f; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_720 = btb_wr_addr == 8'h30; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_723 = btb_wr_addr == 8'h31; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_726 = btb_wr_addr == 8'h32; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_729 = btb_wr_addr == 8'h33; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_732 = btb_wr_addr == 8'h34; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_735 = btb_wr_addr == 8'h35; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_738 = btb_wr_addr == 8'h36; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_741 = btb_wr_addr == 8'h37; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_744 = btb_wr_addr == 8'h38; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_747 = btb_wr_addr == 8'h39; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_750 = btb_wr_addr == 8'h3a; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_753 = btb_wr_addr == 8'h3b; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_756 = btb_wr_addr == 8'h3c; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_759 = btb_wr_addr == 8'h3d; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_762 = btb_wr_addr == 8'h3e; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_765 = btb_wr_addr == 8'h3f; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_768 = btb_wr_addr == 8'h40; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_771 = btb_wr_addr == 8'h41; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_774 = btb_wr_addr == 8'h42; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_777 = btb_wr_addr == 8'h43; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_780 = btb_wr_addr == 8'h44; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_783 = btb_wr_addr == 8'h45; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_786 = btb_wr_addr == 8'h46; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_789 = btb_wr_addr == 8'h47; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_792 = btb_wr_addr == 8'h48; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_795 = btb_wr_addr == 8'h49; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_798 = btb_wr_addr == 8'h4a; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_801 = btb_wr_addr == 8'h4b; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_804 = btb_wr_addr == 8'h4c; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_807 = btb_wr_addr == 8'h4d; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_810 = btb_wr_addr == 8'h4e; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_813 = btb_wr_addr == 8'h4f; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_816 = btb_wr_addr == 8'h50; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_819 = btb_wr_addr == 8'h51; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_822 = btb_wr_addr == 8'h52; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_825 = btb_wr_addr == 8'h53; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_828 = btb_wr_addr == 8'h54; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_831 = btb_wr_addr == 8'h55; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_834 = btb_wr_addr == 8'h56; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_837 = btb_wr_addr == 8'h57; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_840 = btb_wr_addr == 8'h58; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_843 = btb_wr_addr == 8'h59; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_846 = btb_wr_addr == 8'h5a; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_849 = btb_wr_addr == 8'h5b; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_852 = btb_wr_addr == 8'h5c; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_855 = btb_wr_addr == 8'h5d; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_858 = btb_wr_addr == 8'h5e; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_861 = btb_wr_addr == 8'h5f; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_864 = btb_wr_addr == 8'h60; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_867 = btb_wr_addr == 8'h61; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_870 = btb_wr_addr == 8'h62; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_873 = btb_wr_addr == 8'h63; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_876 = btb_wr_addr == 8'h64; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_879 = btb_wr_addr == 8'h65; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_882 = btb_wr_addr == 8'h66; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_885 = btb_wr_addr == 8'h67; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_888 = btb_wr_addr == 8'h68; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_891 = btb_wr_addr == 8'h69; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_894 = btb_wr_addr == 8'h6a; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_897 = btb_wr_addr == 8'h6b; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_900 = btb_wr_addr == 8'h6c; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_903 = btb_wr_addr == 8'h6d; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_906 = btb_wr_addr == 8'h6e; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_909 = btb_wr_addr == 8'h6f; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_912 = btb_wr_addr == 8'h70; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_915 = btb_wr_addr == 8'h71; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_918 = btb_wr_addr == 8'h72; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_921 = btb_wr_addr == 8'h73; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_924 = btb_wr_addr == 8'h74; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_927 = btb_wr_addr == 8'h75; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_930 = btb_wr_addr == 8'h76; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_933 = btb_wr_addr == 8'h77; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_936 = btb_wr_addr == 8'h78; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_939 = btb_wr_addr == 8'h79; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_942 = btb_wr_addr == 8'h7a; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_945 = btb_wr_addr == 8'h7b; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_948 = btb_wr_addr == 8'h7c; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_951 = btb_wr_addr == 8'h7d; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_954 = btb_wr_addr == 8'h7e; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_957 = btb_wr_addr == 8'h7f; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_960 = btb_wr_addr == 8'h80; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_963 = btb_wr_addr == 8'h81; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_966 = btb_wr_addr == 8'h82; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_969 = btb_wr_addr == 8'h83; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_972 = btb_wr_addr == 8'h84; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_975 = btb_wr_addr == 8'h85; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_978 = btb_wr_addr == 8'h86; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_981 = btb_wr_addr == 8'h87; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_984 = btb_wr_addr == 8'h88; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_987 = btb_wr_addr == 8'h89; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_990 = btb_wr_addr == 8'h8a; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_993 = btb_wr_addr == 8'h8b; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_996 = btb_wr_addr == 8'h8c; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_999 = btb_wr_addr == 8'h8d; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1002 = btb_wr_addr == 8'h8e; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1005 = btb_wr_addr == 8'h8f; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1008 = btb_wr_addr == 8'h90; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1011 = btb_wr_addr == 8'h91; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1014 = btb_wr_addr == 8'h92; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1017 = btb_wr_addr == 8'h93; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1020 = btb_wr_addr == 8'h94; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1023 = btb_wr_addr == 8'h95; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1026 = btb_wr_addr == 8'h96; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1029 = btb_wr_addr == 8'h97; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1032 = btb_wr_addr == 8'h98; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1035 = btb_wr_addr == 8'h99; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1038 = btb_wr_addr == 8'h9a; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1041 = btb_wr_addr == 8'h9b; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1044 = btb_wr_addr == 8'h9c; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1047 = btb_wr_addr == 8'h9d; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1050 = btb_wr_addr == 8'h9e; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1053 = btb_wr_addr == 8'h9f; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1056 = btb_wr_addr == 8'ha0; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1059 = btb_wr_addr == 8'ha1; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1062 = btb_wr_addr == 8'ha2; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1065 = btb_wr_addr == 8'ha3; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1068 = btb_wr_addr == 8'ha4; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1071 = btb_wr_addr == 8'ha5; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1074 = btb_wr_addr == 8'ha6; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1077 = btb_wr_addr == 8'ha7; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1080 = btb_wr_addr == 8'ha8; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1083 = btb_wr_addr == 8'ha9; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1086 = btb_wr_addr == 8'haa; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1089 = btb_wr_addr == 8'hab; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1092 = btb_wr_addr == 8'hac; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1095 = btb_wr_addr == 8'had; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1098 = btb_wr_addr == 8'hae; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1101 = btb_wr_addr == 8'haf; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1104 = btb_wr_addr == 8'hb0; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1107 = btb_wr_addr == 8'hb1; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1110 = btb_wr_addr == 8'hb2; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1113 = btb_wr_addr == 8'hb3; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1116 = btb_wr_addr == 8'hb4; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1119 = btb_wr_addr == 8'hb5; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1122 = btb_wr_addr == 8'hb6; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1125 = btb_wr_addr == 8'hb7; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1128 = btb_wr_addr == 8'hb8; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1131 = btb_wr_addr == 8'hb9; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1134 = btb_wr_addr == 8'hba; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1137 = btb_wr_addr == 8'hbb; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1140 = btb_wr_addr == 8'hbc; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1143 = btb_wr_addr == 8'hbd; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1146 = btb_wr_addr == 8'hbe; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1149 = btb_wr_addr == 8'hbf; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1152 = btb_wr_addr == 8'hc0; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1155 = btb_wr_addr == 8'hc1; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1158 = btb_wr_addr == 8'hc2; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1161 = btb_wr_addr == 8'hc3; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1164 = btb_wr_addr == 8'hc4; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1167 = btb_wr_addr == 8'hc5; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1170 = btb_wr_addr == 8'hc6; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1173 = btb_wr_addr == 8'hc7; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1176 = btb_wr_addr == 8'hc8; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1179 = btb_wr_addr == 8'hc9; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1182 = btb_wr_addr == 8'hca; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1185 = btb_wr_addr == 8'hcb; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1188 = btb_wr_addr == 8'hcc; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1191 = btb_wr_addr == 8'hcd; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1194 = btb_wr_addr == 8'hce; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1197 = btb_wr_addr == 8'hcf; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1200 = btb_wr_addr == 8'hd0; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1203 = btb_wr_addr == 8'hd1; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1206 = btb_wr_addr == 8'hd2; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1209 = btb_wr_addr == 8'hd3; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1212 = btb_wr_addr == 8'hd4; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1215 = btb_wr_addr == 8'hd5; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1218 = btb_wr_addr == 8'hd6; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1221 = btb_wr_addr == 8'hd7; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1224 = btb_wr_addr == 8'hd8; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1227 = btb_wr_addr == 8'hd9; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1230 = btb_wr_addr == 8'hda; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1233 = btb_wr_addr == 8'hdb; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1236 = btb_wr_addr == 8'hdc; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1239 = btb_wr_addr == 8'hdd; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1242 = btb_wr_addr == 8'hde; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1245 = btb_wr_addr == 8'hdf; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1248 = btb_wr_addr == 8'he0; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1251 = btb_wr_addr == 8'he1; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1254 = btb_wr_addr == 8'he2; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1257 = btb_wr_addr == 8'he3; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1260 = btb_wr_addr == 8'he4; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1263 = btb_wr_addr == 8'he5; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1266 = btb_wr_addr == 8'he6; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1269 = btb_wr_addr == 8'he7; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1272 = btb_wr_addr == 8'he8; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1275 = btb_wr_addr == 8'he9; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1278 = btb_wr_addr == 8'hea; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1281 = btb_wr_addr == 8'heb; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1284 = btb_wr_addr == 8'hec; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1287 = btb_wr_addr == 8'hed; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1290 = btb_wr_addr == 8'hee; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1293 = btb_wr_addr == 8'hef; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1296 = btb_wr_addr == 8'hf0; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1299 = btb_wr_addr == 8'hf1; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1302 = btb_wr_addr == 8'hf2; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1305 = btb_wr_addr == 8'hf3; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1308 = btb_wr_addr == 8'hf4; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1311 = btb_wr_addr == 8'hf5; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1314 = btb_wr_addr == 8'hf6; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1317 = btb_wr_addr == 8'hf7; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1320 = btb_wr_addr == 8'hf8; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1323 = btb_wr_addr == 8'hf9; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1326 = btb_wr_addr == 8'hfa; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1329 = btb_wr_addr == 8'hfb; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1332 = btb_wr_addr == 8'hfc; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1335 = btb_wr_addr == 8'hfd; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1338 = btb_wr_addr == 8'hfe; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1341 = btb_wr_addr == 8'hff; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_6210 = bht_wr_addr0[7:4] == 4'h0; // @[ifu_bp_ctl.scala 429:109]
  wire  _T_6212 = bht_wr_en0[0] & _T_6210; // @[ifu_bp_ctl.scala 429:44]
  wire  _T_6215 = bht_wr_addr2[7:4] == 4'h0; // @[ifu_bp_ctl.scala 430:109]
  wire  _T_6217 = bht_wr_en2[0] & _T_6215; // @[ifu_bp_ctl.scala 430:44]
  wire  _T_6221 = bht_wr_addr0[7:4] == 4'h1; // @[ifu_bp_ctl.scala 429:109]
  wire  _T_6223 = bht_wr_en0[0] & _T_6221; // @[ifu_bp_ctl.scala 429:44]
  wire  _T_6226 = bht_wr_addr2[7:4] == 4'h1; // @[ifu_bp_ctl.scala 430:109]
  wire  _T_6228 = bht_wr_en2[0] & _T_6226; // @[ifu_bp_ctl.scala 430:44]
  wire  _T_6232 = bht_wr_addr0[7:4] == 4'h2; // @[ifu_bp_ctl.scala 429:109]
  wire  _T_6234 = bht_wr_en0[0] & _T_6232; // @[ifu_bp_ctl.scala 429:44]
  wire  _T_6237 = bht_wr_addr2[7:4] == 4'h2; // @[ifu_bp_ctl.scala 430:109]
  wire  _T_6239 = bht_wr_en2[0] & _T_6237; // @[ifu_bp_ctl.scala 430:44]
  wire  _T_6243 = bht_wr_addr0[7:4] == 4'h3; // @[ifu_bp_ctl.scala 429:109]
  wire  _T_6245 = bht_wr_en0[0] & _T_6243; // @[ifu_bp_ctl.scala 429:44]
  wire  _T_6248 = bht_wr_addr2[7:4] == 4'h3; // @[ifu_bp_ctl.scala 430:109]
  wire  _T_6250 = bht_wr_en2[0] & _T_6248; // @[ifu_bp_ctl.scala 430:44]
  wire  _T_6254 = bht_wr_addr0[7:4] == 4'h4; // @[ifu_bp_ctl.scala 429:109]
  wire  _T_6256 = bht_wr_en0[0] & _T_6254; // @[ifu_bp_ctl.scala 429:44]
  wire  _T_6259 = bht_wr_addr2[7:4] == 4'h4; // @[ifu_bp_ctl.scala 430:109]
  wire  _T_6261 = bht_wr_en2[0] & _T_6259; // @[ifu_bp_ctl.scala 430:44]
  wire  _T_6265 = bht_wr_addr0[7:4] == 4'h5; // @[ifu_bp_ctl.scala 429:109]
  wire  _T_6267 = bht_wr_en0[0] & _T_6265; // @[ifu_bp_ctl.scala 429:44]
  wire  _T_6270 = bht_wr_addr2[7:4] == 4'h5; // @[ifu_bp_ctl.scala 430:109]
  wire  _T_6272 = bht_wr_en2[0] & _T_6270; // @[ifu_bp_ctl.scala 430:44]
  wire  _T_6276 = bht_wr_addr0[7:4] == 4'h6; // @[ifu_bp_ctl.scala 429:109]
  wire  _T_6278 = bht_wr_en0[0] & _T_6276; // @[ifu_bp_ctl.scala 429:44]
  wire  _T_6281 = bht_wr_addr2[7:4] == 4'h6; // @[ifu_bp_ctl.scala 430:109]
  wire  _T_6283 = bht_wr_en2[0] & _T_6281; // @[ifu_bp_ctl.scala 430:44]
  wire  _T_6287 = bht_wr_addr0[7:4] == 4'h7; // @[ifu_bp_ctl.scala 429:109]
  wire  _T_6289 = bht_wr_en0[0] & _T_6287; // @[ifu_bp_ctl.scala 429:44]
  wire  _T_6292 = bht_wr_addr2[7:4] == 4'h7; // @[ifu_bp_ctl.scala 430:109]
  wire  _T_6294 = bht_wr_en2[0] & _T_6292; // @[ifu_bp_ctl.scala 430:44]
  wire  _T_6298 = bht_wr_addr0[7:4] == 4'h8; // @[ifu_bp_ctl.scala 429:109]
  wire  _T_6300 = bht_wr_en0[0] & _T_6298; // @[ifu_bp_ctl.scala 429:44]
  wire  _T_6303 = bht_wr_addr2[7:4] == 4'h8; // @[ifu_bp_ctl.scala 430:109]
  wire  _T_6305 = bht_wr_en2[0] & _T_6303; // @[ifu_bp_ctl.scala 430:44]
  wire  _T_6309 = bht_wr_addr0[7:4] == 4'h9; // @[ifu_bp_ctl.scala 429:109]
  wire  _T_6311 = bht_wr_en0[0] & _T_6309; // @[ifu_bp_ctl.scala 429:44]
  wire  _T_6314 = bht_wr_addr2[7:4] == 4'h9; // @[ifu_bp_ctl.scala 430:109]
  wire  _T_6316 = bht_wr_en2[0] & _T_6314; // @[ifu_bp_ctl.scala 430:44]
  wire  _T_6320 = bht_wr_addr0[7:4] == 4'ha; // @[ifu_bp_ctl.scala 429:109]
  wire  _T_6322 = bht_wr_en0[0] & _T_6320; // @[ifu_bp_ctl.scala 429:44]
  wire  _T_6325 = bht_wr_addr2[7:4] == 4'ha; // @[ifu_bp_ctl.scala 430:109]
  wire  _T_6327 = bht_wr_en2[0] & _T_6325; // @[ifu_bp_ctl.scala 430:44]
  wire  _T_6331 = bht_wr_addr0[7:4] == 4'hb; // @[ifu_bp_ctl.scala 429:109]
  wire  _T_6333 = bht_wr_en0[0] & _T_6331; // @[ifu_bp_ctl.scala 429:44]
  wire  _T_6336 = bht_wr_addr2[7:4] == 4'hb; // @[ifu_bp_ctl.scala 430:109]
  wire  _T_6338 = bht_wr_en2[0] & _T_6336; // @[ifu_bp_ctl.scala 430:44]
  wire  _T_6342 = bht_wr_addr0[7:4] == 4'hc; // @[ifu_bp_ctl.scala 429:109]
  wire  _T_6344 = bht_wr_en0[0] & _T_6342; // @[ifu_bp_ctl.scala 429:44]
  wire  _T_6347 = bht_wr_addr2[7:4] == 4'hc; // @[ifu_bp_ctl.scala 430:109]
  wire  _T_6349 = bht_wr_en2[0] & _T_6347; // @[ifu_bp_ctl.scala 430:44]
  wire  _T_6353 = bht_wr_addr0[7:4] == 4'hd; // @[ifu_bp_ctl.scala 429:109]
  wire  _T_6355 = bht_wr_en0[0] & _T_6353; // @[ifu_bp_ctl.scala 429:44]
  wire  _T_6358 = bht_wr_addr2[7:4] == 4'hd; // @[ifu_bp_ctl.scala 430:109]
  wire  _T_6360 = bht_wr_en2[0] & _T_6358; // @[ifu_bp_ctl.scala 430:44]
  wire  _T_6364 = bht_wr_addr0[7:4] == 4'he; // @[ifu_bp_ctl.scala 429:109]
  wire  _T_6366 = bht_wr_en0[0] & _T_6364; // @[ifu_bp_ctl.scala 429:44]
  wire  _T_6369 = bht_wr_addr2[7:4] == 4'he; // @[ifu_bp_ctl.scala 430:109]
  wire  _T_6371 = bht_wr_en2[0] & _T_6369; // @[ifu_bp_ctl.scala 430:44]
  wire  _T_6375 = bht_wr_addr0[7:4] == 4'hf; // @[ifu_bp_ctl.scala 429:109]
  wire  _T_6377 = bht_wr_en0[0] & _T_6375; // @[ifu_bp_ctl.scala 429:44]
  wire  _T_6380 = bht_wr_addr2[7:4] == 4'hf; // @[ifu_bp_ctl.scala 430:109]
  wire  _T_6382 = bht_wr_en2[0] & _T_6380; // @[ifu_bp_ctl.scala 430:44]
  wire  _T_6388 = bht_wr_en0[1] & _T_6210; // @[ifu_bp_ctl.scala 429:44]
  wire  _T_6393 = bht_wr_en2[1] & _T_6215; // @[ifu_bp_ctl.scala 430:44]
  wire  _T_6399 = bht_wr_en0[1] & _T_6221; // @[ifu_bp_ctl.scala 429:44]
  wire  _T_6404 = bht_wr_en2[1] & _T_6226; // @[ifu_bp_ctl.scala 430:44]
  wire  _T_6410 = bht_wr_en0[1] & _T_6232; // @[ifu_bp_ctl.scala 429:44]
  wire  _T_6415 = bht_wr_en2[1] & _T_6237; // @[ifu_bp_ctl.scala 430:44]
  wire  _T_6421 = bht_wr_en0[1] & _T_6243; // @[ifu_bp_ctl.scala 429:44]
  wire  _T_6426 = bht_wr_en2[1] & _T_6248; // @[ifu_bp_ctl.scala 430:44]
  wire  _T_6432 = bht_wr_en0[1] & _T_6254; // @[ifu_bp_ctl.scala 429:44]
  wire  _T_6437 = bht_wr_en2[1] & _T_6259; // @[ifu_bp_ctl.scala 430:44]
  wire  _T_6443 = bht_wr_en0[1] & _T_6265; // @[ifu_bp_ctl.scala 429:44]
  wire  _T_6448 = bht_wr_en2[1] & _T_6270; // @[ifu_bp_ctl.scala 430:44]
  wire  _T_6454 = bht_wr_en0[1] & _T_6276; // @[ifu_bp_ctl.scala 429:44]
  wire  _T_6459 = bht_wr_en2[1] & _T_6281; // @[ifu_bp_ctl.scala 430:44]
  wire  _T_6465 = bht_wr_en0[1] & _T_6287; // @[ifu_bp_ctl.scala 429:44]
  wire  _T_6470 = bht_wr_en2[1] & _T_6292; // @[ifu_bp_ctl.scala 430:44]
  wire  _T_6476 = bht_wr_en0[1] & _T_6298; // @[ifu_bp_ctl.scala 429:44]
  wire  _T_6481 = bht_wr_en2[1] & _T_6303; // @[ifu_bp_ctl.scala 430:44]
  wire  _T_6487 = bht_wr_en0[1] & _T_6309; // @[ifu_bp_ctl.scala 429:44]
  wire  _T_6492 = bht_wr_en2[1] & _T_6314; // @[ifu_bp_ctl.scala 430:44]
  wire  _T_6498 = bht_wr_en0[1] & _T_6320; // @[ifu_bp_ctl.scala 429:44]
  wire  _T_6503 = bht_wr_en2[1] & _T_6325; // @[ifu_bp_ctl.scala 430:44]
  wire  _T_6509 = bht_wr_en0[1] & _T_6331; // @[ifu_bp_ctl.scala 429:44]
  wire  _T_6514 = bht_wr_en2[1] & _T_6336; // @[ifu_bp_ctl.scala 430:44]
  wire  _T_6520 = bht_wr_en0[1] & _T_6342; // @[ifu_bp_ctl.scala 429:44]
  wire  _T_6525 = bht_wr_en2[1] & _T_6347; // @[ifu_bp_ctl.scala 430:44]
  wire  _T_6531 = bht_wr_en0[1] & _T_6353; // @[ifu_bp_ctl.scala 429:44]
  wire  _T_6536 = bht_wr_en2[1] & _T_6358; // @[ifu_bp_ctl.scala 430:44]
  wire  _T_6542 = bht_wr_en0[1] & _T_6364; // @[ifu_bp_ctl.scala 429:44]
  wire  _T_6547 = bht_wr_en2[1] & _T_6369; // @[ifu_bp_ctl.scala 430:44]
  wire  _T_6553 = bht_wr_en0[1] & _T_6375; // @[ifu_bp_ctl.scala 429:44]
  wire  _T_6558 = bht_wr_en2[1] & _T_6380; // @[ifu_bp_ctl.scala 430:44]
  wire  _T_6562 = bht_wr_addr2[3:0] == 4'h0; // @[ifu_bp_ctl.scala 435:74]
  wire  _T_6563 = bht_wr_en2[0] & _T_6562; // @[ifu_bp_ctl.scala 435:23]
  wire  _T_6566 = _T_6563 & _T_6215; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_6571 = bht_wr_addr2[3:0] == 4'h1; // @[ifu_bp_ctl.scala 435:74]
  wire  _T_6572 = bht_wr_en2[0] & _T_6571; // @[ifu_bp_ctl.scala 435:23]
  wire  _T_6575 = _T_6572 & _T_6215; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_6580 = bht_wr_addr2[3:0] == 4'h2; // @[ifu_bp_ctl.scala 435:74]
  wire  _T_6581 = bht_wr_en2[0] & _T_6580; // @[ifu_bp_ctl.scala 435:23]
  wire  _T_6584 = _T_6581 & _T_6215; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_6589 = bht_wr_addr2[3:0] == 4'h3; // @[ifu_bp_ctl.scala 435:74]
  wire  _T_6590 = bht_wr_en2[0] & _T_6589; // @[ifu_bp_ctl.scala 435:23]
  wire  _T_6593 = _T_6590 & _T_6215; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_6598 = bht_wr_addr2[3:0] == 4'h4; // @[ifu_bp_ctl.scala 435:74]
  wire  _T_6599 = bht_wr_en2[0] & _T_6598; // @[ifu_bp_ctl.scala 435:23]
  wire  _T_6602 = _T_6599 & _T_6215; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_6607 = bht_wr_addr2[3:0] == 4'h5; // @[ifu_bp_ctl.scala 435:74]
  wire  _T_6608 = bht_wr_en2[0] & _T_6607; // @[ifu_bp_ctl.scala 435:23]
  wire  _T_6611 = _T_6608 & _T_6215; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_6616 = bht_wr_addr2[3:0] == 4'h6; // @[ifu_bp_ctl.scala 435:74]
  wire  _T_6617 = bht_wr_en2[0] & _T_6616; // @[ifu_bp_ctl.scala 435:23]
  wire  _T_6620 = _T_6617 & _T_6215; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_6625 = bht_wr_addr2[3:0] == 4'h7; // @[ifu_bp_ctl.scala 435:74]
  wire  _T_6626 = bht_wr_en2[0] & _T_6625; // @[ifu_bp_ctl.scala 435:23]
  wire  _T_6629 = _T_6626 & _T_6215; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_6634 = bht_wr_addr2[3:0] == 4'h8; // @[ifu_bp_ctl.scala 435:74]
  wire  _T_6635 = bht_wr_en2[0] & _T_6634; // @[ifu_bp_ctl.scala 435:23]
  wire  _T_6638 = _T_6635 & _T_6215; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_6643 = bht_wr_addr2[3:0] == 4'h9; // @[ifu_bp_ctl.scala 435:74]
  wire  _T_6644 = bht_wr_en2[0] & _T_6643; // @[ifu_bp_ctl.scala 435:23]
  wire  _T_6647 = _T_6644 & _T_6215; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_6652 = bht_wr_addr2[3:0] == 4'ha; // @[ifu_bp_ctl.scala 435:74]
  wire  _T_6653 = bht_wr_en2[0] & _T_6652; // @[ifu_bp_ctl.scala 435:23]
  wire  _T_6656 = _T_6653 & _T_6215; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_6661 = bht_wr_addr2[3:0] == 4'hb; // @[ifu_bp_ctl.scala 435:74]
  wire  _T_6662 = bht_wr_en2[0] & _T_6661; // @[ifu_bp_ctl.scala 435:23]
  wire  _T_6665 = _T_6662 & _T_6215; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_6670 = bht_wr_addr2[3:0] == 4'hc; // @[ifu_bp_ctl.scala 435:74]
  wire  _T_6671 = bht_wr_en2[0] & _T_6670; // @[ifu_bp_ctl.scala 435:23]
  wire  _T_6674 = _T_6671 & _T_6215; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_6679 = bht_wr_addr2[3:0] == 4'hd; // @[ifu_bp_ctl.scala 435:74]
  wire  _T_6680 = bht_wr_en2[0] & _T_6679; // @[ifu_bp_ctl.scala 435:23]
  wire  _T_6683 = _T_6680 & _T_6215; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_6688 = bht_wr_addr2[3:0] == 4'he; // @[ifu_bp_ctl.scala 435:74]
  wire  _T_6689 = bht_wr_en2[0] & _T_6688; // @[ifu_bp_ctl.scala 435:23]
  wire  _T_6692 = _T_6689 & _T_6215; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_6697 = bht_wr_addr2[3:0] == 4'hf; // @[ifu_bp_ctl.scala 435:74]
  wire  _T_6698 = bht_wr_en2[0] & _T_6697; // @[ifu_bp_ctl.scala 435:23]
  wire  _T_6701 = _T_6698 & _T_6215; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_6710 = _T_6563 & _T_6226; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_6719 = _T_6572 & _T_6226; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_6728 = _T_6581 & _T_6226; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_6737 = _T_6590 & _T_6226; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_6746 = _T_6599 & _T_6226; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_6755 = _T_6608 & _T_6226; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_6764 = _T_6617 & _T_6226; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_6773 = _T_6626 & _T_6226; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_6782 = _T_6635 & _T_6226; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_6791 = _T_6644 & _T_6226; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_6800 = _T_6653 & _T_6226; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_6809 = _T_6662 & _T_6226; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_6818 = _T_6671 & _T_6226; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_6827 = _T_6680 & _T_6226; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_6836 = _T_6689 & _T_6226; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_6845 = _T_6698 & _T_6226; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_6854 = _T_6563 & _T_6237; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_6863 = _T_6572 & _T_6237; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_6872 = _T_6581 & _T_6237; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_6881 = _T_6590 & _T_6237; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_6890 = _T_6599 & _T_6237; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_6899 = _T_6608 & _T_6237; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_6908 = _T_6617 & _T_6237; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_6917 = _T_6626 & _T_6237; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_6926 = _T_6635 & _T_6237; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_6935 = _T_6644 & _T_6237; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_6944 = _T_6653 & _T_6237; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_6953 = _T_6662 & _T_6237; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_6962 = _T_6671 & _T_6237; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_6971 = _T_6680 & _T_6237; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_6980 = _T_6689 & _T_6237; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_6989 = _T_6698 & _T_6237; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_6998 = _T_6563 & _T_6248; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7007 = _T_6572 & _T_6248; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7016 = _T_6581 & _T_6248; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7025 = _T_6590 & _T_6248; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7034 = _T_6599 & _T_6248; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7043 = _T_6608 & _T_6248; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7052 = _T_6617 & _T_6248; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7061 = _T_6626 & _T_6248; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7070 = _T_6635 & _T_6248; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7079 = _T_6644 & _T_6248; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7088 = _T_6653 & _T_6248; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7097 = _T_6662 & _T_6248; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7106 = _T_6671 & _T_6248; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7115 = _T_6680 & _T_6248; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7124 = _T_6689 & _T_6248; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7133 = _T_6698 & _T_6248; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7142 = _T_6563 & _T_6259; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7151 = _T_6572 & _T_6259; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7160 = _T_6581 & _T_6259; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7169 = _T_6590 & _T_6259; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7178 = _T_6599 & _T_6259; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7187 = _T_6608 & _T_6259; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7196 = _T_6617 & _T_6259; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7205 = _T_6626 & _T_6259; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7214 = _T_6635 & _T_6259; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7223 = _T_6644 & _T_6259; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7232 = _T_6653 & _T_6259; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7241 = _T_6662 & _T_6259; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7250 = _T_6671 & _T_6259; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7259 = _T_6680 & _T_6259; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7268 = _T_6689 & _T_6259; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7277 = _T_6698 & _T_6259; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7286 = _T_6563 & _T_6270; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7295 = _T_6572 & _T_6270; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7304 = _T_6581 & _T_6270; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7313 = _T_6590 & _T_6270; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7322 = _T_6599 & _T_6270; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7331 = _T_6608 & _T_6270; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7340 = _T_6617 & _T_6270; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7349 = _T_6626 & _T_6270; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7358 = _T_6635 & _T_6270; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7367 = _T_6644 & _T_6270; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7376 = _T_6653 & _T_6270; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7385 = _T_6662 & _T_6270; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7394 = _T_6671 & _T_6270; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7403 = _T_6680 & _T_6270; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7412 = _T_6689 & _T_6270; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7421 = _T_6698 & _T_6270; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7430 = _T_6563 & _T_6281; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7439 = _T_6572 & _T_6281; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7448 = _T_6581 & _T_6281; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7457 = _T_6590 & _T_6281; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7466 = _T_6599 & _T_6281; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7475 = _T_6608 & _T_6281; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7484 = _T_6617 & _T_6281; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7493 = _T_6626 & _T_6281; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7502 = _T_6635 & _T_6281; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7511 = _T_6644 & _T_6281; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7520 = _T_6653 & _T_6281; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7529 = _T_6662 & _T_6281; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7538 = _T_6671 & _T_6281; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7547 = _T_6680 & _T_6281; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7556 = _T_6689 & _T_6281; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7565 = _T_6698 & _T_6281; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7574 = _T_6563 & _T_6292; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7583 = _T_6572 & _T_6292; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7592 = _T_6581 & _T_6292; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7601 = _T_6590 & _T_6292; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7610 = _T_6599 & _T_6292; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7619 = _T_6608 & _T_6292; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7628 = _T_6617 & _T_6292; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7637 = _T_6626 & _T_6292; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7646 = _T_6635 & _T_6292; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7655 = _T_6644 & _T_6292; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7664 = _T_6653 & _T_6292; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7673 = _T_6662 & _T_6292; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7682 = _T_6671 & _T_6292; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7691 = _T_6680 & _T_6292; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7700 = _T_6689 & _T_6292; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7709 = _T_6698 & _T_6292; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7718 = _T_6563 & _T_6303; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7727 = _T_6572 & _T_6303; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7736 = _T_6581 & _T_6303; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7745 = _T_6590 & _T_6303; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7754 = _T_6599 & _T_6303; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7763 = _T_6608 & _T_6303; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7772 = _T_6617 & _T_6303; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7781 = _T_6626 & _T_6303; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7790 = _T_6635 & _T_6303; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7799 = _T_6644 & _T_6303; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7808 = _T_6653 & _T_6303; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7817 = _T_6662 & _T_6303; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7826 = _T_6671 & _T_6303; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7835 = _T_6680 & _T_6303; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7844 = _T_6689 & _T_6303; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7853 = _T_6698 & _T_6303; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7862 = _T_6563 & _T_6314; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7871 = _T_6572 & _T_6314; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7880 = _T_6581 & _T_6314; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7889 = _T_6590 & _T_6314; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7898 = _T_6599 & _T_6314; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7907 = _T_6608 & _T_6314; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7916 = _T_6617 & _T_6314; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7925 = _T_6626 & _T_6314; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7934 = _T_6635 & _T_6314; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7943 = _T_6644 & _T_6314; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7952 = _T_6653 & _T_6314; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7961 = _T_6662 & _T_6314; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7970 = _T_6671 & _T_6314; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7979 = _T_6680 & _T_6314; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7988 = _T_6689 & _T_6314; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7997 = _T_6698 & _T_6314; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8006 = _T_6563 & _T_6325; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8015 = _T_6572 & _T_6325; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8024 = _T_6581 & _T_6325; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8033 = _T_6590 & _T_6325; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8042 = _T_6599 & _T_6325; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8051 = _T_6608 & _T_6325; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8060 = _T_6617 & _T_6325; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8069 = _T_6626 & _T_6325; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8078 = _T_6635 & _T_6325; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8087 = _T_6644 & _T_6325; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8096 = _T_6653 & _T_6325; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8105 = _T_6662 & _T_6325; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8114 = _T_6671 & _T_6325; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8123 = _T_6680 & _T_6325; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8132 = _T_6689 & _T_6325; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8141 = _T_6698 & _T_6325; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8150 = _T_6563 & _T_6336; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8159 = _T_6572 & _T_6336; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8168 = _T_6581 & _T_6336; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8177 = _T_6590 & _T_6336; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8186 = _T_6599 & _T_6336; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8195 = _T_6608 & _T_6336; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8204 = _T_6617 & _T_6336; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8213 = _T_6626 & _T_6336; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8222 = _T_6635 & _T_6336; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8231 = _T_6644 & _T_6336; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8240 = _T_6653 & _T_6336; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8249 = _T_6662 & _T_6336; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8258 = _T_6671 & _T_6336; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8267 = _T_6680 & _T_6336; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8276 = _T_6689 & _T_6336; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8285 = _T_6698 & _T_6336; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8294 = _T_6563 & _T_6347; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8303 = _T_6572 & _T_6347; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8312 = _T_6581 & _T_6347; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8321 = _T_6590 & _T_6347; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8330 = _T_6599 & _T_6347; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8339 = _T_6608 & _T_6347; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8348 = _T_6617 & _T_6347; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8357 = _T_6626 & _T_6347; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8366 = _T_6635 & _T_6347; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8375 = _T_6644 & _T_6347; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8384 = _T_6653 & _T_6347; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8393 = _T_6662 & _T_6347; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8402 = _T_6671 & _T_6347; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8411 = _T_6680 & _T_6347; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8420 = _T_6689 & _T_6347; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8429 = _T_6698 & _T_6347; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8438 = _T_6563 & _T_6358; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8447 = _T_6572 & _T_6358; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8456 = _T_6581 & _T_6358; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8465 = _T_6590 & _T_6358; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8474 = _T_6599 & _T_6358; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8483 = _T_6608 & _T_6358; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8492 = _T_6617 & _T_6358; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8501 = _T_6626 & _T_6358; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8510 = _T_6635 & _T_6358; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8519 = _T_6644 & _T_6358; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8528 = _T_6653 & _T_6358; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8537 = _T_6662 & _T_6358; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8546 = _T_6671 & _T_6358; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8555 = _T_6680 & _T_6358; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8564 = _T_6689 & _T_6358; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8573 = _T_6698 & _T_6358; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8582 = _T_6563 & _T_6369; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8591 = _T_6572 & _T_6369; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8600 = _T_6581 & _T_6369; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8609 = _T_6590 & _T_6369; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8618 = _T_6599 & _T_6369; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8627 = _T_6608 & _T_6369; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8636 = _T_6617 & _T_6369; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8645 = _T_6626 & _T_6369; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8654 = _T_6635 & _T_6369; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8663 = _T_6644 & _T_6369; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8672 = _T_6653 & _T_6369; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8681 = _T_6662 & _T_6369; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8690 = _T_6671 & _T_6369; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8699 = _T_6680 & _T_6369; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8708 = _T_6689 & _T_6369; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8717 = _T_6698 & _T_6369; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8726 = _T_6563 & _T_6380; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8735 = _T_6572 & _T_6380; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8744 = _T_6581 & _T_6380; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8753 = _T_6590 & _T_6380; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8762 = _T_6599 & _T_6380; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8771 = _T_6608 & _T_6380; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8780 = _T_6617 & _T_6380; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8789 = _T_6626 & _T_6380; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8798 = _T_6635 & _T_6380; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8807 = _T_6644 & _T_6380; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8816 = _T_6653 & _T_6380; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8825 = _T_6662 & _T_6380; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8834 = _T_6671 & _T_6380; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8843 = _T_6680 & _T_6380; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8852 = _T_6689 & _T_6380; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8861 = _T_6698 & _T_6380; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8867 = bht_wr_en2[1] & _T_6562; // @[ifu_bp_ctl.scala 435:23]
  wire  _T_8870 = _T_8867 & _T_6215; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8876 = bht_wr_en2[1] & _T_6571; // @[ifu_bp_ctl.scala 435:23]
  wire  _T_8879 = _T_8876 & _T_6215; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8885 = bht_wr_en2[1] & _T_6580; // @[ifu_bp_ctl.scala 435:23]
  wire  _T_8888 = _T_8885 & _T_6215; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8894 = bht_wr_en2[1] & _T_6589; // @[ifu_bp_ctl.scala 435:23]
  wire  _T_8897 = _T_8894 & _T_6215; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8903 = bht_wr_en2[1] & _T_6598; // @[ifu_bp_ctl.scala 435:23]
  wire  _T_8906 = _T_8903 & _T_6215; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8912 = bht_wr_en2[1] & _T_6607; // @[ifu_bp_ctl.scala 435:23]
  wire  _T_8915 = _T_8912 & _T_6215; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8921 = bht_wr_en2[1] & _T_6616; // @[ifu_bp_ctl.scala 435:23]
  wire  _T_8924 = _T_8921 & _T_6215; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8930 = bht_wr_en2[1] & _T_6625; // @[ifu_bp_ctl.scala 435:23]
  wire  _T_8933 = _T_8930 & _T_6215; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8939 = bht_wr_en2[1] & _T_6634; // @[ifu_bp_ctl.scala 435:23]
  wire  _T_8942 = _T_8939 & _T_6215; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8948 = bht_wr_en2[1] & _T_6643; // @[ifu_bp_ctl.scala 435:23]
  wire  _T_8951 = _T_8948 & _T_6215; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8957 = bht_wr_en2[1] & _T_6652; // @[ifu_bp_ctl.scala 435:23]
  wire  _T_8960 = _T_8957 & _T_6215; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8966 = bht_wr_en2[1] & _T_6661; // @[ifu_bp_ctl.scala 435:23]
  wire  _T_8969 = _T_8966 & _T_6215; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8975 = bht_wr_en2[1] & _T_6670; // @[ifu_bp_ctl.scala 435:23]
  wire  _T_8978 = _T_8975 & _T_6215; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8984 = bht_wr_en2[1] & _T_6679; // @[ifu_bp_ctl.scala 435:23]
  wire  _T_8987 = _T_8984 & _T_6215; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8993 = bht_wr_en2[1] & _T_6688; // @[ifu_bp_ctl.scala 435:23]
  wire  _T_8996 = _T_8993 & _T_6215; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9002 = bht_wr_en2[1] & _T_6697; // @[ifu_bp_ctl.scala 435:23]
  wire  _T_9005 = _T_9002 & _T_6215; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9014 = _T_8867 & _T_6226; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9023 = _T_8876 & _T_6226; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9032 = _T_8885 & _T_6226; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9041 = _T_8894 & _T_6226; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9050 = _T_8903 & _T_6226; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9059 = _T_8912 & _T_6226; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9068 = _T_8921 & _T_6226; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9077 = _T_8930 & _T_6226; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9086 = _T_8939 & _T_6226; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9095 = _T_8948 & _T_6226; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9104 = _T_8957 & _T_6226; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9113 = _T_8966 & _T_6226; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9122 = _T_8975 & _T_6226; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9131 = _T_8984 & _T_6226; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9140 = _T_8993 & _T_6226; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9149 = _T_9002 & _T_6226; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9158 = _T_8867 & _T_6237; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9167 = _T_8876 & _T_6237; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9176 = _T_8885 & _T_6237; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9185 = _T_8894 & _T_6237; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9194 = _T_8903 & _T_6237; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9203 = _T_8912 & _T_6237; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9212 = _T_8921 & _T_6237; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9221 = _T_8930 & _T_6237; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9230 = _T_8939 & _T_6237; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9239 = _T_8948 & _T_6237; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9248 = _T_8957 & _T_6237; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9257 = _T_8966 & _T_6237; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9266 = _T_8975 & _T_6237; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9275 = _T_8984 & _T_6237; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9284 = _T_8993 & _T_6237; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9293 = _T_9002 & _T_6237; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9302 = _T_8867 & _T_6248; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9311 = _T_8876 & _T_6248; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9320 = _T_8885 & _T_6248; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9329 = _T_8894 & _T_6248; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9338 = _T_8903 & _T_6248; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9347 = _T_8912 & _T_6248; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9356 = _T_8921 & _T_6248; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9365 = _T_8930 & _T_6248; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9374 = _T_8939 & _T_6248; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9383 = _T_8948 & _T_6248; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9392 = _T_8957 & _T_6248; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9401 = _T_8966 & _T_6248; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9410 = _T_8975 & _T_6248; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9419 = _T_8984 & _T_6248; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9428 = _T_8993 & _T_6248; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9437 = _T_9002 & _T_6248; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9446 = _T_8867 & _T_6259; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9455 = _T_8876 & _T_6259; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9464 = _T_8885 & _T_6259; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9473 = _T_8894 & _T_6259; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9482 = _T_8903 & _T_6259; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9491 = _T_8912 & _T_6259; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9500 = _T_8921 & _T_6259; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9509 = _T_8930 & _T_6259; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9518 = _T_8939 & _T_6259; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9527 = _T_8948 & _T_6259; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9536 = _T_8957 & _T_6259; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9545 = _T_8966 & _T_6259; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9554 = _T_8975 & _T_6259; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9563 = _T_8984 & _T_6259; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9572 = _T_8993 & _T_6259; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9581 = _T_9002 & _T_6259; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9590 = _T_8867 & _T_6270; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9599 = _T_8876 & _T_6270; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9608 = _T_8885 & _T_6270; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9617 = _T_8894 & _T_6270; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9626 = _T_8903 & _T_6270; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9635 = _T_8912 & _T_6270; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9644 = _T_8921 & _T_6270; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9653 = _T_8930 & _T_6270; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9662 = _T_8939 & _T_6270; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9671 = _T_8948 & _T_6270; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9680 = _T_8957 & _T_6270; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9689 = _T_8966 & _T_6270; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9698 = _T_8975 & _T_6270; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9707 = _T_8984 & _T_6270; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9716 = _T_8993 & _T_6270; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9725 = _T_9002 & _T_6270; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9734 = _T_8867 & _T_6281; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9743 = _T_8876 & _T_6281; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9752 = _T_8885 & _T_6281; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9761 = _T_8894 & _T_6281; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9770 = _T_8903 & _T_6281; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9779 = _T_8912 & _T_6281; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9788 = _T_8921 & _T_6281; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9797 = _T_8930 & _T_6281; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9806 = _T_8939 & _T_6281; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9815 = _T_8948 & _T_6281; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9824 = _T_8957 & _T_6281; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9833 = _T_8966 & _T_6281; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9842 = _T_8975 & _T_6281; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9851 = _T_8984 & _T_6281; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9860 = _T_8993 & _T_6281; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9869 = _T_9002 & _T_6281; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9878 = _T_8867 & _T_6292; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9887 = _T_8876 & _T_6292; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9896 = _T_8885 & _T_6292; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9905 = _T_8894 & _T_6292; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9914 = _T_8903 & _T_6292; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9923 = _T_8912 & _T_6292; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9932 = _T_8921 & _T_6292; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9941 = _T_8930 & _T_6292; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9950 = _T_8939 & _T_6292; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9959 = _T_8948 & _T_6292; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9968 = _T_8957 & _T_6292; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9977 = _T_8966 & _T_6292; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9986 = _T_8975 & _T_6292; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9995 = _T_8984 & _T_6292; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10004 = _T_8993 & _T_6292; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10013 = _T_9002 & _T_6292; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10022 = _T_8867 & _T_6303; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10031 = _T_8876 & _T_6303; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10040 = _T_8885 & _T_6303; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10049 = _T_8894 & _T_6303; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10058 = _T_8903 & _T_6303; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10067 = _T_8912 & _T_6303; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10076 = _T_8921 & _T_6303; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10085 = _T_8930 & _T_6303; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10094 = _T_8939 & _T_6303; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10103 = _T_8948 & _T_6303; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10112 = _T_8957 & _T_6303; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10121 = _T_8966 & _T_6303; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10130 = _T_8975 & _T_6303; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10139 = _T_8984 & _T_6303; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10148 = _T_8993 & _T_6303; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10157 = _T_9002 & _T_6303; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10166 = _T_8867 & _T_6314; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10175 = _T_8876 & _T_6314; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10184 = _T_8885 & _T_6314; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10193 = _T_8894 & _T_6314; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10202 = _T_8903 & _T_6314; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10211 = _T_8912 & _T_6314; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10220 = _T_8921 & _T_6314; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10229 = _T_8930 & _T_6314; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10238 = _T_8939 & _T_6314; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10247 = _T_8948 & _T_6314; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10256 = _T_8957 & _T_6314; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10265 = _T_8966 & _T_6314; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10274 = _T_8975 & _T_6314; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10283 = _T_8984 & _T_6314; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10292 = _T_8993 & _T_6314; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10301 = _T_9002 & _T_6314; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10310 = _T_8867 & _T_6325; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10319 = _T_8876 & _T_6325; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10328 = _T_8885 & _T_6325; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10337 = _T_8894 & _T_6325; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10346 = _T_8903 & _T_6325; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10355 = _T_8912 & _T_6325; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10364 = _T_8921 & _T_6325; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10373 = _T_8930 & _T_6325; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10382 = _T_8939 & _T_6325; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10391 = _T_8948 & _T_6325; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10400 = _T_8957 & _T_6325; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10409 = _T_8966 & _T_6325; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10418 = _T_8975 & _T_6325; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10427 = _T_8984 & _T_6325; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10436 = _T_8993 & _T_6325; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10445 = _T_9002 & _T_6325; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10454 = _T_8867 & _T_6336; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10463 = _T_8876 & _T_6336; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10472 = _T_8885 & _T_6336; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10481 = _T_8894 & _T_6336; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10490 = _T_8903 & _T_6336; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10499 = _T_8912 & _T_6336; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10508 = _T_8921 & _T_6336; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10517 = _T_8930 & _T_6336; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10526 = _T_8939 & _T_6336; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10535 = _T_8948 & _T_6336; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10544 = _T_8957 & _T_6336; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10553 = _T_8966 & _T_6336; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10562 = _T_8975 & _T_6336; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10571 = _T_8984 & _T_6336; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10580 = _T_8993 & _T_6336; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10589 = _T_9002 & _T_6336; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10598 = _T_8867 & _T_6347; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10607 = _T_8876 & _T_6347; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10616 = _T_8885 & _T_6347; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10625 = _T_8894 & _T_6347; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10634 = _T_8903 & _T_6347; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10643 = _T_8912 & _T_6347; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10652 = _T_8921 & _T_6347; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10661 = _T_8930 & _T_6347; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10670 = _T_8939 & _T_6347; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10679 = _T_8948 & _T_6347; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10688 = _T_8957 & _T_6347; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10697 = _T_8966 & _T_6347; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10706 = _T_8975 & _T_6347; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10715 = _T_8984 & _T_6347; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10724 = _T_8993 & _T_6347; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10733 = _T_9002 & _T_6347; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10742 = _T_8867 & _T_6358; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10751 = _T_8876 & _T_6358; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10760 = _T_8885 & _T_6358; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10769 = _T_8894 & _T_6358; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10778 = _T_8903 & _T_6358; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10787 = _T_8912 & _T_6358; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10796 = _T_8921 & _T_6358; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10805 = _T_8930 & _T_6358; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10814 = _T_8939 & _T_6358; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10823 = _T_8948 & _T_6358; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10832 = _T_8957 & _T_6358; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10841 = _T_8966 & _T_6358; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10850 = _T_8975 & _T_6358; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10859 = _T_8984 & _T_6358; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10868 = _T_8993 & _T_6358; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10877 = _T_9002 & _T_6358; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10886 = _T_8867 & _T_6369; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10895 = _T_8876 & _T_6369; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10904 = _T_8885 & _T_6369; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10913 = _T_8894 & _T_6369; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10922 = _T_8903 & _T_6369; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10931 = _T_8912 & _T_6369; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10940 = _T_8921 & _T_6369; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10949 = _T_8930 & _T_6369; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10958 = _T_8939 & _T_6369; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10967 = _T_8948 & _T_6369; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10976 = _T_8957 & _T_6369; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10985 = _T_8966 & _T_6369; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10994 = _T_8975 & _T_6369; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_11003 = _T_8984 & _T_6369; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_11012 = _T_8993 & _T_6369; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_11021 = _T_9002 & _T_6369; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_11030 = _T_8867 & _T_6380; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_11039 = _T_8876 & _T_6380; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_11048 = _T_8885 & _T_6380; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_11057 = _T_8894 & _T_6380; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_11066 = _T_8903 & _T_6380; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_11075 = _T_8912 & _T_6380; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_11084 = _T_8921 & _T_6380; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_11093 = _T_8930 & _T_6380; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_11102 = _T_8939 & _T_6380; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_11111 = _T_8948 & _T_6380; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_11120 = _T_8957 & _T_6380; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_11129 = _T_8966 & _T_6380; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_11138 = _T_8975 & _T_6380; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_11147 = _T_8984 & _T_6380; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_11156 = _T_8993 & _T_6380; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_11165 = _T_9002 & _T_6380; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_11170 = bht_wr_addr0[3:0] == 4'h0; // @[ifu_bp_ctl.scala 443:97]
  wire  _T_11171 = bht_wr_en0[0] & _T_11170; // @[ifu_bp_ctl.scala 443:45]
  wire  _T_11175 = _T_11171 & _T_6210; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_0_0 = _T_11175 | _T_6566; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_11187 = bht_wr_addr0[3:0] == 4'h1; // @[ifu_bp_ctl.scala 443:97]
  wire  _T_11188 = bht_wr_en0[0] & _T_11187; // @[ifu_bp_ctl.scala 443:45]
  wire  _T_11192 = _T_11188 & _T_6210; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_0_1 = _T_11192 | _T_6575; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_11204 = bht_wr_addr0[3:0] == 4'h2; // @[ifu_bp_ctl.scala 443:97]
  wire  _T_11205 = bht_wr_en0[0] & _T_11204; // @[ifu_bp_ctl.scala 443:45]
  wire  _T_11209 = _T_11205 & _T_6210; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_0_2 = _T_11209 | _T_6584; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_11221 = bht_wr_addr0[3:0] == 4'h3; // @[ifu_bp_ctl.scala 443:97]
  wire  _T_11222 = bht_wr_en0[0] & _T_11221; // @[ifu_bp_ctl.scala 443:45]
  wire  _T_11226 = _T_11222 & _T_6210; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_0_3 = _T_11226 | _T_6593; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_11238 = bht_wr_addr0[3:0] == 4'h4; // @[ifu_bp_ctl.scala 443:97]
  wire  _T_11239 = bht_wr_en0[0] & _T_11238; // @[ifu_bp_ctl.scala 443:45]
  wire  _T_11243 = _T_11239 & _T_6210; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_0_4 = _T_11243 | _T_6602; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_11255 = bht_wr_addr0[3:0] == 4'h5; // @[ifu_bp_ctl.scala 443:97]
  wire  _T_11256 = bht_wr_en0[0] & _T_11255; // @[ifu_bp_ctl.scala 443:45]
  wire  _T_11260 = _T_11256 & _T_6210; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_0_5 = _T_11260 | _T_6611; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_11272 = bht_wr_addr0[3:0] == 4'h6; // @[ifu_bp_ctl.scala 443:97]
  wire  _T_11273 = bht_wr_en0[0] & _T_11272; // @[ifu_bp_ctl.scala 443:45]
  wire  _T_11277 = _T_11273 & _T_6210; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_0_6 = _T_11277 | _T_6620; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_11289 = bht_wr_addr0[3:0] == 4'h7; // @[ifu_bp_ctl.scala 443:97]
  wire  _T_11290 = bht_wr_en0[0] & _T_11289; // @[ifu_bp_ctl.scala 443:45]
  wire  _T_11294 = _T_11290 & _T_6210; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_0_7 = _T_11294 | _T_6629; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_11306 = bht_wr_addr0[3:0] == 4'h8; // @[ifu_bp_ctl.scala 443:97]
  wire  _T_11307 = bht_wr_en0[0] & _T_11306; // @[ifu_bp_ctl.scala 443:45]
  wire  _T_11311 = _T_11307 & _T_6210; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_0_8 = _T_11311 | _T_6638; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_11323 = bht_wr_addr0[3:0] == 4'h9; // @[ifu_bp_ctl.scala 443:97]
  wire  _T_11324 = bht_wr_en0[0] & _T_11323; // @[ifu_bp_ctl.scala 443:45]
  wire  _T_11328 = _T_11324 & _T_6210; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_0_9 = _T_11328 | _T_6647; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_11340 = bht_wr_addr0[3:0] == 4'ha; // @[ifu_bp_ctl.scala 443:97]
  wire  _T_11341 = bht_wr_en0[0] & _T_11340; // @[ifu_bp_ctl.scala 443:45]
  wire  _T_11345 = _T_11341 & _T_6210; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_0_10 = _T_11345 | _T_6656; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_11357 = bht_wr_addr0[3:0] == 4'hb; // @[ifu_bp_ctl.scala 443:97]
  wire  _T_11358 = bht_wr_en0[0] & _T_11357; // @[ifu_bp_ctl.scala 443:45]
  wire  _T_11362 = _T_11358 & _T_6210; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_0_11 = _T_11362 | _T_6665; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_11374 = bht_wr_addr0[3:0] == 4'hc; // @[ifu_bp_ctl.scala 443:97]
  wire  _T_11375 = bht_wr_en0[0] & _T_11374; // @[ifu_bp_ctl.scala 443:45]
  wire  _T_11379 = _T_11375 & _T_6210; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_0_12 = _T_11379 | _T_6674; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_11391 = bht_wr_addr0[3:0] == 4'hd; // @[ifu_bp_ctl.scala 443:97]
  wire  _T_11392 = bht_wr_en0[0] & _T_11391; // @[ifu_bp_ctl.scala 443:45]
  wire  _T_11396 = _T_11392 & _T_6210; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_0_13 = _T_11396 | _T_6683; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_11408 = bht_wr_addr0[3:0] == 4'he; // @[ifu_bp_ctl.scala 443:97]
  wire  _T_11409 = bht_wr_en0[0] & _T_11408; // @[ifu_bp_ctl.scala 443:45]
  wire  _T_11413 = _T_11409 & _T_6210; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_0_14 = _T_11413 | _T_6692; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_11425 = bht_wr_addr0[3:0] == 4'hf; // @[ifu_bp_ctl.scala 443:97]
  wire  _T_11426 = bht_wr_en0[0] & _T_11425; // @[ifu_bp_ctl.scala 443:45]
  wire  _T_11430 = _T_11426 & _T_6210; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_0_15 = _T_11430 | _T_6701; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_11447 = _T_11171 & _T_6221; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_1_0 = _T_11447 | _T_6710; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_11464 = _T_11188 & _T_6221; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_1_1 = _T_11464 | _T_6719; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_11481 = _T_11205 & _T_6221; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_1_2 = _T_11481 | _T_6728; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_11498 = _T_11222 & _T_6221; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_1_3 = _T_11498 | _T_6737; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_11515 = _T_11239 & _T_6221; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_1_4 = _T_11515 | _T_6746; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_11532 = _T_11256 & _T_6221; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_1_5 = _T_11532 | _T_6755; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_11549 = _T_11273 & _T_6221; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_1_6 = _T_11549 | _T_6764; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_11566 = _T_11290 & _T_6221; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_1_7 = _T_11566 | _T_6773; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_11583 = _T_11307 & _T_6221; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_1_8 = _T_11583 | _T_6782; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_11600 = _T_11324 & _T_6221; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_1_9 = _T_11600 | _T_6791; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_11617 = _T_11341 & _T_6221; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_1_10 = _T_11617 | _T_6800; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_11634 = _T_11358 & _T_6221; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_1_11 = _T_11634 | _T_6809; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_11651 = _T_11375 & _T_6221; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_1_12 = _T_11651 | _T_6818; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_11668 = _T_11392 & _T_6221; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_1_13 = _T_11668 | _T_6827; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_11685 = _T_11409 & _T_6221; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_1_14 = _T_11685 | _T_6836; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_11702 = _T_11426 & _T_6221; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_1_15 = _T_11702 | _T_6845; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_11719 = _T_11171 & _T_6232; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_2_0 = _T_11719 | _T_6854; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_11736 = _T_11188 & _T_6232; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_2_1 = _T_11736 | _T_6863; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_11753 = _T_11205 & _T_6232; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_2_2 = _T_11753 | _T_6872; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_11770 = _T_11222 & _T_6232; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_2_3 = _T_11770 | _T_6881; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_11787 = _T_11239 & _T_6232; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_2_4 = _T_11787 | _T_6890; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_11804 = _T_11256 & _T_6232; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_2_5 = _T_11804 | _T_6899; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_11821 = _T_11273 & _T_6232; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_2_6 = _T_11821 | _T_6908; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_11838 = _T_11290 & _T_6232; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_2_7 = _T_11838 | _T_6917; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_11855 = _T_11307 & _T_6232; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_2_8 = _T_11855 | _T_6926; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_11872 = _T_11324 & _T_6232; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_2_9 = _T_11872 | _T_6935; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_11889 = _T_11341 & _T_6232; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_2_10 = _T_11889 | _T_6944; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_11906 = _T_11358 & _T_6232; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_2_11 = _T_11906 | _T_6953; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_11923 = _T_11375 & _T_6232; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_2_12 = _T_11923 | _T_6962; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_11940 = _T_11392 & _T_6232; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_2_13 = _T_11940 | _T_6971; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_11957 = _T_11409 & _T_6232; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_2_14 = _T_11957 | _T_6980; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_11974 = _T_11426 & _T_6232; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_2_15 = _T_11974 | _T_6989; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_11991 = _T_11171 & _T_6243; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_3_0 = _T_11991 | _T_6998; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12008 = _T_11188 & _T_6243; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_3_1 = _T_12008 | _T_7007; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12025 = _T_11205 & _T_6243; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_3_2 = _T_12025 | _T_7016; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12042 = _T_11222 & _T_6243; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_3_3 = _T_12042 | _T_7025; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12059 = _T_11239 & _T_6243; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_3_4 = _T_12059 | _T_7034; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12076 = _T_11256 & _T_6243; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_3_5 = _T_12076 | _T_7043; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12093 = _T_11273 & _T_6243; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_3_6 = _T_12093 | _T_7052; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12110 = _T_11290 & _T_6243; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_3_7 = _T_12110 | _T_7061; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12127 = _T_11307 & _T_6243; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_3_8 = _T_12127 | _T_7070; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12144 = _T_11324 & _T_6243; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_3_9 = _T_12144 | _T_7079; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12161 = _T_11341 & _T_6243; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_3_10 = _T_12161 | _T_7088; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12178 = _T_11358 & _T_6243; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_3_11 = _T_12178 | _T_7097; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12195 = _T_11375 & _T_6243; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_3_12 = _T_12195 | _T_7106; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12212 = _T_11392 & _T_6243; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_3_13 = _T_12212 | _T_7115; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12229 = _T_11409 & _T_6243; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_3_14 = _T_12229 | _T_7124; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12246 = _T_11426 & _T_6243; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_3_15 = _T_12246 | _T_7133; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12263 = _T_11171 & _T_6254; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_4_0 = _T_12263 | _T_7142; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12280 = _T_11188 & _T_6254; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_4_1 = _T_12280 | _T_7151; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12297 = _T_11205 & _T_6254; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_4_2 = _T_12297 | _T_7160; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12314 = _T_11222 & _T_6254; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_4_3 = _T_12314 | _T_7169; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12331 = _T_11239 & _T_6254; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_4_4 = _T_12331 | _T_7178; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12348 = _T_11256 & _T_6254; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_4_5 = _T_12348 | _T_7187; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12365 = _T_11273 & _T_6254; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_4_6 = _T_12365 | _T_7196; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12382 = _T_11290 & _T_6254; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_4_7 = _T_12382 | _T_7205; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12399 = _T_11307 & _T_6254; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_4_8 = _T_12399 | _T_7214; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12416 = _T_11324 & _T_6254; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_4_9 = _T_12416 | _T_7223; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12433 = _T_11341 & _T_6254; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_4_10 = _T_12433 | _T_7232; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12450 = _T_11358 & _T_6254; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_4_11 = _T_12450 | _T_7241; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12467 = _T_11375 & _T_6254; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_4_12 = _T_12467 | _T_7250; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12484 = _T_11392 & _T_6254; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_4_13 = _T_12484 | _T_7259; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12501 = _T_11409 & _T_6254; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_4_14 = _T_12501 | _T_7268; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12518 = _T_11426 & _T_6254; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_4_15 = _T_12518 | _T_7277; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12535 = _T_11171 & _T_6265; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_5_0 = _T_12535 | _T_7286; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12552 = _T_11188 & _T_6265; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_5_1 = _T_12552 | _T_7295; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12569 = _T_11205 & _T_6265; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_5_2 = _T_12569 | _T_7304; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12586 = _T_11222 & _T_6265; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_5_3 = _T_12586 | _T_7313; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12603 = _T_11239 & _T_6265; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_5_4 = _T_12603 | _T_7322; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12620 = _T_11256 & _T_6265; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_5_5 = _T_12620 | _T_7331; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12637 = _T_11273 & _T_6265; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_5_6 = _T_12637 | _T_7340; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12654 = _T_11290 & _T_6265; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_5_7 = _T_12654 | _T_7349; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12671 = _T_11307 & _T_6265; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_5_8 = _T_12671 | _T_7358; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12688 = _T_11324 & _T_6265; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_5_9 = _T_12688 | _T_7367; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12705 = _T_11341 & _T_6265; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_5_10 = _T_12705 | _T_7376; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12722 = _T_11358 & _T_6265; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_5_11 = _T_12722 | _T_7385; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12739 = _T_11375 & _T_6265; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_5_12 = _T_12739 | _T_7394; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12756 = _T_11392 & _T_6265; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_5_13 = _T_12756 | _T_7403; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12773 = _T_11409 & _T_6265; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_5_14 = _T_12773 | _T_7412; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12790 = _T_11426 & _T_6265; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_5_15 = _T_12790 | _T_7421; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12807 = _T_11171 & _T_6276; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_6_0 = _T_12807 | _T_7430; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12824 = _T_11188 & _T_6276; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_6_1 = _T_12824 | _T_7439; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12841 = _T_11205 & _T_6276; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_6_2 = _T_12841 | _T_7448; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12858 = _T_11222 & _T_6276; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_6_3 = _T_12858 | _T_7457; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12875 = _T_11239 & _T_6276; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_6_4 = _T_12875 | _T_7466; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12892 = _T_11256 & _T_6276; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_6_5 = _T_12892 | _T_7475; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12909 = _T_11273 & _T_6276; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_6_6 = _T_12909 | _T_7484; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12926 = _T_11290 & _T_6276; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_6_7 = _T_12926 | _T_7493; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12943 = _T_11307 & _T_6276; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_6_8 = _T_12943 | _T_7502; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12960 = _T_11324 & _T_6276; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_6_9 = _T_12960 | _T_7511; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12977 = _T_11341 & _T_6276; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_6_10 = _T_12977 | _T_7520; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12994 = _T_11358 & _T_6276; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_6_11 = _T_12994 | _T_7529; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13011 = _T_11375 & _T_6276; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_6_12 = _T_13011 | _T_7538; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13028 = _T_11392 & _T_6276; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_6_13 = _T_13028 | _T_7547; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13045 = _T_11409 & _T_6276; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_6_14 = _T_13045 | _T_7556; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13062 = _T_11426 & _T_6276; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_6_15 = _T_13062 | _T_7565; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13079 = _T_11171 & _T_6287; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_7_0 = _T_13079 | _T_7574; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13096 = _T_11188 & _T_6287; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_7_1 = _T_13096 | _T_7583; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13113 = _T_11205 & _T_6287; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_7_2 = _T_13113 | _T_7592; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13130 = _T_11222 & _T_6287; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_7_3 = _T_13130 | _T_7601; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13147 = _T_11239 & _T_6287; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_7_4 = _T_13147 | _T_7610; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13164 = _T_11256 & _T_6287; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_7_5 = _T_13164 | _T_7619; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13181 = _T_11273 & _T_6287; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_7_6 = _T_13181 | _T_7628; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13198 = _T_11290 & _T_6287; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_7_7 = _T_13198 | _T_7637; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13215 = _T_11307 & _T_6287; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_7_8 = _T_13215 | _T_7646; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13232 = _T_11324 & _T_6287; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_7_9 = _T_13232 | _T_7655; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13249 = _T_11341 & _T_6287; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_7_10 = _T_13249 | _T_7664; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13266 = _T_11358 & _T_6287; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_7_11 = _T_13266 | _T_7673; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13283 = _T_11375 & _T_6287; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_7_12 = _T_13283 | _T_7682; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13300 = _T_11392 & _T_6287; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_7_13 = _T_13300 | _T_7691; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13317 = _T_11409 & _T_6287; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_7_14 = _T_13317 | _T_7700; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13334 = _T_11426 & _T_6287; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_7_15 = _T_13334 | _T_7709; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13351 = _T_11171 & _T_6298; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_8_0 = _T_13351 | _T_7718; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13368 = _T_11188 & _T_6298; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_8_1 = _T_13368 | _T_7727; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13385 = _T_11205 & _T_6298; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_8_2 = _T_13385 | _T_7736; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13402 = _T_11222 & _T_6298; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_8_3 = _T_13402 | _T_7745; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13419 = _T_11239 & _T_6298; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_8_4 = _T_13419 | _T_7754; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13436 = _T_11256 & _T_6298; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_8_5 = _T_13436 | _T_7763; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13453 = _T_11273 & _T_6298; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_8_6 = _T_13453 | _T_7772; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13470 = _T_11290 & _T_6298; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_8_7 = _T_13470 | _T_7781; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13487 = _T_11307 & _T_6298; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_8_8 = _T_13487 | _T_7790; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13504 = _T_11324 & _T_6298; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_8_9 = _T_13504 | _T_7799; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13521 = _T_11341 & _T_6298; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_8_10 = _T_13521 | _T_7808; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13538 = _T_11358 & _T_6298; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_8_11 = _T_13538 | _T_7817; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13555 = _T_11375 & _T_6298; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_8_12 = _T_13555 | _T_7826; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13572 = _T_11392 & _T_6298; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_8_13 = _T_13572 | _T_7835; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13589 = _T_11409 & _T_6298; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_8_14 = _T_13589 | _T_7844; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13606 = _T_11426 & _T_6298; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_8_15 = _T_13606 | _T_7853; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13623 = _T_11171 & _T_6309; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_9_0 = _T_13623 | _T_7862; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13640 = _T_11188 & _T_6309; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_9_1 = _T_13640 | _T_7871; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13657 = _T_11205 & _T_6309; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_9_2 = _T_13657 | _T_7880; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13674 = _T_11222 & _T_6309; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_9_3 = _T_13674 | _T_7889; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13691 = _T_11239 & _T_6309; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_9_4 = _T_13691 | _T_7898; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13708 = _T_11256 & _T_6309; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_9_5 = _T_13708 | _T_7907; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13725 = _T_11273 & _T_6309; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_9_6 = _T_13725 | _T_7916; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13742 = _T_11290 & _T_6309; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_9_7 = _T_13742 | _T_7925; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13759 = _T_11307 & _T_6309; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_9_8 = _T_13759 | _T_7934; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13776 = _T_11324 & _T_6309; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_9_9 = _T_13776 | _T_7943; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13793 = _T_11341 & _T_6309; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_9_10 = _T_13793 | _T_7952; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13810 = _T_11358 & _T_6309; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_9_11 = _T_13810 | _T_7961; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13827 = _T_11375 & _T_6309; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_9_12 = _T_13827 | _T_7970; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13844 = _T_11392 & _T_6309; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_9_13 = _T_13844 | _T_7979; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13861 = _T_11409 & _T_6309; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_9_14 = _T_13861 | _T_7988; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13878 = _T_11426 & _T_6309; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_9_15 = _T_13878 | _T_7997; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13895 = _T_11171 & _T_6320; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_10_0 = _T_13895 | _T_8006; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13912 = _T_11188 & _T_6320; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_10_1 = _T_13912 | _T_8015; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13929 = _T_11205 & _T_6320; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_10_2 = _T_13929 | _T_8024; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13946 = _T_11222 & _T_6320; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_10_3 = _T_13946 | _T_8033; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13963 = _T_11239 & _T_6320; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_10_4 = _T_13963 | _T_8042; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13980 = _T_11256 & _T_6320; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_10_5 = _T_13980 | _T_8051; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13997 = _T_11273 & _T_6320; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_10_6 = _T_13997 | _T_8060; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14014 = _T_11290 & _T_6320; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_10_7 = _T_14014 | _T_8069; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14031 = _T_11307 & _T_6320; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_10_8 = _T_14031 | _T_8078; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14048 = _T_11324 & _T_6320; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_10_9 = _T_14048 | _T_8087; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14065 = _T_11341 & _T_6320; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_10_10 = _T_14065 | _T_8096; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14082 = _T_11358 & _T_6320; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_10_11 = _T_14082 | _T_8105; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14099 = _T_11375 & _T_6320; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_10_12 = _T_14099 | _T_8114; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14116 = _T_11392 & _T_6320; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_10_13 = _T_14116 | _T_8123; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14133 = _T_11409 & _T_6320; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_10_14 = _T_14133 | _T_8132; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14150 = _T_11426 & _T_6320; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_10_15 = _T_14150 | _T_8141; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14167 = _T_11171 & _T_6331; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_11_0 = _T_14167 | _T_8150; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14184 = _T_11188 & _T_6331; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_11_1 = _T_14184 | _T_8159; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14201 = _T_11205 & _T_6331; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_11_2 = _T_14201 | _T_8168; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14218 = _T_11222 & _T_6331; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_11_3 = _T_14218 | _T_8177; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14235 = _T_11239 & _T_6331; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_11_4 = _T_14235 | _T_8186; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14252 = _T_11256 & _T_6331; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_11_5 = _T_14252 | _T_8195; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14269 = _T_11273 & _T_6331; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_11_6 = _T_14269 | _T_8204; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14286 = _T_11290 & _T_6331; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_11_7 = _T_14286 | _T_8213; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14303 = _T_11307 & _T_6331; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_11_8 = _T_14303 | _T_8222; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14320 = _T_11324 & _T_6331; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_11_9 = _T_14320 | _T_8231; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14337 = _T_11341 & _T_6331; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_11_10 = _T_14337 | _T_8240; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14354 = _T_11358 & _T_6331; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_11_11 = _T_14354 | _T_8249; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14371 = _T_11375 & _T_6331; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_11_12 = _T_14371 | _T_8258; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14388 = _T_11392 & _T_6331; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_11_13 = _T_14388 | _T_8267; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14405 = _T_11409 & _T_6331; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_11_14 = _T_14405 | _T_8276; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14422 = _T_11426 & _T_6331; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_11_15 = _T_14422 | _T_8285; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14439 = _T_11171 & _T_6342; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_12_0 = _T_14439 | _T_8294; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14456 = _T_11188 & _T_6342; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_12_1 = _T_14456 | _T_8303; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14473 = _T_11205 & _T_6342; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_12_2 = _T_14473 | _T_8312; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14490 = _T_11222 & _T_6342; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_12_3 = _T_14490 | _T_8321; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14507 = _T_11239 & _T_6342; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_12_4 = _T_14507 | _T_8330; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14524 = _T_11256 & _T_6342; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_12_5 = _T_14524 | _T_8339; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14541 = _T_11273 & _T_6342; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_12_6 = _T_14541 | _T_8348; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14558 = _T_11290 & _T_6342; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_12_7 = _T_14558 | _T_8357; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14575 = _T_11307 & _T_6342; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_12_8 = _T_14575 | _T_8366; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14592 = _T_11324 & _T_6342; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_12_9 = _T_14592 | _T_8375; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14609 = _T_11341 & _T_6342; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_12_10 = _T_14609 | _T_8384; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14626 = _T_11358 & _T_6342; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_12_11 = _T_14626 | _T_8393; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14643 = _T_11375 & _T_6342; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_12_12 = _T_14643 | _T_8402; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14660 = _T_11392 & _T_6342; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_12_13 = _T_14660 | _T_8411; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14677 = _T_11409 & _T_6342; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_12_14 = _T_14677 | _T_8420; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14694 = _T_11426 & _T_6342; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_12_15 = _T_14694 | _T_8429; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14711 = _T_11171 & _T_6353; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_13_0 = _T_14711 | _T_8438; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14728 = _T_11188 & _T_6353; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_13_1 = _T_14728 | _T_8447; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14745 = _T_11205 & _T_6353; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_13_2 = _T_14745 | _T_8456; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14762 = _T_11222 & _T_6353; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_13_3 = _T_14762 | _T_8465; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14779 = _T_11239 & _T_6353; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_13_4 = _T_14779 | _T_8474; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14796 = _T_11256 & _T_6353; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_13_5 = _T_14796 | _T_8483; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14813 = _T_11273 & _T_6353; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_13_6 = _T_14813 | _T_8492; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14830 = _T_11290 & _T_6353; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_13_7 = _T_14830 | _T_8501; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14847 = _T_11307 & _T_6353; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_13_8 = _T_14847 | _T_8510; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14864 = _T_11324 & _T_6353; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_13_9 = _T_14864 | _T_8519; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14881 = _T_11341 & _T_6353; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_13_10 = _T_14881 | _T_8528; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14898 = _T_11358 & _T_6353; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_13_11 = _T_14898 | _T_8537; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14915 = _T_11375 & _T_6353; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_13_12 = _T_14915 | _T_8546; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14932 = _T_11392 & _T_6353; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_13_13 = _T_14932 | _T_8555; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14949 = _T_11409 & _T_6353; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_13_14 = _T_14949 | _T_8564; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14966 = _T_11426 & _T_6353; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_13_15 = _T_14966 | _T_8573; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14983 = _T_11171 & _T_6364; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_14_0 = _T_14983 | _T_8582; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15000 = _T_11188 & _T_6364; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_14_1 = _T_15000 | _T_8591; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15017 = _T_11205 & _T_6364; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_14_2 = _T_15017 | _T_8600; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15034 = _T_11222 & _T_6364; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_14_3 = _T_15034 | _T_8609; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15051 = _T_11239 & _T_6364; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_14_4 = _T_15051 | _T_8618; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15068 = _T_11256 & _T_6364; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_14_5 = _T_15068 | _T_8627; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15085 = _T_11273 & _T_6364; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_14_6 = _T_15085 | _T_8636; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15102 = _T_11290 & _T_6364; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_14_7 = _T_15102 | _T_8645; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15119 = _T_11307 & _T_6364; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_14_8 = _T_15119 | _T_8654; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15136 = _T_11324 & _T_6364; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_14_9 = _T_15136 | _T_8663; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15153 = _T_11341 & _T_6364; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_14_10 = _T_15153 | _T_8672; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15170 = _T_11358 & _T_6364; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_14_11 = _T_15170 | _T_8681; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15187 = _T_11375 & _T_6364; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_14_12 = _T_15187 | _T_8690; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15204 = _T_11392 & _T_6364; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_14_13 = _T_15204 | _T_8699; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15221 = _T_11409 & _T_6364; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_14_14 = _T_15221 | _T_8708; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15238 = _T_11426 & _T_6364; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_14_15 = _T_15238 | _T_8717; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15255 = _T_11171 & _T_6375; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_15_0 = _T_15255 | _T_8726; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15272 = _T_11188 & _T_6375; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_15_1 = _T_15272 | _T_8735; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15289 = _T_11205 & _T_6375; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_15_2 = _T_15289 | _T_8744; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15306 = _T_11222 & _T_6375; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_15_3 = _T_15306 | _T_8753; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15323 = _T_11239 & _T_6375; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_15_4 = _T_15323 | _T_8762; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15340 = _T_11256 & _T_6375; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_15_5 = _T_15340 | _T_8771; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15357 = _T_11273 & _T_6375; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_15_6 = _T_15357 | _T_8780; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15374 = _T_11290 & _T_6375; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_15_7 = _T_15374 | _T_8789; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15391 = _T_11307 & _T_6375; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_15_8 = _T_15391 | _T_8798; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15408 = _T_11324 & _T_6375; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_15_9 = _T_15408 | _T_8807; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15425 = _T_11341 & _T_6375; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_15_10 = _T_15425 | _T_8816; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15442 = _T_11358 & _T_6375; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_15_11 = _T_15442 | _T_8825; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15459 = _T_11375 & _T_6375; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_15_12 = _T_15459 | _T_8834; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15476 = _T_11392 & _T_6375; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_15_13 = _T_15476 | _T_8843; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15493 = _T_11409 & _T_6375; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_15_14 = _T_15493 | _T_8852; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15510 = _T_11426 & _T_6375; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_15_15 = _T_15510 | _T_8861; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15523 = bht_wr_en0[1] & _T_11170; // @[ifu_bp_ctl.scala 443:45]
  wire  _T_15527 = _T_15523 & _T_6210; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_0_0 = _T_15527 | _T_8870; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15540 = bht_wr_en0[1] & _T_11187; // @[ifu_bp_ctl.scala 443:45]
  wire  _T_15544 = _T_15540 & _T_6210; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_0_1 = _T_15544 | _T_8879; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15557 = bht_wr_en0[1] & _T_11204; // @[ifu_bp_ctl.scala 443:45]
  wire  _T_15561 = _T_15557 & _T_6210; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_0_2 = _T_15561 | _T_8888; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15574 = bht_wr_en0[1] & _T_11221; // @[ifu_bp_ctl.scala 443:45]
  wire  _T_15578 = _T_15574 & _T_6210; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_0_3 = _T_15578 | _T_8897; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15591 = bht_wr_en0[1] & _T_11238; // @[ifu_bp_ctl.scala 443:45]
  wire  _T_15595 = _T_15591 & _T_6210; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_0_4 = _T_15595 | _T_8906; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15608 = bht_wr_en0[1] & _T_11255; // @[ifu_bp_ctl.scala 443:45]
  wire  _T_15612 = _T_15608 & _T_6210; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_0_5 = _T_15612 | _T_8915; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15625 = bht_wr_en0[1] & _T_11272; // @[ifu_bp_ctl.scala 443:45]
  wire  _T_15629 = _T_15625 & _T_6210; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_0_6 = _T_15629 | _T_8924; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15642 = bht_wr_en0[1] & _T_11289; // @[ifu_bp_ctl.scala 443:45]
  wire  _T_15646 = _T_15642 & _T_6210; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_0_7 = _T_15646 | _T_8933; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15659 = bht_wr_en0[1] & _T_11306; // @[ifu_bp_ctl.scala 443:45]
  wire  _T_15663 = _T_15659 & _T_6210; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_0_8 = _T_15663 | _T_8942; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15676 = bht_wr_en0[1] & _T_11323; // @[ifu_bp_ctl.scala 443:45]
  wire  _T_15680 = _T_15676 & _T_6210; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_0_9 = _T_15680 | _T_8951; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15693 = bht_wr_en0[1] & _T_11340; // @[ifu_bp_ctl.scala 443:45]
  wire  _T_15697 = _T_15693 & _T_6210; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_0_10 = _T_15697 | _T_8960; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15710 = bht_wr_en0[1] & _T_11357; // @[ifu_bp_ctl.scala 443:45]
  wire  _T_15714 = _T_15710 & _T_6210; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_0_11 = _T_15714 | _T_8969; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15727 = bht_wr_en0[1] & _T_11374; // @[ifu_bp_ctl.scala 443:45]
  wire  _T_15731 = _T_15727 & _T_6210; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_0_12 = _T_15731 | _T_8978; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15744 = bht_wr_en0[1] & _T_11391; // @[ifu_bp_ctl.scala 443:45]
  wire  _T_15748 = _T_15744 & _T_6210; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_0_13 = _T_15748 | _T_8987; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15761 = bht_wr_en0[1] & _T_11408; // @[ifu_bp_ctl.scala 443:45]
  wire  _T_15765 = _T_15761 & _T_6210; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_0_14 = _T_15765 | _T_8996; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15778 = bht_wr_en0[1] & _T_11425; // @[ifu_bp_ctl.scala 443:45]
  wire  _T_15782 = _T_15778 & _T_6210; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_0_15 = _T_15782 | _T_9005; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15799 = _T_15523 & _T_6221; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_1_0 = _T_15799 | _T_9014; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15816 = _T_15540 & _T_6221; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_1_1 = _T_15816 | _T_9023; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15833 = _T_15557 & _T_6221; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_1_2 = _T_15833 | _T_9032; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15850 = _T_15574 & _T_6221; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_1_3 = _T_15850 | _T_9041; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15867 = _T_15591 & _T_6221; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_1_4 = _T_15867 | _T_9050; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15884 = _T_15608 & _T_6221; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_1_5 = _T_15884 | _T_9059; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15901 = _T_15625 & _T_6221; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_1_6 = _T_15901 | _T_9068; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15918 = _T_15642 & _T_6221; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_1_7 = _T_15918 | _T_9077; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15935 = _T_15659 & _T_6221; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_1_8 = _T_15935 | _T_9086; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15952 = _T_15676 & _T_6221; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_1_9 = _T_15952 | _T_9095; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15969 = _T_15693 & _T_6221; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_1_10 = _T_15969 | _T_9104; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15986 = _T_15710 & _T_6221; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_1_11 = _T_15986 | _T_9113; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16003 = _T_15727 & _T_6221; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_1_12 = _T_16003 | _T_9122; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16020 = _T_15744 & _T_6221; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_1_13 = _T_16020 | _T_9131; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16037 = _T_15761 & _T_6221; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_1_14 = _T_16037 | _T_9140; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16054 = _T_15778 & _T_6221; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_1_15 = _T_16054 | _T_9149; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16071 = _T_15523 & _T_6232; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_2_0 = _T_16071 | _T_9158; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16088 = _T_15540 & _T_6232; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_2_1 = _T_16088 | _T_9167; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16105 = _T_15557 & _T_6232; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_2_2 = _T_16105 | _T_9176; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16122 = _T_15574 & _T_6232; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_2_3 = _T_16122 | _T_9185; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16139 = _T_15591 & _T_6232; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_2_4 = _T_16139 | _T_9194; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16156 = _T_15608 & _T_6232; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_2_5 = _T_16156 | _T_9203; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16173 = _T_15625 & _T_6232; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_2_6 = _T_16173 | _T_9212; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16190 = _T_15642 & _T_6232; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_2_7 = _T_16190 | _T_9221; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16207 = _T_15659 & _T_6232; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_2_8 = _T_16207 | _T_9230; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16224 = _T_15676 & _T_6232; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_2_9 = _T_16224 | _T_9239; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16241 = _T_15693 & _T_6232; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_2_10 = _T_16241 | _T_9248; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16258 = _T_15710 & _T_6232; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_2_11 = _T_16258 | _T_9257; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16275 = _T_15727 & _T_6232; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_2_12 = _T_16275 | _T_9266; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16292 = _T_15744 & _T_6232; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_2_13 = _T_16292 | _T_9275; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16309 = _T_15761 & _T_6232; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_2_14 = _T_16309 | _T_9284; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16326 = _T_15778 & _T_6232; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_2_15 = _T_16326 | _T_9293; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16343 = _T_15523 & _T_6243; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_3_0 = _T_16343 | _T_9302; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16360 = _T_15540 & _T_6243; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_3_1 = _T_16360 | _T_9311; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16377 = _T_15557 & _T_6243; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_3_2 = _T_16377 | _T_9320; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16394 = _T_15574 & _T_6243; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_3_3 = _T_16394 | _T_9329; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16411 = _T_15591 & _T_6243; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_3_4 = _T_16411 | _T_9338; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16428 = _T_15608 & _T_6243; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_3_5 = _T_16428 | _T_9347; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16445 = _T_15625 & _T_6243; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_3_6 = _T_16445 | _T_9356; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16462 = _T_15642 & _T_6243; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_3_7 = _T_16462 | _T_9365; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16479 = _T_15659 & _T_6243; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_3_8 = _T_16479 | _T_9374; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16496 = _T_15676 & _T_6243; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_3_9 = _T_16496 | _T_9383; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16513 = _T_15693 & _T_6243; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_3_10 = _T_16513 | _T_9392; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16530 = _T_15710 & _T_6243; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_3_11 = _T_16530 | _T_9401; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16547 = _T_15727 & _T_6243; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_3_12 = _T_16547 | _T_9410; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16564 = _T_15744 & _T_6243; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_3_13 = _T_16564 | _T_9419; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16581 = _T_15761 & _T_6243; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_3_14 = _T_16581 | _T_9428; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16598 = _T_15778 & _T_6243; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_3_15 = _T_16598 | _T_9437; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16615 = _T_15523 & _T_6254; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_4_0 = _T_16615 | _T_9446; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16632 = _T_15540 & _T_6254; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_4_1 = _T_16632 | _T_9455; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16649 = _T_15557 & _T_6254; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_4_2 = _T_16649 | _T_9464; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16666 = _T_15574 & _T_6254; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_4_3 = _T_16666 | _T_9473; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16683 = _T_15591 & _T_6254; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_4_4 = _T_16683 | _T_9482; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16700 = _T_15608 & _T_6254; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_4_5 = _T_16700 | _T_9491; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16717 = _T_15625 & _T_6254; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_4_6 = _T_16717 | _T_9500; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16734 = _T_15642 & _T_6254; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_4_7 = _T_16734 | _T_9509; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16751 = _T_15659 & _T_6254; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_4_8 = _T_16751 | _T_9518; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16768 = _T_15676 & _T_6254; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_4_9 = _T_16768 | _T_9527; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16785 = _T_15693 & _T_6254; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_4_10 = _T_16785 | _T_9536; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16802 = _T_15710 & _T_6254; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_4_11 = _T_16802 | _T_9545; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16819 = _T_15727 & _T_6254; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_4_12 = _T_16819 | _T_9554; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16836 = _T_15744 & _T_6254; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_4_13 = _T_16836 | _T_9563; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16853 = _T_15761 & _T_6254; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_4_14 = _T_16853 | _T_9572; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16870 = _T_15778 & _T_6254; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_4_15 = _T_16870 | _T_9581; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16887 = _T_15523 & _T_6265; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_5_0 = _T_16887 | _T_9590; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16904 = _T_15540 & _T_6265; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_5_1 = _T_16904 | _T_9599; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16921 = _T_15557 & _T_6265; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_5_2 = _T_16921 | _T_9608; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16938 = _T_15574 & _T_6265; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_5_3 = _T_16938 | _T_9617; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16955 = _T_15591 & _T_6265; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_5_4 = _T_16955 | _T_9626; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16972 = _T_15608 & _T_6265; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_5_5 = _T_16972 | _T_9635; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16989 = _T_15625 & _T_6265; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_5_6 = _T_16989 | _T_9644; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17006 = _T_15642 & _T_6265; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_5_7 = _T_17006 | _T_9653; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17023 = _T_15659 & _T_6265; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_5_8 = _T_17023 | _T_9662; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17040 = _T_15676 & _T_6265; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_5_9 = _T_17040 | _T_9671; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17057 = _T_15693 & _T_6265; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_5_10 = _T_17057 | _T_9680; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17074 = _T_15710 & _T_6265; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_5_11 = _T_17074 | _T_9689; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17091 = _T_15727 & _T_6265; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_5_12 = _T_17091 | _T_9698; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17108 = _T_15744 & _T_6265; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_5_13 = _T_17108 | _T_9707; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17125 = _T_15761 & _T_6265; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_5_14 = _T_17125 | _T_9716; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17142 = _T_15778 & _T_6265; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_5_15 = _T_17142 | _T_9725; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17159 = _T_15523 & _T_6276; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_6_0 = _T_17159 | _T_9734; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17176 = _T_15540 & _T_6276; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_6_1 = _T_17176 | _T_9743; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17193 = _T_15557 & _T_6276; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_6_2 = _T_17193 | _T_9752; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17210 = _T_15574 & _T_6276; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_6_3 = _T_17210 | _T_9761; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17227 = _T_15591 & _T_6276; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_6_4 = _T_17227 | _T_9770; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17244 = _T_15608 & _T_6276; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_6_5 = _T_17244 | _T_9779; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17261 = _T_15625 & _T_6276; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_6_6 = _T_17261 | _T_9788; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17278 = _T_15642 & _T_6276; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_6_7 = _T_17278 | _T_9797; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17295 = _T_15659 & _T_6276; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_6_8 = _T_17295 | _T_9806; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17312 = _T_15676 & _T_6276; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_6_9 = _T_17312 | _T_9815; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17329 = _T_15693 & _T_6276; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_6_10 = _T_17329 | _T_9824; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17346 = _T_15710 & _T_6276; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_6_11 = _T_17346 | _T_9833; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17363 = _T_15727 & _T_6276; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_6_12 = _T_17363 | _T_9842; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17380 = _T_15744 & _T_6276; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_6_13 = _T_17380 | _T_9851; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17397 = _T_15761 & _T_6276; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_6_14 = _T_17397 | _T_9860; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17414 = _T_15778 & _T_6276; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_6_15 = _T_17414 | _T_9869; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17431 = _T_15523 & _T_6287; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_7_0 = _T_17431 | _T_9878; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17448 = _T_15540 & _T_6287; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_7_1 = _T_17448 | _T_9887; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17465 = _T_15557 & _T_6287; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_7_2 = _T_17465 | _T_9896; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17482 = _T_15574 & _T_6287; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_7_3 = _T_17482 | _T_9905; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17499 = _T_15591 & _T_6287; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_7_4 = _T_17499 | _T_9914; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17516 = _T_15608 & _T_6287; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_7_5 = _T_17516 | _T_9923; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17533 = _T_15625 & _T_6287; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_7_6 = _T_17533 | _T_9932; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17550 = _T_15642 & _T_6287; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_7_7 = _T_17550 | _T_9941; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17567 = _T_15659 & _T_6287; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_7_8 = _T_17567 | _T_9950; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17584 = _T_15676 & _T_6287; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_7_9 = _T_17584 | _T_9959; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17601 = _T_15693 & _T_6287; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_7_10 = _T_17601 | _T_9968; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17618 = _T_15710 & _T_6287; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_7_11 = _T_17618 | _T_9977; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17635 = _T_15727 & _T_6287; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_7_12 = _T_17635 | _T_9986; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17652 = _T_15744 & _T_6287; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_7_13 = _T_17652 | _T_9995; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17669 = _T_15761 & _T_6287; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_7_14 = _T_17669 | _T_10004; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17686 = _T_15778 & _T_6287; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_7_15 = _T_17686 | _T_10013; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17703 = _T_15523 & _T_6298; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_8_0 = _T_17703 | _T_10022; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17720 = _T_15540 & _T_6298; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_8_1 = _T_17720 | _T_10031; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17737 = _T_15557 & _T_6298; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_8_2 = _T_17737 | _T_10040; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17754 = _T_15574 & _T_6298; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_8_3 = _T_17754 | _T_10049; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17771 = _T_15591 & _T_6298; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_8_4 = _T_17771 | _T_10058; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17788 = _T_15608 & _T_6298; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_8_5 = _T_17788 | _T_10067; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17805 = _T_15625 & _T_6298; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_8_6 = _T_17805 | _T_10076; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17822 = _T_15642 & _T_6298; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_8_7 = _T_17822 | _T_10085; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17839 = _T_15659 & _T_6298; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_8_8 = _T_17839 | _T_10094; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17856 = _T_15676 & _T_6298; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_8_9 = _T_17856 | _T_10103; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17873 = _T_15693 & _T_6298; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_8_10 = _T_17873 | _T_10112; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17890 = _T_15710 & _T_6298; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_8_11 = _T_17890 | _T_10121; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17907 = _T_15727 & _T_6298; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_8_12 = _T_17907 | _T_10130; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17924 = _T_15744 & _T_6298; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_8_13 = _T_17924 | _T_10139; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17941 = _T_15761 & _T_6298; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_8_14 = _T_17941 | _T_10148; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17958 = _T_15778 & _T_6298; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_8_15 = _T_17958 | _T_10157; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17975 = _T_15523 & _T_6309; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_9_0 = _T_17975 | _T_10166; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17992 = _T_15540 & _T_6309; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_9_1 = _T_17992 | _T_10175; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18009 = _T_15557 & _T_6309; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_9_2 = _T_18009 | _T_10184; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18026 = _T_15574 & _T_6309; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_9_3 = _T_18026 | _T_10193; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18043 = _T_15591 & _T_6309; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_9_4 = _T_18043 | _T_10202; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18060 = _T_15608 & _T_6309; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_9_5 = _T_18060 | _T_10211; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18077 = _T_15625 & _T_6309; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_9_6 = _T_18077 | _T_10220; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18094 = _T_15642 & _T_6309; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_9_7 = _T_18094 | _T_10229; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18111 = _T_15659 & _T_6309; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_9_8 = _T_18111 | _T_10238; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18128 = _T_15676 & _T_6309; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_9_9 = _T_18128 | _T_10247; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18145 = _T_15693 & _T_6309; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_9_10 = _T_18145 | _T_10256; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18162 = _T_15710 & _T_6309; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_9_11 = _T_18162 | _T_10265; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18179 = _T_15727 & _T_6309; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_9_12 = _T_18179 | _T_10274; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18196 = _T_15744 & _T_6309; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_9_13 = _T_18196 | _T_10283; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18213 = _T_15761 & _T_6309; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_9_14 = _T_18213 | _T_10292; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18230 = _T_15778 & _T_6309; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_9_15 = _T_18230 | _T_10301; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18247 = _T_15523 & _T_6320; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_10_0 = _T_18247 | _T_10310; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18264 = _T_15540 & _T_6320; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_10_1 = _T_18264 | _T_10319; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18281 = _T_15557 & _T_6320; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_10_2 = _T_18281 | _T_10328; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18298 = _T_15574 & _T_6320; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_10_3 = _T_18298 | _T_10337; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18315 = _T_15591 & _T_6320; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_10_4 = _T_18315 | _T_10346; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18332 = _T_15608 & _T_6320; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_10_5 = _T_18332 | _T_10355; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18349 = _T_15625 & _T_6320; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_10_6 = _T_18349 | _T_10364; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18366 = _T_15642 & _T_6320; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_10_7 = _T_18366 | _T_10373; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18383 = _T_15659 & _T_6320; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_10_8 = _T_18383 | _T_10382; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18400 = _T_15676 & _T_6320; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_10_9 = _T_18400 | _T_10391; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18417 = _T_15693 & _T_6320; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_10_10 = _T_18417 | _T_10400; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18434 = _T_15710 & _T_6320; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_10_11 = _T_18434 | _T_10409; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18451 = _T_15727 & _T_6320; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_10_12 = _T_18451 | _T_10418; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18468 = _T_15744 & _T_6320; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_10_13 = _T_18468 | _T_10427; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18485 = _T_15761 & _T_6320; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_10_14 = _T_18485 | _T_10436; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18502 = _T_15778 & _T_6320; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_10_15 = _T_18502 | _T_10445; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18519 = _T_15523 & _T_6331; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_11_0 = _T_18519 | _T_10454; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18536 = _T_15540 & _T_6331; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_11_1 = _T_18536 | _T_10463; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18553 = _T_15557 & _T_6331; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_11_2 = _T_18553 | _T_10472; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18570 = _T_15574 & _T_6331; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_11_3 = _T_18570 | _T_10481; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18587 = _T_15591 & _T_6331; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_11_4 = _T_18587 | _T_10490; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18604 = _T_15608 & _T_6331; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_11_5 = _T_18604 | _T_10499; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18621 = _T_15625 & _T_6331; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_11_6 = _T_18621 | _T_10508; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18638 = _T_15642 & _T_6331; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_11_7 = _T_18638 | _T_10517; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18655 = _T_15659 & _T_6331; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_11_8 = _T_18655 | _T_10526; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18672 = _T_15676 & _T_6331; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_11_9 = _T_18672 | _T_10535; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18689 = _T_15693 & _T_6331; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_11_10 = _T_18689 | _T_10544; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18706 = _T_15710 & _T_6331; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_11_11 = _T_18706 | _T_10553; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18723 = _T_15727 & _T_6331; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_11_12 = _T_18723 | _T_10562; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18740 = _T_15744 & _T_6331; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_11_13 = _T_18740 | _T_10571; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18757 = _T_15761 & _T_6331; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_11_14 = _T_18757 | _T_10580; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18774 = _T_15778 & _T_6331; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_11_15 = _T_18774 | _T_10589; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18791 = _T_15523 & _T_6342; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_12_0 = _T_18791 | _T_10598; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18808 = _T_15540 & _T_6342; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_12_1 = _T_18808 | _T_10607; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18825 = _T_15557 & _T_6342; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_12_2 = _T_18825 | _T_10616; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18842 = _T_15574 & _T_6342; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_12_3 = _T_18842 | _T_10625; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18859 = _T_15591 & _T_6342; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_12_4 = _T_18859 | _T_10634; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18876 = _T_15608 & _T_6342; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_12_5 = _T_18876 | _T_10643; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18893 = _T_15625 & _T_6342; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_12_6 = _T_18893 | _T_10652; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18910 = _T_15642 & _T_6342; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_12_7 = _T_18910 | _T_10661; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18927 = _T_15659 & _T_6342; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_12_8 = _T_18927 | _T_10670; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18944 = _T_15676 & _T_6342; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_12_9 = _T_18944 | _T_10679; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18961 = _T_15693 & _T_6342; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_12_10 = _T_18961 | _T_10688; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18978 = _T_15710 & _T_6342; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_12_11 = _T_18978 | _T_10697; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18995 = _T_15727 & _T_6342; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_12_12 = _T_18995 | _T_10706; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_19012 = _T_15744 & _T_6342; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_12_13 = _T_19012 | _T_10715; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_19029 = _T_15761 & _T_6342; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_12_14 = _T_19029 | _T_10724; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_19046 = _T_15778 & _T_6342; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_12_15 = _T_19046 | _T_10733; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_19063 = _T_15523 & _T_6353; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_13_0 = _T_19063 | _T_10742; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_19080 = _T_15540 & _T_6353; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_13_1 = _T_19080 | _T_10751; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_19097 = _T_15557 & _T_6353; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_13_2 = _T_19097 | _T_10760; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_19114 = _T_15574 & _T_6353; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_13_3 = _T_19114 | _T_10769; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_19131 = _T_15591 & _T_6353; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_13_4 = _T_19131 | _T_10778; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_19148 = _T_15608 & _T_6353; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_13_5 = _T_19148 | _T_10787; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_19165 = _T_15625 & _T_6353; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_13_6 = _T_19165 | _T_10796; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_19182 = _T_15642 & _T_6353; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_13_7 = _T_19182 | _T_10805; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_19199 = _T_15659 & _T_6353; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_13_8 = _T_19199 | _T_10814; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_19216 = _T_15676 & _T_6353; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_13_9 = _T_19216 | _T_10823; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_19233 = _T_15693 & _T_6353; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_13_10 = _T_19233 | _T_10832; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_19250 = _T_15710 & _T_6353; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_13_11 = _T_19250 | _T_10841; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_19267 = _T_15727 & _T_6353; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_13_12 = _T_19267 | _T_10850; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_19284 = _T_15744 & _T_6353; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_13_13 = _T_19284 | _T_10859; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_19301 = _T_15761 & _T_6353; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_13_14 = _T_19301 | _T_10868; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_19318 = _T_15778 & _T_6353; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_13_15 = _T_19318 | _T_10877; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_19335 = _T_15523 & _T_6364; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_14_0 = _T_19335 | _T_10886; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_19352 = _T_15540 & _T_6364; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_14_1 = _T_19352 | _T_10895; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_19369 = _T_15557 & _T_6364; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_14_2 = _T_19369 | _T_10904; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_19386 = _T_15574 & _T_6364; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_14_3 = _T_19386 | _T_10913; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_19403 = _T_15591 & _T_6364; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_14_4 = _T_19403 | _T_10922; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_19420 = _T_15608 & _T_6364; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_14_5 = _T_19420 | _T_10931; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_19437 = _T_15625 & _T_6364; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_14_6 = _T_19437 | _T_10940; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_19454 = _T_15642 & _T_6364; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_14_7 = _T_19454 | _T_10949; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_19471 = _T_15659 & _T_6364; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_14_8 = _T_19471 | _T_10958; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_19488 = _T_15676 & _T_6364; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_14_9 = _T_19488 | _T_10967; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_19505 = _T_15693 & _T_6364; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_14_10 = _T_19505 | _T_10976; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_19522 = _T_15710 & _T_6364; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_14_11 = _T_19522 | _T_10985; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_19539 = _T_15727 & _T_6364; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_14_12 = _T_19539 | _T_10994; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_19556 = _T_15744 & _T_6364; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_14_13 = _T_19556 | _T_11003; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_19573 = _T_15761 & _T_6364; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_14_14 = _T_19573 | _T_11012; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_19590 = _T_15778 & _T_6364; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_14_15 = _T_19590 | _T_11021; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_19607 = _T_15523 & _T_6375; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_15_0 = _T_19607 | _T_11030; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_19624 = _T_15540 & _T_6375; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_15_1 = _T_19624 | _T_11039; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_19641 = _T_15557 & _T_6375; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_15_2 = _T_19641 | _T_11048; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_19658 = _T_15574 & _T_6375; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_15_3 = _T_19658 | _T_11057; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_19675 = _T_15591 & _T_6375; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_15_4 = _T_19675 | _T_11066; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_19692 = _T_15608 & _T_6375; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_15_5 = _T_19692 | _T_11075; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_19709 = _T_15625 & _T_6375; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_15_6 = _T_19709 | _T_11084; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_19726 = _T_15642 & _T_6375; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_15_7 = _T_19726 | _T_11093; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_19743 = _T_15659 & _T_6375; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_15_8 = _T_19743 | _T_11102; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_19760 = _T_15676 & _T_6375; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_15_9 = _T_19760 | _T_11111; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_19777 = _T_15693 & _T_6375; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_15_10 = _T_19777 | _T_11120; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_19794 = _T_15710 & _T_6375; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_15_11 = _T_19794 | _T_11129; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_19811 = _T_15727 & _T_6375; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_15_12 = _T_19811 | _T_11138; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_19828 = _T_15744 & _T_6375; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_15_13 = _T_19828 | _T_11147; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_19845 = _T_15761 & _T_6375; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_15_14 = _T_19845 | _T_11156; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_19862 = _T_15778 & _T_6375; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_15_15 = _T_19862 | _T_11165; // @[ifu_bp_ctl.scala 443:223]
  rvclkhdr rvclkhdr ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_io_l1clk),
    .io_clk(rvclkhdr_io_clk),
    .io_en(rvclkhdr_io_en),
    .io_scan_mode(rvclkhdr_io_scan_mode)
  );
  rvclkhdr rvclkhdr_1 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_1_io_l1clk),
    .io_clk(rvclkhdr_1_io_clk),
    .io_en(rvclkhdr_1_io_en),
    .io_scan_mode(rvclkhdr_1_io_scan_mode)
  );
  rvclkhdr rvclkhdr_2 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_2_io_l1clk),
    .io_clk(rvclkhdr_2_io_clk),
    .io_en(rvclkhdr_2_io_en),
    .io_scan_mode(rvclkhdr_2_io_scan_mode)
  );
  rvclkhdr rvclkhdr_3 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_3_io_l1clk),
    .io_clk(rvclkhdr_3_io_clk),
    .io_en(rvclkhdr_3_io_en),
    .io_scan_mode(rvclkhdr_3_io_scan_mode)
  );
  rvclkhdr rvclkhdr_4 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_4_io_l1clk),
    .io_clk(rvclkhdr_4_io_clk),
    .io_en(rvclkhdr_4_io_en),
    .io_scan_mode(rvclkhdr_4_io_scan_mode)
  );
  rvclkhdr rvclkhdr_5 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_5_io_l1clk),
    .io_clk(rvclkhdr_5_io_clk),
    .io_en(rvclkhdr_5_io_en),
    .io_scan_mode(rvclkhdr_5_io_scan_mode)
  );
  rvclkhdr rvclkhdr_6 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_6_io_l1clk),
    .io_clk(rvclkhdr_6_io_clk),
    .io_en(rvclkhdr_6_io_en),
    .io_scan_mode(rvclkhdr_6_io_scan_mode)
  );
  rvclkhdr rvclkhdr_7 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_7_io_l1clk),
    .io_clk(rvclkhdr_7_io_clk),
    .io_en(rvclkhdr_7_io_en),
    .io_scan_mode(rvclkhdr_7_io_scan_mode)
  );
  rvclkhdr rvclkhdr_8 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_8_io_l1clk),
    .io_clk(rvclkhdr_8_io_clk),
    .io_en(rvclkhdr_8_io_en),
    .io_scan_mode(rvclkhdr_8_io_scan_mode)
  );
  rvclkhdr rvclkhdr_9 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_9_io_l1clk),
    .io_clk(rvclkhdr_9_io_clk),
    .io_en(rvclkhdr_9_io_en),
    .io_scan_mode(rvclkhdr_9_io_scan_mode)
  );
  rvclkhdr rvclkhdr_10 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_10_io_l1clk),
    .io_clk(rvclkhdr_10_io_clk),
    .io_en(rvclkhdr_10_io_en),
    .io_scan_mode(rvclkhdr_10_io_scan_mode)
  );
  rvclkhdr rvclkhdr_11 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_11_io_l1clk),
    .io_clk(rvclkhdr_11_io_clk),
    .io_en(rvclkhdr_11_io_en),
    .io_scan_mode(rvclkhdr_11_io_scan_mode)
  );
  rvclkhdr rvclkhdr_12 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_12_io_l1clk),
    .io_clk(rvclkhdr_12_io_clk),
    .io_en(rvclkhdr_12_io_en),
    .io_scan_mode(rvclkhdr_12_io_scan_mode)
  );
  rvclkhdr rvclkhdr_13 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_13_io_l1clk),
    .io_clk(rvclkhdr_13_io_clk),
    .io_en(rvclkhdr_13_io_en),
    .io_scan_mode(rvclkhdr_13_io_scan_mode)
  );
  rvclkhdr rvclkhdr_14 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_14_io_l1clk),
    .io_clk(rvclkhdr_14_io_clk),
    .io_en(rvclkhdr_14_io_en),
    .io_scan_mode(rvclkhdr_14_io_scan_mode)
  );
  rvclkhdr rvclkhdr_15 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_15_io_l1clk),
    .io_clk(rvclkhdr_15_io_clk),
    .io_en(rvclkhdr_15_io_en),
    .io_scan_mode(rvclkhdr_15_io_scan_mode)
  );
  rvclkhdr rvclkhdr_16 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_16_io_l1clk),
    .io_clk(rvclkhdr_16_io_clk),
    .io_en(rvclkhdr_16_io_en),
    .io_scan_mode(rvclkhdr_16_io_scan_mode)
  );
  rvclkhdr rvclkhdr_17 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_17_io_l1clk),
    .io_clk(rvclkhdr_17_io_clk),
    .io_en(rvclkhdr_17_io_en),
    .io_scan_mode(rvclkhdr_17_io_scan_mode)
  );
  rvclkhdr rvclkhdr_18 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_18_io_l1clk),
    .io_clk(rvclkhdr_18_io_clk),
    .io_en(rvclkhdr_18_io_en),
    .io_scan_mode(rvclkhdr_18_io_scan_mode)
  );
  rvclkhdr rvclkhdr_19 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_19_io_l1clk),
    .io_clk(rvclkhdr_19_io_clk),
    .io_en(rvclkhdr_19_io_en),
    .io_scan_mode(rvclkhdr_19_io_scan_mode)
  );
  rvclkhdr rvclkhdr_20 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_20_io_l1clk),
    .io_clk(rvclkhdr_20_io_clk),
    .io_en(rvclkhdr_20_io_en),
    .io_scan_mode(rvclkhdr_20_io_scan_mode)
  );
  rvclkhdr rvclkhdr_21 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_21_io_l1clk),
    .io_clk(rvclkhdr_21_io_clk),
    .io_en(rvclkhdr_21_io_en),
    .io_scan_mode(rvclkhdr_21_io_scan_mode)
  );
  rvclkhdr rvclkhdr_22 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_22_io_l1clk),
    .io_clk(rvclkhdr_22_io_clk),
    .io_en(rvclkhdr_22_io_en),
    .io_scan_mode(rvclkhdr_22_io_scan_mode)
  );
  rvclkhdr rvclkhdr_23 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_23_io_l1clk),
    .io_clk(rvclkhdr_23_io_clk),
    .io_en(rvclkhdr_23_io_en),
    .io_scan_mode(rvclkhdr_23_io_scan_mode)
  );
  rvclkhdr rvclkhdr_24 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_24_io_l1clk),
    .io_clk(rvclkhdr_24_io_clk),
    .io_en(rvclkhdr_24_io_en),
    .io_scan_mode(rvclkhdr_24_io_scan_mode)
  );
  rvclkhdr rvclkhdr_25 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_25_io_l1clk),
    .io_clk(rvclkhdr_25_io_clk),
    .io_en(rvclkhdr_25_io_en),
    .io_scan_mode(rvclkhdr_25_io_scan_mode)
  );
  rvclkhdr rvclkhdr_26 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_26_io_l1clk),
    .io_clk(rvclkhdr_26_io_clk),
    .io_en(rvclkhdr_26_io_en),
    .io_scan_mode(rvclkhdr_26_io_scan_mode)
  );
  rvclkhdr rvclkhdr_27 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_27_io_l1clk),
    .io_clk(rvclkhdr_27_io_clk),
    .io_en(rvclkhdr_27_io_en),
    .io_scan_mode(rvclkhdr_27_io_scan_mode)
  );
  rvclkhdr rvclkhdr_28 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_28_io_l1clk),
    .io_clk(rvclkhdr_28_io_clk),
    .io_en(rvclkhdr_28_io_en),
    .io_scan_mode(rvclkhdr_28_io_scan_mode)
  );
  rvclkhdr rvclkhdr_29 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_29_io_l1clk),
    .io_clk(rvclkhdr_29_io_clk),
    .io_en(rvclkhdr_29_io_en),
    .io_scan_mode(rvclkhdr_29_io_scan_mode)
  );
  rvclkhdr rvclkhdr_30 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_30_io_l1clk),
    .io_clk(rvclkhdr_30_io_clk),
    .io_en(rvclkhdr_30_io_en),
    .io_scan_mode(rvclkhdr_30_io_scan_mode)
  );
  rvclkhdr rvclkhdr_31 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_31_io_l1clk),
    .io_clk(rvclkhdr_31_io_clk),
    .io_en(rvclkhdr_31_io_en),
    .io_scan_mode(rvclkhdr_31_io_scan_mode)
  );
  rvclkhdr rvclkhdr_32 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_32_io_l1clk),
    .io_clk(rvclkhdr_32_io_clk),
    .io_en(rvclkhdr_32_io_en),
    .io_scan_mode(rvclkhdr_32_io_scan_mode)
  );
  rvclkhdr rvclkhdr_33 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_33_io_l1clk),
    .io_clk(rvclkhdr_33_io_clk),
    .io_en(rvclkhdr_33_io_en),
    .io_scan_mode(rvclkhdr_33_io_scan_mode)
  );
  rvclkhdr rvclkhdr_34 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_34_io_l1clk),
    .io_clk(rvclkhdr_34_io_clk),
    .io_en(rvclkhdr_34_io_en),
    .io_scan_mode(rvclkhdr_34_io_scan_mode)
  );
  rvclkhdr rvclkhdr_35 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_35_io_l1clk),
    .io_clk(rvclkhdr_35_io_clk),
    .io_en(rvclkhdr_35_io_en),
    .io_scan_mode(rvclkhdr_35_io_scan_mode)
  );
  rvclkhdr rvclkhdr_36 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_36_io_l1clk),
    .io_clk(rvclkhdr_36_io_clk),
    .io_en(rvclkhdr_36_io_en),
    .io_scan_mode(rvclkhdr_36_io_scan_mode)
  );
  rvclkhdr rvclkhdr_37 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_37_io_l1clk),
    .io_clk(rvclkhdr_37_io_clk),
    .io_en(rvclkhdr_37_io_en),
    .io_scan_mode(rvclkhdr_37_io_scan_mode)
  );
  rvclkhdr rvclkhdr_38 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_38_io_l1clk),
    .io_clk(rvclkhdr_38_io_clk),
    .io_en(rvclkhdr_38_io_en),
    .io_scan_mode(rvclkhdr_38_io_scan_mode)
  );
  rvclkhdr rvclkhdr_39 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_39_io_l1clk),
    .io_clk(rvclkhdr_39_io_clk),
    .io_en(rvclkhdr_39_io_en),
    .io_scan_mode(rvclkhdr_39_io_scan_mode)
  );
  rvclkhdr rvclkhdr_40 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_40_io_l1clk),
    .io_clk(rvclkhdr_40_io_clk),
    .io_en(rvclkhdr_40_io_en),
    .io_scan_mode(rvclkhdr_40_io_scan_mode)
  );
  rvclkhdr rvclkhdr_41 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_41_io_l1clk),
    .io_clk(rvclkhdr_41_io_clk),
    .io_en(rvclkhdr_41_io_en),
    .io_scan_mode(rvclkhdr_41_io_scan_mode)
  );
  rvclkhdr rvclkhdr_42 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_42_io_l1clk),
    .io_clk(rvclkhdr_42_io_clk),
    .io_en(rvclkhdr_42_io_en),
    .io_scan_mode(rvclkhdr_42_io_scan_mode)
  );
  rvclkhdr rvclkhdr_43 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_43_io_l1clk),
    .io_clk(rvclkhdr_43_io_clk),
    .io_en(rvclkhdr_43_io_en),
    .io_scan_mode(rvclkhdr_43_io_scan_mode)
  );
  rvclkhdr rvclkhdr_44 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_44_io_l1clk),
    .io_clk(rvclkhdr_44_io_clk),
    .io_en(rvclkhdr_44_io_en),
    .io_scan_mode(rvclkhdr_44_io_scan_mode)
  );
  rvclkhdr rvclkhdr_45 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_45_io_l1clk),
    .io_clk(rvclkhdr_45_io_clk),
    .io_en(rvclkhdr_45_io_en),
    .io_scan_mode(rvclkhdr_45_io_scan_mode)
  );
  rvclkhdr rvclkhdr_46 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_46_io_l1clk),
    .io_clk(rvclkhdr_46_io_clk),
    .io_en(rvclkhdr_46_io_en),
    .io_scan_mode(rvclkhdr_46_io_scan_mode)
  );
  rvclkhdr rvclkhdr_47 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_47_io_l1clk),
    .io_clk(rvclkhdr_47_io_clk),
    .io_en(rvclkhdr_47_io_en),
    .io_scan_mode(rvclkhdr_47_io_scan_mode)
  );
  rvclkhdr rvclkhdr_48 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_48_io_l1clk),
    .io_clk(rvclkhdr_48_io_clk),
    .io_en(rvclkhdr_48_io_en),
    .io_scan_mode(rvclkhdr_48_io_scan_mode)
  );
  rvclkhdr rvclkhdr_49 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_49_io_l1clk),
    .io_clk(rvclkhdr_49_io_clk),
    .io_en(rvclkhdr_49_io_en),
    .io_scan_mode(rvclkhdr_49_io_scan_mode)
  );
  rvclkhdr rvclkhdr_50 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_50_io_l1clk),
    .io_clk(rvclkhdr_50_io_clk),
    .io_en(rvclkhdr_50_io_en),
    .io_scan_mode(rvclkhdr_50_io_scan_mode)
  );
  rvclkhdr rvclkhdr_51 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_51_io_l1clk),
    .io_clk(rvclkhdr_51_io_clk),
    .io_en(rvclkhdr_51_io_en),
    .io_scan_mode(rvclkhdr_51_io_scan_mode)
  );
  rvclkhdr rvclkhdr_52 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_52_io_l1clk),
    .io_clk(rvclkhdr_52_io_clk),
    .io_en(rvclkhdr_52_io_en),
    .io_scan_mode(rvclkhdr_52_io_scan_mode)
  );
  rvclkhdr rvclkhdr_53 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_53_io_l1clk),
    .io_clk(rvclkhdr_53_io_clk),
    .io_en(rvclkhdr_53_io_en),
    .io_scan_mode(rvclkhdr_53_io_scan_mode)
  );
  rvclkhdr rvclkhdr_54 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_54_io_l1clk),
    .io_clk(rvclkhdr_54_io_clk),
    .io_en(rvclkhdr_54_io_en),
    .io_scan_mode(rvclkhdr_54_io_scan_mode)
  );
  rvclkhdr rvclkhdr_55 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_55_io_l1clk),
    .io_clk(rvclkhdr_55_io_clk),
    .io_en(rvclkhdr_55_io_en),
    .io_scan_mode(rvclkhdr_55_io_scan_mode)
  );
  rvclkhdr rvclkhdr_56 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_56_io_l1clk),
    .io_clk(rvclkhdr_56_io_clk),
    .io_en(rvclkhdr_56_io_en),
    .io_scan_mode(rvclkhdr_56_io_scan_mode)
  );
  rvclkhdr rvclkhdr_57 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_57_io_l1clk),
    .io_clk(rvclkhdr_57_io_clk),
    .io_en(rvclkhdr_57_io_en),
    .io_scan_mode(rvclkhdr_57_io_scan_mode)
  );
  rvclkhdr rvclkhdr_58 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_58_io_l1clk),
    .io_clk(rvclkhdr_58_io_clk),
    .io_en(rvclkhdr_58_io_en),
    .io_scan_mode(rvclkhdr_58_io_scan_mode)
  );
  rvclkhdr rvclkhdr_59 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_59_io_l1clk),
    .io_clk(rvclkhdr_59_io_clk),
    .io_en(rvclkhdr_59_io_en),
    .io_scan_mode(rvclkhdr_59_io_scan_mode)
  );
  rvclkhdr rvclkhdr_60 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_60_io_l1clk),
    .io_clk(rvclkhdr_60_io_clk),
    .io_en(rvclkhdr_60_io_en),
    .io_scan_mode(rvclkhdr_60_io_scan_mode)
  );
  rvclkhdr rvclkhdr_61 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_61_io_l1clk),
    .io_clk(rvclkhdr_61_io_clk),
    .io_en(rvclkhdr_61_io_en),
    .io_scan_mode(rvclkhdr_61_io_scan_mode)
  );
  rvclkhdr rvclkhdr_62 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_62_io_l1clk),
    .io_clk(rvclkhdr_62_io_clk),
    .io_en(rvclkhdr_62_io_en),
    .io_scan_mode(rvclkhdr_62_io_scan_mode)
  );
  rvclkhdr rvclkhdr_63 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_63_io_l1clk),
    .io_clk(rvclkhdr_63_io_clk),
    .io_en(rvclkhdr_63_io_en),
    .io_scan_mode(rvclkhdr_63_io_scan_mode)
  );
  rvclkhdr rvclkhdr_64 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_64_io_l1clk),
    .io_clk(rvclkhdr_64_io_clk),
    .io_en(rvclkhdr_64_io_en),
    .io_scan_mode(rvclkhdr_64_io_scan_mode)
  );
  rvclkhdr rvclkhdr_65 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_65_io_l1clk),
    .io_clk(rvclkhdr_65_io_clk),
    .io_en(rvclkhdr_65_io_en),
    .io_scan_mode(rvclkhdr_65_io_scan_mode)
  );
  rvclkhdr rvclkhdr_66 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_66_io_l1clk),
    .io_clk(rvclkhdr_66_io_clk),
    .io_en(rvclkhdr_66_io_en),
    .io_scan_mode(rvclkhdr_66_io_scan_mode)
  );
  rvclkhdr rvclkhdr_67 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_67_io_l1clk),
    .io_clk(rvclkhdr_67_io_clk),
    .io_en(rvclkhdr_67_io_en),
    .io_scan_mode(rvclkhdr_67_io_scan_mode)
  );
  rvclkhdr rvclkhdr_68 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_68_io_l1clk),
    .io_clk(rvclkhdr_68_io_clk),
    .io_en(rvclkhdr_68_io_en),
    .io_scan_mode(rvclkhdr_68_io_scan_mode)
  );
  rvclkhdr rvclkhdr_69 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_69_io_l1clk),
    .io_clk(rvclkhdr_69_io_clk),
    .io_en(rvclkhdr_69_io_en),
    .io_scan_mode(rvclkhdr_69_io_scan_mode)
  );
  rvclkhdr rvclkhdr_70 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_70_io_l1clk),
    .io_clk(rvclkhdr_70_io_clk),
    .io_en(rvclkhdr_70_io_en),
    .io_scan_mode(rvclkhdr_70_io_scan_mode)
  );
  rvclkhdr rvclkhdr_71 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_71_io_l1clk),
    .io_clk(rvclkhdr_71_io_clk),
    .io_en(rvclkhdr_71_io_en),
    .io_scan_mode(rvclkhdr_71_io_scan_mode)
  );
  rvclkhdr rvclkhdr_72 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_72_io_l1clk),
    .io_clk(rvclkhdr_72_io_clk),
    .io_en(rvclkhdr_72_io_en),
    .io_scan_mode(rvclkhdr_72_io_scan_mode)
  );
  rvclkhdr rvclkhdr_73 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_73_io_l1clk),
    .io_clk(rvclkhdr_73_io_clk),
    .io_en(rvclkhdr_73_io_en),
    .io_scan_mode(rvclkhdr_73_io_scan_mode)
  );
  rvclkhdr rvclkhdr_74 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_74_io_l1clk),
    .io_clk(rvclkhdr_74_io_clk),
    .io_en(rvclkhdr_74_io_en),
    .io_scan_mode(rvclkhdr_74_io_scan_mode)
  );
  rvclkhdr rvclkhdr_75 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_75_io_l1clk),
    .io_clk(rvclkhdr_75_io_clk),
    .io_en(rvclkhdr_75_io_en),
    .io_scan_mode(rvclkhdr_75_io_scan_mode)
  );
  rvclkhdr rvclkhdr_76 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_76_io_l1clk),
    .io_clk(rvclkhdr_76_io_clk),
    .io_en(rvclkhdr_76_io_en),
    .io_scan_mode(rvclkhdr_76_io_scan_mode)
  );
  rvclkhdr rvclkhdr_77 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_77_io_l1clk),
    .io_clk(rvclkhdr_77_io_clk),
    .io_en(rvclkhdr_77_io_en),
    .io_scan_mode(rvclkhdr_77_io_scan_mode)
  );
  rvclkhdr rvclkhdr_78 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_78_io_l1clk),
    .io_clk(rvclkhdr_78_io_clk),
    .io_en(rvclkhdr_78_io_en),
    .io_scan_mode(rvclkhdr_78_io_scan_mode)
  );
  rvclkhdr rvclkhdr_79 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_79_io_l1clk),
    .io_clk(rvclkhdr_79_io_clk),
    .io_en(rvclkhdr_79_io_en),
    .io_scan_mode(rvclkhdr_79_io_scan_mode)
  );
  rvclkhdr rvclkhdr_80 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_80_io_l1clk),
    .io_clk(rvclkhdr_80_io_clk),
    .io_en(rvclkhdr_80_io_en),
    .io_scan_mode(rvclkhdr_80_io_scan_mode)
  );
  rvclkhdr rvclkhdr_81 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_81_io_l1clk),
    .io_clk(rvclkhdr_81_io_clk),
    .io_en(rvclkhdr_81_io_en),
    .io_scan_mode(rvclkhdr_81_io_scan_mode)
  );
  rvclkhdr rvclkhdr_82 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_82_io_l1clk),
    .io_clk(rvclkhdr_82_io_clk),
    .io_en(rvclkhdr_82_io_en),
    .io_scan_mode(rvclkhdr_82_io_scan_mode)
  );
  rvclkhdr rvclkhdr_83 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_83_io_l1clk),
    .io_clk(rvclkhdr_83_io_clk),
    .io_en(rvclkhdr_83_io_en),
    .io_scan_mode(rvclkhdr_83_io_scan_mode)
  );
  rvclkhdr rvclkhdr_84 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_84_io_l1clk),
    .io_clk(rvclkhdr_84_io_clk),
    .io_en(rvclkhdr_84_io_en),
    .io_scan_mode(rvclkhdr_84_io_scan_mode)
  );
  rvclkhdr rvclkhdr_85 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_85_io_l1clk),
    .io_clk(rvclkhdr_85_io_clk),
    .io_en(rvclkhdr_85_io_en),
    .io_scan_mode(rvclkhdr_85_io_scan_mode)
  );
  rvclkhdr rvclkhdr_86 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_86_io_l1clk),
    .io_clk(rvclkhdr_86_io_clk),
    .io_en(rvclkhdr_86_io_en),
    .io_scan_mode(rvclkhdr_86_io_scan_mode)
  );
  rvclkhdr rvclkhdr_87 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_87_io_l1clk),
    .io_clk(rvclkhdr_87_io_clk),
    .io_en(rvclkhdr_87_io_en),
    .io_scan_mode(rvclkhdr_87_io_scan_mode)
  );
  rvclkhdr rvclkhdr_88 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_88_io_l1clk),
    .io_clk(rvclkhdr_88_io_clk),
    .io_en(rvclkhdr_88_io_en),
    .io_scan_mode(rvclkhdr_88_io_scan_mode)
  );
  rvclkhdr rvclkhdr_89 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_89_io_l1clk),
    .io_clk(rvclkhdr_89_io_clk),
    .io_en(rvclkhdr_89_io_en),
    .io_scan_mode(rvclkhdr_89_io_scan_mode)
  );
  rvclkhdr rvclkhdr_90 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_90_io_l1clk),
    .io_clk(rvclkhdr_90_io_clk),
    .io_en(rvclkhdr_90_io_en),
    .io_scan_mode(rvclkhdr_90_io_scan_mode)
  );
  rvclkhdr rvclkhdr_91 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_91_io_l1clk),
    .io_clk(rvclkhdr_91_io_clk),
    .io_en(rvclkhdr_91_io_en),
    .io_scan_mode(rvclkhdr_91_io_scan_mode)
  );
  rvclkhdr rvclkhdr_92 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_92_io_l1clk),
    .io_clk(rvclkhdr_92_io_clk),
    .io_en(rvclkhdr_92_io_en),
    .io_scan_mode(rvclkhdr_92_io_scan_mode)
  );
  rvclkhdr rvclkhdr_93 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_93_io_l1clk),
    .io_clk(rvclkhdr_93_io_clk),
    .io_en(rvclkhdr_93_io_en),
    .io_scan_mode(rvclkhdr_93_io_scan_mode)
  );
  rvclkhdr rvclkhdr_94 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_94_io_l1clk),
    .io_clk(rvclkhdr_94_io_clk),
    .io_en(rvclkhdr_94_io_en),
    .io_scan_mode(rvclkhdr_94_io_scan_mode)
  );
  rvclkhdr rvclkhdr_95 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_95_io_l1clk),
    .io_clk(rvclkhdr_95_io_clk),
    .io_en(rvclkhdr_95_io_en),
    .io_scan_mode(rvclkhdr_95_io_scan_mode)
  );
  rvclkhdr rvclkhdr_96 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_96_io_l1clk),
    .io_clk(rvclkhdr_96_io_clk),
    .io_en(rvclkhdr_96_io_en),
    .io_scan_mode(rvclkhdr_96_io_scan_mode)
  );
  rvclkhdr rvclkhdr_97 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_97_io_l1clk),
    .io_clk(rvclkhdr_97_io_clk),
    .io_en(rvclkhdr_97_io_en),
    .io_scan_mode(rvclkhdr_97_io_scan_mode)
  );
  rvclkhdr rvclkhdr_98 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_98_io_l1clk),
    .io_clk(rvclkhdr_98_io_clk),
    .io_en(rvclkhdr_98_io_en),
    .io_scan_mode(rvclkhdr_98_io_scan_mode)
  );
  rvclkhdr rvclkhdr_99 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_99_io_l1clk),
    .io_clk(rvclkhdr_99_io_clk),
    .io_en(rvclkhdr_99_io_en),
    .io_scan_mode(rvclkhdr_99_io_scan_mode)
  );
  rvclkhdr rvclkhdr_100 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_100_io_l1clk),
    .io_clk(rvclkhdr_100_io_clk),
    .io_en(rvclkhdr_100_io_en),
    .io_scan_mode(rvclkhdr_100_io_scan_mode)
  );
  rvclkhdr rvclkhdr_101 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_101_io_l1clk),
    .io_clk(rvclkhdr_101_io_clk),
    .io_en(rvclkhdr_101_io_en),
    .io_scan_mode(rvclkhdr_101_io_scan_mode)
  );
  rvclkhdr rvclkhdr_102 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_102_io_l1clk),
    .io_clk(rvclkhdr_102_io_clk),
    .io_en(rvclkhdr_102_io_en),
    .io_scan_mode(rvclkhdr_102_io_scan_mode)
  );
  rvclkhdr rvclkhdr_103 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_103_io_l1clk),
    .io_clk(rvclkhdr_103_io_clk),
    .io_en(rvclkhdr_103_io_en),
    .io_scan_mode(rvclkhdr_103_io_scan_mode)
  );
  rvclkhdr rvclkhdr_104 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_104_io_l1clk),
    .io_clk(rvclkhdr_104_io_clk),
    .io_en(rvclkhdr_104_io_en),
    .io_scan_mode(rvclkhdr_104_io_scan_mode)
  );
  rvclkhdr rvclkhdr_105 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_105_io_l1clk),
    .io_clk(rvclkhdr_105_io_clk),
    .io_en(rvclkhdr_105_io_en),
    .io_scan_mode(rvclkhdr_105_io_scan_mode)
  );
  rvclkhdr rvclkhdr_106 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_106_io_l1clk),
    .io_clk(rvclkhdr_106_io_clk),
    .io_en(rvclkhdr_106_io_en),
    .io_scan_mode(rvclkhdr_106_io_scan_mode)
  );
  rvclkhdr rvclkhdr_107 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_107_io_l1clk),
    .io_clk(rvclkhdr_107_io_clk),
    .io_en(rvclkhdr_107_io_en),
    .io_scan_mode(rvclkhdr_107_io_scan_mode)
  );
  rvclkhdr rvclkhdr_108 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_108_io_l1clk),
    .io_clk(rvclkhdr_108_io_clk),
    .io_en(rvclkhdr_108_io_en),
    .io_scan_mode(rvclkhdr_108_io_scan_mode)
  );
  rvclkhdr rvclkhdr_109 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_109_io_l1clk),
    .io_clk(rvclkhdr_109_io_clk),
    .io_en(rvclkhdr_109_io_en),
    .io_scan_mode(rvclkhdr_109_io_scan_mode)
  );
  rvclkhdr rvclkhdr_110 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_110_io_l1clk),
    .io_clk(rvclkhdr_110_io_clk),
    .io_en(rvclkhdr_110_io_en),
    .io_scan_mode(rvclkhdr_110_io_scan_mode)
  );
  rvclkhdr rvclkhdr_111 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_111_io_l1clk),
    .io_clk(rvclkhdr_111_io_clk),
    .io_en(rvclkhdr_111_io_en),
    .io_scan_mode(rvclkhdr_111_io_scan_mode)
  );
  rvclkhdr rvclkhdr_112 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_112_io_l1clk),
    .io_clk(rvclkhdr_112_io_clk),
    .io_en(rvclkhdr_112_io_en),
    .io_scan_mode(rvclkhdr_112_io_scan_mode)
  );
  rvclkhdr rvclkhdr_113 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_113_io_l1clk),
    .io_clk(rvclkhdr_113_io_clk),
    .io_en(rvclkhdr_113_io_en),
    .io_scan_mode(rvclkhdr_113_io_scan_mode)
  );
  rvclkhdr rvclkhdr_114 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_114_io_l1clk),
    .io_clk(rvclkhdr_114_io_clk),
    .io_en(rvclkhdr_114_io_en),
    .io_scan_mode(rvclkhdr_114_io_scan_mode)
  );
  rvclkhdr rvclkhdr_115 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_115_io_l1clk),
    .io_clk(rvclkhdr_115_io_clk),
    .io_en(rvclkhdr_115_io_en),
    .io_scan_mode(rvclkhdr_115_io_scan_mode)
  );
  rvclkhdr rvclkhdr_116 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_116_io_l1clk),
    .io_clk(rvclkhdr_116_io_clk),
    .io_en(rvclkhdr_116_io_en),
    .io_scan_mode(rvclkhdr_116_io_scan_mode)
  );
  rvclkhdr rvclkhdr_117 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_117_io_l1clk),
    .io_clk(rvclkhdr_117_io_clk),
    .io_en(rvclkhdr_117_io_en),
    .io_scan_mode(rvclkhdr_117_io_scan_mode)
  );
  rvclkhdr rvclkhdr_118 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_118_io_l1clk),
    .io_clk(rvclkhdr_118_io_clk),
    .io_en(rvclkhdr_118_io_en),
    .io_scan_mode(rvclkhdr_118_io_scan_mode)
  );
  rvclkhdr rvclkhdr_119 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_119_io_l1clk),
    .io_clk(rvclkhdr_119_io_clk),
    .io_en(rvclkhdr_119_io_en),
    .io_scan_mode(rvclkhdr_119_io_scan_mode)
  );
  rvclkhdr rvclkhdr_120 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_120_io_l1clk),
    .io_clk(rvclkhdr_120_io_clk),
    .io_en(rvclkhdr_120_io_en),
    .io_scan_mode(rvclkhdr_120_io_scan_mode)
  );
  rvclkhdr rvclkhdr_121 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_121_io_l1clk),
    .io_clk(rvclkhdr_121_io_clk),
    .io_en(rvclkhdr_121_io_en),
    .io_scan_mode(rvclkhdr_121_io_scan_mode)
  );
  rvclkhdr rvclkhdr_122 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_122_io_l1clk),
    .io_clk(rvclkhdr_122_io_clk),
    .io_en(rvclkhdr_122_io_en),
    .io_scan_mode(rvclkhdr_122_io_scan_mode)
  );
  rvclkhdr rvclkhdr_123 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_123_io_l1clk),
    .io_clk(rvclkhdr_123_io_clk),
    .io_en(rvclkhdr_123_io_en),
    .io_scan_mode(rvclkhdr_123_io_scan_mode)
  );
  rvclkhdr rvclkhdr_124 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_124_io_l1clk),
    .io_clk(rvclkhdr_124_io_clk),
    .io_en(rvclkhdr_124_io_en),
    .io_scan_mode(rvclkhdr_124_io_scan_mode)
  );
  rvclkhdr rvclkhdr_125 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_125_io_l1clk),
    .io_clk(rvclkhdr_125_io_clk),
    .io_en(rvclkhdr_125_io_en),
    .io_scan_mode(rvclkhdr_125_io_scan_mode)
  );
  rvclkhdr rvclkhdr_126 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_126_io_l1clk),
    .io_clk(rvclkhdr_126_io_clk),
    .io_en(rvclkhdr_126_io_en),
    .io_scan_mode(rvclkhdr_126_io_scan_mode)
  );
  rvclkhdr rvclkhdr_127 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_127_io_l1clk),
    .io_clk(rvclkhdr_127_io_clk),
    .io_en(rvclkhdr_127_io_en),
    .io_scan_mode(rvclkhdr_127_io_scan_mode)
  );
  rvclkhdr rvclkhdr_128 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_128_io_l1clk),
    .io_clk(rvclkhdr_128_io_clk),
    .io_en(rvclkhdr_128_io_en),
    .io_scan_mode(rvclkhdr_128_io_scan_mode)
  );
  rvclkhdr rvclkhdr_129 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_129_io_l1clk),
    .io_clk(rvclkhdr_129_io_clk),
    .io_en(rvclkhdr_129_io_en),
    .io_scan_mode(rvclkhdr_129_io_scan_mode)
  );
  rvclkhdr rvclkhdr_130 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_130_io_l1clk),
    .io_clk(rvclkhdr_130_io_clk),
    .io_en(rvclkhdr_130_io_en),
    .io_scan_mode(rvclkhdr_130_io_scan_mode)
  );
  rvclkhdr rvclkhdr_131 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_131_io_l1clk),
    .io_clk(rvclkhdr_131_io_clk),
    .io_en(rvclkhdr_131_io_en),
    .io_scan_mode(rvclkhdr_131_io_scan_mode)
  );
  rvclkhdr rvclkhdr_132 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_132_io_l1clk),
    .io_clk(rvclkhdr_132_io_clk),
    .io_en(rvclkhdr_132_io_en),
    .io_scan_mode(rvclkhdr_132_io_scan_mode)
  );
  rvclkhdr rvclkhdr_133 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_133_io_l1clk),
    .io_clk(rvclkhdr_133_io_clk),
    .io_en(rvclkhdr_133_io_en),
    .io_scan_mode(rvclkhdr_133_io_scan_mode)
  );
  rvclkhdr rvclkhdr_134 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_134_io_l1clk),
    .io_clk(rvclkhdr_134_io_clk),
    .io_en(rvclkhdr_134_io_en),
    .io_scan_mode(rvclkhdr_134_io_scan_mode)
  );
  rvclkhdr rvclkhdr_135 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_135_io_l1clk),
    .io_clk(rvclkhdr_135_io_clk),
    .io_en(rvclkhdr_135_io_en),
    .io_scan_mode(rvclkhdr_135_io_scan_mode)
  );
  rvclkhdr rvclkhdr_136 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_136_io_l1clk),
    .io_clk(rvclkhdr_136_io_clk),
    .io_en(rvclkhdr_136_io_en),
    .io_scan_mode(rvclkhdr_136_io_scan_mode)
  );
  rvclkhdr rvclkhdr_137 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_137_io_l1clk),
    .io_clk(rvclkhdr_137_io_clk),
    .io_en(rvclkhdr_137_io_en),
    .io_scan_mode(rvclkhdr_137_io_scan_mode)
  );
  rvclkhdr rvclkhdr_138 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_138_io_l1clk),
    .io_clk(rvclkhdr_138_io_clk),
    .io_en(rvclkhdr_138_io_en),
    .io_scan_mode(rvclkhdr_138_io_scan_mode)
  );
  rvclkhdr rvclkhdr_139 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_139_io_l1clk),
    .io_clk(rvclkhdr_139_io_clk),
    .io_en(rvclkhdr_139_io_en),
    .io_scan_mode(rvclkhdr_139_io_scan_mode)
  );
  rvclkhdr rvclkhdr_140 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_140_io_l1clk),
    .io_clk(rvclkhdr_140_io_clk),
    .io_en(rvclkhdr_140_io_en),
    .io_scan_mode(rvclkhdr_140_io_scan_mode)
  );
  rvclkhdr rvclkhdr_141 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_141_io_l1clk),
    .io_clk(rvclkhdr_141_io_clk),
    .io_en(rvclkhdr_141_io_en),
    .io_scan_mode(rvclkhdr_141_io_scan_mode)
  );
  rvclkhdr rvclkhdr_142 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_142_io_l1clk),
    .io_clk(rvclkhdr_142_io_clk),
    .io_en(rvclkhdr_142_io_en),
    .io_scan_mode(rvclkhdr_142_io_scan_mode)
  );
  rvclkhdr rvclkhdr_143 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_143_io_l1clk),
    .io_clk(rvclkhdr_143_io_clk),
    .io_en(rvclkhdr_143_io_en),
    .io_scan_mode(rvclkhdr_143_io_scan_mode)
  );
  rvclkhdr rvclkhdr_144 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_144_io_l1clk),
    .io_clk(rvclkhdr_144_io_clk),
    .io_en(rvclkhdr_144_io_en),
    .io_scan_mode(rvclkhdr_144_io_scan_mode)
  );
  rvclkhdr rvclkhdr_145 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_145_io_l1clk),
    .io_clk(rvclkhdr_145_io_clk),
    .io_en(rvclkhdr_145_io_en),
    .io_scan_mode(rvclkhdr_145_io_scan_mode)
  );
  rvclkhdr rvclkhdr_146 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_146_io_l1clk),
    .io_clk(rvclkhdr_146_io_clk),
    .io_en(rvclkhdr_146_io_en),
    .io_scan_mode(rvclkhdr_146_io_scan_mode)
  );
  rvclkhdr rvclkhdr_147 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_147_io_l1clk),
    .io_clk(rvclkhdr_147_io_clk),
    .io_en(rvclkhdr_147_io_en),
    .io_scan_mode(rvclkhdr_147_io_scan_mode)
  );
  rvclkhdr rvclkhdr_148 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_148_io_l1clk),
    .io_clk(rvclkhdr_148_io_clk),
    .io_en(rvclkhdr_148_io_en),
    .io_scan_mode(rvclkhdr_148_io_scan_mode)
  );
  rvclkhdr rvclkhdr_149 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_149_io_l1clk),
    .io_clk(rvclkhdr_149_io_clk),
    .io_en(rvclkhdr_149_io_en),
    .io_scan_mode(rvclkhdr_149_io_scan_mode)
  );
  rvclkhdr rvclkhdr_150 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_150_io_l1clk),
    .io_clk(rvclkhdr_150_io_clk),
    .io_en(rvclkhdr_150_io_en),
    .io_scan_mode(rvclkhdr_150_io_scan_mode)
  );
  rvclkhdr rvclkhdr_151 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_151_io_l1clk),
    .io_clk(rvclkhdr_151_io_clk),
    .io_en(rvclkhdr_151_io_en),
    .io_scan_mode(rvclkhdr_151_io_scan_mode)
  );
  rvclkhdr rvclkhdr_152 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_152_io_l1clk),
    .io_clk(rvclkhdr_152_io_clk),
    .io_en(rvclkhdr_152_io_en),
    .io_scan_mode(rvclkhdr_152_io_scan_mode)
  );
  rvclkhdr rvclkhdr_153 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_153_io_l1clk),
    .io_clk(rvclkhdr_153_io_clk),
    .io_en(rvclkhdr_153_io_en),
    .io_scan_mode(rvclkhdr_153_io_scan_mode)
  );
  rvclkhdr rvclkhdr_154 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_154_io_l1clk),
    .io_clk(rvclkhdr_154_io_clk),
    .io_en(rvclkhdr_154_io_en),
    .io_scan_mode(rvclkhdr_154_io_scan_mode)
  );
  rvclkhdr rvclkhdr_155 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_155_io_l1clk),
    .io_clk(rvclkhdr_155_io_clk),
    .io_en(rvclkhdr_155_io_en),
    .io_scan_mode(rvclkhdr_155_io_scan_mode)
  );
  rvclkhdr rvclkhdr_156 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_156_io_l1clk),
    .io_clk(rvclkhdr_156_io_clk),
    .io_en(rvclkhdr_156_io_en),
    .io_scan_mode(rvclkhdr_156_io_scan_mode)
  );
  rvclkhdr rvclkhdr_157 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_157_io_l1clk),
    .io_clk(rvclkhdr_157_io_clk),
    .io_en(rvclkhdr_157_io_en),
    .io_scan_mode(rvclkhdr_157_io_scan_mode)
  );
  rvclkhdr rvclkhdr_158 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_158_io_l1clk),
    .io_clk(rvclkhdr_158_io_clk),
    .io_en(rvclkhdr_158_io_en),
    .io_scan_mode(rvclkhdr_158_io_scan_mode)
  );
  rvclkhdr rvclkhdr_159 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_159_io_l1clk),
    .io_clk(rvclkhdr_159_io_clk),
    .io_en(rvclkhdr_159_io_en),
    .io_scan_mode(rvclkhdr_159_io_scan_mode)
  );
  rvclkhdr rvclkhdr_160 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_160_io_l1clk),
    .io_clk(rvclkhdr_160_io_clk),
    .io_en(rvclkhdr_160_io_en),
    .io_scan_mode(rvclkhdr_160_io_scan_mode)
  );
  rvclkhdr rvclkhdr_161 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_161_io_l1clk),
    .io_clk(rvclkhdr_161_io_clk),
    .io_en(rvclkhdr_161_io_en),
    .io_scan_mode(rvclkhdr_161_io_scan_mode)
  );
  rvclkhdr rvclkhdr_162 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_162_io_l1clk),
    .io_clk(rvclkhdr_162_io_clk),
    .io_en(rvclkhdr_162_io_en),
    .io_scan_mode(rvclkhdr_162_io_scan_mode)
  );
  rvclkhdr rvclkhdr_163 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_163_io_l1clk),
    .io_clk(rvclkhdr_163_io_clk),
    .io_en(rvclkhdr_163_io_en),
    .io_scan_mode(rvclkhdr_163_io_scan_mode)
  );
  rvclkhdr rvclkhdr_164 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_164_io_l1clk),
    .io_clk(rvclkhdr_164_io_clk),
    .io_en(rvclkhdr_164_io_en),
    .io_scan_mode(rvclkhdr_164_io_scan_mode)
  );
  rvclkhdr rvclkhdr_165 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_165_io_l1clk),
    .io_clk(rvclkhdr_165_io_clk),
    .io_en(rvclkhdr_165_io_en),
    .io_scan_mode(rvclkhdr_165_io_scan_mode)
  );
  rvclkhdr rvclkhdr_166 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_166_io_l1clk),
    .io_clk(rvclkhdr_166_io_clk),
    .io_en(rvclkhdr_166_io_en),
    .io_scan_mode(rvclkhdr_166_io_scan_mode)
  );
  rvclkhdr rvclkhdr_167 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_167_io_l1clk),
    .io_clk(rvclkhdr_167_io_clk),
    .io_en(rvclkhdr_167_io_en),
    .io_scan_mode(rvclkhdr_167_io_scan_mode)
  );
  rvclkhdr rvclkhdr_168 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_168_io_l1clk),
    .io_clk(rvclkhdr_168_io_clk),
    .io_en(rvclkhdr_168_io_en),
    .io_scan_mode(rvclkhdr_168_io_scan_mode)
  );
  rvclkhdr rvclkhdr_169 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_169_io_l1clk),
    .io_clk(rvclkhdr_169_io_clk),
    .io_en(rvclkhdr_169_io_en),
    .io_scan_mode(rvclkhdr_169_io_scan_mode)
  );
  rvclkhdr rvclkhdr_170 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_170_io_l1clk),
    .io_clk(rvclkhdr_170_io_clk),
    .io_en(rvclkhdr_170_io_en),
    .io_scan_mode(rvclkhdr_170_io_scan_mode)
  );
  rvclkhdr rvclkhdr_171 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_171_io_l1clk),
    .io_clk(rvclkhdr_171_io_clk),
    .io_en(rvclkhdr_171_io_en),
    .io_scan_mode(rvclkhdr_171_io_scan_mode)
  );
  rvclkhdr rvclkhdr_172 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_172_io_l1clk),
    .io_clk(rvclkhdr_172_io_clk),
    .io_en(rvclkhdr_172_io_en),
    .io_scan_mode(rvclkhdr_172_io_scan_mode)
  );
  rvclkhdr rvclkhdr_173 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_173_io_l1clk),
    .io_clk(rvclkhdr_173_io_clk),
    .io_en(rvclkhdr_173_io_en),
    .io_scan_mode(rvclkhdr_173_io_scan_mode)
  );
  rvclkhdr rvclkhdr_174 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_174_io_l1clk),
    .io_clk(rvclkhdr_174_io_clk),
    .io_en(rvclkhdr_174_io_en),
    .io_scan_mode(rvclkhdr_174_io_scan_mode)
  );
  rvclkhdr rvclkhdr_175 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_175_io_l1clk),
    .io_clk(rvclkhdr_175_io_clk),
    .io_en(rvclkhdr_175_io_en),
    .io_scan_mode(rvclkhdr_175_io_scan_mode)
  );
  rvclkhdr rvclkhdr_176 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_176_io_l1clk),
    .io_clk(rvclkhdr_176_io_clk),
    .io_en(rvclkhdr_176_io_en),
    .io_scan_mode(rvclkhdr_176_io_scan_mode)
  );
  rvclkhdr rvclkhdr_177 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_177_io_l1clk),
    .io_clk(rvclkhdr_177_io_clk),
    .io_en(rvclkhdr_177_io_en),
    .io_scan_mode(rvclkhdr_177_io_scan_mode)
  );
  rvclkhdr rvclkhdr_178 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_178_io_l1clk),
    .io_clk(rvclkhdr_178_io_clk),
    .io_en(rvclkhdr_178_io_en),
    .io_scan_mode(rvclkhdr_178_io_scan_mode)
  );
  rvclkhdr rvclkhdr_179 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_179_io_l1clk),
    .io_clk(rvclkhdr_179_io_clk),
    .io_en(rvclkhdr_179_io_en),
    .io_scan_mode(rvclkhdr_179_io_scan_mode)
  );
  rvclkhdr rvclkhdr_180 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_180_io_l1clk),
    .io_clk(rvclkhdr_180_io_clk),
    .io_en(rvclkhdr_180_io_en),
    .io_scan_mode(rvclkhdr_180_io_scan_mode)
  );
  rvclkhdr rvclkhdr_181 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_181_io_l1clk),
    .io_clk(rvclkhdr_181_io_clk),
    .io_en(rvclkhdr_181_io_en),
    .io_scan_mode(rvclkhdr_181_io_scan_mode)
  );
  rvclkhdr rvclkhdr_182 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_182_io_l1clk),
    .io_clk(rvclkhdr_182_io_clk),
    .io_en(rvclkhdr_182_io_en),
    .io_scan_mode(rvclkhdr_182_io_scan_mode)
  );
  rvclkhdr rvclkhdr_183 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_183_io_l1clk),
    .io_clk(rvclkhdr_183_io_clk),
    .io_en(rvclkhdr_183_io_en),
    .io_scan_mode(rvclkhdr_183_io_scan_mode)
  );
  rvclkhdr rvclkhdr_184 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_184_io_l1clk),
    .io_clk(rvclkhdr_184_io_clk),
    .io_en(rvclkhdr_184_io_en),
    .io_scan_mode(rvclkhdr_184_io_scan_mode)
  );
  rvclkhdr rvclkhdr_185 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_185_io_l1clk),
    .io_clk(rvclkhdr_185_io_clk),
    .io_en(rvclkhdr_185_io_en),
    .io_scan_mode(rvclkhdr_185_io_scan_mode)
  );
  rvclkhdr rvclkhdr_186 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_186_io_l1clk),
    .io_clk(rvclkhdr_186_io_clk),
    .io_en(rvclkhdr_186_io_en),
    .io_scan_mode(rvclkhdr_186_io_scan_mode)
  );
  rvclkhdr rvclkhdr_187 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_187_io_l1clk),
    .io_clk(rvclkhdr_187_io_clk),
    .io_en(rvclkhdr_187_io_en),
    .io_scan_mode(rvclkhdr_187_io_scan_mode)
  );
  rvclkhdr rvclkhdr_188 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_188_io_l1clk),
    .io_clk(rvclkhdr_188_io_clk),
    .io_en(rvclkhdr_188_io_en),
    .io_scan_mode(rvclkhdr_188_io_scan_mode)
  );
  rvclkhdr rvclkhdr_189 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_189_io_l1clk),
    .io_clk(rvclkhdr_189_io_clk),
    .io_en(rvclkhdr_189_io_en),
    .io_scan_mode(rvclkhdr_189_io_scan_mode)
  );
  rvclkhdr rvclkhdr_190 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_190_io_l1clk),
    .io_clk(rvclkhdr_190_io_clk),
    .io_en(rvclkhdr_190_io_en),
    .io_scan_mode(rvclkhdr_190_io_scan_mode)
  );
  rvclkhdr rvclkhdr_191 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_191_io_l1clk),
    .io_clk(rvclkhdr_191_io_clk),
    .io_en(rvclkhdr_191_io_en),
    .io_scan_mode(rvclkhdr_191_io_scan_mode)
  );
  rvclkhdr rvclkhdr_192 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_192_io_l1clk),
    .io_clk(rvclkhdr_192_io_clk),
    .io_en(rvclkhdr_192_io_en),
    .io_scan_mode(rvclkhdr_192_io_scan_mode)
  );
  rvclkhdr rvclkhdr_193 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_193_io_l1clk),
    .io_clk(rvclkhdr_193_io_clk),
    .io_en(rvclkhdr_193_io_en),
    .io_scan_mode(rvclkhdr_193_io_scan_mode)
  );
  rvclkhdr rvclkhdr_194 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_194_io_l1clk),
    .io_clk(rvclkhdr_194_io_clk),
    .io_en(rvclkhdr_194_io_en),
    .io_scan_mode(rvclkhdr_194_io_scan_mode)
  );
  rvclkhdr rvclkhdr_195 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_195_io_l1clk),
    .io_clk(rvclkhdr_195_io_clk),
    .io_en(rvclkhdr_195_io_en),
    .io_scan_mode(rvclkhdr_195_io_scan_mode)
  );
  rvclkhdr rvclkhdr_196 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_196_io_l1clk),
    .io_clk(rvclkhdr_196_io_clk),
    .io_en(rvclkhdr_196_io_en),
    .io_scan_mode(rvclkhdr_196_io_scan_mode)
  );
  rvclkhdr rvclkhdr_197 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_197_io_l1clk),
    .io_clk(rvclkhdr_197_io_clk),
    .io_en(rvclkhdr_197_io_en),
    .io_scan_mode(rvclkhdr_197_io_scan_mode)
  );
  rvclkhdr rvclkhdr_198 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_198_io_l1clk),
    .io_clk(rvclkhdr_198_io_clk),
    .io_en(rvclkhdr_198_io_en),
    .io_scan_mode(rvclkhdr_198_io_scan_mode)
  );
  rvclkhdr rvclkhdr_199 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_199_io_l1clk),
    .io_clk(rvclkhdr_199_io_clk),
    .io_en(rvclkhdr_199_io_en),
    .io_scan_mode(rvclkhdr_199_io_scan_mode)
  );
  rvclkhdr rvclkhdr_200 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_200_io_l1clk),
    .io_clk(rvclkhdr_200_io_clk),
    .io_en(rvclkhdr_200_io_en),
    .io_scan_mode(rvclkhdr_200_io_scan_mode)
  );
  rvclkhdr rvclkhdr_201 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_201_io_l1clk),
    .io_clk(rvclkhdr_201_io_clk),
    .io_en(rvclkhdr_201_io_en),
    .io_scan_mode(rvclkhdr_201_io_scan_mode)
  );
  rvclkhdr rvclkhdr_202 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_202_io_l1clk),
    .io_clk(rvclkhdr_202_io_clk),
    .io_en(rvclkhdr_202_io_en),
    .io_scan_mode(rvclkhdr_202_io_scan_mode)
  );
  rvclkhdr rvclkhdr_203 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_203_io_l1clk),
    .io_clk(rvclkhdr_203_io_clk),
    .io_en(rvclkhdr_203_io_en),
    .io_scan_mode(rvclkhdr_203_io_scan_mode)
  );
  rvclkhdr rvclkhdr_204 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_204_io_l1clk),
    .io_clk(rvclkhdr_204_io_clk),
    .io_en(rvclkhdr_204_io_en),
    .io_scan_mode(rvclkhdr_204_io_scan_mode)
  );
  rvclkhdr rvclkhdr_205 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_205_io_l1clk),
    .io_clk(rvclkhdr_205_io_clk),
    .io_en(rvclkhdr_205_io_en),
    .io_scan_mode(rvclkhdr_205_io_scan_mode)
  );
  rvclkhdr rvclkhdr_206 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_206_io_l1clk),
    .io_clk(rvclkhdr_206_io_clk),
    .io_en(rvclkhdr_206_io_en),
    .io_scan_mode(rvclkhdr_206_io_scan_mode)
  );
  rvclkhdr rvclkhdr_207 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_207_io_l1clk),
    .io_clk(rvclkhdr_207_io_clk),
    .io_en(rvclkhdr_207_io_en),
    .io_scan_mode(rvclkhdr_207_io_scan_mode)
  );
  rvclkhdr rvclkhdr_208 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_208_io_l1clk),
    .io_clk(rvclkhdr_208_io_clk),
    .io_en(rvclkhdr_208_io_en),
    .io_scan_mode(rvclkhdr_208_io_scan_mode)
  );
  rvclkhdr rvclkhdr_209 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_209_io_l1clk),
    .io_clk(rvclkhdr_209_io_clk),
    .io_en(rvclkhdr_209_io_en),
    .io_scan_mode(rvclkhdr_209_io_scan_mode)
  );
  rvclkhdr rvclkhdr_210 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_210_io_l1clk),
    .io_clk(rvclkhdr_210_io_clk),
    .io_en(rvclkhdr_210_io_en),
    .io_scan_mode(rvclkhdr_210_io_scan_mode)
  );
  rvclkhdr rvclkhdr_211 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_211_io_l1clk),
    .io_clk(rvclkhdr_211_io_clk),
    .io_en(rvclkhdr_211_io_en),
    .io_scan_mode(rvclkhdr_211_io_scan_mode)
  );
  rvclkhdr rvclkhdr_212 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_212_io_l1clk),
    .io_clk(rvclkhdr_212_io_clk),
    .io_en(rvclkhdr_212_io_en),
    .io_scan_mode(rvclkhdr_212_io_scan_mode)
  );
  rvclkhdr rvclkhdr_213 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_213_io_l1clk),
    .io_clk(rvclkhdr_213_io_clk),
    .io_en(rvclkhdr_213_io_en),
    .io_scan_mode(rvclkhdr_213_io_scan_mode)
  );
  rvclkhdr rvclkhdr_214 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_214_io_l1clk),
    .io_clk(rvclkhdr_214_io_clk),
    .io_en(rvclkhdr_214_io_en),
    .io_scan_mode(rvclkhdr_214_io_scan_mode)
  );
  rvclkhdr rvclkhdr_215 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_215_io_l1clk),
    .io_clk(rvclkhdr_215_io_clk),
    .io_en(rvclkhdr_215_io_en),
    .io_scan_mode(rvclkhdr_215_io_scan_mode)
  );
  rvclkhdr rvclkhdr_216 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_216_io_l1clk),
    .io_clk(rvclkhdr_216_io_clk),
    .io_en(rvclkhdr_216_io_en),
    .io_scan_mode(rvclkhdr_216_io_scan_mode)
  );
  rvclkhdr rvclkhdr_217 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_217_io_l1clk),
    .io_clk(rvclkhdr_217_io_clk),
    .io_en(rvclkhdr_217_io_en),
    .io_scan_mode(rvclkhdr_217_io_scan_mode)
  );
  rvclkhdr rvclkhdr_218 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_218_io_l1clk),
    .io_clk(rvclkhdr_218_io_clk),
    .io_en(rvclkhdr_218_io_en),
    .io_scan_mode(rvclkhdr_218_io_scan_mode)
  );
  rvclkhdr rvclkhdr_219 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_219_io_l1clk),
    .io_clk(rvclkhdr_219_io_clk),
    .io_en(rvclkhdr_219_io_en),
    .io_scan_mode(rvclkhdr_219_io_scan_mode)
  );
  rvclkhdr rvclkhdr_220 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_220_io_l1clk),
    .io_clk(rvclkhdr_220_io_clk),
    .io_en(rvclkhdr_220_io_en),
    .io_scan_mode(rvclkhdr_220_io_scan_mode)
  );
  rvclkhdr rvclkhdr_221 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_221_io_l1clk),
    .io_clk(rvclkhdr_221_io_clk),
    .io_en(rvclkhdr_221_io_en),
    .io_scan_mode(rvclkhdr_221_io_scan_mode)
  );
  rvclkhdr rvclkhdr_222 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_222_io_l1clk),
    .io_clk(rvclkhdr_222_io_clk),
    .io_en(rvclkhdr_222_io_en),
    .io_scan_mode(rvclkhdr_222_io_scan_mode)
  );
  rvclkhdr rvclkhdr_223 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_223_io_l1clk),
    .io_clk(rvclkhdr_223_io_clk),
    .io_en(rvclkhdr_223_io_en),
    .io_scan_mode(rvclkhdr_223_io_scan_mode)
  );
  rvclkhdr rvclkhdr_224 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_224_io_l1clk),
    .io_clk(rvclkhdr_224_io_clk),
    .io_en(rvclkhdr_224_io_en),
    .io_scan_mode(rvclkhdr_224_io_scan_mode)
  );
  rvclkhdr rvclkhdr_225 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_225_io_l1clk),
    .io_clk(rvclkhdr_225_io_clk),
    .io_en(rvclkhdr_225_io_en),
    .io_scan_mode(rvclkhdr_225_io_scan_mode)
  );
  rvclkhdr rvclkhdr_226 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_226_io_l1clk),
    .io_clk(rvclkhdr_226_io_clk),
    .io_en(rvclkhdr_226_io_en),
    .io_scan_mode(rvclkhdr_226_io_scan_mode)
  );
  rvclkhdr rvclkhdr_227 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_227_io_l1clk),
    .io_clk(rvclkhdr_227_io_clk),
    .io_en(rvclkhdr_227_io_en),
    .io_scan_mode(rvclkhdr_227_io_scan_mode)
  );
  rvclkhdr rvclkhdr_228 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_228_io_l1clk),
    .io_clk(rvclkhdr_228_io_clk),
    .io_en(rvclkhdr_228_io_en),
    .io_scan_mode(rvclkhdr_228_io_scan_mode)
  );
  rvclkhdr rvclkhdr_229 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_229_io_l1clk),
    .io_clk(rvclkhdr_229_io_clk),
    .io_en(rvclkhdr_229_io_en),
    .io_scan_mode(rvclkhdr_229_io_scan_mode)
  );
  rvclkhdr rvclkhdr_230 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_230_io_l1clk),
    .io_clk(rvclkhdr_230_io_clk),
    .io_en(rvclkhdr_230_io_en),
    .io_scan_mode(rvclkhdr_230_io_scan_mode)
  );
  rvclkhdr rvclkhdr_231 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_231_io_l1clk),
    .io_clk(rvclkhdr_231_io_clk),
    .io_en(rvclkhdr_231_io_en),
    .io_scan_mode(rvclkhdr_231_io_scan_mode)
  );
  rvclkhdr rvclkhdr_232 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_232_io_l1clk),
    .io_clk(rvclkhdr_232_io_clk),
    .io_en(rvclkhdr_232_io_en),
    .io_scan_mode(rvclkhdr_232_io_scan_mode)
  );
  rvclkhdr rvclkhdr_233 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_233_io_l1clk),
    .io_clk(rvclkhdr_233_io_clk),
    .io_en(rvclkhdr_233_io_en),
    .io_scan_mode(rvclkhdr_233_io_scan_mode)
  );
  rvclkhdr rvclkhdr_234 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_234_io_l1clk),
    .io_clk(rvclkhdr_234_io_clk),
    .io_en(rvclkhdr_234_io_en),
    .io_scan_mode(rvclkhdr_234_io_scan_mode)
  );
  rvclkhdr rvclkhdr_235 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_235_io_l1clk),
    .io_clk(rvclkhdr_235_io_clk),
    .io_en(rvclkhdr_235_io_en),
    .io_scan_mode(rvclkhdr_235_io_scan_mode)
  );
  rvclkhdr rvclkhdr_236 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_236_io_l1clk),
    .io_clk(rvclkhdr_236_io_clk),
    .io_en(rvclkhdr_236_io_en),
    .io_scan_mode(rvclkhdr_236_io_scan_mode)
  );
  rvclkhdr rvclkhdr_237 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_237_io_l1clk),
    .io_clk(rvclkhdr_237_io_clk),
    .io_en(rvclkhdr_237_io_en),
    .io_scan_mode(rvclkhdr_237_io_scan_mode)
  );
  rvclkhdr rvclkhdr_238 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_238_io_l1clk),
    .io_clk(rvclkhdr_238_io_clk),
    .io_en(rvclkhdr_238_io_en),
    .io_scan_mode(rvclkhdr_238_io_scan_mode)
  );
  rvclkhdr rvclkhdr_239 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_239_io_l1clk),
    .io_clk(rvclkhdr_239_io_clk),
    .io_en(rvclkhdr_239_io_en),
    .io_scan_mode(rvclkhdr_239_io_scan_mode)
  );
  rvclkhdr rvclkhdr_240 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_240_io_l1clk),
    .io_clk(rvclkhdr_240_io_clk),
    .io_en(rvclkhdr_240_io_en),
    .io_scan_mode(rvclkhdr_240_io_scan_mode)
  );
  rvclkhdr rvclkhdr_241 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_241_io_l1clk),
    .io_clk(rvclkhdr_241_io_clk),
    .io_en(rvclkhdr_241_io_en),
    .io_scan_mode(rvclkhdr_241_io_scan_mode)
  );
  rvclkhdr rvclkhdr_242 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_242_io_l1clk),
    .io_clk(rvclkhdr_242_io_clk),
    .io_en(rvclkhdr_242_io_en),
    .io_scan_mode(rvclkhdr_242_io_scan_mode)
  );
  rvclkhdr rvclkhdr_243 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_243_io_l1clk),
    .io_clk(rvclkhdr_243_io_clk),
    .io_en(rvclkhdr_243_io_en),
    .io_scan_mode(rvclkhdr_243_io_scan_mode)
  );
  rvclkhdr rvclkhdr_244 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_244_io_l1clk),
    .io_clk(rvclkhdr_244_io_clk),
    .io_en(rvclkhdr_244_io_en),
    .io_scan_mode(rvclkhdr_244_io_scan_mode)
  );
  rvclkhdr rvclkhdr_245 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_245_io_l1clk),
    .io_clk(rvclkhdr_245_io_clk),
    .io_en(rvclkhdr_245_io_en),
    .io_scan_mode(rvclkhdr_245_io_scan_mode)
  );
  rvclkhdr rvclkhdr_246 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_246_io_l1clk),
    .io_clk(rvclkhdr_246_io_clk),
    .io_en(rvclkhdr_246_io_en),
    .io_scan_mode(rvclkhdr_246_io_scan_mode)
  );
  rvclkhdr rvclkhdr_247 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_247_io_l1clk),
    .io_clk(rvclkhdr_247_io_clk),
    .io_en(rvclkhdr_247_io_en),
    .io_scan_mode(rvclkhdr_247_io_scan_mode)
  );
  rvclkhdr rvclkhdr_248 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_248_io_l1clk),
    .io_clk(rvclkhdr_248_io_clk),
    .io_en(rvclkhdr_248_io_en),
    .io_scan_mode(rvclkhdr_248_io_scan_mode)
  );
  rvclkhdr rvclkhdr_249 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_249_io_l1clk),
    .io_clk(rvclkhdr_249_io_clk),
    .io_en(rvclkhdr_249_io_en),
    .io_scan_mode(rvclkhdr_249_io_scan_mode)
  );
  rvclkhdr rvclkhdr_250 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_250_io_l1clk),
    .io_clk(rvclkhdr_250_io_clk),
    .io_en(rvclkhdr_250_io_en),
    .io_scan_mode(rvclkhdr_250_io_scan_mode)
  );
  rvclkhdr rvclkhdr_251 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_251_io_l1clk),
    .io_clk(rvclkhdr_251_io_clk),
    .io_en(rvclkhdr_251_io_en),
    .io_scan_mode(rvclkhdr_251_io_scan_mode)
  );
  rvclkhdr rvclkhdr_252 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_252_io_l1clk),
    .io_clk(rvclkhdr_252_io_clk),
    .io_en(rvclkhdr_252_io_en),
    .io_scan_mode(rvclkhdr_252_io_scan_mode)
  );
  rvclkhdr rvclkhdr_253 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_253_io_l1clk),
    .io_clk(rvclkhdr_253_io_clk),
    .io_en(rvclkhdr_253_io_en),
    .io_scan_mode(rvclkhdr_253_io_scan_mode)
  );
  rvclkhdr rvclkhdr_254 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_254_io_l1clk),
    .io_clk(rvclkhdr_254_io_clk),
    .io_en(rvclkhdr_254_io_en),
    .io_scan_mode(rvclkhdr_254_io_scan_mode)
  );
  rvclkhdr rvclkhdr_255 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_255_io_l1clk),
    .io_clk(rvclkhdr_255_io_clk),
    .io_en(rvclkhdr_255_io_en),
    .io_scan_mode(rvclkhdr_255_io_scan_mode)
  );
  rvclkhdr rvclkhdr_256 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_256_io_l1clk),
    .io_clk(rvclkhdr_256_io_clk),
    .io_en(rvclkhdr_256_io_en),
    .io_scan_mode(rvclkhdr_256_io_scan_mode)
  );
  rvclkhdr rvclkhdr_257 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_257_io_l1clk),
    .io_clk(rvclkhdr_257_io_clk),
    .io_en(rvclkhdr_257_io_en),
    .io_scan_mode(rvclkhdr_257_io_scan_mode)
  );
  rvclkhdr rvclkhdr_258 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_258_io_l1clk),
    .io_clk(rvclkhdr_258_io_clk),
    .io_en(rvclkhdr_258_io_en),
    .io_scan_mode(rvclkhdr_258_io_scan_mode)
  );
  rvclkhdr rvclkhdr_259 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_259_io_l1clk),
    .io_clk(rvclkhdr_259_io_clk),
    .io_en(rvclkhdr_259_io_en),
    .io_scan_mode(rvclkhdr_259_io_scan_mode)
  );
  rvclkhdr rvclkhdr_260 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_260_io_l1clk),
    .io_clk(rvclkhdr_260_io_clk),
    .io_en(rvclkhdr_260_io_en),
    .io_scan_mode(rvclkhdr_260_io_scan_mode)
  );
  rvclkhdr rvclkhdr_261 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_261_io_l1clk),
    .io_clk(rvclkhdr_261_io_clk),
    .io_en(rvclkhdr_261_io_en),
    .io_scan_mode(rvclkhdr_261_io_scan_mode)
  );
  rvclkhdr rvclkhdr_262 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_262_io_l1clk),
    .io_clk(rvclkhdr_262_io_clk),
    .io_en(rvclkhdr_262_io_en),
    .io_scan_mode(rvclkhdr_262_io_scan_mode)
  );
  rvclkhdr rvclkhdr_263 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_263_io_l1clk),
    .io_clk(rvclkhdr_263_io_clk),
    .io_en(rvclkhdr_263_io_en),
    .io_scan_mode(rvclkhdr_263_io_scan_mode)
  );
  rvclkhdr rvclkhdr_264 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_264_io_l1clk),
    .io_clk(rvclkhdr_264_io_clk),
    .io_en(rvclkhdr_264_io_en),
    .io_scan_mode(rvclkhdr_264_io_scan_mode)
  );
  rvclkhdr rvclkhdr_265 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_265_io_l1clk),
    .io_clk(rvclkhdr_265_io_clk),
    .io_en(rvclkhdr_265_io_en),
    .io_scan_mode(rvclkhdr_265_io_scan_mode)
  );
  rvclkhdr rvclkhdr_266 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_266_io_l1clk),
    .io_clk(rvclkhdr_266_io_clk),
    .io_en(rvclkhdr_266_io_en),
    .io_scan_mode(rvclkhdr_266_io_scan_mode)
  );
  rvclkhdr rvclkhdr_267 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_267_io_l1clk),
    .io_clk(rvclkhdr_267_io_clk),
    .io_en(rvclkhdr_267_io_en),
    .io_scan_mode(rvclkhdr_267_io_scan_mode)
  );
  rvclkhdr rvclkhdr_268 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_268_io_l1clk),
    .io_clk(rvclkhdr_268_io_clk),
    .io_en(rvclkhdr_268_io_en),
    .io_scan_mode(rvclkhdr_268_io_scan_mode)
  );
  rvclkhdr rvclkhdr_269 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_269_io_l1clk),
    .io_clk(rvclkhdr_269_io_clk),
    .io_en(rvclkhdr_269_io_en),
    .io_scan_mode(rvclkhdr_269_io_scan_mode)
  );
  rvclkhdr rvclkhdr_270 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_270_io_l1clk),
    .io_clk(rvclkhdr_270_io_clk),
    .io_en(rvclkhdr_270_io_en),
    .io_scan_mode(rvclkhdr_270_io_scan_mode)
  );
  rvclkhdr rvclkhdr_271 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_271_io_l1clk),
    .io_clk(rvclkhdr_271_io_clk),
    .io_en(rvclkhdr_271_io_en),
    .io_scan_mode(rvclkhdr_271_io_scan_mode)
  );
  rvclkhdr rvclkhdr_272 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_272_io_l1clk),
    .io_clk(rvclkhdr_272_io_clk),
    .io_en(rvclkhdr_272_io_en),
    .io_scan_mode(rvclkhdr_272_io_scan_mode)
  );
  rvclkhdr rvclkhdr_273 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_273_io_l1clk),
    .io_clk(rvclkhdr_273_io_clk),
    .io_en(rvclkhdr_273_io_en),
    .io_scan_mode(rvclkhdr_273_io_scan_mode)
  );
  rvclkhdr rvclkhdr_274 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_274_io_l1clk),
    .io_clk(rvclkhdr_274_io_clk),
    .io_en(rvclkhdr_274_io_en),
    .io_scan_mode(rvclkhdr_274_io_scan_mode)
  );
  rvclkhdr rvclkhdr_275 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_275_io_l1clk),
    .io_clk(rvclkhdr_275_io_clk),
    .io_en(rvclkhdr_275_io_en),
    .io_scan_mode(rvclkhdr_275_io_scan_mode)
  );
  rvclkhdr rvclkhdr_276 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_276_io_l1clk),
    .io_clk(rvclkhdr_276_io_clk),
    .io_en(rvclkhdr_276_io_en),
    .io_scan_mode(rvclkhdr_276_io_scan_mode)
  );
  rvclkhdr rvclkhdr_277 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_277_io_l1clk),
    .io_clk(rvclkhdr_277_io_clk),
    .io_en(rvclkhdr_277_io_en),
    .io_scan_mode(rvclkhdr_277_io_scan_mode)
  );
  rvclkhdr rvclkhdr_278 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_278_io_l1clk),
    .io_clk(rvclkhdr_278_io_clk),
    .io_en(rvclkhdr_278_io_en),
    .io_scan_mode(rvclkhdr_278_io_scan_mode)
  );
  rvclkhdr rvclkhdr_279 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_279_io_l1clk),
    .io_clk(rvclkhdr_279_io_clk),
    .io_en(rvclkhdr_279_io_en),
    .io_scan_mode(rvclkhdr_279_io_scan_mode)
  );
  rvclkhdr rvclkhdr_280 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_280_io_l1clk),
    .io_clk(rvclkhdr_280_io_clk),
    .io_en(rvclkhdr_280_io_en),
    .io_scan_mode(rvclkhdr_280_io_scan_mode)
  );
  rvclkhdr rvclkhdr_281 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_281_io_l1clk),
    .io_clk(rvclkhdr_281_io_clk),
    .io_en(rvclkhdr_281_io_en),
    .io_scan_mode(rvclkhdr_281_io_scan_mode)
  );
  rvclkhdr rvclkhdr_282 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_282_io_l1clk),
    .io_clk(rvclkhdr_282_io_clk),
    .io_en(rvclkhdr_282_io_en),
    .io_scan_mode(rvclkhdr_282_io_scan_mode)
  );
  rvclkhdr rvclkhdr_283 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_283_io_l1clk),
    .io_clk(rvclkhdr_283_io_clk),
    .io_en(rvclkhdr_283_io_en),
    .io_scan_mode(rvclkhdr_283_io_scan_mode)
  );
  rvclkhdr rvclkhdr_284 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_284_io_l1clk),
    .io_clk(rvclkhdr_284_io_clk),
    .io_en(rvclkhdr_284_io_en),
    .io_scan_mode(rvclkhdr_284_io_scan_mode)
  );
  rvclkhdr rvclkhdr_285 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_285_io_l1clk),
    .io_clk(rvclkhdr_285_io_clk),
    .io_en(rvclkhdr_285_io_en),
    .io_scan_mode(rvclkhdr_285_io_scan_mode)
  );
  rvclkhdr rvclkhdr_286 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_286_io_l1clk),
    .io_clk(rvclkhdr_286_io_clk),
    .io_en(rvclkhdr_286_io_en),
    .io_scan_mode(rvclkhdr_286_io_scan_mode)
  );
  rvclkhdr rvclkhdr_287 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_287_io_l1clk),
    .io_clk(rvclkhdr_287_io_clk),
    .io_en(rvclkhdr_287_io_en),
    .io_scan_mode(rvclkhdr_287_io_scan_mode)
  );
  rvclkhdr rvclkhdr_288 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_288_io_l1clk),
    .io_clk(rvclkhdr_288_io_clk),
    .io_en(rvclkhdr_288_io_en),
    .io_scan_mode(rvclkhdr_288_io_scan_mode)
  );
  rvclkhdr rvclkhdr_289 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_289_io_l1clk),
    .io_clk(rvclkhdr_289_io_clk),
    .io_en(rvclkhdr_289_io_en),
    .io_scan_mode(rvclkhdr_289_io_scan_mode)
  );
  rvclkhdr rvclkhdr_290 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_290_io_l1clk),
    .io_clk(rvclkhdr_290_io_clk),
    .io_en(rvclkhdr_290_io_en),
    .io_scan_mode(rvclkhdr_290_io_scan_mode)
  );
  rvclkhdr rvclkhdr_291 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_291_io_l1clk),
    .io_clk(rvclkhdr_291_io_clk),
    .io_en(rvclkhdr_291_io_en),
    .io_scan_mode(rvclkhdr_291_io_scan_mode)
  );
  rvclkhdr rvclkhdr_292 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_292_io_l1clk),
    .io_clk(rvclkhdr_292_io_clk),
    .io_en(rvclkhdr_292_io_en),
    .io_scan_mode(rvclkhdr_292_io_scan_mode)
  );
  rvclkhdr rvclkhdr_293 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_293_io_l1clk),
    .io_clk(rvclkhdr_293_io_clk),
    .io_en(rvclkhdr_293_io_en),
    .io_scan_mode(rvclkhdr_293_io_scan_mode)
  );
  rvclkhdr rvclkhdr_294 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_294_io_l1clk),
    .io_clk(rvclkhdr_294_io_clk),
    .io_en(rvclkhdr_294_io_en),
    .io_scan_mode(rvclkhdr_294_io_scan_mode)
  );
  rvclkhdr rvclkhdr_295 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_295_io_l1clk),
    .io_clk(rvclkhdr_295_io_clk),
    .io_en(rvclkhdr_295_io_en),
    .io_scan_mode(rvclkhdr_295_io_scan_mode)
  );
  rvclkhdr rvclkhdr_296 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_296_io_l1clk),
    .io_clk(rvclkhdr_296_io_clk),
    .io_en(rvclkhdr_296_io_en),
    .io_scan_mode(rvclkhdr_296_io_scan_mode)
  );
  rvclkhdr rvclkhdr_297 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_297_io_l1clk),
    .io_clk(rvclkhdr_297_io_clk),
    .io_en(rvclkhdr_297_io_en),
    .io_scan_mode(rvclkhdr_297_io_scan_mode)
  );
  rvclkhdr rvclkhdr_298 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_298_io_l1clk),
    .io_clk(rvclkhdr_298_io_clk),
    .io_en(rvclkhdr_298_io_en),
    .io_scan_mode(rvclkhdr_298_io_scan_mode)
  );
  rvclkhdr rvclkhdr_299 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_299_io_l1clk),
    .io_clk(rvclkhdr_299_io_clk),
    .io_en(rvclkhdr_299_io_en),
    .io_scan_mode(rvclkhdr_299_io_scan_mode)
  );
  rvclkhdr rvclkhdr_300 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_300_io_l1clk),
    .io_clk(rvclkhdr_300_io_clk),
    .io_en(rvclkhdr_300_io_en),
    .io_scan_mode(rvclkhdr_300_io_scan_mode)
  );
  rvclkhdr rvclkhdr_301 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_301_io_l1clk),
    .io_clk(rvclkhdr_301_io_clk),
    .io_en(rvclkhdr_301_io_en),
    .io_scan_mode(rvclkhdr_301_io_scan_mode)
  );
  rvclkhdr rvclkhdr_302 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_302_io_l1clk),
    .io_clk(rvclkhdr_302_io_clk),
    .io_en(rvclkhdr_302_io_en),
    .io_scan_mode(rvclkhdr_302_io_scan_mode)
  );
  rvclkhdr rvclkhdr_303 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_303_io_l1clk),
    .io_clk(rvclkhdr_303_io_clk),
    .io_en(rvclkhdr_303_io_en),
    .io_scan_mode(rvclkhdr_303_io_scan_mode)
  );
  rvclkhdr rvclkhdr_304 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_304_io_l1clk),
    .io_clk(rvclkhdr_304_io_clk),
    .io_en(rvclkhdr_304_io_en),
    .io_scan_mode(rvclkhdr_304_io_scan_mode)
  );
  rvclkhdr rvclkhdr_305 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_305_io_l1clk),
    .io_clk(rvclkhdr_305_io_clk),
    .io_en(rvclkhdr_305_io_en),
    .io_scan_mode(rvclkhdr_305_io_scan_mode)
  );
  rvclkhdr rvclkhdr_306 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_306_io_l1clk),
    .io_clk(rvclkhdr_306_io_clk),
    .io_en(rvclkhdr_306_io_en),
    .io_scan_mode(rvclkhdr_306_io_scan_mode)
  );
  rvclkhdr rvclkhdr_307 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_307_io_l1clk),
    .io_clk(rvclkhdr_307_io_clk),
    .io_en(rvclkhdr_307_io_en),
    .io_scan_mode(rvclkhdr_307_io_scan_mode)
  );
  rvclkhdr rvclkhdr_308 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_308_io_l1clk),
    .io_clk(rvclkhdr_308_io_clk),
    .io_en(rvclkhdr_308_io_en),
    .io_scan_mode(rvclkhdr_308_io_scan_mode)
  );
  rvclkhdr rvclkhdr_309 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_309_io_l1clk),
    .io_clk(rvclkhdr_309_io_clk),
    .io_en(rvclkhdr_309_io_en),
    .io_scan_mode(rvclkhdr_309_io_scan_mode)
  );
  rvclkhdr rvclkhdr_310 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_310_io_l1clk),
    .io_clk(rvclkhdr_310_io_clk),
    .io_en(rvclkhdr_310_io_en),
    .io_scan_mode(rvclkhdr_310_io_scan_mode)
  );
  rvclkhdr rvclkhdr_311 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_311_io_l1clk),
    .io_clk(rvclkhdr_311_io_clk),
    .io_en(rvclkhdr_311_io_en),
    .io_scan_mode(rvclkhdr_311_io_scan_mode)
  );
  rvclkhdr rvclkhdr_312 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_312_io_l1clk),
    .io_clk(rvclkhdr_312_io_clk),
    .io_en(rvclkhdr_312_io_en),
    .io_scan_mode(rvclkhdr_312_io_scan_mode)
  );
  rvclkhdr rvclkhdr_313 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_313_io_l1clk),
    .io_clk(rvclkhdr_313_io_clk),
    .io_en(rvclkhdr_313_io_en),
    .io_scan_mode(rvclkhdr_313_io_scan_mode)
  );
  rvclkhdr rvclkhdr_314 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_314_io_l1clk),
    .io_clk(rvclkhdr_314_io_clk),
    .io_en(rvclkhdr_314_io_en),
    .io_scan_mode(rvclkhdr_314_io_scan_mode)
  );
  rvclkhdr rvclkhdr_315 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_315_io_l1clk),
    .io_clk(rvclkhdr_315_io_clk),
    .io_en(rvclkhdr_315_io_en),
    .io_scan_mode(rvclkhdr_315_io_scan_mode)
  );
  rvclkhdr rvclkhdr_316 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_316_io_l1clk),
    .io_clk(rvclkhdr_316_io_clk),
    .io_en(rvclkhdr_316_io_en),
    .io_scan_mode(rvclkhdr_316_io_scan_mode)
  );
  rvclkhdr rvclkhdr_317 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_317_io_l1clk),
    .io_clk(rvclkhdr_317_io_clk),
    .io_en(rvclkhdr_317_io_en),
    .io_scan_mode(rvclkhdr_317_io_scan_mode)
  );
  rvclkhdr rvclkhdr_318 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_318_io_l1clk),
    .io_clk(rvclkhdr_318_io_clk),
    .io_en(rvclkhdr_318_io_en),
    .io_scan_mode(rvclkhdr_318_io_scan_mode)
  );
  rvclkhdr rvclkhdr_319 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_319_io_l1clk),
    .io_clk(rvclkhdr_319_io_clk),
    .io_en(rvclkhdr_319_io_en),
    .io_scan_mode(rvclkhdr_319_io_scan_mode)
  );
  rvclkhdr rvclkhdr_320 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_320_io_l1clk),
    .io_clk(rvclkhdr_320_io_clk),
    .io_en(rvclkhdr_320_io_en),
    .io_scan_mode(rvclkhdr_320_io_scan_mode)
  );
  rvclkhdr rvclkhdr_321 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_321_io_l1clk),
    .io_clk(rvclkhdr_321_io_clk),
    .io_en(rvclkhdr_321_io_en),
    .io_scan_mode(rvclkhdr_321_io_scan_mode)
  );
  rvclkhdr rvclkhdr_322 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_322_io_l1clk),
    .io_clk(rvclkhdr_322_io_clk),
    .io_en(rvclkhdr_322_io_en),
    .io_scan_mode(rvclkhdr_322_io_scan_mode)
  );
  rvclkhdr rvclkhdr_323 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_323_io_l1clk),
    .io_clk(rvclkhdr_323_io_clk),
    .io_en(rvclkhdr_323_io_en),
    .io_scan_mode(rvclkhdr_323_io_scan_mode)
  );
  rvclkhdr rvclkhdr_324 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_324_io_l1clk),
    .io_clk(rvclkhdr_324_io_clk),
    .io_en(rvclkhdr_324_io_en),
    .io_scan_mode(rvclkhdr_324_io_scan_mode)
  );
  rvclkhdr rvclkhdr_325 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_325_io_l1clk),
    .io_clk(rvclkhdr_325_io_clk),
    .io_en(rvclkhdr_325_io_en),
    .io_scan_mode(rvclkhdr_325_io_scan_mode)
  );
  rvclkhdr rvclkhdr_326 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_326_io_l1clk),
    .io_clk(rvclkhdr_326_io_clk),
    .io_en(rvclkhdr_326_io_en),
    .io_scan_mode(rvclkhdr_326_io_scan_mode)
  );
  rvclkhdr rvclkhdr_327 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_327_io_l1clk),
    .io_clk(rvclkhdr_327_io_clk),
    .io_en(rvclkhdr_327_io_en),
    .io_scan_mode(rvclkhdr_327_io_scan_mode)
  );
  rvclkhdr rvclkhdr_328 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_328_io_l1clk),
    .io_clk(rvclkhdr_328_io_clk),
    .io_en(rvclkhdr_328_io_en),
    .io_scan_mode(rvclkhdr_328_io_scan_mode)
  );
  rvclkhdr rvclkhdr_329 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_329_io_l1clk),
    .io_clk(rvclkhdr_329_io_clk),
    .io_en(rvclkhdr_329_io_en),
    .io_scan_mode(rvclkhdr_329_io_scan_mode)
  );
  rvclkhdr rvclkhdr_330 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_330_io_l1clk),
    .io_clk(rvclkhdr_330_io_clk),
    .io_en(rvclkhdr_330_io_en),
    .io_scan_mode(rvclkhdr_330_io_scan_mode)
  );
  rvclkhdr rvclkhdr_331 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_331_io_l1clk),
    .io_clk(rvclkhdr_331_io_clk),
    .io_en(rvclkhdr_331_io_en),
    .io_scan_mode(rvclkhdr_331_io_scan_mode)
  );
  rvclkhdr rvclkhdr_332 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_332_io_l1clk),
    .io_clk(rvclkhdr_332_io_clk),
    .io_en(rvclkhdr_332_io_en),
    .io_scan_mode(rvclkhdr_332_io_scan_mode)
  );
  rvclkhdr rvclkhdr_333 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_333_io_l1clk),
    .io_clk(rvclkhdr_333_io_clk),
    .io_en(rvclkhdr_333_io_en),
    .io_scan_mode(rvclkhdr_333_io_scan_mode)
  );
  rvclkhdr rvclkhdr_334 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_334_io_l1clk),
    .io_clk(rvclkhdr_334_io_clk),
    .io_en(rvclkhdr_334_io_en),
    .io_scan_mode(rvclkhdr_334_io_scan_mode)
  );
  rvclkhdr rvclkhdr_335 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_335_io_l1clk),
    .io_clk(rvclkhdr_335_io_clk),
    .io_en(rvclkhdr_335_io_en),
    .io_scan_mode(rvclkhdr_335_io_scan_mode)
  );
  rvclkhdr rvclkhdr_336 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_336_io_l1clk),
    .io_clk(rvclkhdr_336_io_clk),
    .io_en(rvclkhdr_336_io_en),
    .io_scan_mode(rvclkhdr_336_io_scan_mode)
  );
  rvclkhdr rvclkhdr_337 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_337_io_l1clk),
    .io_clk(rvclkhdr_337_io_clk),
    .io_en(rvclkhdr_337_io_en),
    .io_scan_mode(rvclkhdr_337_io_scan_mode)
  );
  rvclkhdr rvclkhdr_338 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_338_io_l1clk),
    .io_clk(rvclkhdr_338_io_clk),
    .io_en(rvclkhdr_338_io_en),
    .io_scan_mode(rvclkhdr_338_io_scan_mode)
  );
  rvclkhdr rvclkhdr_339 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_339_io_l1clk),
    .io_clk(rvclkhdr_339_io_clk),
    .io_en(rvclkhdr_339_io_en),
    .io_scan_mode(rvclkhdr_339_io_scan_mode)
  );
  rvclkhdr rvclkhdr_340 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_340_io_l1clk),
    .io_clk(rvclkhdr_340_io_clk),
    .io_en(rvclkhdr_340_io_en),
    .io_scan_mode(rvclkhdr_340_io_scan_mode)
  );
  rvclkhdr rvclkhdr_341 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_341_io_l1clk),
    .io_clk(rvclkhdr_341_io_clk),
    .io_en(rvclkhdr_341_io_en),
    .io_scan_mode(rvclkhdr_341_io_scan_mode)
  );
  rvclkhdr rvclkhdr_342 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_342_io_l1clk),
    .io_clk(rvclkhdr_342_io_clk),
    .io_en(rvclkhdr_342_io_en),
    .io_scan_mode(rvclkhdr_342_io_scan_mode)
  );
  rvclkhdr rvclkhdr_343 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_343_io_l1clk),
    .io_clk(rvclkhdr_343_io_clk),
    .io_en(rvclkhdr_343_io_en),
    .io_scan_mode(rvclkhdr_343_io_scan_mode)
  );
  rvclkhdr rvclkhdr_344 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_344_io_l1clk),
    .io_clk(rvclkhdr_344_io_clk),
    .io_en(rvclkhdr_344_io_en),
    .io_scan_mode(rvclkhdr_344_io_scan_mode)
  );
  rvclkhdr rvclkhdr_345 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_345_io_l1clk),
    .io_clk(rvclkhdr_345_io_clk),
    .io_en(rvclkhdr_345_io_en),
    .io_scan_mode(rvclkhdr_345_io_scan_mode)
  );
  rvclkhdr rvclkhdr_346 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_346_io_l1clk),
    .io_clk(rvclkhdr_346_io_clk),
    .io_en(rvclkhdr_346_io_en),
    .io_scan_mode(rvclkhdr_346_io_scan_mode)
  );
  rvclkhdr rvclkhdr_347 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_347_io_l1clk),
    .io_clk(rvclkhdr_347_io_clk),
    .io_en(rvclkhdr_347_io_en),
    .io_scan_mode(rvclkhdr_347_io_scan_mode)
  );
  rvclkhdr rvclkhdr_348 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_348_io_l1clk),
    .io_clk(rvclkhdr_348_io_clk),
    .io_en(rvclkhdr_348_io_en),
    .io_scan_mode(rvclkhdr_348_io_scan_mode)
  );
  rvclkhdr rvclkhdr_349 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_349_io_l1clk),
    .io_clk(rvclkhdr_349_io_clk),
    .io_en(rvclkhdr_349_io_en),
    .io_scan_mode(rvclkhdr_349_io_scan_mode)
  );
  rvclkhdr rvclkhdr_350 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_350_io_l1clk),
    .io_clk(rvclkhdr_350_io_clk),
    .io_en(rvclkhdr_350_io_en),
    .io_scan_mode(rvclkhdr_350_io_scan_mode)
  );
  rvclkhdr rvclkhdr_351 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_351_io_l1clk),
    .io_clk(rvclkhdr_351_io_clk),
    .io_en(rvclkhdr_351_io_en),
    .io_scan_mode(rvclkhdr_351_io_scan_mode)
  );
  rvclkhdr rvclkhdr_352 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_352_io_l1clk),
    .io_clk(rvclkhdr_352_io_clk),
    .io_en(rvclkhdr_352_io_en),
    .io_scan_mode(rvclkhdr_352_io_scan_mode)
  );
  rvclkhdr rvclkhdr_353 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_353_io_l1clk),
    .io_clk(rvclkhdr_353_io_clk),
    .io_en(rvclkhdr_353_io_en),
    .io_scan_mode(rvclkhdr_353_io_scan_mode)
  );
  rvclkhdr rvclkhdr_354 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_354_io_l1clk),
    .io_clk(rvclkhdr_354_io_clk),
    .io_en(rvclkhdr_354_io_en),
    .io_scan_mode(rvclkhdr_354_io_scan_mode)
  );
  rvclkhdr rvclkhdr_355 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_355_io_l1clk),
    .io_clk(rvclkhdr_355_io_clk),
    .io_en(rvclkhdr_355_io_en),
    .io_scan_mode(rvclkhdr_355_io_scan_mode)
  );
  rvclkhdr rvclkhdr_356 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_356_io_l1clk),
    .io_clk(rvclkhdr_356_io_clk),
    .io_en(rvclkhdr_356_io_en),
    .io_scan_mode(rvclkhdr_356_io_scan_mode)
  );
  rvclkhdr rvclkhdr_357 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_357_io_l1clk),
    .io_clk(rvclkhdr_357_io_clk),
    .io_en(rvclkhdr_357_io_en),
    .io_scan_mode(rvclkhdr_357_io_scan_mode)
  );
  rvclkhdr rvclkhdr_358 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_358_io_l1clk),
    .io_clk(rvclkhdr_358_io_clk),
    .io_en(rvclkhdr_358_io_en),
    .io_scan_mode(rvclkhdr_358_io_scan_mode)
  );
  rvclkhdr rvclkhdr_359 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_359_io_l1clk),
    .io_clk(rvclkhdr_359_io_clk),
    .io_en(rvclkhdr_359_io_en),
    .io_scan_mode(rvclkhdr_359_io_scan_mode)
  );
  rvclkhdr rvclkhdr_360 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_360_io_l1clk),
    .io_clk(rvclkhdr_360_io_clk),
    .io_en(rvclkhdr_360_io_en),
    .io_scan_mode(rvclkhdr_360_io_scan_mode)
  );
  rvclkhdr rvclkhdr_361 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_361_io_l1clk),
    .io_clk(rvclkhdr_361_io_clk),
    .io_en(rvclkhdr_361_io_en),
    .io_scan_mode(rvclkhdr_361_io_scan_mode)
  );
  rvclkhdr rvclkhdr_362 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_362_io_l1clk),
    .io_clk(rvclkhdr_362_io_clk),
    .io_en(rvclkhdr_362_io_en),
    .io_scan_mode(rvclkhdr_362_io_scan_mode)
  );
  rvclkhdr rvclkhdr_363 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_363_io_l1clk),
    .io_clk(rvclkhdr_363_io_clk),
    .io_en(rvclkhdr_363_io_en),
    .io_scan_mode(rvclkhdr_363_io_scan_mode)
  );
  rvclkhdr rvclkhdr_364 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_364_io_l1clk),
    .io_clk(rvclkhdr_364_io_clk),
    .io_en(rvclkhdr_364_io_en),
    .io_scan_mode(rvclkhdr_364_io_scan_mode)
  );
  rvclkhdr rvclkhdr_365 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_365_io_l1clk),
    .io_clk(rvclkhdr_365_io_clk),
    .io_en(rvclkhdr_365_io_en),
    .io_scan_mode(rvclkhdr_365_io_scan_mode)
  );
  rvclkhdr rvclkhdr_366 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_366_io_l1clk),
    .io_clk(rvclkhdr_366_io_clk),
    .io_en(rvclkhdr_366_io_en),
    .io_scan_mode(rvclkhdr_366_io_scan_mode)
  );
  rvclkhdr rvclkhdr_367 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_367_io_l1clk),
    .io_clk(rvclkhdr_367_io_clk),
    .io_en(rvclkhdr_367_io_en),
    .io_scan_mode(rvclkhdr_367_io_scan_mode)
  );
  rvclkhdr rvclkhdr_368 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_368_io_l1clk),
    .io_clk(rvclkhdr_368_io_clk),
    .io_en(rvclkhdr_368_io_en),
    .io_scan_mode(rvclkhdr_368_io_scan_mode)
  );
  rvclkhdr rvclkhdr_369 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_369_io_l1clk),
    .io_clk(rvclkhdr_369_io_clk),
    .io_en(rvclkhdr_369_io_en),
    .io_scan_mode(rvclkhdr_369_io_scan_mode)
  );
  rvclkhdr rvclkhdr_370 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_370_io_l1clk),
    .io_clk(rvclkhdr_370_io_clk),
    .io_en(rvclkhdr_370_io_en),
    .io_scan_mode(rvclkhdr_370_io_scan_mode)
  );
  rvclkhdr rvclkhdr_371 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_371_io_l1clk),
    .io_clk(rvclkhdr_371_io_clk),
    .io_en(rvclkhdr_371_io_en),
    .io_scan_mode(rvclkhdr_371_io_scan_mode)
  );
  rvclkhdr rvclkhdr_372 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_372_io_l1clk),
    .io_clk(rvclkhdr_372_io_clk),
    .io_en(rvclkhdr_372_io_en),
    .io_scan_mode(rvclkhdr_372_io_scan_mode)
  );
  rvclkhdr rvclkhdr_373 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_373_io_l1clk),
    .io_clk(rvclkhdr_373_io_clk),
    .io_en(rvclkhdr_373_io_en),
    .io_scan_mode(rvclkhdr_373_io_scan_mode)
  );
  rvclkhdr rvclkhdr_374 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_374_io_l1clk),
    .io_clk(rvclkhdr_374_io_clk),
    .io_en(rvclkhdr_374_io_en),
    .io_scan_mode(rvclkhdr_374_io_scan_mode)
  );
  rvclkhdr rvclkhdr_375 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_375_io_l1clk),
    .io_clk(rvclkhdr_375_io_clk),
    .io_en(rvclkhdr_375_io_en),
    .io_scan_mode(rvclkhdr_375_io_scan_mode)
  );
  rvclkhdr rvclkhdr_376 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_376_io_l1clk),
    .io_clk(rvclkhdr_376_io_clk),
    .io_en(rvclkhdr_376_io_en),
    .io_scan_mode(rvclkhdr_376_io_scan_mode)
  );
  rvclkhdr rvclkhdr_377 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_377_io_l1clk),
    .io_clk(rvclkhdr_377_io_clk),
    .io_en(rvclkhdr_377_io_en),
    .io_scan_mode(rvclkhdr_377_io_scan_mode)
  );
  rvclkhdr rvclkhdr_378 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_378_io_l1clk),
    .io_clk(rvclkhdr_378_io_clk),
    .io_en(rvclkhdr_378_io_en),
    .io_scan_mode(rvclkhdr_378_io_scan_mode)
  );
  rvclkhdr rvclkhdr_379 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_379_io_l1clk),
    .io_clk(rvclkhdr_379_io_clk),
    .io_en(rvclkhdr_379_io_en),
    .io_scan_mode(rvclkhdr_379_io_scan_mode)
  );
  rvclkhdr rvclkhdr_380 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_380_io_l1clk),
    .io_clk(rvclkhdr_380_io_clk),
    .io_en(rvclkhdr_380_io_en),
    .io_scan_mode(rvclkhdr_380_io_scan_mode)
  );
  rvclkhdr rvclkhdr_381 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_381_io_l1clk),
    .io_clk(rvclkhdr_381_io_clk),
    .io_en(rvclkhdr_381_io_en),
    .io_scan_mode(rvclkhdr_381_io_scan_mode)
  );
  rvclkhdr rvclkhdr_382 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_382_io_l1clk),
    .io_clk(rvclkhdr_382_io_clk),
    .io_en(rvclkhdr_382_io_en),
    .io_scan_mode(rvclkhdr_382_io_scan_mode)
  );
  rvclkhdr rvclkhdr_383 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_383_io_l1clk),
    .io_clk(rvclkhdr_383_io_clk),
    .io_en(rvclkhdr_383_io_en),
    .io_scan_mode(rvclkhdr_383_io_scan_mode)
  );
  rvclkhdr rvclkhdr_384 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_384_io_l1clk),
    .io_clk(rvclkhdr_384_io_clk),
    .io_en(rvclkhdr_384_io_en),
    .io_scan_mode(rvclkhdr_384_io_scan_mode)
  );
  rvclkhdr rvclkhdr_385 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_385_io_l1clk),
    .io_clk(rvclkhdr_385_io_clk),
    .io_en(rvclkhdr_385_io_en),
    .io_scan_mode(rvclkhdr_385_io_scan_mode)
  );
  rvclkhdr rvclkhdr_386 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_386_io_l1clk),
    .io_clk(rvclkhdr_386_io_clk),
    .io_en(rvclkhdr_386_io_en),
    .io_scan_mode(rvclkhdr_386_io_scan_mode)
  );
  rvclkhdr rvclkhdr_387 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_387_io_l1clk),
    .io_clk(rvclkhdr_387_io_clk),
    .io_en(rvclkhdr_387_io_en),
    .io_scan_mode(rvclkhdr_387_io_scan_mode)
  );
  rvclkhdr rvclkhdr_388 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_388_io_l1clk),
    .io_clk(rvclkhdr_388_io_clk),
    .io_en(rvclkhdr_388_io_en),
    .io_scan_mode(rvclkhdr_388_io_scan_mode)
  );
  rvclkhdr rvclkhdr_389 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_389_io_l1clk),
    .io_clk(rvclkhdr_389_io_clk),
    .io_en(rvclkhdr_389_io_en),
    .io_scan_mode(rvclkhdr_389_io_scan_mode)
  );
  rvclkhdr rvclkhdr_390 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_390_io_l1clk),
    .io_clk(rvclkhdr_390_io_clk),
    .io_en(rvclkhdr_390_io_en),
    .io_scan_mode(rvclkhdr_390_io_scan_mode)
  );
  rvclkhdr rvclkhdr_391 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_391_io_l1clk),
    .io_clk(rvclkhdr_391_io_clk),
    .io_en(rvclkhdr_391_io_en),
    .io_scan_mode(rvclkhdr_391_io_scan_mode)
  );
  rvclkhdr rvclkhdr_392 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_392_io_l1clk),
    .io_clk(rvclkhdr_392_io_clk),
    .io_en(rvclkhdr_392_io_en),
    .io_scan_mode(rvclkhdr_392_io_scan_mode)
  );
  rvclkhdr rvclkhdr_393 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_393_io_l1clk),
    .io_clk(rvclkhdr_393_io_clk),
    .io_en(rvclkhdr_393_io_en),
    .io_scan_mode(rvclkhdr_393_io_scan_mode)
  );
  rvclkhdr rvclkhdr_394 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_394_io_l1clk),
    .io_clk(rvclkhdr_394_io_clk),
    .io_en(rvclkhdr_394_io_en),
    .io_scan_mode(rvclkhdr_394_io_scan_mode)
  );
  rvclkhdr rvclkhdr_395 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_395_io_l1clk),
    .io_clk(rvclkhdr_395_io_clk),
    .io_en(rvclkhdr_395_io_en),
    .io_scan_mode(rvclkhdr_395_io_scan_mode)
  );
  rvclkhdr rvclkhdr_396 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_396_io_l1clk),
    .io_clk(rvclkhdr_396_io_clk),
    .io_en(rvclkhdr_396_io_en),
    .io_scan_mode(rvclkhdr_396_io_scan_mode)
  );
  rvclkhdr rvclkhdr_397 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_397_io_l1clk),
    .io_clk(rvclkhdr_397_io_clk),
    .io_en(rvclkhdr_397_io_en),
    .io_scan_mode(rvclkhdr_397_io_scan_mode)
  );
  rvclkhdr rvclkhdr_398 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_398_io_l1clk),
    .io_clk(rvclkhdr_398_io_clk),
    .io_en(rvclkhdr_398_io_en),
    .io_scan_mode(rvclkhdr_398_io_scan_mode)
  );
  rvclkhdr rvclkhdr_399 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_399_io_l1clk),
    .io_clk(rvclkhdr_399_io_clk),
    .io_en(rvclkhdr_399_io_en),
    .io_scan_mode(rvclkhdr_399_io_scan_mode)
  );
  rvclkhdr rvclkhdr_400 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_400_io_l1clk),
    .io_clk(rvclkhdr_400_io_clk),
    .io_en(rvclkhdr_400_io_en),
    .io_scan_mode(rvclkhdr_400_io_scan_mode)
  );
  rvclkhdr rvclkhdr_401 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_401_io_l1clk),
    .io_clk(rvclkhdr_401_io_clk),
    .io_en(rvclkhdr_401_io_en),
    .io_scan_mode(rvclkhdr_401_io_scan_mode)
  );
  rvclkhdr rvclkhdr_402 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_402_io_l1clk),
    .io_clk(rvclkhdr_402_io_clk),
    .io_en(rvclkhdr_402_io_en),
    .io_scan_mode(rvclkhdr_402_io_scan_mode)
  );
  rvclkhdr rvclkhdr_403 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_403_io_l1clk),
    .io_clk(rvclkhdr_403_io_clk),
    .io_en(rvclkhdr_403_io_en),
    .io_scan_mode(rvclkhdr_403_io_scan_mode)
  );
  rvclkhdr rvclkhdr_404 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_404_io_l1clk),
    .io_clk(rvclkhdr_404_io_clk),
    .io_en(rvclkhdr_404_io_en),
    .io_scan_mode(rvclkhdr_404_io_scan_mode)
  );
  rvclkhdr rvclkhdr_405 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_405_io_l1clk),
    .io_clk(rvclkhdr_405_io_clk),
    .io_en(rvclkhdr_405_io_en),
    .io_scan_mode(rvclkhdr_405_io_scan_mode)
  );
  rvclkhdr rvclkhdr_406 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_406_io_l1clk),
    .io_clk(rvclkhdr_406_io_clk),
    .io_en(rvclkhdr_406_io_en),
    .io_scan_mode(rvclkhdr_406_io_scan_mode)
  );
  rvclkhdr rvclkhdr_407 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_407_io_l1clk),
    .io_clk(rvclkhdr_407_io_clk),
    .io_en(rvclkhdr_407_io_en),
    .io_scan_mode(rvclkhdr_407_io_scan_mode)
  );
  rvclkhdr rvclkhdr_408 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_408_io_l1clk),
    .io_clk(rvclkhdr_408_io_clk),
    .io_en(rvclkhdr_408_io_en),
    .io_scan_mode(rvclkhdr_408_io_scan_mode)
  );
  rvclkhdr rvclkhdr_409 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_409_io_l1clk),
    .io_clk(rvclkhdr_409_io_clk),
    .io_en(rvclkhdr_409_io_en),
    .io_scan_mode(rvclkhdr_409_io_scan_mode)
  );
  rvclkhdr rvclkhdr_410 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_410_io_l1clk),
    .io_clk(rvclkhdr_410_io_clk),
    .io_en(rvclkhdr_410_io_en),
    .io_scan_mode(rvclkhdr_410_io_scan_mode)
  );
  rvclkhdr rvclkhdr_411 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_411_io_l1clk),
    .io_clk(rvclkhdr_411_io_clk),
    .io_en(rvclkhdr_411_io_en),
    .io_scan_mode(rvclkhdr_411_io_scan_mode)
  );
  rvclkhdr rvclkhdr_412 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_412_io_l1clk),
    .io_clk(rvclkhdr_412_io_clk),
    .io_en(rvclkhdr_412_io_en),
    .io_scan_mode(rvclkhdr_412_io_scan_mode)
  );
  rvclkhdr rvclkhdr_413 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_413_io_l1clk),
    .io_clk(rvclkhdr_413_io_clk),
    .io_en(rvclkhdr_413_io_en),
    .io_scan_mode(rvclkhdr_413_io_scan_mode)
  );
  rvclkhdr rvclkhdr_414 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_414_io_l1clk),
    .io_clk(rvclkhdr_414_io_clk),
    .io_en(rvclkhdr_414_io_en),
    .io_scan_mode(rvclkhdr_414_io_scan_mode)
  );
  rvclkhdr rvclkhdr_415 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_415_io_l1clk),
    .io_clk(rvclkhdr_415_io_clk),
    .io_en(rvclkhdr_415_io_en),
    .io_scan_mode(rvclkhdr_415_io_scan_mode)
  );
  rvclkhdr rvclkhdr_416 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_416_io_l1clk),
    .io_clk(rvclkhdr_416_io_clk),
    .io_en(rvclkhdr_416_io_en),
    .io_scan_mode(rvclkhdr_416_io_scan_mode)
  );
  rvclkhdr rvclkhdr_417 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_417_io_l1clk),
    .io_clk(rvclkhdr_417_io_clk),
    .io_en(rvclkhdr_417_io_en),
    .io_scan_mode(rvclkhdr_417_io_scan_mode)
  );
  rvclkhdr rvclkhdr_418 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_418_io_l1clk),
    .io_clk(rvclkhdr_418_io_clk),
    .io_en(rvclkhdr_418_io_en),
    .io_scan_mode(rvclkhdr_418_io_scan_mode)
  );
  rvclkhdr rvclkhdr_419 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_419_io_l1clk),
    .io_clk(rvclkhdr_419_io_clk),
    .io_en(rvclkhdr_419_io_en),
    .io_scan_mode(rvclkhdr_419_io_scan_mode)
  );
  rvclkhdr rvclkhdr_420 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_420_io_l1clk),
    .io_clk(rvclkhdr_420_io_clk),
    .io_en(rvclkhdr_420_io_en),
    .io_scan_mode(rvclkhdr_420_io_scan_mode)
  );
  rvclkhdr rvclkhdr_421 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_421_io_l1clk),
    .io_clk(rvclkhdr_421_io_clk),
    .io_en(rvclkhdr_421_io_en),
    .io_scan_mode(rvclkhdr_421_io_scan_mode)
  );
  rvclkhdr rvclkhdr_422 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_422_io_l1clk),
    .io_clk(rvclkhdr_422_io_clk),
    .io_en(rvclkhdr_422_io_en),
    .io_scan_mode(rvclkhdr_422_io_scan_mode)
  );
  rvclkhdr rvclkhdr_423 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_423_io_l1clk),
    .io_clk(rvclkhdr_423_io_clk),
    .io_en(rvclkhdr_423_io_en),
    .io_scan_mode(rvclkhdr_423_io_scan_mode)
  );
  rvclkhdr rvclkhdr_424 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_424_io_l1clk),
    .io_clk(rvclkhdr_424_io_clk),
    .io_en(rvclkhdr_424_io_en),
    .io_scan_mode(rvclkhdr_424_io_scan_mode)
  );
  rvclkhdr rvclkhdr_425 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_425_io_l1clk),
    .io_clk(rvclkhdr_425_io_clk),
    .io_en(rvclkhdr_425_io_en),
    .io_scan_mode(rvclkhdr_425_io_scan_mode)
  );
  rvclkhdr rvclkhdr_426 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_426_io_l1clk),
    .io_clk(rvclkhdr_426_io_clk),
    .io_en(rvclkhdr_426_io_en),
    .io_scan_mode(rvclkhdr_426_io_scan_mode)
  );
  rvclkhdr rvclkhdr_427 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_427_io_l1clk),
    .io_clk(rvclkhdr_427_io_clk),
    .io_en(rvclkhdr_427_io_en),
    .io_scan_mode(rvclkhdr_427_io_scan_mode)
  );
  rvclkhdr rvclkhdr_428 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_428_io_l1clk),
    .io_clk(rvclkhdr_428_io_clk),
    .io_en(rvclkhdr_428_io_en),
    .io_scan_mode(rvclkhdr_428_io_scan_mode)
  );
  rvclkhdr rvclkhdr_429 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_429_io_l1clk),
    .io_clk(rvclkhdr_429_io_clk),
    .io_en(rvclkhdr_429_io_en),
    .io_scan_mode(rvclkhdr_429_io_scan_mode)
  );
  rvclkhdr rvclkhdr_430 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_430_io_l1clk),
    .io_clk(rvclkhdr_430_io_clk),
    .io_en(rvclkhdr_430_io_en),
    .io_scan_mode(rvclkhdr_430_io_scan_mode)
  );
  rvclkhdr rvclkhdr_431 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_431_io_l1clk),
    .io_clk(rvclkhdr_431_io_clk),
    .io_en(rvclkhdr_431_io_en),
    .io_scan_mode(rvclkhdr_431_io_scan_mode)
  );
  rvclkhdr rvclkhdr_432 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_432_io_l1clk),
    .io_clk(rvclkhdr_432_io_clk),
    .io_en(rvclkhdr_432_io_en),
    .io_scan_mode(rvclkhdr_432_io_scan_mode)
  );
  rvclkhdr rvclkhdr_433 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_433_io_l1clk),
    .io_clk(rvclkhdr_433_io_clk),
    .io_en(rvclkhdr_433_io_en),
    .io_scan_mode(rvclkhdr_433_io_scan_mode)
  );
  rvclkhdr rvclkhdr_434 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_434_io_l1clk),
    .io_clk(rvclkhdr_434_io_clk),
    .io_en(rvclkhdr_434_io_en),
    .io_scan_mode(rvclkhdr_434_io_scan_mode)
  );
  rvclkhdr rvclkhdr_435 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_435_io_l1clk),
    .io_clk(rvclkhdr_435_io_clk),
    .io_en(rvclkhdr_435_io_en),
    .io_scan_mode(rvclkhdr_435_io_scan_mode)
  );
  rvclkhdr rvclkhdr_436 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_436_io_l1clk),
    .io_clk(rvclkhdr_436_io_clk),
    .io_en(rvclkhdr_436_io_en),
    .io_scan_mode(rvclkhdr_436_io_scan_mode)
  );
  rvclkhdr rvclkhdr_437 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_437_io_l1clk),
    .io_clk(rvclkhdr_437_io_clk),
    .io_en(rvclkhdr_437_io_en),
    .io_scan_mode(rvclkhdr_437_io_scan_mode)
  );
  rvclkhdr rvclkhdr_438 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_438_io_l1clk),
    .io_clk(rvclkhdr_438_io_clk),
    .io_en(rvclkhdr_438_io_en),
    .io_scan_mode(rvclkhdr_438_io_scan_mode)
  );
  rvclkhdr rvclkhdr_439 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_439_io_l1clk),
    .io_clk(rvclkhdr_439_io_clk),
    .io_en(rvclkhdr_439_io_en),
    .io_scan_mode(rvclkhdr_439_io_scan_mode)
  );
  rvclkhdr rvclkhdr_440 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_440_io_l1clk),
    .io_clk(rvclkhdr_440_io_clk),
    .io_en(rvclkhdr_440_io_en),
    .io_scan_mode(rvclkhdr_440_io_scan_mode)
  );
  rvclkhdr rvclkhdr_441 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_441_io_l1clk),
    .io_clk(rvclkhdr_441_io_clk),
    .io_en(rvclkhdr_441_io_en),
    .io_scan_mode(rvclkhdr_441_io_scan_mode)
  );
  rvclkhdr rvclkhdr_442 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_442_io_l1clk),
    .io_clk(rvclkhdr_442_io_clk),
    .io_en(rvclkhdr_442_io_en),
    .io_scan_mode(rvclkhdr_442_io_scan_mode)
  );
  rvclkhdr rvclkhdr_443 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_443_io_l1clk),
    .io_clk(rvclkhdr_443_io_clk),
    .io_en(rvclkhdr_443_io_en),
    .io_scan_mode(rvclkhdr_443_io_scan_mode)
  );
  rvclkhdr rvclkhdr_444 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_444_io_l1clk),
    .io_clk(rvclkhdr_444_io_clk),
    .io_en(rvclkhdr_444_io_en),
    .io_scan_mode(rvclkhdr_444_io_scan_mode)
  );
  rvclkhdr rvclkhdr_445 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_445_io_l1clk),
    .io_clk(rvclkhdr_445_io_clk),
    .io_en(rvclkhdr_445_io_en),
    .io_scan_mode(rvclkhdr_445_io_scan_mode)
  );
  rvclkhdr rvclkhdr_446 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_446_io_l1clk),
    .io_clk(rvclkhdr_446_io_clk),
    .io_en(rvclkhdr_446_io_en),
    .io_scan_mode(rvclkhdr_446_io_scan_mode)
  );
  rvclkhdr rvclkhdr_447 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_447_io_l1clk),
    .io_clk(rvclkhdr_447_io_clk),
    .io_en(rvclkhdr_447_io_en),
    .io_scan_mode(rvclkhdr_447_io_scan_mode)
  );
  rvclkhdr rvclkhdr_448 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_448_io_l1clk),
    .io_clk(rvclkhdr_448_io_clk),
    .io_en(rvclkhdr_448_io_en),
    .io_scan_mode(rvclkhdr_448_io_scan_mode)
  );
  rvclkhdr rvclkhdr_449 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_449_io_l1clk),
    .io_clk(rvclkhdr_449_io_clk),
    .io_en(rvclkhdr_449_io_en),
    .io_scan_mode(rvclkhdr_449_io_scan_mode)
  );
  rvclkhdr rvclkhdr_450 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_450_io_l1clk),
    .io_clk(rvclkhdr_450_io_clk),
    .io_en(rvclkhdr_450_io_en),
    .io_scan_mode(rvclkhdr_450_io_scan_mode)
  );
  rvclkhdr rvclkhdr_451 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_451_io_l1clk),
    .io_clk(rvclkhdr_451_io_clk),
    .io_en(rvclkhdr_451_io_en),
    .io_scan_mode(rvclkhdr_451_io_scan_mode)
  );
  rvclkhdr rvclkhdr_452 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_452_io_l1clk),
    .io_clk(rvclkhdr_452_io_clk),
    .io_en(rvclkhdr_452_io_en),
    .io_scan_mode(rvclkhdr_452_io_scan_mode)
  );
  rvclkhdr rvclkhdr_453 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_453_io_l1clk),
    .io_clk(rvclkhdr_453_io_clk),
    .io_en(rvclkhdr_453_io_en),
    .io_scan_mode(rvclkhdr_453_io_scan_mode)
  );
  rvclkhdr rvclkhdr_454 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_454_io_l1clk),
    .io_clk(rvclkhdr_454_io_clk),
    .io_en(rvclkhdr_454_io_en),
    .io_scan_mode(rvclkhdr_454_io_scan_mode)
  );
  rvclkhdr rvclkhdr_455 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_455_io_l1clk),
    .io_clk(rvclkhdr_455_io_clk),
    .io_en(rvclkhdr_455_io_en),
    .io_scan_mode(rvclkhdr_455_io_scan_mode)
  );
  rvclkhdr rvclkhdr_456 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_456_io_l1clk),
    .io_clk(rvclkhdr_456_io_clk),
    .io_en(rvclkhdr_456_io_en),
    .io_scan_mode(rvclkhdr_456_io_scan_mode)
  );
  rvclkhdr rvclkhdr_457 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_457_io_l1clk),
    .io_clk(rvclkhdr_457_io_clk),
    .io_en(rvclkhdr_457_io_en),
    .io_scan_mode(rvclkhdr_457_io_scan_mode)
  );
  rvclkhdr rvclkhdr_458 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_458_io_l1clk),
    .io_clk(rvclkhdr_458_io_clk),
    .io_en(rvclkhdr_458_io_en),
    .io_scan_mode(rvclkhdr_458_io_scan_mode)
  );
  rvclkhdr rvclkhdr_459 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_459_io_l1clk),
    .io_clk(rvclkhdr_459_io_clk),
    .io_en(rvclkhdr_459_io_en),
    .io_scan_mode(rvclkhdr_459_io_scan_mode)
  );
  rvclkhdr rvclkhdr_460 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_460_io_l1clk),
    .io_clk(rvclkhdr_460_io_clk),
    .io_en(rvclkhdr_460_io_en),
    .io_scan_mode(rvclkhdr_460_io_scan_mode)
  );
  rvclkhdr rvclkhdr_461 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_461_io_l1clk),
    .io_clk(rvclkhdr_461_io_clk),
    .io_en(rvclkhdr_461_io_en),
    .io_scan_mode(rvclkhdr_461_io_scan_mode)
  );
  rvclkhdr rvclkhdr_462 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_462_io_l1clk),
    .io_clk(rvclkhdr_462_io_clk),
    .io_en(rvclkhdr_462_io_en),
    .io_scan_mode(rvclkhdr_462_io_scan_mode)
  );
  rvclkhdr rvclkhdr_463 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_463_io_l1clk),
    .io_clk(rvclkhdr_463_io_clk),
    .io_en(rvclkhdr_463_io_en),
    .io_scan_mode(rvclkhdr_463_io_scan_mode)
  );
  rvclkhdr rvclkhdr_464 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_464_io_l1clk),
    .io_clk(rvclkhdr_464_io_clk),
    .io_en(rvclkhdr_464_io_en),
    .io_scan_mode(rvclkhdr_464_io_scan_mode)
  );
  rvclkhdr rvclkhdr_465 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_465_io_l1clk),
    .io_clk(rvclkhdr_465_io_clk),
    .io_en(rvclkhdr_465_io_en),
    .io_scan_mode(rvclkhdr_465_io_scan_mode)
  );
  rvclkhdr rvclkhdr_466 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_466_io_l1clk),
    .io_clk(rvclkhdr_466_io_clk),
    .io_en(rvclkhdr_466_io_en),
    .io_scan_mode(rvclkhdr_466_io_scan_mode)
  );
  rvclkhdr rvclkhdr_467 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_467_io_l1clk),
    .io_clk(rvclkhdr_467_io_clk),
    .io_en(rvclkhdr_467_io_en),
    .io_scan_mode(rvclkhdr_467_io_scan_mode)
  );
  rvclkhdr rvclkhdr_468 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_468_io_l1clk),
    .io_clk(rvclkhdr_468_io_clk),
    .io_en(rvclkhdr_468_io_en),
    .io_scan_mode(rvclkhdr_468_io_scan_mode)
  );
  rvclkhdr rvclkhdr_469 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_469_io_l1clk),
    .io_clk(rvclkhdr_469_io_clk),
    .io_en(rvclkhdr_469_io_en),
    .io_scan_mode(rvclkhdr_469_io_scan_mode)
  );
  rvclkhdr rvclkhdr_470 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_470_io_l1clk),
    .io_clk(rvclkhdr_470_io_clk),
    .io_en(rvclkhdr_470_io_en),
    .io_scan_mode(rvclkhdr_470_io_scan_mode)
  );
  rvclkhdr rvclkhdr_471 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_471_io_l1clk),
    .io_clk(rvclkhdr_471_io_clk),
    .io_en(rvclkhdr_471_io_en),
    .io_scan_mode(rvclkhdr_471_io_scan_mode)
  );
  rvclkhdr rvclkhdr_472 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_472_io_l1clk),
    .io_clk(rvclkhdr_472_io_clk),
    .io_en(rvclkhdr_472_io_en),
    .io_scan_mode(rvclkhdr_472_io_scan_mode)
  );
  rvclkhdr rvclkhdr_473 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_473_io_l1clk),
    .io_clk(rvclkhdr_473_io_clk),
    .io_en(rvclkhdr_473_io_en),
    .io_scan_mode(rvclkhdr_473_io_scan_mode)
  );
  rvclkhdr rvclkhdr_474 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_474_io_l1clk),
    .io_clk(rvclkhdr_474_io_clk),
    .io_en(rvclkhdr_474_io_en),
    .io_scan_mode(rvclkhdr_474_io_scan_mode)
  );
  rvclkhdr rvclkhdr_475 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_475_io_l1clk),
    .io_clk(rvclkhdr_475_io_clk),
    .io_en(rvclkhdr_475_io_en),
    .io_scan_mode(rvclkhdr_475_io_scan_mode)
  );
  rvclkhdr rvclkhdr_476 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_476_io_l1clk),
    .io_clk(rvclkhdr_476_io_clk),
    .io_en(rvclkhdr_476_io_en),
    .io_scan_mode(rvclkhdr_476_io_scan_mode)
  );
  rvclkhdr rvclkhdr_477 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_477_io_l1clk),
    .io_clk(rvclkhdr_477_io_clk),
    .io_en(rvclkhdr_477_io_en),
    .io_scan_mode(rvclkhdr_477_io_scan_mode)
  );
  rvclkhdr rvclkhdr_478 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_478_io_l1clk),
    .io_clk(rvclkhdr_478_io_clk),
    .io_en(rvclkhdr_478_io_en),
    .io_scan_mode(rvclkhdr_478_io_scan_mode)
  );
  rvclkhdr rvclkhdr_479 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_479_io_l1clk),
    .io_clk(rvclkhdr_479_io_clk),
    .io_en(rvclkhdr_479_io_en),
    .io_scan_mode(rvclkhdr_479_io_scan_mode)
  );
  rvclkhdr rvclkhdr_480 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_480_io_l1clk),
    .io_clk(rvclkhdr_480_io_clk),
    .io_en(rvclkhdr_480_io_en),
    .io_scan_mode(rvclkhdr_480_io_scan_mode)
  );
  rvclkhdr rvclkhdr_481 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_481_io_l1clk),
    .io_clk(rvclkhdr_481_io_clk),
    .io_en(rvclkhdr_481_io_en),
    .io_scan_mode(rvclkhdr_481_io_scan_mode)
  );
  rvclkhdr rvclkhdr_482 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_482_io_l1clk),
    .io_clk(rvclkhdr_482_io_clk),
    .io_en(rvclkhdr_482_io_en),
    .io_scan_mode(rvclkhdr_482_io_scan_mode)
  );
  rvclkhdr rvclkhdr_483 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_483_io_l1clk),
    .io_clk(rvclkhdr_483_io_clk),
    .io_en(rvclkhdr_483_io_en),
    .io_scan_mode(rvclkhdr_483_io_scan_mode)
  );
  rvclkhdr rvclkhdr_484 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_484_io_l1clk),
    .io_clk(rvclkhdr_484_io_clk),
    .io_en(rvclkhdr_484_io_en),
    .io_scan_mode(rvclkhdr_484_io_scan_mode)
  );
  rvclkhdr rvclkhdr_485 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_485_io_l1clk),
    .io_clk(rvclkhdr_485_io_clk),
    .io_en(rvclkhdr_485_io_en),
    .io_scan_mode(rvclkhdr_485_io_scan_mode)
  );
  rvclkhdr rvclkhdr_486 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_486_io_l1clk),
    .io_clk(rvclkhdr_486_io_clk),
    .io_en(rvclkhdr_486_io_en),
    .io_scan_mode(rvclkhdr_486_io_scan_mode)
  );
  rvclkhdr rvclkhdr_487 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_487_io_l1clk),
    .io_clk(rvclkhdr_487_io_clk),
    .io_en(rvclkhdr_487_io_en),
    .io_scan_mode(rvclkhdr_487_io_scan_mode)
  );
  rvclkhdr rvclkhdr_488 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_488_io_l1clk),
    .io_clk(rvclkhdr_488_io_clk),
    .io_en(rvclkhdr_488_io_en),
    .io_scan_mode(rvclkhdr_488_io_scan_mode)
  );
  rvclkhdr rvclkhdr_489 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_489_io_l1clk),
    .io_clk(rvclkhdr_489_io_clk),
    .io_en(rvclkhdr_489_io_en),
    .io_scan_mode(rvclkhdr_489_io_scan_mode)
  );
  rvclkhdr rvclkhdr_490 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_490_io_l1clk),
    .io_clk(rvclkhdr_490_io_clk),
    .io_en(rvclkhdr_490_io_en),
    .io_scan_mode(rvclkhdr_490_io_scan_mode)
  );
  rvclkhdr rvclkhdr_491 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_491_io_l1clk),
    .io_clk(rvclkhdr_491_io_clk),
    .io_en(rvclkhdr_491_io_en),
    .io_scan_mode(rvclkhdr_491_io_scan_mode)
  );
  rvclkhdr rvclkhdr_492 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_492_io_l1clk),
    .io_clk(rvclkhdr_492_io_clk),
    .io_en(rvclkhdr_492_io_en),
    .io_scan_mode(rvclkhdr_492_io_scan_mode)
  );
  rvclkhdr rvclkhdr_493 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_493_io_l1clk),
    .io_clk(rvclkhdr_493_io_clk),
    .io_en(rvclkhdr_493_io_en),
    .io_scan_mode(rvclkhdr_493_io_scan_mode)
  );
  rvclkhdr rvclkhdr_494 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_494_io_l1clk),
    .io_clk(rvclkhdr_494_io_clk),
    .io_en(rvclkhdr_494_io_en),
    .io_scan_mode(rvclkhdr_494_io_scan_mode)
  );
  rvclkhdr rvclkhdr_495 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_495_io_l1clk),
    .io_clk(rvclkhdr_495_io_clk),
    .io_en(rvclkhdr_495_io_en),
    .io_scan_mode(rvclkhdr_495_io_scan_mode)
  );
  rvclkhdr rvclkhdr_496 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_496_io_l1clk),
    .io_clk(rvclkhdr_496_io_clk),
    .io_en(rvclkhdr_496_io_en),
    .io_scan_mode(rvclkhdr_496_io_scan_mode)
  );
  rvclkhdr rvclkhdr_497 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_497_io_l1clk),
    .io_clk(rvclkhdr_497_io_clk),
    .io_en(rvclkhdr_497_io_en),
    .io_scan_mode(rvclkhdr_497_io_scan_mode)
  );
  rvclkhdr rvclkhdr_498 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_498_io_l1clk),
    .io_clk(rvclkhdr_498_io_clk),
    .io_en(rvclkhdr_498_io_en),
    .io_scan_mode(rvclkhdr_498_io_scan_mode)
  );
  rvclkhdr rvclkhdr_499 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_499_io_l1clk),
    .io_clk(rvclkhdr_499_io_clk),
    .io_en(rvclkhdr_499_io_en),
    .io_scan_mode(rvclkhdr_499_io_scan_mode)
  );
  rvclkhdr rvclkhdr_500 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_500_io_l1clk),
    .io_clk(rvclkhdr_500_io_clk),
    .io_en(rvclkhdr_500_io_en),
    .io_scan_mode(rvclkhdr_500_io_scan_mode)
  );
  rvclkhdr rvclkhdr_501 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_501_io_l1clk),
    .io_clk(rvclkhdr_501_io_clk),
    .io_en(rvclkhdr_501_io_en),
    .io_scan_mode(rvclkhdr_501_io_scan_mode)
  );
  rvclkhdr rvclkhdr_502 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_502_io_l1clk),
    .io_clk(rvclkhdr_502_io_clk),
    .io_en(rvclkhdr_502_io_en),
    .io_scan_mode(rvclkhdr_502_io_scan_mode)
  );
  rvclkhdr rvclkhdr_503 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_503_io_l1clk),
    .io_clk(rvclkhdr_503_io_clk),
    .io_en(rvclkhdr_503_io_en),
    .io_scan_mode(rvclkhdr_503_io_scan_mode)
  );
  rvclkhdr rvclkhdr_504 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_504_io_l1clk),
    .io_clk(rvclkhdr_504_io_clk),
    .io_en(rvclkhdr_504_io_en),
    .io_scan_mode(rvclkhdr_504_io_scan_mode)
  );
  rvclkhdr rvclkhdr_505 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_505_io_l1clk),
    .io_clk(rvclkhdr_505_io_clk),
    .io_en(rvclkhdr_505_io_en),
    .io_scan_mode(rvclkhdr_505_io_scan_mode)
  );
  rvclkhdr rvclkhdr_506 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_506_io_l1clk),
    .io_clk(rvclkhdr_506_io_clk),
    .io_en(rvclkhdr_506_io_en),
    .io_scan_mode(rvclkhdr_506_io_scan_mode)
  );
  rvclkhdr rvclkhdr_507 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_507_io_l1clk),
    .io_clk(rvclkhdr_507_io_clk),
    .io_en(rvclkhdr_507_io_en),
    .io_scan_mode(rvclkhdr_507_io_scan_mode)
  );
  rvclkhdr rvclkhdr_508 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_508_io_l1clk),
    .io_clk(rvclkhdr_508_io_clk),
    .io_en(rvclkhdr_508_io_en),
    .io_scan_mode(rvclkhdr_508_io_scan_mode)
  );
  rvclkhdr rvclkhdr_509 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_509_io_l1clk),
    .io_clk(rvclkhdr_509_io_clk),
    .io_en(rvclkhdr_509_io_en),
    .io_scan_mode(rvclkhdr_509_io_scan_mode)
  );
  rvclkhdr rvclkhdr_510 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_510_io_l1clk),
    .io_clk(rvclkhdr_510_io_clk),
    .io_en(rvclkhdr_510_io_en),
    .io_scan_mode(rvclkhdr_510_io_scan_mode)
  );
  rvclkhdr rvclkhdr_511 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_511_io_l1clk),
    .io_clk(rvclkhdr_511_io_clk),
    .io_en(rvclkhdr_511_io_en),
    .io_scan_mode(rvclkhdr_511_io_scan_mode)
  );
  rvclkhdr rvclkhdr_512 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_512_io_l1clk),
    .io_clk(rvclkhdr_512_io_clk),
    .io_en(rvclkhdr_512_io_en),
    .io_scan_mode(rvclkhdr_512_io_scan_mode)
  );
  rvclkhdr rvclkhdr_513 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_513_io_l1clk),
    .io_clk(rvclkhdr_513_io_clk),
    .io_en(rvclkhdr_513_io_en),
    .io_scan_mode(rvclkhdr_513_io_scan_mode)
  );
  rvclkhdr rvclkhdr_514 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_514_io_l1clk),
    .io_clk(rvclkhdr_514_io_clk),
    .io_en(rvclkhdr_514_io_en),
    .io_scan_mode(rvclkhdr_514_io_scan_mode)
  );
  rvclkhdr rvclkhdr_515 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_515_io_l1clk),
    .io_clk(rvclkhdr_515_io_clk),
    .io_en(rvclkhdr_515_io_en),
    .io_scan_mode(rvclkhdr_515_io_scan_mode)
  );
  rvclkhdr rvclkhdr_516 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_516_io_l1clk),
    .io_clk(rvclkhdr_516_io_clk),
    .io_en(rvclkhdr_516_io_en),
    .io_scan_mode(rvclkhdr_516_io_scan_mode)
  );
  rvclkhdr rvclkhdr_517 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_517_io_l1clk),
    .io_clk(rvclkhdr_517_io_clk),
    .io_en(rvclkhdr_517_io_en),
    .io_scan_mode(rvclkhdr_517_io_scan_mode)
  );
  rvclkhdr rvclkhdr_518 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_518_io_l1clk),
    .io_clk(rvclkhdr_518_io_clk),
    .io_en(rvclkhdr_518_io_en),
    .io_scan_mode(rvclkhdr_518_io_scan_mode)
  );
  rvclkhdr rvclkhdr_519 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_519_io_l1clk),
    .io_clk(rvclkhdr_519_io_clk),
    .io_en(rvclkhdr_519_io_en),
    .io_scan_mode(rvclkhdr_519_io_scan_mode)
  );
  rvclkhdr rvclkhdr_520 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_520_io_l1clk),
    .io_clk(rvclkhdr_520_io_clk),
    .io_en(rvclkhdr_520_io_en),
    .io_scan_mode(rvclkhdr_520_io_scan_mode)
  );
  rvclkhdr rvclkhdr_521 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_521_io_l1clk),
    .io_clk(rvclkhdr_521_io_clk),
    .io_en(rvclkhdr_521_io_en),
    .io_scan_mode(rvclkhdr_521_io_scan_mode)
  );
  rvclkhdr rvclkhdr_522 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_522_io_l1clk),
    .io_clk(rvclkhdr_522_io_clk),
    .io_en(rvclkhdr_522_io_en),
    .io_scan_mode(rvclkhdr_522_io_scan_mode)
  );
  rvclkhdr rvclkhdr_523 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_523_io_l1clk),
    .io_clk(rvclkhdr_523_io_clk),
    .io_en(rvclkhdr_523_io_en),
    .io_scan_mode(rvclkhdr_523_io_scan_mode)
  );
  rvclkhdr rvclkhdr_524 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_524_io_l1clk),
    .io_clk(rvclkhdr_524_io_clk),
    .io_en(rvclkhdr_524_io_en),
    .io_scan_mode(rvclkhdr_524_io_scan_mode)
  );
  rvclkhdr rvclkhdr_525 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_525_io_l1clk),
    .io_clk(rvclkhdr_525_io_clk),
    .io_en(rvclkhdr_525_io_en),
    .io_scan_mode(rvclkhdr_525_io_scan_mode)
  );
  rvclkhdr rvclkhdr_526 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_526_io_l1clk),
    .io_clk(rvclkhdr_526_io_clk),
    .io_en(rvclkhdr_526_io_en),
    .io_scan_mode(rvclkhdr_526_io_scan_mode)
  );
  rvclkhdr rvclkhdr_527 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_527_io_l1clk),
    .io_clk(rvclkhdr_527_io_clk),
    .io_en(rvclkhdr_527_io_en),
    .io_scan_mode(rvclkhdr_527_io_scan_mode)
  );
  rvclkhdr rvclkhdr_528 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_528_io_l1clk),
    .io_clk(rvclkhdr_528_io_clk),
    .io_en(rvclkhdr_528_io_en),
    .io_scan_mode(rvclkhdr_528_io_scan_mode)
  );
  rvclkhdr rvclkhdr_529 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_529_io_l1clk),
    .io_clk(rvclkhdr_529_io_clk),
    .io_en(rvclkhdr_529_io_en),
    .io_scan_mode(rvclkhdr_529_io_scan_mode)
  );
  rvclkhdr rvclkhdr_530 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_530_io_l1clk),
    .io_clk(rvclkhdr_530_io_clk),
    .io_en(rvclkhdr_530_io_en),
    .io_scan_mode(rvclkhdr_530_io_scan_mode)
  );
  rvclkhdr rvclkhdr_531 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_531_io_l1clk),
    .io_clk(rvclkhdr_531_io_clk),
    .io_en(rvclkhdr_531_io_en),
    .io_scan_mode(rvclkhdr_531_io_scan_mode)
  );
  rvclkhdr rvclkhdr_532 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_532_io_l1clk),
    .io_clk(rvclkhdr_532_io_clk),
    .io_en(rvclkhdr_532_io_en),
    .io_scan_mode(rvclkhdr_532_io_scan_mode)
  );
  rvclkhdr rvclkhdr_533 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_533_io_l1clk),
    .io_clk(rvclkhdr_533_io_clk),
    .io_en(rvclkhdr_533_io_en),
    .io_scan_mode(rvclkhdr_533_io_scan_mode)
  );
  rvclkhdr rvclkhdr_534 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_534_io_l1clk),
    .io_clk(rvclkhdr_534_io_clk),
    .io_en(rvclkhdr_534_io_en),
    .io_scan_mode(rvclkhdr_534_io_scan_mode)
  );
  rvclkhdr rvclkhdr_535 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_535_io_l1clk),
    .io_clk(rvclkhdr_535_io_clk),
    .io_en(rvclkhdr_535_io_en),
    .io_scan_mode(rvclkhdr_535_io_scan_mode)
  );
  rvclkhdr rvclkhdr_536 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_536_io_l1clk),
    .io_clk(rvclkhdr_536_io_clk),
    .io_en(rvclkhdr_536_io_en),
    .io_scan_mode(rvclkhdr_536_io_scan_mode)
  );
  rvclkhdr rvclkhdr_537 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_537_io_l1clk),
    .io_clk(rvclkhdr_537_io_clk),
    .io_en(rvclkhdr_537_io_en),
    .io_scan_mode(rvclkhdr_537_io_scan_mode)
  );
  rvclkhdr rvclkhdr_538 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_538_io_l1clk),
    .io_clk(rvclkhdr_538_io_clk),
    .io_en(rvclkhdr_538_io_en),
    .io_scan_mode(rvclkhdr_538_io_scan_mode)
  );
  rvclkhdr rvclkhdr_539 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_539_io_l1clk),
    .io_clk(rvclkhdr_539_io_clk),
    .io_en(rvclkhdr_539_io_en),
    .io_scan_mode(rvclkhdr_539_io_scan_mode)
  );
  rvclkhdr rvclkhdr_540 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_540_io_l1clk),
    .io_clk(rvclkhdr_540_io_clk),
    .io_en(rvclkhdr_540_io_en),
    .io_scan_mode(rvclkhdr_540_io_scan_mode)
  );
  rvclkhdr rvclkhdr_541 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_541_io_l1clk),
    .io_clk(rvclkhdr_541_io_clk),
    .io_en(rvclkhdr_541_io_en),
    .io_scan_mode(rvclkhdr_541_io_scan_mode)
  );
  rvclkhdr rvclkhdr_542 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_542_io_l1clk),
    .io_clk(rvclkhdr_542_io_clk),
    .io_en(rvclkhdr_542_io_en),
    .io_scan_mode(rvclkhdr_542_io_scan_mode)
  );
  rvclkhdr rvclkhdr_543 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_543_io_l1clk),
    .io_clk(rvclkhdr_543_io_clk),
    .io_en(rvclkhdr_543_io_en),
    .io_scan_mode(rvclkhdr_543_io_scan_mode)
  );
  rvclkhdr rvclkhdr_544 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_544_io_l1clk),
    .io_clk(rvclkhdr_544_io_clk),
    .io_en(rvclkhdr_544_io_en),
    .io_scan_mode(rvclkhdr_544_io_scan_mode)
  );
  rvclkhdr rvclkhdr_545 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_545_io_l1clk),
    .io_clk(rvclkhdr_545_io_clk),
    .io_en(rvclkhdr_545_io_en),
    .io_scan_mode(rvclkhdr_545_io_scan_mode)
  );
  rvclkhdr rvclkhdr_546 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_546_io_l1clk),
    .io_clk(rvclkhdr_546_io_clk),
    .io_en(rvclkhdr_546_io_en),
    .io_scan_mode(rvclkhdr_546_io_scan_mode)
  );
  rvclkhdr rvclkhdr_547 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_547_io_l1clk),
    .io_clk(rvclkhdr_547_io_clk),
    .io_en(rvclkhdr_547_io_en),
    .io_scan_mode(rvclkhdr_547_io_scan_mode)
  );
  rvclkhdr rvclkhdr_548 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_548_io_l1clk),
    .io_clk(rvclkhdr_548_io_clk),
    .io_en(rvclkhdr_548_io_en),
    .io_scan_mode(rvclkhdr_548_io_scan_mode)
  );
  rvclkhdr rvclkhdr_549 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_549_io_l1clk),
    .io_clk(rvclkhdr_549_io_clk),
    .io_en(rvclkhdr_549_io_en),
    .io_scan_mode(rvclkhdr_549_io_scan_mode)
  );
  rvclkhdr rvclkhdr_550 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_550_io_l1clk),
    .io_clk(rvclkhdr_550_io_clk),
    .io_en(rvclkhdr_550_io_en),
    .io_scan_mode(rvclkhdr_550_io_scan_mode)
  );
  rvclkhdr rvclkhdr_551 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_551_io_l1clk),
    .io_clk(rvclkhdr_551_io_clk),
    .io_en(rvclkhdr_551_io_en),
    .io_scan_mode(rvclkhdr_551_io_scan_mode)
  );
  rvclkhdr rvclkhdr_552 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_552_io_l1clk),
    .io_clk(rvclkhdr_552_io_clk),
    .io_en(rvclkhdr_552_io_en),
    .io_scan_mode(rvclkhdr_552_io_scan_mode)
  );
  rvclkhdr rvclkhdr_553 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_553_io_l1clk),
    .io_clk(rvclkhdr_553_io_clk),
    .io_en(rvclkhdr_553_io_en),
    .io_scan_mode(rvclkhdr_553_io_scan_mode)
  );
  assign io_ifu_bp_hit_taken_f = _T_238 & _T_239; // @[ifu_bp_ctl.scala 261:25]
  assign io_ifu_bp_btb_target_f = _T_429 ? rets_out_0[31:1] : bp_btb_target_adder_f[31:1]; // @[ifu_bp_ctl.scala 357:26]
  assign io_ifu_bp_inst_mask_f = _T_275 | _T_276; // @[ifu_bp_ctl.scala 285:25]
  assign io_ifu_bp_fghr_f = fghr; // @[ifu_bp_ctl.scala 325:20]
  assign io_ifu_bp_way_f = tag_match_vway1_expanded_f | _T_213; // @[ifu_bp_ctl.scala 235:19]
  assign io_ifu_bp_ret_f = {_T_295,_T_301}; // @[ifu_bp_ctl.scala 331:19]
  assign io_ifu_bp_hist1_f = bht_force_taken_f | _T_280; // @[ifu_bp_ctl.scala 326:21]
  assign io_ifu_bp_hist0_f = {bht_vbank1_rd_data_f[0],bht_vbank0_rd_data_f[0]}; // @[ifu_bp_ctl.scala 327:21]
  assign io_ifu_bp_pc4_f = {_T_286,_T_289}; // @[ifu_bp_ctl.scala 328:19]
  assign io_ifu_bp_valid_f = bht_valid_f & _T_345; // @[ifu_bp_ctl.scala 330:21]
  assign io_ifu_bp_poffset_f = btb_sel_data_f[15:4]; // @[ifu_bp_ctl.scala 344:23]
  assign rvclkhdr_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_io_en = io_ifc_fetch_req_f | exu_mp_valid; // @[lib.scala 371:17]
  assign rvclkhdr_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_1_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_1_io_en = _T_376 & io_ic_hit_f; // @[lib.scala 371:17]
  assign rvclkhdr_1_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_2_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_2_io_en = ~rs_hold; // @[lib.scala 371:17]
  assign rvclkhdr_2_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_3_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_3_io_en = rs_push | rs_pop; // @[lib.scala 371:17]
  assign rvclkhdr_3_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_4_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_4_io_en = rs_push | rs_pop; // @[lib.scala 371:17]
  assign rvclkhdr_4_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_5_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_5_io_en = rs_push | rs_pop; // @[lib.scala 371:17]
  assign rvclkhdr_5_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_6_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_6_io_en = rs_push | rs_pop; // @[lib.scala 371:17]
  assign rvclkhdr_6_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_7_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_7_io_en = rs_push | rs_pop; // @[lib.scala 371:17]
  assign rvclkhdr_7_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_8_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_8_io_en = rs_push | rs_pop; // @[lib.scala 371:17]
  assign rvclkhdr_8_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_9_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_9_io_en = _T_473 & io_ifu_bp_hit_taken_f; // @[lib.scala 371:17]
  assign rvclkhdr_9_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_10_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_10_io_en = _T_576 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_10_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_11_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_11_io_en = _T_579 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_11_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_12_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_12_io_en = _T_582 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_12_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_13_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_13_io_en = _T_585 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_13_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_14_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_14_io_en = _T_588 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_14_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_15_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_15_io_en = _T_591 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_15_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_16_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_16_io_en = _T_594 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_16_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_17_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_17_io_en = _T_597 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_17_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_18_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_18_io_en = _T_600 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_18_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_19_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_19_io_en = _T_603 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_19_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_20_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_20_io_en = _T_606 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_20_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_21_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_21_io_en = _T_609 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_21_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_22_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_22_io_en = _T_612 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_22_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_23_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_23_io_en = _T_615 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_23_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_24_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_24_io_en = _T_618 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_24_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_25_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_25_io_en = _T_621 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_25_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_26_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_26_io_en = _T_624 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_26_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_27_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_27_io_en = _T_627 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_27_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_28_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_28_io_en = _T_630 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_28_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_29_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_29_io_en = _T_633 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_29_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_30_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_30_io_en = _T_636 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_30_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_31_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_31_io_en = _T_639 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_31_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_32_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_32_io_en = _T_642 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_32_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_33_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_33_io_en = _T_645 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_33_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_34_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_34_io_en = _T_648 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_34_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_35_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_35_io_en = _T_651 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_35_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_36_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_36_io_en = _T_654 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_36_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_37_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_37_io_en = _T_657 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_37_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_38_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_38_io_en = _T_660 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_38_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_39_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_39_io_en = _T_663 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_39_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_40_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_40_io_en = _T_666 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_40_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_41_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_41_io_en = _T_669 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_41_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_42_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_42_io_en = _T_672 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_42_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_43_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_43_io_en = _T_675 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_43_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_44_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_44_io_en = _T_678 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_44_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_45_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_45_io_en = _T_681 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_45_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_46_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_46_io_en = _T_684 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_46_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_47_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_47_io_en = _T_687 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_47_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_48_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_48_io_en = _T_690 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_48_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_49_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_49_io_en = _T_693 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_49_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_50_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_50_io_en = _T_696 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_50_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_51_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_51_io_en = _T_699 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_51_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_52_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_52_io_en = _T_702 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_52_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_53_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_53_io_en = _T_705 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_53_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_54_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_54_io_en = _T_708 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_54_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_55_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_55_io_en = _T_711 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_55_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_56_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_56_io_en = _T_714 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_56_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_57_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_57_io_en = _T_717 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_57_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_58_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_58_io_en = _T_720 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_58_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_59_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_59_io_en = _T_723 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_59_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_60_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_60_io_en = _T_726 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_60_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_61_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_61_io_en = _T_729 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_61_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_62_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_62_io_en = _T_732 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_62_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_63_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_63_io_en = _T_735 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_63_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_64_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_64_io_en = _T_738 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_64_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_65_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_65_io_en = _T_741 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_65_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_66_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_66_io_en = _T_744 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_66_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_67_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_67_io_en = _T_747 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_67_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_68_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_68_io_en = _T_750 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_68_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_69_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_69_io_en = _T_753 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_69_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_70_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_70_io_en = _T_756 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_70_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_71_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_71_io_en = _T_759 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_71_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_72_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_72_io_en = _T_762 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_72_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_73_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_73_io_en = _T_765 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_73_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_74_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_74_io_en = _T_768 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_74_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_75_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_75_io_en = _T_771 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_75_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_76_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_76_io_en = _T_774 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_76_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_77_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_77_io_en = _T_777 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_77_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_78_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_78_io_en = _T_780 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_78_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_79_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_79_io_en = _T_783 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_79_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_80_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_80_io_en = _T_786 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_80_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_81_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_81_io_en = _T_789 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_81_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_82_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_82_io_en = _T_792 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_82_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_83_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_83_io_en = _T_795 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_83_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_84_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_84_io_en = _T_798 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_84_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_85_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_85_io_en = _T_801 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_85_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_86_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_86_io_en = _T_804 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_86_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_87_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_87_io_en = _T_807 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_87_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_88_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_88_io_en = _T_810 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_88_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_89_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_89_io_en = _T_813 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_89_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_90_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_90_io_en = _T_816 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_90_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_91_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_91_io_en = _T_819 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_91_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_92_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_92_io_en = _T_822 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_92_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_93_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_93_io_en = _T_825 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_93_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_94_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_94_io_en = _T_828 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_94_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_95_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_95_io_en = _T_831 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_95_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_96_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_96_io_en = _T_834 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_96_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_97_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_97_io_en = _T_837 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_97_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_98_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_98_io_en = _T_840 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_98_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_99_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_99_io_en = _T_843 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_99_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_100_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_100_io_en = _T_846 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_100_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_101_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_101_io_en = _T_849 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_101_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_102_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_102_io_en = _T_852 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_102_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_103_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_103_io_en = _T_855 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_103_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_104_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_104_io_en = _T_858 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_104_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_105_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_105_io_en = _T_861 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_105_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_106_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_106_io_en = _T_864 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_106_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_107_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_107_io_en = _T_867 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_107_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_108_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_108_io_en = _T_870 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_108_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_109_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_109_io_en = _T_873 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_109_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_110_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_110_io_en = _T_876 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_110_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_111_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_111_io_en = _T_879 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_111_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_112_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_112_io_en = _T_882 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_112_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_113_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_113_io_en = _T_885 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_113_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_114_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_114_io_en = _T_888 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_114_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_115_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_115_io_en = _T_891 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_115_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_116_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_116_io_en = _T_894 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_116_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_117_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_117_io_en = _T_897 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_117_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_118_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_118_io_en = _T_900 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_118_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_119_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_119_io_en = _T_903 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_119_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_120_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_120_io_en = _T_906 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_120_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_121_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_121_io_en = _T_909 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_121_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_122_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_122_io_en = _T_912 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_122_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_123_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_123_io_en = _T_915 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_123_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_124_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_124_io_en = _T_918 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_124_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_125_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_125_io_en = _T_921 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_125_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_126_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_126_io_en = _T_924 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_126_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_127_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_127_io_en = _T_927 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_127_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_128_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_128_io_en = _T_930 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_128_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_129_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_129_io_en = _T_933 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_129_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_130_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_130_io_en = _T_936 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_130_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_131_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_131_io_en = _T_939 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_131_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_132_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_132_io_en = _T_942 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_132_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_133_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_133_io_en = _T_945 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_133_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_134_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_134_io_en = _T_948 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_134_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_135_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_135_io_en = _T_951 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_135_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_136_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_136_io_en = _T_954 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_136_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_137_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_137_io_en = _T_957 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_137_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_138_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_138_io_en = _T_960 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_138_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_139_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_139_io_en = _T_963 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_139_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_140_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_140_io_en = _T_966 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_140_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_141_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_141_io_en = _T_969 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_141_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_142_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_142_io_en = _T_972 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_142_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_143_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_143_io_en = _T_975 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_143_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_144_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_144_io_en = _T_978 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_144_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_145_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_145_io_en = _T_981 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_145_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_146_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_146_io_en = _T_984 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_146_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_147_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_147_io_en = _T_987 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_147_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_148_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_148_io_en = _T_990 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_148_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_149_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_149_io_en = _T_993 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_149_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_150_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_150_io_en = _T_996 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_150_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_151_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_151_io_en = _T_999 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_151_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_152_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_152_io_en = _T_1002 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_152_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_153_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_153_io_en = _T_1005 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_153_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_154_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_154_io_en = _T_1008 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_154_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_155_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_155_io_en = _T_1011 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_155_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_156_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_156_io_en = _T_1014 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_156_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_157_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_157_io_en = _T_1017 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_157_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_158_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_158_io_en = _T_1020 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_158_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_159_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_159_io_en = _T_1023 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_159_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_160_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_160_io_en = _T_1026 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_160_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_161_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_161_io_en = _T_1029 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_161_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_162_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_162_io_en = _T_1032 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_162_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_163_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_163_io_en = _T_1035 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_163_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_164_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_164_io_en = _T_1038 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_164_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_165_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_165_io_en = _T_1041 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_165_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_166_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_166_io_en = _T_1044 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_166_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_167_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_167_io_en = _T_1047 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_167_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_168_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_168_io_en = _T_1050 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_168_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_169_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_169_io_en = _T_1053 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_169_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_170_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_170_io_en = _T_1056 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_170_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_171_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_171_io_en = _T_1059 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_171_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_172_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_172_io_en = _T_1062 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_172_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_173_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_173_io_en = _T_1065 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_173_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_174_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_174_io_en = _T_1068 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_174_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_175_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_175_io_en = _T_1071 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_175_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_176_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_176_io_en = _T_1074 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_176_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_177_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_177_io_en = _T_1077 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_177_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_178_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_178_io_en = _T_1080 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_178_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_179_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_179_io_en = _T_1083 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_179_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_180_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_180_io_en = _T_1086 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_180_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_181_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_181_io_en = _T_1089 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_181_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_182_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_182_io_en = _T_1092 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_182_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_183_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_183_io_en = _T_1095 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_183_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_184_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_184_io_en = _T_1098 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_184_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_185_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_185_io_en = _T_1101 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_185_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_186_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_186_io_en = _T_1104 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_186_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_187_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_187_io_en = _T_1107 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_187_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_188_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_188_io_en = _T_1110 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_188_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_189_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_189_io_en = _T_1113 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_189_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_190_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_190_io_en = _T_1116 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_190_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_191_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_191_io_en = _T_1119 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_191_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_192_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_192_io_en = _T_1122 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_192_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_193_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_193_io_en = _T_1125 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_193_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_194_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_194_io_en = _T_1128 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_194_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_195_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_195_io_en = _T_1131 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_195_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_196_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_196_io_en = _T_1134 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_196_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_197_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_197_io_en = _T_1137 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_197_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_198_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_198_io_en = _T_1140 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_198_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_199_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_199_io_en = _T_1143 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_199_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_200_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_200_io_en = _T_1146 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_200_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_201_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_201_io_en = _T_1149 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_201_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_202_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_202_io_en = _T_1152 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_202_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_203_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_203_io_en = _T_1155 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_203_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_204_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_204_io_en = _T_1158 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_204_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_205_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_205_io_en = _T_1161 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_205_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_206_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_206_io_en = _T_1164 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_206_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_207_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_207_io_en = _T_1167 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_207_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_208_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_208_io_en = _T_1170 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_208_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_209_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_209_io_en = _T_1173 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_209_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_210_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_210_io_en = _T_1176 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_210_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_211_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_211_io_en = _T_1179 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_211_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_212_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_212_io_en = _T_1182 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_212_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_213_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_213_io_en = _T_1185 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_213_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_214_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_214_io_en = _T_1188 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_214_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_215_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_215_io_en = _T_1191 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_215_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_216_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_216_io_en = _T_1194 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_216_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_217_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_217_io_en = _T_1197 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_217_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_218_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_218_io_en = _T_1200 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_218_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_219_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_219_io_en = _T_1203 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_219_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_220_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_220_io_en = _T_1206 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_220_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_221_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_221_io_en = _T_1209 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_221_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_222_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_222_io_en = _T_1212 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_222_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_223_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_223_io_en = _T_1215 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_223_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_224_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_224_io_en = _T_1218 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_224_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_225_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_225_io_en = _T_1221 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_225_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_226_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_226_io_en = _T_1224 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_226_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_227_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_227_io_en = _T_1227 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_227_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_228_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_228_io_en = _T_1230 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_228_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_229_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_229_io_en = _T_1233 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_229_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_230_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_230_io_en = _T_1236 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_230_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_231_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_231_io_en = _T_1239 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_231_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_232_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_232_io_en = _T_1242 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_232_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_233_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_233_io_en = _T_1245 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_233_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_234_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_234_io_en = _T_1248 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_234_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_235_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_235_io_en = _T_1251 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_235_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_236_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_236_io_en = _T_1254 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_236_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_237_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_237_io_en = _T_1257 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_237_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_238_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_238_io_en = _T_1260 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_238_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_239_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_239_io_en = _T_1263 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_239_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_240_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_240_io_en = _T_1266 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_240_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_241_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_241_io_en = _T_1269 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_241_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_242_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_242_io_en = _T_1272 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_242_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_243_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_243_io_en = _T_1275 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_243_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_244_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_244_io_en = _T_1278 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_244_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_245_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_245_io_en = _T_1281 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_245_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_246_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_246_io_en = _T_1284 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_246_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_247_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_247_io_en = _T_1287 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_247_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_248_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_248_io_en = _T_1290 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_248_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_249_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_249_io_en = _T_1293 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_249_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_250_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_250_io_en = _T_1296 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_250_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_251_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_251_io_en = _T_1299 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_251_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_252_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_252_io_en = _T_1302 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_252_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_253_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_253_io_en = _T_1305 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_253_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_254_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_254_io_en = _T_1308 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_254_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_255_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_255_io_en = _T_1311 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_255_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_256_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_256_io_en = _T_1314 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_256_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_257_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_257_io_en = _T_1317 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_257_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_258_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_258_io_en = _T_1320 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_258_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_259_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_259_io_en = _T_1323 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_259_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_260_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_260_io_en = _T_1326 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_260_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_261_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_261_io_en = _T_1329 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_261_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_262_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_262_io_en = _T_1332 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_262_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_263_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_263_io_en = _T_1335 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_263_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_264_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_264_io_en = _T_1338 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_264_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_265_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_265_io_en = _T_1341 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_265_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_266_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_266_io_en = _T_576 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_266_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_267_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_267_io_en = _T_579 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_267_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_268_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_268_io_en = _T_582 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_268_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_269_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_269_io_en = _T_585 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_269_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_270_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_270_io_en = _T_588 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_270_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_271_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_271_io_en = _T_591 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_271_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_272_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_272_io_en = _T_594 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_272_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_273_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_273_io_en = _T_597 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_273_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_274_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_274_io_en = _T_600 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_274_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_275_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_275_io_en = _T_603 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_275_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_276_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_276_io_en = _T_606 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_276_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_277_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_277_io_en = _T_609 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_277_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_278_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_278_io_en = _T_612 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_278_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_279_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_279_io_en = _T_615 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_279_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_280_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_280_io_en = _T_618 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_280_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_281_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_281_io_en = _T_621 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_281_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_282_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_282_io_en = _T_624 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_282_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_283_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_283_io_en = _T_627 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_283_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_284_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_284_io_en = _T_630 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_284_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_285_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_285_io_en = _T_633 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_285_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_286_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_286_io_en = _T_636 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_286_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_287_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_287_io_en = _T_639 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_287_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_288_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_288_io_en = _T_642 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_288_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_289_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_289_io_en = _T_645 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_289_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_290_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_290_io_en = _T_648 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_290_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_291_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_291_io_en = _T_651 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_291_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_292_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_292_io_en = _T_654 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_292_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_293_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_293_io_en = _T_657 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_293_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_294_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_294_io_en = _T_660 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_294_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_295_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_295_io_en = _T_663 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_295_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_296_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_296_io_en = _T_666 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_296_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_297_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_297_io_en = _T_669 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_297_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_298_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_298_io_en = _T_672 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_298_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_299_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_299_io_en = _T_675 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_299_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_300_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_300_io_en = _T_678 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_300_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_301_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_301_io_en = _T_681 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_301_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_302_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_302_io_en = _T_684 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_302_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_303_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_303_io_en = _T_687 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_303_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_304_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_304_io_en = _T_690 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_304_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_305_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_305_io_en = _T_693 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_305_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_306_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_306_io_en = _T_696 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_306_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_307_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_307_io_en = _T_699 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_307_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_308_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_308_io_en = _T_702 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_308_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_309_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_309_io_en = _T_705 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_309_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_310_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_310_io_en = _T_708 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_310_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_311_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_311_io_en = _T_711 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_311_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_312_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_312_io_en = _T_714 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_312_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_313_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_313_io_en = _T_717 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_313_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_314_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_314_io_en = _T_720 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_314_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_315_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_315_io_en = _T_723 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_315_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_316_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_316_io_en = _T_726 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_316_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_317_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_317_io_en = _T_729 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_317_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_318_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_318_io_en = _T_732 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_318_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_319_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_319_io_en = _T_735 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_319_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_320_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_320_io_en = _T_738 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_320_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_321_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_321_io_en = _T_741 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_321_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_322_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_322_io_en = _T_744 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_322_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_323_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_323_io_en = _T_747 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_323_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_324_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_324_io_en = _T_750 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_324_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_325_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_325_io_en = _T_753 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_325_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_326_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_326_io_en = _T_756 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_326_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_327_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_327_io_en = _T_759 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_327_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_328_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_328_io_en = _T_762 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_328_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_329_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_329_io_en = _T_765 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_329_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_330_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_330_io_en = _T_768 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_330_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_331_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_331_io_en = _T_771 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_331_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_332_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_332_io_en = _T_774 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_332_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_333_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_333_io_en = _T_777 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_333_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_334_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_334_io_en = _T_780 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_334_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_335_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_335_io_en = _T_783 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_335_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_336_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_336_io_en = _T_786 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_336_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_337_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_337_io_en = _T_789 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_337_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_338_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_338_io_en = _T_792 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_338_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_339_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_339_io_en = _T_795 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_339_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_340_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_340_io_en = _T_798 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_340_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_341_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_341_io_en = _T_801 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_341_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_342_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_342_io_en = _T_804 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_342_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_343_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_343_io_en = _T_807 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_343_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_344_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_344_io_en = _T_810 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_344_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_345_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_345_io_en = _T_813 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_345_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_346_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_346_io_en = _T_816 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_346_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_347_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_347_io_en = _T_819 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_347_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_348_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_348_io_en = _T_822 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_348_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_349_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_349_io_en = _T_825 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_349_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_350_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_350_io_en = _T_828 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_350_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_351_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_351_io_en = _T_831 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_351_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_352_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_352_io_en = _T_834 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_352_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_353_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_353_io_en = _T_837 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_353_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_354_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_354_io_en = _T_840 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_354_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_355_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_355_io_en = _T_843 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_355_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_356_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_356_io_en = _T_846 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_356_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_357_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_357_io_en = _T_849 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_357_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_358_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_358_io_en = _T_852 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_358_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_359_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_359_io_en = _T_855 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_359_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_360_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_360_io_en = _T_858 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_360_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_361_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_361_io_en = _T_861 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_361_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_362_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_362_io_en = _T_864 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_362_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_363_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_363_io_en = _T_867 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_363_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_364_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_364_io_en = _T_870 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_364_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_365_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_365_io_en = _T_873 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_365_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_366_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_366_io_en = _T_876 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_366_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_367_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_367_io_en = _T_879 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_367_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_368_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_368_io_en = _T_882 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_368_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_369_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_369_io_en = _T_885 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_369_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_370_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_370_io_en = _T_888 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_370_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_371_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_371_io_en = _T_891 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_371_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_372_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_372_io_en = _T_894 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_372_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_373_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_373_io_en = _T_897 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_373_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_374_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_374_io_en = _T_900 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_374_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_375_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_375_io_en = _T_903 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_375_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_376_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_376_io_en = _T_906 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_376_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_377_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_377_io_en = _T_909 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_377_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_378_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_378_io_en = _T_912 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_378_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_379_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_379_io_en = _T_915 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_379_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_380_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_380_io_en = _T_918 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_380_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_381_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_381_io_en = _T_921 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_381_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_382_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_382_io_en = _T_924 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_382_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_383_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_383_io_en = _T_927 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_383_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_384_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_384_io_en = _T_930 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_384_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_385_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_385_io_en = _T_933 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_385_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_386_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_386_io_en = _T_936 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_386_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_387_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_387_io_en = _T_939 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_387_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_388_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_388_io_en = _T_942 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_388_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_389_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_389_io_en = _T_945 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_389_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_390_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_390_io_en = _T_948 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_390_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_391_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_391_io_en = _T_951 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_391_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_392_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_392_io_en = _T_954 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_392_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_393_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_393_io_en = _T_957 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_393_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_394_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_394_io_en = _T_960 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_394_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_395_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_395_io_en = _T_963 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_395_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_396_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_396_io_en = _T_966 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_396_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_397_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_397_io_en = _T_969 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_397_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_398_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_398_io_en = _T_972 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_398_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_399_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_399_io_en = _T_975 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_399_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_400_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_400_io_en = _T_978 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_400_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_401_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_401_io_en = _T_981 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_401_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_402_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_402_io_en = _T_984 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_402_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_403_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_403_io_en = _T_987 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_403_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_404_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_404_io_en = _T_990 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_404_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_405_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_405_io_en = _T_993 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_405_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_406_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_406_io_en = _T_996 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_406_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_407_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_407_io_en = _T_999 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_407_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_408_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_408_io_en = _T_1002 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_408_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_409_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_409_io_en = _T_1005 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_409_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_410_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_410_io_en = _T_1008 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_410_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_411_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_411_io_en = _T_1011 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_411_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_412_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_412_io_en = _T_1014 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_412_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_413_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_413_io_en = _T_1017 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_413_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_414_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_414_io_en = _T_1020 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_414_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_415_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_415_io_en = _T_1023 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_415_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_416_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_416_io_en = _T_1026 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_416_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_417_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_417_io_en = _T_1029 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_417_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_418_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_418_io_en = _T_1032 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_418_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_419_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_419_io_en = _T_1035 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_419_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_420_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_420_io_en = _T_1038 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_420_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_421_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_421_io_en = _T_1041 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_421_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_422_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_422_io_en = _T_1044 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_422_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_423_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_423_io_en = _T_1047 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_423_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_424_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_424_io_en = _T_1050 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_424_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_425_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_425_io_en = _T_1053 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_425_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_426_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_426_io_en = _T_1056 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_426_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_427_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_427_io_en = _T_1059 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_427_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_428_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_428_io_en = _T_1062 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_428_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_429_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_429_io_en = _T_1065 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_429_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_430_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_430_io_en = _T_1068 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_430_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_431_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_431_io_en = _T_1071 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_431_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_432_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_432_io_en = _T_1074 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_432_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_433_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_433_io_en = _T_1077 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_433_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_434_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_434_io_en = _T_1080 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_434_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_435_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_435_io_en = _T_1083 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_435_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_436_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_436_io_en = _T_1086 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_436_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_437_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_437_io_en = _T_1089 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_437_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_438_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_438_io_en = _T_1092 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_438_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_439_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_439_io_en = _T_1095 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_439_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_440_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_440_io_en = _T_1098 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_440_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_441_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_441_io_en = _T_1101 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_441_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_442_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_442_io_en = _T_1104 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_442_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_443_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_443_io_en = _T_1107 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_443_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_444_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_444_io_en = _T_1110 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_444_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_445_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_445_io_en = _T_1113 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_445_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_446_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_446_io_en = _T_1116 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_446_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_447_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_447_io_en = _T_1119 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_447_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_448_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_448_io_en = _T_1122 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_448_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_449_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_449_io_en = _T_1125 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_449_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_450_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_450_io_en = _T_1128 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_450_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_451_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_451_io_en = _T_1131 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_451_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_452_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_452_io_en = _T_1134 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_452_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_453_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_453_io_en = _T_1137 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_453_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_454_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_454_io_en = _T_1140 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_454_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_455_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_455_io_en = _T_1143 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_455_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_456_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_456_io_en = _T_1146 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_456_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_457_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_457_io_en = _T_1149 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_457_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_458_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_458_io_en = _T_1152 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_458_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_459_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_459_io_en = _T_1155 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_459_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_460_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_460_io_en = _T_1158 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_460_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_461_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_461_io_en = _T_1161 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_461_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_462_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_462_io_en = _T_1164 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_462_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_463_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_463_io_en = _T_1167 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_463_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_464_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_464_io_en = _T_1170 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_464_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_465_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_465_io_en = _T_1173 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_465_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_466_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_466_io_en = _T_1176 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_466_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_467_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_467_io_en = _T_1179 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_467_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_468_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_468_io_en = _T_1182 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_468_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_469_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_469_io_en = _T_1185 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_469_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_470_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_470_io_en = _T_1188 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_470_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_471_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_471_io_en = _T_1191 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_471_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_472_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_472_io_en = _T_1194 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_472_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_473_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_473_io_en = _T_1197 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_473_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_474_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_474_io_en = _T_1200 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_474_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_475_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_475_io_en = _T_1203 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_475_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_476_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_476_io_en = _T_1206 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_476_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_477_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_477_io_en = _T_1209 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_477_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_478_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_478_io_en = _T_1212 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_478_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_479_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_479_io_en = _T_1215 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_479_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_480_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_480_io_en = _T_1218 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_480_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_481_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_481_io_en = _T_1221 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_481_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_482_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_482_io_en = _T_1224 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_482_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_483_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_483_io_en = _T_1227 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_483_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_484_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_484_io_en = _T_1230 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_484_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_485_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_485_io_en = _T_1233 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_485_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_486_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_486_io_en = _T_1236 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_486_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_487_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_487_io_en = _T_1239 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_487_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_488_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_488_io_en = _T_1242 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_488_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_489_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_489_io_en = _T_1245 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_489_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_490_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_490_io_en = _T_1248 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_490_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_491_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_491_io_en = _T_1251 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_491_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_492_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_492_io_en = _T_1254 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_492_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_493_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_493_io_en = _T_1257 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_493_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_494_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_494_io_en = _T_1260 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_494_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_495_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_495_io_en = _T_1263 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_495_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_496_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_496_io_en = _T_1266 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_496_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_497_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_497_io_en = _T_1269 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_497_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_498_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_498_io_en = _T_1272 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_498_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_499_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_499_io_en = _T_1275 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_499_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_500_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_500_io_en = _T_1278 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_500_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_501_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_501_io_en = _T_1281 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_501_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_502_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_502_io_en = _T_1284 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_502_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_503_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_503_io_en = _T_1287 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_503_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_504_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_504_io_en = _T_1290 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_504_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_505_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_505_io_en = _T_1293 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_505_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_506_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_506_io_en = _T_1296 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_506_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_507_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_507_io_en = _T_1299 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_507_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_508_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_508_io_en = _T_1302 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_508_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_509_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_509_io_en = _T_1305 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_509_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_510_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_510_io_en = _T_1308 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_510_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_511_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_511_io_en = _T_1311 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_511_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_512_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_512_io_en = _T_1314 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_512_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_513_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_513_io_en = _T_1317 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_513_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_514_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_514_io_en = _T_1320 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_514_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_515_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_515_io_en = _T_1323 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_515_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_516_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_516_io_en = _T_1326 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_516_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_517_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_517_io_en = _T_1329 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_517_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_518_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_518_io_en = _T_1332 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_518_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_519_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_519_io_en = _T_1335 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_519_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_520_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_520_io_en = _T_1338 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_520_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_521_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_521_io_en = _T_1341 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_521_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_522_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_522_io_en = _T_6212 | _T_6217; // @[lib.scala 345:16]
  assign rvclkhdr_522_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_523_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_523_io_en = _T_6223 | _T_6228; // @[lib.scala 345:16]
  assign rvclkhdr_523_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_524_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_524_io_en = _T_6234 | _T_6239; // @[lib.scala 345:16]
  assign rvclkhdr_524_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_525_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_525_io_en = _T_6245 | _T_6250; // @[lib.scala 345:16]
  assign rvclkhdr_525_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_526_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_526_io_en = _T_6256 | _T_6261; // @[lib.scala 345:16]
  assign rvclkhdr_526_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_527_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_527_io_en = _T_6267 | _T_6272; // @[lib.scala 345:16]
  assign rvclkhdr_527_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_528_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_528_io_en = _T_6278 | _T_6283; // @[lib.scala 345:16]
  assign rvclkhdr_528_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_529_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_529_io_en = _T_6289 | _T_6294; // @[lib.scala 345:16]
  assign rvclkhdr_529_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_530_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_530_io_en = _T_6300 | _T_6305; // @[lib.scala 345:16]
  assign rvclkhdr_530_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_531_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_531_io_en = _T_6311 | _T_6316; // @[lib.scala 345:16]
  assign rvclkhdr_531_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_532_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_532_io_en = _T_6322 | _T_6327; // @[lib.scala 345:16]
  assign rvclkhdr_532_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_533_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_533_io_en = _T_6333 | _T_6338; // @[lib.scala 345:16]
  assign rvclkhdr_533_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_534_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_534_io_en = _T_6344 | _T_6349; // @[lib.scala 345:16]
  assign rvclkhdr_534_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_535_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_535_io_en = _T_6355 | _T_6360; // @[lib.scala 345:16]
  assign rvclkhdr_535_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_536_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_536_io_en = _T_6366 | _T_6371; // @[lib.scala 345:16]
  assign rvclkhdr_536_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_537_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_537_io_en = _T_6377 | _T_6382; // @[lib.scala 345:16]
  assign rvclkhdr_537_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_538_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_538_io_en = _T_6388 | _T_6393; // @[lib.scala 345:16]
  assign rvclkhdr_538_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_539_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_539_io_en = _T_6399 | _T_6404; // @[lib.scala 345:16]
  assign rvclkhdr_539_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_540_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_540_io_en = _T_6410 | _T_6415; // @[lib.scala 345:16]
  assign rvclkhdr_540_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_541_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_541_io_en = _T_6421 | _T_6426; // @[lib.scala 345:16]
  assign rvclkhdr_541_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_542_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_542_io_en = _T_6432 | _T_6437; // @[lib.scala 345:16]
  assign rvclkhdr_542_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_543_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_543_io_en = _T_6443 | _T_6448; // @[lib.scala 345:16]
  assign rvclkhdr_543_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_544_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_544_io_en = _T_6454 | _T_6459; // @[lib.scala 345:16]
  assign rvclkhdr_544_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_545_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_545_io_en = _T_6465 | _T_6470; // @[lib.scala 345:16]
  assign rvclkhdr_545_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_546_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_546_io_en = _T_6476 | _T_6481; // @[lib.scala 345:16]
  assign rvclkhdr_546_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_547_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_547_io_en = _T_6487 | _T_6492; // @[lib.scala 345:16]
  assign rvclkhdr_547_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_548_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_548_io_en = _T_6498 | _T_6503; // @[lib.scala 345:16]
  assign rvclkhdr_548_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_549_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_549_io_en = _T_6509 | _T_6514; // @[lib.scala 345:16]
  assign rvclkhdr_549_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_550_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_550_io_en = _T_6520 | _T_6525; // @[lib.scala 345:16]
  assign rvclkhdr_550_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_551_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_551_io_en = _T_6531 | _T_6536; // @[lib.scala 345:16]
  assign rvclkhdr_551_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_552_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_552_io_en = _T_6542 | _T_6547; // @[lib.scala 345:16]
  assign rvclkhdr_552_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_553_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_553_io_en = _T_6553 | _T_6558; // @[lib.scala 345:16]
  assign rvclkhdr_553_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  leak_one_f_d1 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_0 = _RAND_1[21:0];
  _RAND_2 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_1 = _RAND_2[21:0];
  _RAND_3 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_2 = _RAND_3[21:0];
  _RAND_4 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_3 = _RAND_4[21:0];
  _RAND_5 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_4 = _RAND_5[21:0];
  _RAND_6 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_5 = _RAND_6[21:0];
  _RAND_7 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_6 = _RAND_7[21:0];
  _RAND_8 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_7 = _RAND_8[21:0];
  _RAND_9 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_8 = _RAND_9[21:0];
  _RAND_10 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_9 = _RAND_10[21:0];
  _RAND_11 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_10 = _RAND_11[21:0];
  _RAND_12 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_11 = _RAND_12[21:0];
  _RAND_13 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_12 = _RAND_13[21:0];
  _RAND_14 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_13 = _RAND_14[21:0];
  _RAND_15 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_14 = _RAND_15[21:0];
  _RAND_16 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_15 = _RAND_16[21:0];
  _RAND_17 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_16 = _RAND_17[21:0];
  _RAND_18 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_17 = _RAND_18[21:0];
  _RAND_19 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_18 = _RAND_19[21:0];
  _RAND_20 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_19 = _RAND_20[21:0];
  _RAND_21 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_20 = _RAND_21[21:0];
  _RAND_22 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_21 = _RAND_22[21:0];
  _RAND_23 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_22 = _RAND_23[21:0];
  _RAND_24 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_23 = _RAND_24[21:0];
  _RAND_25 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_24 = _RAND_25[21:0];
  _RAND_26 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_25 = _RAND_26[21:0];
  _RAND_27 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_26 = _RAND_27[21:0];
  _RAND_28 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_27 = _RAND_28[21:0];
  _RAND_29 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_28 = _RAND_29[21:0];
  _RAND_30 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_29 = _RAND_30[21:0];
  _RAND_31 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_30 = _RAND_31[21:0];
  _RAND_32 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_31 = _RAND_32[21:0];
  _RAND_33 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_32 = _RAND_33[21:0];
  _RAND_34 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_33 = _RAND_34[21:0];
  _RAND_35 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_34 = _RAND_35[21:0];
  _RAND_36 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_35 = _RAND_36[21:0];
  _RAND_37 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_36 = _RAND_37[21:0];
  _RAND_38 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_37 = _RAND_38[21:0];
  _RAND_39 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_38 = _RAND_39[21:0];
  _RAND_40 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_39 = _RAND_40[21:0];
  _RAND_41 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_40 = _RAND_41[21:0];
  _RAND_42 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_41 = _RAND_42[21:0];
  _RAND_43 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_42 = _RAND_43[21:0];
  _RAND_44 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_43 = _RAND_44[21:0];
  _RAND_45 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_44 = _RAND_45[21:0];
  _RAND_46 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_45 = _RAND_46[21:0];
  _RAND_47 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_46 = _RAND_47[21:0];
  _RAND_48 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_47 = _RAND_48[21:0];
  _RAND_49 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_48 = _RAND_49[21:0];
  _RAND_50 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_49 = _RAND_50[21:0];
  _RAND_51 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_50 = _RAND_51[21:0];
  _RAND_52 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_51 = _RAND_52[21:0];
  _RAND_53 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_52 = _RAND_53[21:0];
  _RAND_54 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_53 = _RAND_54[21:0];
  _RAND_55 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_54 = _RAND_55[21:0];
  _RAND_56 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_55 = _RAND_56[21:0];
  _RAND_57 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_56 = _RAND_57[21:0];
  _RAND_58 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_57 = _RAND_58[21:0];
  _RAND_59 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_58 = _RAND_59[21:0];
  _RAND_60 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_59 = _RAND_60[21:0];
  _RAND_61 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_60 = _RAND_61[21:0];
  _RAND_62 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_61 = _RAND_62[21:0];
  _RAND_63 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_62 = _RAND_63[21:0];
  _RAND_64 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_63 = _RAND_64[21:0];
  _RAND_65 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_64 = _RAND_65[21:0];
  _RAND_66 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_65 = _RAND_66[21:0];
  _RAND_67 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_66 = _RAND_67[21:0];
  _RAND_68 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_67 = _RAND_68[21:0];
  _RAND_69 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_68 = _RAND_69[21:0];
  _RAND_70 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_69 = _RAND_70[21:0];
  _RAND_71 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_70 = _RAND_71[21:0];
  _RAND_72 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_71 = _RAND_72[21:0];
  _RAND_73 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_72 = _RAND_73[21:0];
  _RAND_74 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_73 = _RAND_74[21:0];
  _RAND_75 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_74 = _RAND_75[21:0];
  _RAND_76 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_75 = _RAND_76[21:0];
  _RAND_77 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_76 = _RAND_77[21:0];
  _RAND_78 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_77 = _RAND_78[21:0];
  _RAND_79 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_78 = _RAND_79[21:0];
  _RAND_80 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_79 = _RAND_80[21:0];
  _RAND_81 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_80 = _RAND_81[21:0];
  _RAND_82 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_81 = _RAND_82[21:0];
  _RAND_83 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_82 = _RAND_83[21:0];
  _RAND_84 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_83 = _RAND_84[21:0];
  _RAND_85 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_84 = _RAND_85[21:0];
  _RAND_86 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_85 = _RAND_86[21:0];
  _RAND_87 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_86 = _RAND_87[21:0];
  _RAND_88 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_87 = _RAND_88[21:0];
  _RAND_89 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_88 = _RAND_89[21:0];
  _RAND_90 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_89 = _RAND_90[21:0];
  _RAND_91 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_90 = _RAND_91[21:0];
  _RAND_92 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_91 = _RAND_92[21:0];
  _RAND_93 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_92 = _RAND_93[21:0];
  _RAND_94 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_93 = _RAND_94[21:0];
  _RAND_95 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_94 = _RAND_95[21:0];
  _RAND_96 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_95 = _RAND_96[21:0];
  _RAND_97 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_96 = _RAND_97[21:0];
  _RAND_98 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_97 = _RAND_98[21:0];
  _RAND_99 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_98 = _RAND_99[21:0];
  _RAND_100 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_99 = _RAND_100[21:0];
  _RAND_101 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_100 = _RAND_101[21:0];
  _RAND_102 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_101 = _RAND_102[21:0];
  _RAND_103 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_102 = _RAND_103[21:0];
  _RAND_104 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_103 = _RAND_104[21:0];
  _RAND_105 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_104 = _RAND_105[21:0];
  _RAND_106 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_105 = _RAND_106[21:0];
  _RAND_107 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_106 = _RAND_107[21:0];
  _RAND_108 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_107 = _RAND_108[21:0];
  _RAND_109 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_108 = _RAND_109[21:0];
  _RAND_110 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_109 = _RAND_110[21:0];
  _RAND_111 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_110 = _RAND_111[21:0];
  _RAND_112 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_111 = _RAND_112[21:0];
  _RAND_113 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_112 = _RAND_113[21:0];
  _RAND_114 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_113 = _RAND_114[21:0];
  _RAND_115 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_114 = _RAND_115[21:0];
  _RAND_116 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_115 = _RAND_116[21:0];
  _RAND_117 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_116 = _RAND_117[21:0];
  _RAND_118 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_117 = _RAND_118[21:0];
  _RAND_119 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_118 = _RAND_119[21:0];
  _RAND_120 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_119 = _RAND_120[21:0];
  _RAND_121 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_120 = _RAND_121[21:0];
  _RAND_122 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_121 = _RAND_122[21:0];
  _RAND_123 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_122 = _RAND_123[21:0];
  _RAND_124 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_123 = _RAND_124[21:0];
  _RAND_125 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_124 = _RAND_125[21:0];
  _RAND_126 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_125 = _RAND_126[21:0];
  _RAND_127 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_126 = _RAND_127[21:0];
  _RAND_128 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_127 = _RAND_128[21:0];
  _RAND_129 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_128 = _RAND_129[21:0];
  _RAND_130 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_129 = _RAND_130[21:0];
  _RAND_131 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_130 = _RAND_131[21:0];
  _RAND_132 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_131 = _RAND_132[21:0];
  _RAND_133 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_132 = _RAND_133[21:0];
  _RAND_134 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_133 = _RAND_134[21:0];
  _RAND_135 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_134 = _RAND_135[21:0];
  _RAND_136 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_135 = _RAND_136[21:0];
  _RAND_137 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_136 = _RAND_137[21:0];
  _RAND_138 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_137 = _RAND_138[21:0];
  _RAND_139 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_138 = _RAND_139[21:0];
  _RAND_140 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_139 = _RAND_140[21:0];
  _RAND_141 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_140 = _RAND_141[21:0];
  _RAND_142 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_141 = _RAND_142[21:0];
  _RAND_143 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_142 = _RAND_143[21:0];
  _RAND_144 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_143 = _RAND_144[21:0];
  _RAND_145 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_144 = _RAND_145[21:0];
  _RAND_146 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_145 = _RAND_146[21:0];
  _RAND_147 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_146 = _RAND_147[21:0];
  _RAND_148 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_147 = _RAND_148[21:0];
  _RAND_149 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_148 = _RAND_149[21:0];
  _RAND_150 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_149 = _RAND_150[21:0];
  _RAND_151 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_150 = _RAND_151[21:0];
  _RAND_152 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_151 = _RAND_152[21:0];
  _RAND_153 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_152 = _RAND_153[21:0];
  _RAND_154 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_153 = _RAND_154[21:0];
  _RAND_155 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_154 = _RAND_155[21:0];
  _RAND_156 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_155 = _RAND_156[21:0];
  _RAND_157 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_156 = _RAND_157[21:0];
  _RAND_158 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_157 = _RAND_158[21:0];
  _RAND_159 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_158 = _RAND_159[21:0];
  _RAND_160 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_159 = _RAND_160[21:0];
  _RAND_161 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_160 = _RAND_161[21:0];
  _RAND_162 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_161 = _RAND_162[21:0];
  _RAND_163 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_162 = _RAND_163[21:0];
  _RAND_164 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_163 = _RAND_164[21:0];
  _RAND_165 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_164 = _RAND_165[21:0];
  _RAND_166 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_165 = _RAND_166[21:0];
  _RAND_167 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_166 = _RAND_167[21:0];
  _RAND_168 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_167 = _RAND_168[21:0];
  _RAND_169 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_168 = _RAND_169[21:0];
  _RAND_170 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_169 = _RAND_170[21:0];
  _RAND_171 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_170 = _RAND_171[21:0];
  _RAND_172 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_171 = _RAND_172[21:0];
  _RAND_173 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_172 = _RAND_173[21:0];
  _RAND_174 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_173 = _RAND_174[21:0];
  _RAND_175 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_174 = _RAND_175[21:0];
  _RAND_176 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_175 = _RAND_176[21:0];
  _RAND_177 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_176 = _RAND_177[21:0];
  _RAND_178 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_177 = _RAND_178[21:0];
  _RAND_179 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_178 = _RAND_179[21:0];
  _RAND_180 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_179 = _RAND_180[21:0];
  _RAND_181 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_180 = _RAND_181[21:0];
  _RAND_182 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_181 = _RAND_182[21:0];
  _RAND_183 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_182 = _RAND_183[21:0];
  _RAND_184 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_183 = _RAND_184[21:0];
  _RAND_185 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_184 = _RAND_185[21:0];
  _RAND_186 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_185 = _RAND_186[21:0];
  _RAND_187 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_186 = _RAND_187[21:0];
  _RAND_188 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_187 = _RAND_188[21:0];
  _RAND_189 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_188 = _RAND_189[21:0];
  _RAND_190 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_189 = _RAND_190[21:0];
  _RAND_191 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_190 = _RAND_191[21:0];
  _RAND_192 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_191 = _RAND_192[21:0];
  _RAND_193 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_192 = _RAND_193[21:0];
  _RAND_194 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_193 = _RAND_194[21:0];
  _RAND_195 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_194 = _RAND_195[21:0];
  _RAND_196 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_195 = _RAND_196[21:0];
  _RAND_197 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_196 = _RAND_197[21:0];
  _RAND_198 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_197 = _RAND_198[21:0];
  _RAND_199 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_198 = _RAND_199[21:0];
  _RAND_200 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_199 = _RAND_200[21:0];
  _RAND_201 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_200 = _RAND_201[21:0];
  _RAND_202 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_201 = _RAND_202[21:0];
  _RAND_203 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_202 = _RAND_203[21:0];
  _RAND_204 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_203 = _RAND_204[21:0];
  _RAND_205 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_204 = _RAND_205[21:0];
  _RAND_206 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_205 = _RAND_206[21:0];
  _RAND_207 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_206 = _RAND_207[21:0];
  _RAND_208 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_207 = _RAND_208[21:0];
  _RAND_209 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_208 = _RAND_209[21:0];
  _RAND_210 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_209 = _RAND_210[21:0];
  _RAND_211 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_210 = _RAND_211[21:0];
  _RAND_212 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_211 = _RAND_212[21:0];
  _RAND_213 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_212 = _RAND_213[21:0];
  _RAND_214 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_213 = _RAND_214[21:0];
  _RAND_215 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_214 = _RAND_215[21:0];
  _RAND_216 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_215 = _RAND_216[21:0];
  _RAND_217 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_216 = _RAND_217[21:0];
  _RAND_218 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_217 = _RAND_218[21:0];
  _RAND_219 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_218 = _RAND_219[21:0];
  _RAND_220 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_219 = _RAND_220[21:0];
  _RAND_221 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_220 = _RAND_221[21:0];
  _RAND_222 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_221 = _RAND_222[21:0];
  _RAND_223 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_222 = _RAND_223[21:0];
  _RAND_224 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_223 = _RAND_224[21:0];
  _RAND_225 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_224 = _RAND_225[21:0];
  _RAND_226 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_225 = _RAND_226[21:0];
  _RAND_227 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_226 = _RAND_227[21:0];
  _RAND_228 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_227 = _RAND_228[21:0];
  _RAND_229 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_228 = _RAND_229[21:0];
  _RAND_230 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_229 = _RAND_230[21:0];
  _RAND_231 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_230 = _RAND_231[21:0];
  _RAND_232 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_231 = _RAND_232[21:0];
  _RAND_233 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_232 = _RAND_233[21:0];
  _RAND_234 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_233 = _RAND_234[21:0];
  _RAND_235 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_234 = _RAND_235[21:0];
  _RAND_236 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_235 = _RAND_236[21:0];
  _RAND_237 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_236 = _RAND_237[21:0];
  _RAND_238 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_237 = _RAND_238[21:0];
  _RAND_239 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_238 = _RAND_239[21:0];
  _RAND_240 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_239 = _RAND_240[21:0];
  _RAND_241 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_240 = _RAND_241[21:0];
  _RAND_242 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_241 = _RAND_242[21:0];
  _RAND_243 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_242 = _RAND_243[21:0];
  _RAND_244 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_243 = _RAND_244[21:0];
  _RAND_245 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_244 = _RAND_245[21:0];
  _RAND_246 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_245 = _RAND_246[21:0];
  _RAND_247 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_246 = _RAND_247[21:0];
  _RAND_248 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_247 = _RAND_248[21:0];
  _RAND_249 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_248 = _RAND_249[21:0];
  _RAND_250 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_249 = _RAND_250[21:0];
  _RAND_251 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_250 = _RAND_251[21:0];
  _RAND_252 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_251 = _RAND_252[21:0];
  _RAND_253 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_252 = _RAND_253[21:0];
  _RAND_254 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_253 = _RAND_254[21:0];
  _RAND_255 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_254 = _RAND_255[21:0];
  _RAND_256 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_255 = _RAND_256[21:0];
  _RAND_257 = {1{`RANDOM}};
  dec_tlu_way_wb_f = _RAND_257[0:0];
  _RAND_258 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_0 = _RAND_258[21:0];
  _RAND_259 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_1 = _RAND_259[21:0];
  _RAND_260 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_2 = _RAND_260[21:0];
  _RAND_261 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_3 = _RAND_261[21:0];
  _RAND_262 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_4 = _RAND_262[21:0];
  _RAND_263 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_5 = _RAND_263[21:0];
  _RAND_264 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_6 = _RAND_264[21:0];
  _RAND_265 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_7 = _RAND_265[21:0];
  _RAND_266 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_8 = _RAND_266[21:0];
  _RAND_267 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_9 = _RAND_267[21:0];
  _RAND_268 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_10 = _RAND_268[21:0];
  _RAND_269 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_11 = _RAND_269[21:0];
  _RAND_270 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_12 = _RAND_270[21:0];
  _RAND_271 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_13 = _RAND_271[21:0];
  _RAND_272 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_14 = _RAND_272[21:0];
  _RAND_273 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_15 = _RAND_273[21:0];
  _RAND_274 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_16 = _RAND_274[21:0];
  _RAND_275 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_17 = _RAND_275[21:0];
  _RAND_276 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_18 = _RAND_276[21:0];
  _RAND_277 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_19 = _RAND_277[21:0];
  _RAND_278 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_20 = _RAND_278[21:0];
  _RAND_279 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_21 = _RAND_279[21:0];
  _RAND_280 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_22 = _RAND_280[21:0];
  _RAND_281 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_23 = _RAND_281[21:0];
  _RAND_282 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_24 = _RAND_282[21:0];
  _RAND_283 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_25 = _RAND_283[21:0];
  _RAND_284 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_26 = _RAND_284[21:0];
  _RAND_285 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_27 = _RAND_285[21:0];
  _RAND_286 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_28 = _RAND_286[21:0];
  _RAND_287 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_29 = _RAND_287[21:0];
  _RAND_288 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_30 = _RAND_288[21:0];
  _RAND_289 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_31 = _RAND_289[21:0];
  _RAND_290 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_32 = _RAND_290[21:0];
  _RAND_291 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_33 = _RAND_291[21:0];
  _RAND_292 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_34 = _RAND_292[21:0];
  _RAND_293 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_35 = _RAND_293[21:0];
  _RAND_294 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_36 = _RAND_294[21:0];
  _RAND_295 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_37 = _RAND_295[21:0];
  _RAND_296 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_38 = _RAND_296[21:0];
  _RAND_297 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_39 = _RAND_297[21:0];
  _RAND_298 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_40 = _RAND_298[21:0];
  _RAND_299 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_41 = _RAND_299[21:0];
  _RAND_300 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_42 = _RAND_300[21:0];
  _RAND_301 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_43 = _RAND_301[21:0];
  _RAND_302 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_44 = _RAND_302[21:0];
  _RAND_303 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_45 = _RAND_303[21:0];
  _RAND_304 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_46 = _RAND_304[21:0];
  _RAND_305 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_47 = _RAND_305[21:0];
  _RAND_306 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_48 = _RAND_306[21:0];
  _RAND_307 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_49 = _RAND_307[21:0];
  _RAND_308 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_50 = _RAND_308[21:0];
  _RAND_309 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_51 = _RAND_309[21:0];
  _RAND_310 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_52 = _RAND_310[21:0];
  _RAND_311 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_53 = _RAND_311[21:0];
  _RAND_312 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_54 = _RAND_312[21:0];
  _RAND_313 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_55 = _RAND_313[21:0];
  _RAND_314 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_56 = _RAND_314[21:0];
  _RAND_315 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_57 = _RAND_315[21:0];
  _RAND_316 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_58 = _RAND_316[21:0];
  _RAND_317 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_59 = _RAND_317[21:0];
  _RAND_318 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_60 = _RAND_318[21:0];
  _RAND_319 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_61 = _RAND_319[21:0];
  _RAND_320 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_62 = _RAND_320[21:0];
  _RAND_321 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_63 = _RAND_321[21:0];
  _RAND_322 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_64 = _RAND_322[21:0];
  _RAND_323 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_65 = _RAND_323[21:0];
  _RAND_324 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_66 = _RAND_324[21:0];
  _RAND_325 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_67 = _RAND_325[21:0];
  _RAND_326 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_68 = _RAND_326[21:0];
  _RAND_327 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_69 = _RAND_327[21:0];
  _RAND_328 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_70 = _RAND_328[21:0];
  _RAND_329 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_71 = _RAND_329[21:0];
  _RAND_330 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_72 = _RAND_330[21:0];
  _RAND_331 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_73 = _RAND_331[21:0];
  _RAND_332 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_74 = _RAND_332[21:0];
  _RAND_333 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_75 = _RAND_333[21:0];
  _RAND_334 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_76 = _RAND_334[21:0];
  _RAND_335 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_77 = _RAND_335[21:0];
  _RAND_336 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_78 = _RAND_336[21:0];
  _RAND_337 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_79 = _RAND_337[21:0];
  _RAND_338 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_80 = _RAND_338[21:0];
  _RAND_339 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_81 = _RAND_339[21:0];
  _RAND_340 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_82 = _RAND_340[21:0];
  _RAND_341 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_83 = _RAND_341[21:0];
  _RAND_342 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_84 = _RAND_342[21:0];
  _RAND_343 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_85 = _RAND_343[21:0];
  _RAND_344 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_86 = _RAND_344[21:0];
  _RAND_345 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_87 = _RAND_345[21:0];
  _RAND_346 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_88 = _RAND_346[21:0];
  _RAND_347 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_89 = _RAND_347[21:0];
  _RAND_348 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_90 = _RAND_348[21:0];
  _RAND_349 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_91 = _RAND_349[21:0];
  _RAND_350 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_92 = _RAND_350[21:0];
  _RAND_351 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_93 = _RAND_351[21:0];
  _RAND_352 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_94 = _RAND_352[21:0];
  _RAND_353 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_95 = _RAND_353[21:0];
  _RAND_354 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_96 = _RAND_354[21:0];
  _RAND_355 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_97 = _RAND_355[21:0];
  _RAND_356 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_98 = _RAND_356[21:0];
  _RAND_357 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_99 = _RAND_357[21:0];
  _RAND_358 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_100 = _RAND_358[21:0];
  _RAND_359 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_101 = _RAND_359[21:0];
  _RAND_360 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_102 = _RAND_360[21:0];
  _RAND_361 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_103 = _RAND_361[21:0];
  _RAND_362 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_104 = _RAND_362[21:0];
  _RAND_363 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_105 = _RAND_363[21:0];
  _RAND_364 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_106 = _RAND_364[21:0];
  _RAND_365 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_107 = _RAND_365[21:0];
  _RAND_366 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_108 = _RAND_366[21:0];
  _RAND_367 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_109 = _RAND_367[21:0];
  _RAND_368 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_110 = _RAND_368[21:0];
  _RAND_369 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_111 = _RAND_369[21:0];
  _RAND_370 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_112 = _RAND_370[21:0];
  _RAND_371 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_113 = _RAND_371[21:0];
  _RAND_372 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_114 = _RAND_372[21:0];
  _RAND_373 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_115 = _RAND_373[21:0];
  _RAND_374 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_116 = _RAND_374[21:0];
  _RAND_375 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_117 = _RAND_375[21:0];
  _RAND_376 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_118 = _RAND_376[21:0];
  _RAND_377 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_119 = _RAND_377[21:0];
  _RAND_378 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_120 = _RAND_378[21:0];
  _RAND_379 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_121 = _RAND_379[21:0];
  _RAND_380 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_122 = _RAND_380[21:0];
  _RAND_381 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_123 = _RAND_381[21:0];
  _RAND_382 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_124 = _RAND_382[21:0];
  _RAND_383 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_125 = _RAND_383[21:0];
  _RAND_384 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_126 = _RAND_384[21:0];
  _RAND_385 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_127 = _RAND_385[21:0];
  _RAND_386 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_128 = _RAND_386[21:0];
  _RAND_387 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_129 = _RAND_387[21:0];
  _RAND_388 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_130 = _RAND_388[21:0];
  _RAND_389 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_131 = _RAND_389[21:0];
  _RAND_390 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_132 = _RAND_390[21:0];
  _RAND_391 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_133 = _RAND_391[21:0];
  _RAND_392 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_134 = _RAND_392[21:0];
  _RAND_393 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_135 = _RAND_393[21:0];
  _RAND_394 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_136 = _RAND_394[21:0];
  _RAND_395 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_137 = _RAND_395[21:0];
  _RAND_396 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_138 = _RAND_396[21:0];
  _RAND_397 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_139 = _RAND_397[21:0];
  _RAND_398 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_140 = _RAND_398[21:0];
  _RAND_399 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_141 = _RAND_399[21:0];
  _RAND_400 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_142 = _RAND_400[21:0];
  _RAND_401 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_143 = _RAND_401[21:0];
  _RAND_402 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_144 = _RAND_402[21:0];
  _RAND_403 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_145 = _RAND_403[21:0];
  _RAND_404 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_146 = _RAND_404[21:0];
  _RAND_405 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_147 = _RAND_405[21:0];
  _RAND_406 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_148 = _RAND_406[21:0];
  _RAND_407 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_149 = _RAND_407[21:0];
  _RAND_408 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_150 = _RAND_408[21:0];
  _RAND_409 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_151 = _RAND_409[21:0];
  _RAND_410 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_152 = _RAND_410[21:0];
  _RAND_411 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_153 = _RAND_411[21:0];
  _RAND_412 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_154 = _RAND_412[21:0];
  _RAND_413 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_155 = _RAND_413[21:0];
  _RAND_414 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_156 = _RAND_414[21:0];
  _RAND_415 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_157 = _RAND_415[21:0];
  _RAND_416 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_158 = _RAND_416[21:0];
  _RAND_417 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_159 = _RAND_417[21:0];
  _RAND_418 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_160 = _RAND_418[21:0];
  _RAND_419 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_161 = _RAND_419[21:0];
  _RAND_420 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_162 = _RAND_420[21:0];
  _RAND_421 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_163 = _RAND_421[21:0];
  _RAND_422 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_164 = _RAND_422[21:0];
  _RAND_423 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_165 = _RAND_423[21:0];
  _RAND_424 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_166 = _RAND_424[21:0];
  _RAND_425 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_167 = _RAND_425[21:0];
  _RAND_426 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_168 = _RAND_426[21:0];
  _RAND_427 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_169 = _RAND_427[21:0];
  _RAND_428 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_170 = _RAND_428[21:0];
  _RAND_429 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_171 = _RAND_429[21:0];
  _RAND_430 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_172 = _RAND_430[21:0];
  _RAND_431 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_173 = _RAND_431[21:0];
  _RAND_432 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_174 = _RAND_432[21:0];
  _RAND_433 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_175 = _RAND_433[21:0];
  _RAND_434 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_176 = _RAND_434[21:0];
  _RAND_435 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_177 = _RAND_435[21:0];
  _RAND_436 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_178 = _RAND_436[21:0];
  _RAND_437 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_179 = _RAND_437[21:0];
  _RAND_438 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_180 = _RAND_438[21:0];
  _RAND_439 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_181 = _RAND_439[21:0];
  _RAND_440 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_182 = _RAND_440[21:0];
  _RAND_441 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_183 = _RAND_441[21:0];
  _RAND_442 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_184 = _RAND_442[21:0];
  _RAND_443 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_185 = _RAND_443[21:0];
  _RAND_444 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_186 = _RAND_444[21:0];
  _RAND_445 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_187 = _RAND_445[21:0];
  _RAND_446 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_188 = _RAND_446[21:0];
  _RAND_447 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_189 = _RAND_447[21:0];
  _RAND_448 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_190 = _RAND_448[21:0];
  _RAND_449 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_191 = _RAND_449[21:0];
  _RAND_450 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_192 = _RAND_450[21:0];
  _RAND_451 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_193 = _RAND_451[21:0];
  _RAND_452 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_194 = _RAND_452[21:0];
  _RAND_453 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_195 = _RAND_453[21:0];
  _RAND_454 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_196 = _RAND_454[21:0];
  _RAND_455 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_197 = _RAND_455[21:0];
  _RAND_456 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_198 = _RAND_456[21:0];
  _RAND_457 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_199 = _RAND_457[21:0];
  _RAND_458 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_200 = _RAND_458[21:0];
  _RAND_459 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_201 = _RAND_459[21:0];
  _RAND_460 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_202 = _RAND_460[21:0];
  _RAND_461 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_203 = _RAND_461[21:0];
  _RAND_462 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_204 = _RAND_462[21:0];
  _RAND_463 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_205 = _RAND_463[21:0];
  _RAND_464 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_206 = _RAND_464[21:0];
  _RAND_465 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_207 = _RAND_465[21:0];
  _RAND_466 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_208 = _RAND_466[21:0];
  _RAND_467 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_209 = _RAND_467[21:0];
  _RAND_468 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_210 = _RAND_468[21:0];
  _RAND_469 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_211 = _RAND_469[21:0];
  _RAND_470 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_212 = _RAND_470[21:0];
  _RAND_471 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_213 = _RAND_471[21:0];
  _RAND_472 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_214 = _RAND_472[21:0];
  _RAND_473 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_215 = _RAND_473[21:0];
  _RAND_474 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_216 = _RAND_474[21:0];
  _RAND_475 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_217 = _RAND_475[21:0];
  _RAND_476 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_218 = _RAND_476[21:0];
  _RAND_477 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_219 = _RAND_477[21:0];
  _RAND_478 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_220 = _RAND_478[21:0];
  _RAND_479 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_221 = _RAND_479[21:0];
  _RAND_480 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_222 = _RAND_480[21:0];
  _RAND_481 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_223 = _RAND_481[21:0];
  _RAND_482 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_224 = _RAND_482[21:0];
  _RAND_483 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_225 = _RAND_483[21:0];
  _RAND_484 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_226 = _RAND_484[21:0];
  _RAND_485 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_227 = _RAND_485[21:0];
  _RAND_486 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_228 = _RAND_486[21:0];
  _RAND_487 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_229 = _RAND_487[21:0];
  _RAND_488 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_230 = _RAND_488[21:0];
  _RAND_489 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_231 = _RAND_489[21:0];
  _RAND_490 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_232 = _RAND_490[21:0];
  _RAND_491 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_233 = _RAND_491[21:0];
  _RAND_492 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_234 = _RAND_492[21:0];
  _RAND_493 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_235 = _RAND_493[21:0];
  _RAND_494 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_236 = _RAND_494[21:0];
  _RAND_495 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_237 = _RAND_495[21:0];
  _RAND_496 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_238 = _RAND_496[21:0];
  _RAND_497 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_239 = _RAND_497[21:0];
  _RAND_498 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_240 = _RAND_498[21:0];
  _RAND_499 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_241 = _RAND_499[21:0];
  _RAND_500 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_242 = _RAND_500[21:0];
  _RAND_501 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_243 = _RAND_501[21:0];
  _RAND_502 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_244 = _RAND_502[21:0];
  _RAND_503 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_245 = _RAND_503[21:0];
  _RAND_504 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_246 = _RAND_504[21:0];
  _RAND_505 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_247 = _RAND_505[21:0];
  _RAND_506 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_248 = _RAND_506[21:0];
  _RAND_507 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_249 = _RAND_507[21:0];
  _RAND_508 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_250 = _RAND_508[21:0];
  _RAND_509 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_251 = _RAND_509[21:0];
  _RAND_510 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_252 = _RAND_510[21:0];
  _RAND_511 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_253 = _RAND_511[21:0];
  _RAND_512 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_254 = _RAND_512[21:0];
  _RAND_513 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_255 = _RAND_513[21:0];
  _RAND_514 = {1{`RANDOM}};
  fghr = _RAND_514[7:0];
  _RAND_515 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_0 = _RAND_515[1:0];
  _RAND_516 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_1 = _RAND_516[1:0];
  _RAND_517 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_2 = _RAND_517[1:0];
  _RAND_518 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_3 = _RAND_518[1:0];
  _RAND_519 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_4 = _RAND_519[1:0];
  _RAND_520 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_5 = _RAND_520[1:0];
  _RAND_521 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_6 = _RAND_521[1:0];
  _RAND_522 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_7 = _RAND_522[1:0];
  _RAND_523 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_8 = _RAND_523[1:0];
  _RAND_524 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_9 = _RAND_524[1:0];
  _RAND_525 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_10 = _RAND_525[1:0];
  _RAND_526 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_11 = _RAND_526[1:0];
  _RAND_527 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_12 = _RAND_527[1:0];
  _RAND_528 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_13 = _RAND_528[1:0];
  _RAND_529 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_14 = _RAND_529[1:0];
  _RAND_530 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_15 = _RAND_530[1:0];
  _RAND_531 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_16 = _RAND_531[1:0];
  _RAND_532 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_17 = _RAND_532[1:0];
  _RAND_533 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_18 = _RAND_533[1:0];
  _RAND_534 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_19 = _RAND_534[1:0];
  _RAND_535 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_20 = _RAND_535[1:0];
  _RAND_536 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_21 = _RAND_536[1:0];
  _RAND_537 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_22 = _RAND_537[1:0];
  _RAND_538 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_23 = _RAND_538[1:0];
  _RAND_539 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_24 = _RAND_539[1:0];
  _RAND_540 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_25 = _RAND_540[1:0];
  _RAND_541 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_26 = _RAND_541[1:0];
  _RAND_542 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_27 = _RAND_542[1:0];
  _RAND_543 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_28 = _RAND_543[1:0];
  _RAND_544 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_29 = _RAND_544[1:0];
  _RAND_545 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_30 = _RAND_545[1:0];
  _RAND_546 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_31 = _RAND_546[1:0];
  _RAND_547 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_32 = _RAND_547[1:0];
  _RAND_548 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_33 = _RAND_548[1:0];
  _RAND_549 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_34 = _RAND_549[1:0];
  _RAND_550 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_35 = _RAND_550[1:0];
  _RAND_551 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_36 = _RAND_551[1:0];
  _RAND_552 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_37 = _RAND_552[1:0];
  _RAND_553 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_38 = _RAND_553[1:0];
  _RAND_554 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_39 = _RAND_554[1:0];
  _RAND_555 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_40 = _RAND_555[1:0];
  _RAND_556 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_41 = _RAND_556[1:0];
  _RAND_557 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_42 = _RAND_557[1:0];
  _RAND_558 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_43 = _RAND_558[1:0];
  _RAND_559 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_44 = _RAND_559[1:0];
  _RAND_560 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_45 = _RAND_560[1:0];
  _RAND_561 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_46 = _RAND_561[1:0];
  _RAND_562 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_47 = _RAND_562[1:0];
  _RAND_563 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_48 = _RAND_563[1:0];
  _RAND_564 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_49 = _RAND_564[1:0];
  _RAND_565 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_50 = _RAND_565[1:0];
  _RAND_566 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_51 = _RAND_566[1:0];
  _RAND_567 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_52 = _RAND_567[1:0];
  _RAND_568 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_53 = _RAND_568[1:0];
  _RAND_569 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_54 = _RAND_569[1:0];
  _RAND_570 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_55 = _RAND_570[1:0];
  _RAND_571 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_56 = _RAND_571[1:0];
  _RAND_572 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_57 = _RAND_572[1:0];
  _RAND_573 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_58 = _RAND_573[1:0];
  _RAND_574 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_59 = _RAND_574[1:0];
  _RAND_575 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_60 = _RAND_575[1:0];
  _RAND_576 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_61 = _RAND_576[1:0];
  _RAND_577 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_62 = _RAND_577[1:0];
  _RAND_578 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_63 = _RAND_578[1:0];
  _RAND_579 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_64 = _RAND_579[1:0];
  _RAND_580 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_65 = _RAND_580[1:0];
  _RAND_581 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_66 = _RAND_581[1:0];
  _RAND_582 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_67 = _RAND_582[1:0];
  _RAND_583 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_68 = _RAND_583[1:0];
  _RAND_584 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_69 = _RAND_584[1:0];
  _RAND_585 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_70 = _RAND_585[1:0];
  _RAND_586 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_71 = _RAND_586[1:0];
  _RAND_587 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_72 = _RAND_587[1:0];
  _RAND_588 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_73 = _RAND_588[1:0];
  _RAND_589 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_74 = _RAND_589[1:0];
  _RAND_590 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_75 = _RAND_590[1:0];
  _RAND_591 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_76 = _RAND_591[1:0];
  _RAND_592 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_77 = _RAND_592[1:0];
  _RAND_593 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_78 = _RAND_593[1:0];
  _RAND_594 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_79 = _RAND_594[1:0];
  _RAND_595 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_80 = _RAND_595[1:0];
  _RAND_596 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_81 = _RAND_596[1:0];
  _RAND_597 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_82 = _RAND_597[1:0];
  _RAND_598 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_83 = _RAND_598[1:0];
  _RAND_599 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_84 = _RAND_599[1:0];
  _RAND_600 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_85 = _RAND_600[1:0];
  _RAND_601 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_86 = _RAND_601[1:0];
  _RAND_602 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_87 = _RAND_602[1:0];
  _RAND_603 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_88 = _RAND_603[1:0];
  _RAND_604 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_89 = _RAND_604[1:0];
  _RAND_605 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_90 = _RAND_605[1:0];
  _RAND_606 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_91 = _RAND_606[1:0];
  _RAND_607 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_92 = _RAND_607[1:0];
  _RAND_608 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_93 = _RAND_608[1:0];
  _RAND_609 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_94 = _RAND_609[1:0];
  _RAND_610 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_95 = _RAND_610[1:0];
  _RAND_611 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_96 = _RAND_611[1:0];
  _RAND_612 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_97 = _RAND_612[1:0];
  _RAND_613 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_98 = _RAND_613[1:0];
  _RAND_614 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_99 = _RAND_614[1:0];
  _RAND_615 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_100 = _RAND_615[1:0];
  _RAND_616 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_101 = _RAND_616[1:0];
  _RAND_617 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_102 = _RAND_617[1:0];
  _RAND_618 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_103 = _RAND_618[1:0];
  _RAND_619 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_104 = _RAND_619[1:0];
  _RAND_620 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_105 = _RAND_620[1:0];
  _RAND_621 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_106 = _RAND_621[1:0];
  _RAND_622 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_107 = _RAND_622[1:0];
  _RAND_623 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_108 = _RAND_623[1:0];
  _RAND_624 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_109 = _RAND_624[1:0];
  _RAND_625 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_110 = _RAND_625[1:0];
  _RAND_626 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_111 = _RAND_626[1:0];
  _RAND_627 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_112 = _RAND_627[1:0];
  _RAND_628 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_113 = _RAND_628[1:0];
  _RAND_629 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_114 = _RAND_629[1:0];
  _RAND_630 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_115 = _RAND_630[1:0];
  _RAND_631 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_116 = _RAND_631[1:0];
  _RAND_632 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_117 = _RAND_632[1:0];
  _RAND_633 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_118 = _RAND_633[1:0];
  _RAND_634 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_119 = _RAND_634[1:0];
  _RAND_635 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_120 = _RAND_635[1:0];
  _RAND_636 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_121 = _RAND_636[1:0];
  _RAND_637 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_122 = _RAND_637[1:0];
  _RAND_638 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_123 = _RAND_638[1:0];
  _RAND_639 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_124 = _RAND_639[1:0];
  _RAND_640 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_125 = _RAND_640[1:0];
  _RAND_641 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_126 = _RAND_641[1:0];
  _RAND_642 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_127 = _RAND_642[1:0];
  _RAND_643 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_128 = _RAND_643[1:0];
  _RAND_644 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_129 = _RAND_644[1:0];
  _RAND_645 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_130 = _RAND_645[1:0];
  _RAND_646 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_131 = _RAND_646[1:0];
  _RAND_647 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_132 = _RAND_647[1:0];
  _RAND_648 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_133 = _RAND_648[1:0];
  _RAND_649 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_134 = _RAND_649[1:0];
  _RAND_650 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_135 = _RAND_650[1:0];
  _RAND_651 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_136 = _RAND_651[1:0];
  _RAND_652 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_137 = _RAND_652[1:0];
  _RAND_653 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_138 = _RAND_653[1:0];
  _RAND_654 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_139 = _RAND_654[1:0];
  _RAND_655 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_140 = _RAND_655[1:0];
  _RAND_656 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_141 = _RAND_656[1:0];
  _RAND_657 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_142 = _RAND_657[1:0];
  _RAND_658 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_143 = _RAND_658[1:0];
  _RAND_659 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_144 = _RAND_659[1:0];
  _RAND_660 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_145 = _RAND_660[1:0];
  _RAND_661 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_146 = _RAND_661[1:0];
  _RAND_662 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_147 = _RAND_662[1:0];
  _RAND_663 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_148 = _RAND_663[1:0];
  _RAND_664 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_149 = _RAND_664[1:0];
  _RAND_665 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_150 = _RAND_665[1:0];
  _RAND_666 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_151 = _RAND_666[1:0];
  _RAND_667 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_152 = _RAND_667[1:0];
  _RAND_668 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_153 = _RAND_668[1:0];
  _RAND_669 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_154 = _RAND_669[1:0];
  _RAND_670 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_155 = _RAND_670[1:0];
  _RAND_671 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_156 = _RAND_671[1:0];
  _RAND_672 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_157 = _RAND_672[1:0];
  _RAND_673 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_158 = _RAND_673[1:0];
  _RAND_674 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_159 = _RAND_674[1:0];
  _RAND_675 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_160 = _RAND_675[1:0];
  _RAND_676 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_161 = _RAND_676[1:0];
  _RAND_677 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_162 = _RAND_677[1:0];
  _RAND_678 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_163 = _RAND_678[1:0];
  _RAND_679 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_164 = _RAND_679[1:0];
  _RAND_680 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_165 = _RAND_680[1:0];
  _RAND_681 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_166 = _RAND_681[1:0];
  _RAND_682 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_167 = _RAND_682[1:0];
  _RAND_683 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_168 = _RAND_683[1:0];
  _RAND_684 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_169 = _RAND_684[1:0];
  _RAND_685 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_170 = _RAND_685[1:0];
  _RAND_686 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_171 = _RAND_686[1:0];
  _RAND_687 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_172 = _RAND_687[1:0];
  _RAND_688 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_173 = _RAND_688[1:0];
  _RAND_689 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_174 = _RAND_689[1:0];
  _RAND_690 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_175 = _RAND_690[1:0];
  _RAND_691 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_176 = _RAND_691[1:0];
  _RAND_692 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_177 = _RAND_692[1:0];
  _RAND_693 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_178 = _RAND_693[1:0];
  _RAND_694 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_179 = _RAND_694[1:0];
  _RAND_695 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_180 = _RAND_695[1:0];
  _RAND_696 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_181 = _RAND_696[1:0];
  _RAND_697 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_182 = _RAND_697[1:0];
  _RAND_698 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_183 = _RAND_698[1:0];
  _RAND_699 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_184 = _RAND_699[1:0];
  _RAND_700 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_185 = _RAND_700[1:0];
  _RAND_701 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_186 = _RAND_701[1:0];
  _RAND_702 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_187 = _RAND_702[1:0];
  _RAND_703 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_188 = _RAND_703[1:0];
  _RAND_704 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_189 = _RAND_704[1:0];
  _RAND_705 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_190 = _RAND_705[1:0];
  _RAND_706 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_191 = _RAND_706[1:0];
  _RAND_707 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_192 = _RAND_707[1:0];
  _RAND_708 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_193 = _RAND_708[1:0];
  _RAND_709 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_194 = _RAND_709[1:0];
  _RAND_710 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_195 = _RAND_710[1:0];
  _RAND_711 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_196 = _RAND_711[1:0];
  _RAND_712 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_197 = _RAND_712[1:0];
  _RAND_713 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_198 = _RAND_713[1:0];
  _RAND_714 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_199 = _RAND_714[1:0];
  _RAND_715 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_200 = _RAND_715[1:0];
  _RAND_716 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_201 = _RAND_716[1:0];
  _RAND_717 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_202 = _RAND_717[1:0];
  _RAND_718 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_203 = _RAND_718[1:0];
  _RAND_719 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_204 = _RAND_719[1:0];
  _RAND_720 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_205 = _RAND_720[1:0];
  _RAND_721 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_206 = _RAND_721[1:0];
  _RAND_722 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_207 = _RAND_722[1:0];
  _RAND_723 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_208 = _RAND_723[1:0];
  _RAND_724 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_209 = _RAND_724[1:0];
  _RAND_725 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_210 = _RAND_725[1:0];
  _RAND_726 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_211 = _RAND_726[1:0];
  _RAND_727 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_212 = _RAND_727[1:0];
  _RAND_728 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_213 = _RAND_728[1:0];
  _RAND_729 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_214 = _RAND_729[1:0];
  _RAND_730 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_215 = _RAND_730[1:0];
  _RAND_731 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_216 = _RAND_731[1:0];
  _RAND_732 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_217 = _RAND_732[1:0];
  _RAND_733 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_218 = _RAND_733[1:0];
  _RAND_734 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_219 = _RAND_734[1:0];
  _RAND_735 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_220 = _RAND_735[1:0];
  _RAND_736 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_221 = _RAND_736[1:0];
  _RAND_737 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_222 = _RAND_737[1:0];
  _RAND_738 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_223 = _RAND_738[1:0];
  _RAND_739 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_224 = _RAND_739[1:0];
  _RAND_740 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_225 = _RAND_740[1:0];
  _RAND_741 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_226 = _RAND_741[1:0];
  _RAND_742 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_227 = _RAND_742[1:0];
  _RAND_743 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_228 = _RAND_743[1:0];
  _RAND_744 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_229 = _RAND_744[1:0];
  _RAND_745 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_230 = _RAND_745[1:0];
  _RAND_746 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_231 = _RAND_746[1:0];
  _RAND_747 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_232 = _RAND_747[1:0];
  _RAND_748 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_233 = _RAND_748[1:0];
  _RAND_749 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_234 = _RAND_749[1:0];
  _RAND_750 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_235 = _RAND_750[1:0];
  _RAND_751 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_236 = _RAND_751[1:0];
  _RAND_752 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_237 = _RAND_752[1:0];
  _RAND_753 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_238 = _RAND_753[1:0];
  _RAND_754 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_239 = _RAND_754[1:0];
  _RAND_755 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_240 = _RAND_755[1:0];
  _RAND_756 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_241 = _RAND_756[1:0];
  _RAND_757 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_242 = _RAND_757[1:0];
  _RAND_758 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_243 = _RAND_758[1:0];
  _RAND_759 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_244 = _RAND_759[1:0];
  _RAND_760 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_245 = _RAND_760[1:0];
  _RAND_761 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_246 = _RAND_761[1:0];
  _RAND_762 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_247 = _RAND_762[1:0];
  _RAND_763 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_248 = _RAND_763[1:0];
  _RAND_764 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_249 = _RAND_764[1:0];
  _RAND_765 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_250 = _RAND_765[1:0];
  _RAND_766 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_251 = _RAND_766[1:0];
  _RAND_767 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_252 = _RAND_767[1:0];
  _RAND_768 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_253 = _RAND_768[1:0];
  _RAND_769 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_254 = _RAND_769[1:0];
  _RAND_770 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_255 = _RAND_770[1:0];
  _RAND_771 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_0 = _RAND_771[1:0];
  _RAND_772 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_1 = _RAND_772[1:0];
  _RAND_773 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_2 = _RAND_773[1:0];
  _RAND_774 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_3 = _RAND_774[1:0];
  _RAND_775 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_4 = _RAND_775[1:0];
  _RAND_776 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_5 = _RAND_776[1:0];
  _RAND_777 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_6 = _RAND_777[1:0];
  _RAND_778 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_7 = _RAND_778[1:0];
  _RAND_779 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_8 = _RAND_779[1:0];
  _RAND_780 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_9 = _RAND_780[1:0];
  _RAND_781 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_10 = _RAND_781[1:0];
  _RAND_782 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_11 = _RAND_782[1:0];
  _RAND_783 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_12 = _RAND_783[1:0];
  _RAND_784 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_13 = _RAND_784[1:0];
  _RAND_785 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_14 = _RAND_785[1:0];
  _RAND_786 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_15 = _RAND_786[1:0];
  _RAND_787 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_16 = _RAND_787[1:0];
  _RAND_788 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_17 = _RAND_788[1:0];
  _RAND_789 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_18 = _RAND_789[1:0];
  _RAND_790 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_19 = _RAND_790[1:0];
  _RAND_791 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_20 = _RAND_791[1:0];
  _RAND_792 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_21 = _RAND_792[1:0];
  _RAND_793 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_22 = _RAND_793[1:0];
  _RAND_794 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_23 = _RAND_794[1:0];
  _RAND_795 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_24 = _RAND_795[1:0];
  _RAND_796 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_25 = _RAND_796[1:0];
  _RAND_797 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_26 = _RAND_797[1:0];
  _RAND_798 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_27 = _RAND_798[1:0];
  _RAND_799 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_28 = _RAND_799[1:0];
  _RAND_800 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_29 = _RAND_800[1:0];
  _RAND_801 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_30 = _RAND_801[1:0];
  _RAND_802 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_31 = _RAND_802[1:0];
  _RAND_803 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_32 = _RAND_803[1:0];
  _RAND_804 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_33 = _RAND_804[1:0];
  _RAND_805 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_34 = _RAND_805[1:0];
  _RAND_806 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_35 = _RAND_806[1:0];
  _RAND_807 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_36 = _RAND_807[1:0];
  _RAND_808 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_37 = _RAND_808[1:0];
  _RAND_809 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_38 = _RAND_809[1:0];
  _RAND_810 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_39 = _RAND_810[1:0];
  _RAND_811 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_40 = _RAND_811[1:0];
  _RAND_812 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_41 = _RAND_812[1:0];
  _RAND_813 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_42 = _RAND_813[1:0];
  _RAND_814 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_43 = _RAND_814[1:0];
  _RAND_815 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_44 = _RAND_815[1:0];
  _RAND_816 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_45 = _RAND_816[1:0];
  _RAND_817 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_46 = _RAND_817[1:0];
  _RAND_818 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_47 = _RAND_818[1:0];
  _RAND_819 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_48 = _RAND_819[1:0];
  _RAND_820 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_49 = _RAND_820[1:0];
  _RAND_821 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_50 = _RAND_821[1:0];
  _RAND_822 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_51 = _RAND_822[1:0];
  _RAND_823 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_52 = _RAND_823[1:0];
  _RAND_824 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_53 = _RAND_824[1:0];
  _RAND_825 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_54 = _RAND_825[1:0];
  _RAND_826 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_55 = _RAND_826[1:0];
  _RAND_827 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_56 = _RAND_827[1:0];
  _RAND_828 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_57 = _RAND_828[1:0];
  _RAND_829 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_58 = _RAND_829[1:0];
  _RAND_830 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_59 = _RAND_830[1:0];
  _RAND_831 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_60 = _RAND_831[1:0];
  _RAND_832 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_61 = _RAND_832[1:0];
  _RAND_833 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_62 = _RAND_833[1:0];
  _RAND_834 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_63 = _RAND_834[1:0];
  _RAND_835 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_64 = _RAND_835[1:0];
  _RAND_836 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_65 = _RAND_836[1:0];
  _RAND_837 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_66 = _RAND_837[1:0];
  _RAND_838 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_67 = _RAND_838[1:0];
  _RAND_839 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_68 = _RAND_839[1:0];
  _RAND_840 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_69 = _RAND_840[1:0];
  _RAND_841 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_70 = _RAND_841[1:0];
  _RAND_842 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_71 = _RAND_842[1:0];
  _RAND_843 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_72 = _RAND_843[1:0];
  _RAND_844 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_73 = _RAND_844[1:0];
  _RAND_845 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_74 = _RAND_845[1:0];
  _RAND_846 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_75 = _RAND_846[1:0];
  _RAND_847 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_76 = _RAND_847[1:0];
  _RAND_848 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_77 = _RAND_848[1:0];
  _RAND_849 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_78 = _RAND_849[1:0];
  _RAND_850 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_79 = _RAND_850[1:0];
  _RAND_851 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_80 = _RAND_851[1:0];
  _RAND_852 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_81 = _RAND_852[1:0];
  _RAND_853 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_82 = _RAND_853[1:0];
  _RAND_854 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_83 = _RAND_854[1:0];
  _RAND_855 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_84 = _RAND_855[1:0];
  _RAND_856 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_85 = _RAND_856[1:0];
  _RAND_857 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_86 = _RAND_857[1:0];
  _RAND_858 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_87 = _RAND_858[1:0];
  _RAND_859 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_88 = _RAND_859[1:0];
  _RAND_860 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_89 = _RAND_860[1:0];
  _RAND_861 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_90 = _RAND_861[1:0];
  _RAND_862 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_91 = _RAND_862[1:0];
  _RAND_863 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_92 = _RAND_863[1:0];
  _RAND_864 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_93 = _RAND_864[1:0];
  _RAND_865 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_94 = _RAND_865[1:0];
  _RAND_866 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_95 = _RAND_866[1:0];
  _RAND_867 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_96 = _RAND_867[1:0];
  _RAND_868 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_97 = _RAND_868[1:0];
  _RAND_869 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_98 = _RAND_869[1:0];
  _RAND_870 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_99 = _RAND_870[1:0];
  _RAND_871 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_100 = _RAND_871[1:0];
  _RAND_872 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_101 = _RAND_872[1:0];
  _RAND_873 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_102 = _RAND_873[1:0];
  _RAND_874 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_103 = _RAND_874[1:0];
  _RAND_875 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_104 = _RAND_875[1:0];
  _RAND_876 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_105 = _RAND_876[1:0];
  _RAND_877 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_106 = _RAND_877[1:0];
  _RAND_878 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_107 = _RAND_878[1:0];
  _RAND_879 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_108 = _RAND_879[1:0];
  _RAND_880 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_109 = _RAND_880[1:0];
  _RAND_881 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_110 = _RAND_881[1:0];
  _RAND_882 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_111 = _RAND_882[1:0];
  _RAND_883 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_112 = _RAND_883[1:0];
  _RAND_884 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_113 = _RAND_884[1:0];
  _RAND_885 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_114 = _RAND_885[1:0];
  _RAND_886 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_115 = _RAND_886[1:0];
  _RAND_887 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_116 = _RAND_887[1:0];
  _RAND_888 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_117 = _RAND_888[1:0];
  _RAND_889 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_118 = _RAND_889[1:0];
  _RAND_890 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_119 = _RAND_890[1:0];
  _RAND_891 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_120 = _RAND_891[1:0];
  _RAND_892 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_121 = _RAND_892[1:0];
  _RAND_893 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_122 = _RAND_893[1:0];
  _RAND_894 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_123 = _RAND_894[1:0];
  _RAND_895 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_124 = _RAND_895[1:0];
  _RAND_896 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_125 = _RAND_896[1:0];
  _RAND_897 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_126 = _RAND_897[1:0];
  _RAND_898 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_127 = _RAND_898[1:0];
  _RAND_899 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_128 = _RAND_899[1:0];
  _RAND_900 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_129 = _RAND_900[1:0];
  _RAND_901 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_130 = _RAND_901[1:0];
  _RAND_902 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_131 = _RAND_902[1:0];
  _RAND_903 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_132 = _RAND_903[1:0];
  _RAND_904 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_133 = _RAND_904[1:0];
  _RAND_905 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_134 = _RAND_905[1:0];
  _RAND_906 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_135 = _RAND_906[1:0];
  _RAND_907 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_136 = _RAND_907[1:0];
  _RAND_908 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_137 = _RAND_908[1:0];
  _RAND_909 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_138 = _RAND_909[1:0];
  _RAND_910 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_139 = _RAND_910[1:0];
  _RAND_911 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_140 = _RAND_911[1:0];
  _RAND_912 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_141 = _RAND_912[1:0];
  _RAND_913 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_142 = _RAND_913[1:0];
  _RAND_914 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_143 = _RAND_914[1:0];
  _RAND_915 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_144 = _RAND_915[1:0];
  _RAND_916 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_145 = _RAND_916[1:0];
  _RAND_917 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_146 = _RAND_917[1:0];
  _RAND_918 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_147 = _RAND_918[1:0];
  _RAND_919 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_148 = _RAND_919[1:0];
  _RAND_920 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_149 = _RAND_920[1:0];
  _RAND_921 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_150 = _RAND_921[1:0];
  _RAND_922 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_151 = _RAND_922[1:0];
  _RAND_923 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_152 = _RAND_923[1:0];
  _RAND_924 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_153 = _RAND_924[1:0];
  _RAND_925 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_154 = _RAND_925[1:0];
  _RAND_926 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_155 = _RAND_926[1:0];
  _RAND_927 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_156 = _RAND_927[1:0];
  _RAND_928 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_157 = _RAND_928[1:0];
  _RAND_929 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_158 = _RAND_929[1:0];
  _RAND_930 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_159 = _RAND_930[1:0];
  _RAND_931 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_160 = _RAND_931[1:0];
  _RAND_932 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_161 = _RAND_932[1:0];
  _RAND_933 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_162 = _RAND_933[1:0];
  _RAND_934 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_163 = _RAND_934[1:0];
  _RAND_935 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_164 = _RAND_935[1:0];
  _RAND_936 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_165 = _RAND_936[1:0];
  _RAND_937 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_166 = _RAND_937[1:0];
  _RAND_938 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_167 = _RAND_938[1:0];
  _RAND_939 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_168 = _RAND_939[1:0];
  _RAND_940 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_169 = _RAND_940[1:0];
  _RAND_941 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_170 = _RAND_941[1:0];
  _RAND_942 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_171 = _RAND_942[1:0];
  _RAND_943 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_172 = _RAND_943[1:0];
  _RAND_944 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_173 = _RAND_944[1:0];
  _RAND_945 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_174 = _RAND_945[1:0];
  _RAND_946 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_175 = _RAND_946[1:0];
  _RAND_947 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_176 = _RAND_947[1:0];
  _RAND_948 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_177 = _RAND_948[1:0];
  _RAND_949 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_178 = _RAND_949[1:0];
  _RAND_950 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_179 = _RAND_950[1:0];
  _RAND_951 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_180 = _RAND_951[1:0];
  _RAND_952 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_181 = _RAND_952[1:0];
  _RAND_953 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_182 = _RAND_953[1:0];
  _RAND_954 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_183 = _RAND_954[1:0];
  _RAND_955 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_184 = _RAND_955[1:0];
  _RAND_956 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_185 = _RAND_956[1:0];
  _RAND_957 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_186 = _RAND_957[1:0];
  _RAND_958 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_187 = _RAND_958[1:0];
  _RAND_959 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_188 = _RAND_959[1:0];
  _RAND_960 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_189 = _RAND_960[1:0];
  _RAND_961 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_190 = _RAND_961[1:0];
  _RAND_962 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_191 = _RAND_962[1:0];
  _RAND_963 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_192 = _RAND_963[1:0];
  _RAND_964 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_193 = _RAND_964[1:0];
  _RAND_965 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_194 = _RAND_965[1:0];
  _RAND_966 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_195 = _RAND_966[1:0];
  _RAND_967 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_196 = _RAND_967[1:0];
  _RAND_968 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_197 = _RAND_968[1:0];
  _RAND_969 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_198 = _RAND_969[1:0];
  _RAND_970 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_199 = _RAND_970[1:0];
  _RAND_971 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_200 = _RAND_971[1:0];
  _RAND_972 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_201 = _RAND_972[1:0];
  _RAND_973 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_202 = _RAND_973[1:0];
  _RAND_974 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_203 = _RAND_974[1:0];
  _RAND_975 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_204 = _RAND_975[1:0];
  _RAND_976 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_205 = _RAND_976[1:0];
  _RAND_977 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_206 = _RAND_977[1:0];
  _RAND_978 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_207 = _RAND_978[1:0];
  _RAND_979 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_208 = _RAND_979[1:0];
  _RAND_980 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_209 = _RAND_980[1:0];
  _RAND_981 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_210 = _RAND_981[1:0];
  _RAND_982 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_211 = _RAND_982[1:0];
  _RAND_983 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_212 = _RAND_983[1:0];
  _RAND_984 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_213 = _RAND_984[1:0];
  _RAND_985 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_214 = _RAND_985[1:0];
  _RAND_986 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_215 = _RAND_986[1:0];
  _RAND_987 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_216 = _RAND_987[1:0];
  _RAND_988 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_217 = _RAND_988[1:0];
  _RAND_989 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_218 = _RAND_989[1:0];
  _RAND_990 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_219 = _RAND_990[1:0];
  _RAND_991 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_220 = _RAND_991[1:0];
  _RAND_992 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_221 = _RAND_992[1:0];
  _RAND_993 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_222 = _RAND_993[1:0];
  _RAND_994 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_223 = _RAND_994[1:0];
  _RAND_995 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_224 = _RAND_995[1:0];
  _RAND_996 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_225 = _RAND_996[1:0];
  _RAND_997 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_226 = _RAND_997[1:0];
  _RAND_998 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_227 = _RAND_998[1:0];
  _RAND_999 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_228 = _RAND_999[1:0];
  _RAND_1000 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_229 = _RAND_1000[1:0];
  _RAND_1001 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_230 = _RAND_1001[1:0];
  _RAND_1002 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_231 = _RAND_1002[1:0];
  _RAND_1003 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_232 = _RAND_1003[1:0];
  _RAND_1004 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_233 = _RAND_1004[1:0];
  _RAND_1005 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_234 = _RAND_1005[1:0];
  _RAND_1006 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_235 = _RAND_1006[1:0];
  _RAND_1007 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_236 = _RAND_1007[1:0];
  _RAND_1008 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_237 = _RAND_1008[1:0];
  _RAND_1009 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_238 = _RAND_1009[1:0];
  _RAND_1010 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_239 = _RAND_1010[1:0];
  _RAND_1011 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_240 = _RAND_1011[1:0];
  _RAND_1012 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_241 = _RAND_1012[1:0];
  _RAND_1013 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_242 = _RAND_1013[1:0];
  _RAND_1014 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_243 = _RAND_1014[1:0];
  _RAND_1015 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_244 = _RAND_1015[1:0];
  _RAND_1016 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_245 = _RAND_1016[1:0];
  _RAND_1017 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_246 = _RAND_1017[1:0];
  _RAND_1018 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_247 = _RAND_1018[1:0];
  _RAND_1019 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_248 = _RAND_1019[1:0];
  _RAND_1020 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_249 = _RAND_1020[1:0];
  _RAND_1021 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_250 = _RAND_1021[1:0];
  _RAND_1022 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_251 = _RAND_1022[1:0];
  _RAND_1023 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_252 = _RAND_1023[1:0];
  _RAND_1024 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_253 = _RAND_1024[1:0];
  _RAND_1025 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_254 = _RAND_1025[1:0];
  _RAND_1026 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_255 = _RAND_1026[1:0];
  _RAND_1027 = {1{`RANDOM}};
  exu_mp_way_f = _RAND_1027[0:0];
  _RAND_1028 = {1{`RANDOM}};
  exu_flush_final_d1 = _RAND_1028[0:0];
  _RAND_1029 = {8{`RANDOM}};
  btb_lru_b0_f = _RAND_1029[255:0];
  _RAND_1030 = {1{`RANDOM}};
  ifc_fetch_adder_prior = _RAND_1030[29:0];
  _RAND_1031 = {1{`RANDOM}};
  rets_out_0 = _RAND_1031[31:0];
  _RAND_1032 = {1{`RANDOM}};
  rets_out_1 = _RAND_1032[31:0];
  _RAND_1033 = {1{`RANDOM}};
  rets_out_2 = _RAND_1033[31:0];
  _RAND_1034 = {1{`RANDOM}};
  rets_out_3 = _RAND_1034[31:0];
  _RAND_1035 = {1{`RANDOM}};
  rets_out_4 = _RAND_1035[31:0];
  _RAND_1036 = {1{`RANDOM}};
  rets_out_5 = _RAND_1036[31:0];
  _RAND_1037 = {1{`RANDOM}};
  rets_out_6 = _RAND_1037[31:0];
  _RAND_1038 = {1{`RANDOM}};
  rets_out_7 = _RAND_1038[31:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    leak_one_f_d1 = 1'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_0 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_1 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_2 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_3 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_4 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_5 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_6 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_7 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_8 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_9 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_10 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_11 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_12 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_13 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_14 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_15 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_16 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_17 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_18 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_19 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_20 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_21 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_22 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_23 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_24 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_25 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_26 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_27 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_28 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_29 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_30 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_31 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_32 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_33 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_34 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_35 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_36 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_37 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_38 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_39 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_40 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_41 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_42 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_43 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_44 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_45 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_46 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_47 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_48 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_49 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_50 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_51 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_52 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_53 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_54 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_55 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_56 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_57 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_58 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_59 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_60 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_61 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_62 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_63 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_64 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_65 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_66 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_67 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_68 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_69 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_70 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_71 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_72 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_73 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_74 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_75 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_76 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_77 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_78 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_79 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_80 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_81 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_82 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_83 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_84 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_85 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_86 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_87 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_88 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_89 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_90 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_91 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_92 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_93 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_94 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_95 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_96 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_97 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_98 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_99 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_100 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_101 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_102 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_103 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_104 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_105 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_106 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_107 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_108 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_109 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_110 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_111 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_112 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_113 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_114 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_115 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_116 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_117 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_118 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_119 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_120 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_121 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_122 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_123 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_124 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_125 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_126 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_127 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_128 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_129 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_130 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_131 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_132 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_133 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_134 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_135 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_136 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_137 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_138 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_139 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_140 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_141 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_142 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_143 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_144 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_145 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_146 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_147 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_148 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_149 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_150 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_151 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_152 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_153 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_154 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_155 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_156 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_157 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_158 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_159 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_160 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_161 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_162 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_163 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_164 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_165 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_166 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_167 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_168 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_169 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_170 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_171 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_172 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_173 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_174 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_175 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_176 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_177 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_178 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_179 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_180 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_181 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_182 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_183 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_184 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_185 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_186 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_187 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_188 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_189 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_190 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_191 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_192 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_193 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_194 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_195 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_196 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_197 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_198 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_199 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_200 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_201 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_202 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_203 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_204 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_205 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_206 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_207 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_208 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_209 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_210 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_211 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_212 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_213 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_214 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_215 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_216 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_217 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_218 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_219 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_220 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_221 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_222 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_223 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_224 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_225 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_226 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_227 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_228 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_229 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_230 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_231 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_232 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_233 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_234 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_235 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_236 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_237 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_238 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_239 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_240 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_241 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_242 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_243 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_244 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_245 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_246 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_247 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_248 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_249 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_250 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_251 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_252 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_253 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_254 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_255 = 22'h0;
  end
  if (reset) begin
    dec_tlu_way_wb_f = 1'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_0 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_1 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_2 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_3 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_4 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_5 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_6 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_7 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_8 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_9 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_10 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_11 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_12 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_13 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_14 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_15 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_16 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_17 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_18 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_19 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_20 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_21 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_22 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_23 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_24 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_25 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_26 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_27 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_28 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_29 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_30 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_31 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_32 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_33 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_34 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_35 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_36 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_37 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_38 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_39 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_40 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_41 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_42 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_43 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_44 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_45 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_46 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_47 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_48 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_49 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_50 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_51 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_52 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_53 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_54 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_55 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_56 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_57 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_58 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_59 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_60 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_61 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_62 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_63 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_64 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_65 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_66 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_67 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_68 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_69 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_70 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_71 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_72 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_73 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_74 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_75 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_76 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_77 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_78 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_79 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_80 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_81 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_82 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_83 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_84 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_85 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_86 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_87 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_88 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_89 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_90 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_91 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_92 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_93 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_94 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_95 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_96 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_97 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_98 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_99 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_100 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_101 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_102 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_103 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_104 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_105 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_106 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_107 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_108 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_109 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_110 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_111 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_112 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_113 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_114 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_115 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_116 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_117 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_118 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_119 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_120 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_121 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_122 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_123 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_124 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_125 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_126 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_127 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_128 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_129 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_130 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_131 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_132 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_133 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_134 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_135 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_136 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_137 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_138 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_139 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_140 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_141 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_142 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_143 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_144 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_145 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_146 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_147 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_148 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_149 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_150 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_151 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_152 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_153 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_154 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_155 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_156 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_157 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_158 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_159 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_160 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_161 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_162 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_163 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_164 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_165 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_166 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_167 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_168 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_169 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_170 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_171 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_172 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_173 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_174 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_175 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_176 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_177 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_178 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_179 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_180 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_181 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_182 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_183 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_184 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_185 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_186 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_187 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_188 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_189 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_190 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_191 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_192 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_193 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_194 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_195 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_196 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_197 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_198 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_199 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_200 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_201 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_202 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_203 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_204 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_205 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_206 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_207 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_208 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_209 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_210 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_211 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_212 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_213 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_214 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_215 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_216 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_217 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_218 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_219 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_220 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_221 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_222 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_223 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_224 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_225 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_226 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_227 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_228 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_229 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_230 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_231 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_232 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_233 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_234 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_235 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_236 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_237 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_238 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_239 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_240 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_241 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_242 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_243 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_244 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_245 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_246 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_247 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_248 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_249 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_250 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_251 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_252 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_253 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_254 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_255 = 22'h0;
  end
  if (reset) begin
    fghr = 8'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_0 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_1 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_2 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_3 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_4 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_5 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_6 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_7 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_8 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_9 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_10 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_11 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_12 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_13 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_14 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_15 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_16 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_17 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_18 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_19 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_20 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_21 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_22 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_23 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_24 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_25 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_26 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_27 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_28 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_29 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_30 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_31 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_32 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_33 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_34 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_35 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_36 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_37 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_38 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_39 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_40 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_41 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_42 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_43 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_44 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_45 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_46 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_47 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_48 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_49 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_50 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_51 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_52 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_53 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_54 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_55 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_56 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_57 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_58 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_59 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_60 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_61 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_62 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_63 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_64 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_65 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_66 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_67 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_68 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_69 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_70 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_71 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_72 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_73 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_74 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_75 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_76 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_77 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_78 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_79 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_80 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_81 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_82 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_83 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_84 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_85 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_86 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_87 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_88 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_89 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_90 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_91 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_92 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_93 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_94 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_95 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_96 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_97 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_98 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_99 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_100 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_101 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_102 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_103 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_104 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_105 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_106 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_107 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_108 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_109 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_110 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_111 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_112 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_113 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_114 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_115 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_116 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_117 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_118 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_119 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_120 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_121 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_122 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_123 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_124 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_125 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_126 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_127 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_128 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_129 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_130 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_131 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_132 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_133 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_134 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_135 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_136 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_137 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_138 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_139 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_140 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_141 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_142 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_143 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_144 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_145 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_146 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_147 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_148 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_149 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_150 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_151 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_152 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_153 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_154 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_155 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_156 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_157 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_158 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_159 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_160 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_161 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_162 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_163 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_164 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_165 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_166 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_167 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_168 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_169 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_170 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_171 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_172 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_173 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_174 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_175 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_176 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_177 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_178 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_179 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_180 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_181 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_182 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_183 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_184 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_185 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_186 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_187 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_188 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_189 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_190 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_191 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_192 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_193 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_194 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_195 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_196 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_197 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_198 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_199 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_200 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_201 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_202 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_203 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_204 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_205 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_206 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_207 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_208 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_209 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_210 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_211 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_212 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_213 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_214 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_215 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_216 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_217 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_218 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_219 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_220 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_221 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_222 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_223 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_224 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_225 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_226 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_227 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_228 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_229 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_230 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_231 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_232 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_233 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_234 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_235 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_236 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_237 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_238 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_239 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_240 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_241 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_242 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_243 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_244 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_245 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_246 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_247 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_248 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_249 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_250 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_251 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_252 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_253 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_254 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_255 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_0 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_1 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_2 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_3 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_4 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_5 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_6 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_7 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_8 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_9 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_10 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_11 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_12 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_13 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_14 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_15 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_16 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_17 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_18 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_19 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_20 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_21 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_22 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_23 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_24 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_25 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_26 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_27 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_28 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_29 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_30 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_31 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_32 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_33 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_34 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_35 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_36 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_37 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_38 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_39 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_40 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_41 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_42 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_43 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_44 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_45 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_46 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_47 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_48 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_49 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_50 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_51 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_52 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_53 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_54 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_55 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_56 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_57 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_58 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_59 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_60 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_61 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_62 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_63 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_64 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_65 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_66 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_67 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_68 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_69 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_70 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_71 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_72 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_73 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_74 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_75 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_76 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_77 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_78 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_79 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_80 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_81 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_82 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_83 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_84 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_85 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_86 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_87 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_88 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_89 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_90 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_91 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_92 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_93 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_94 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_95 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_96 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_97 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_98 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_99 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_100 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_101 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_102 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_103 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_104 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_105 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_106 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_107 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_108 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_109 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_110 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_111 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_112 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_113 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_114 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_115 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_116 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_117 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_118 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_119 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_120 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_121 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_122 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_123 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_124 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_125 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_126 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_127 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_128 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_129 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_130 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_131 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_132 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_133 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_134 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_135 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_136 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_137 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_138 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_139 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_140 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_141 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_142 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_143 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_144 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_145 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_146 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_147 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_148 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_149 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_150 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_151 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_152 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_153 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_154 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_155 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_156 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_157 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_158 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_159 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_160 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_161 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_162 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_163 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_164 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_165 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_166 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_167 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_168 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_169 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_170 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_171 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_172 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_173 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_174 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_175 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_176 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_177 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_178 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_179 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_180 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_181 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_182 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_183 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_184 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_185 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_186 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_187 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_188 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_189 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_190 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_191 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_192 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_193 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_194 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_195 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_196 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_197 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_198 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_199 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_200 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_201 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_202 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_203 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_204 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_205 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_206 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_207 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_208 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_209 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_210 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_211 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_212 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_213 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_214 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_215 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_216 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_217 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_218 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_219 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_220 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_221 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_222 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_223 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_224 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_225 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_226 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_227 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_228 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_229 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_230 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_231 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_232 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_233 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_234 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_235 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_236 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_237 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_238 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_239 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_240 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_241 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_242 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_243 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_244 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_245 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_246 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_247 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_248 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_249 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_250 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_251 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_252 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_253 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_254 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_255 = 2'h0;
  end
  if (reset) begin
    exu_mp_way_f = 1'h0;
  end
  if (reset) begin
    exu_flush_final_d1 = 1'h0;
  end
  if (reset) begin
    btb_lru_b0_f = 256'h0;
  end
  if (reset) begin
    ifc_fetch_adder_prior = 30'h0;
  end
  if (reset) begin
    rets_out_0 = 32'h0;
  end
  if (reset) begin
    rets_out_1 = 32'h0;
  end
  if (reset) begin
    rets_out_2 = 32'h0;
  end
  if (reset) begin
    rets_out_3 = 32'h0;
  end
  if (reset) begin
    rets_out_4 = 32'h0;
  end
  if (reset) begin
    rets_out_5 = 32'h0;
  end
  if (reset) begin
    rets_out_6 = 32'h0;
  end
  if (reset) begin
    rets_out_7 = 32'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      leak_one_f_d1 <= 1'h0;
    end else begin
      leak_one_f_d1 <= _T_40 | _T_42;
    end
  end
  always @(posedge rvclkhdr_10_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_0 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_0 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_11_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_1 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_1 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_12_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_2 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_2 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_13_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_3 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_3 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_14_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_4 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_4 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_15_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_5 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_5 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_16_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_6 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_6 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_17_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_7 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_7 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_18_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_8 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_8 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_19_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_9 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_9 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_20_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_10 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_10 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_21_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_11 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_11 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_22_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_12 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_12 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_23_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_13 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_13 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_24_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_14 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_14 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_25_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_15 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_15 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_26_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_16 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_16 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_27_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_17 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_17 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_28_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_18 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_18 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_29_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_19 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_19 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_30_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_20 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_20 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_31_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_21 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_21 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_32_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_22 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_22 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_33_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_23 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_23 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_34_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_24 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_24 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_35_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_25 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_25 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_36_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_26 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_26 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_37_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_27 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_27 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_38_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_28 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_28 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_39_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_29 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_29 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_40_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_30 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_30 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_41_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_31 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_31 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_42_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_32 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_32 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_43_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_33 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_33 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_44_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_34 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_34 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_45_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_35 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_35 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_46_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_36 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_36 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_47_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_37 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_37 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_48_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_38 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_38 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_49_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_39 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_39 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_50_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_40 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_40 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_51_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_41 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_41 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_52_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_42 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_42 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_53_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_43 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_43 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_54_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_44 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_44 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_55_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_45 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_45 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_56_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_46 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_46 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_57_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_47 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_47 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_58_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_48 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_48 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_59_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_49 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_49 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_60_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_50 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_50 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_61_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_51 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_51 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_62_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_52 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_52 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_63_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_53 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_53 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_64_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_54 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_54 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_65_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_55 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_55 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_66_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_56 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_56 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_67_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_57 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_57 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_68_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_58 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_58 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_69_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_59 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_59 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_70_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_60 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_60 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_71_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_61 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_61 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_72_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_62 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_62 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_73_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_63 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_63 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_74_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_64 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_64 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_75_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_65 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_65 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_76_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_66 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_66 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_77_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_67 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_67 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_78_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_68 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_68 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_79_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_69 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_69 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_80_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_70 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_70 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_81_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_71 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_71 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_82_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_72 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_72 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_83_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_73 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_73 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_84_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_74 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_74 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_85_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_75 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_75 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_76 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_76 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_77 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_77 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_78 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_78 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_79 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_79 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_80 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_80 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_81 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_81 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_82 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_82 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_83 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_83 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_94_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_84 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_84 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_95_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_85 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_85 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_96_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_86 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_86 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_97_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_87 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_87 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_98_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_88 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_88 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_99_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_89 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_89 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_100_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_90 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_90 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_101_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_91 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_91 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_102_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_92 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_92 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_103_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_93 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_93 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_104_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_94 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_94 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_105_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_95 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_95 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_106_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_96 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_96 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_107_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_97 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_97 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_108_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_98 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_98 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_109_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_99 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_99 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_110_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_100 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_100 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_111_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_101 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_101 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_112_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_102 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_102 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_113_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_103 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_103 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_114_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_104 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_104 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_115_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_105 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_105 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_116_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_106 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_106 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_117_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_107 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_107 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_118_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_108 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_108 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_119_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_109 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_109 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_120_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_110 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_110 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_121_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_111 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_111 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_122_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_112 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_112 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_123_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_113 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_113 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_124_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_114 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_114 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_125_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_115 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_115 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_126_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_116 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_116 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_127_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_117 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_117 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_128_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_118 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_118 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_129_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_119 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_119 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_130_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_120 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_120 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_131_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_121 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_121 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_132_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_122 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_122 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_133_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_123 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_123 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_134_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_124 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_124 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_135_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_125 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_125 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_136_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_126 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_126 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_137_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_127 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_127 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_138_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_128 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_128 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_139_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_129 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_129 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_140_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_130 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_130 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_141_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_131 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_131 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_142_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_132 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_132 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_143_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_133 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_133 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_144_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_134 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_134 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_145_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_135 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_135 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_146_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_136 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_136 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_147_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_137 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_137 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_148_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_138 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_138 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_149_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_139 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_139 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_150_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_140 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_140 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_151_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_141 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_141 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_152_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_142 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_142 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_153_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_143 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_143 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_154_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_144 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_144 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_155_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_145 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_145 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_156_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_146 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_146 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_157_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_147 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_147 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_158_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_148 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_148 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_159_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_149 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_149 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_160_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_150 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_150 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_161_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_151 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_151 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_162_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_152 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_152 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_163_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_153 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_153 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_164_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_154 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_154 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_165_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_155 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_155 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_166_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_156 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_156 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_167_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_157 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_157 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_168_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_158 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_158 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_169_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_159 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_159 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_170_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_160 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_160 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_171_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_161 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_161 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_172_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_162 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_162 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_173_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_163 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_163 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_174_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_164 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_164 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_175_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_165 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_165 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_176_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_166 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_166 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_177_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_167 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_167 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_178_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_168 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_168 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_179_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_169 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_169 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_180_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_170 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_170 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_181_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_171 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_171 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_182_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_172 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_172 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_183_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_173 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_173 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_184_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_174 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_174 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_185_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_175 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_175 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_186_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_176 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_176 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_187_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_177 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_177 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_188_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_178 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_178 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_189_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_179 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_179 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_190_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_180 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_180 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_191_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_181 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_181 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_192_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_182 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_182 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_193_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_183 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_183 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_194_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_184 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_184 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_195_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_185 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_185 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_196_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_186 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_186 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_197_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_187 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_187 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_198_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_188 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_188 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_199_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_189 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_189 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_200_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_190 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_190 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_201_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_191 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_191 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_202_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_192 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_192 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_203_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_193 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_193 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_204_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_194 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_194 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_205_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_195 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_195 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_206_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_196 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_196 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_207_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_197 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_197 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_208_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_198 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_198 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_209_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_199 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_199 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_210_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_200 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_200 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_211_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_201 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_201 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_212_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_202 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_202 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_213_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_203 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_203 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_214_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_204 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_204 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_215_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_205 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_205 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_216_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_206 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_206 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_217_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_207 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_207 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_218_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_208 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_208 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_219_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_209 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_209 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_220_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_210 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_210 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_221_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_211 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_211 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_222_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_212 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_212 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_223_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_213 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_213 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_224_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_214 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_214 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_225_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_215 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_215 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_226_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_216 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_216 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_227_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_217 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_217 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_228_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_218 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_218 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_229_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_219 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_219 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_230_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_220 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_220 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_231_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_221 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_221 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_232_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_222 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_222 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_233_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_223 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_223 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_234_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_224 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_224 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_235_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_225 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_225 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_236_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_226 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_226 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_237_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_227 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_227 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_238_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_228 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_228 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_239_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_229 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_229 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_240_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_230 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_230 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_241_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_231 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_231 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_242_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_232 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_232 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_243_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_233 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_233 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_244_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_234 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_234 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_245_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_235 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_235 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_246_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_236 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_236 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_247_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_237 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_237 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_248_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_238 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_238 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_249_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_239 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_239 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_250_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_240 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_240 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_251_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_241 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_241 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_252_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_242 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_242 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_253_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_243 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_243 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_254_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_244 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_244 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_255_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_245 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_245 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_256_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_246 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_246 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_257_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_247 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_247 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_258_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_248 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_248 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_259_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_249 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_249 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_260_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_250 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_250 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_261_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_251 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_251 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_262_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_252 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_252 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_263_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_253 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_253 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_264_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_254 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_254 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_265_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_255 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_255 <= {_T_538,_T_535};
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      dec_tlu_way_wb_f <= 1'h0;
    end else begin
      dec_tlu_way_wb_f <= io_dec_bp_dec_tlu_br0_r_pkt_bits_way;
    end
  end
  always @(posedge rvclkhdr_266_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_0 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_0 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_267_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_1 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_1 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_268_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_2 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_2 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_269_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_3 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_3 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_270_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_4 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_4 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_271_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_5 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_5 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_272_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_6 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_6 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_273_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_7 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_7 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_274_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_8 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_8 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_275_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_9 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_9 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_276_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_10 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_10 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_277_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_11 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_11 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_278_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_12 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_12 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_279_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_13 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_13 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_280_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_14 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_14 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_281_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_15 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_15 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_282_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_16 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_16 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_283_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_17 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_17 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_284_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_18 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_18 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_285_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_19 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_19 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_286_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_20 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_20 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_287_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_21 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_21 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_288_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_22 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_22 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_289_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_23 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_23 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_290_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_24 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_24 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_291_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_25 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_25 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_292_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_26 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_26 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_293_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_27 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_27 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_294_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_28 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_28 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_295_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_29 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_29 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_296_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_30 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_30 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_297_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_31 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_31 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_298_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_32 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_32 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_299_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_33 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_33 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_300_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_34 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_34 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_301_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_35 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_35 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_302_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_36 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_36 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_303_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_37 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_37 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_304_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_38 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_38 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_305_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_39 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_39 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_306_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_40 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_40 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_307_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_41 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_41 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_308_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_42 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_42 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_309_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_43 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_43 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_310_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_44 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_44 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_311_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_45 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_45 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_312_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_46 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_46 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_313_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_47 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_47 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_314_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_48 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_48 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_315_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_49 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_49 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_316_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_50 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_50 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_317_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_51 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_51 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_318_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_52 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_52 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_319_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_53 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_53 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_320_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_54 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_54 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_321_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_55 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_55 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_322_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_56 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_56 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_323_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_57 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_57 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_324_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_58 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_58 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_325_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_59 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_59 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_326_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_60 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_60 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_327_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_61 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_61 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_328_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_62 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_62 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_329_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_63 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_63 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_330_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_64 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_64 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_331_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_65 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_65 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_332_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_66 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_66 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_333_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_67 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_67 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_334_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_68 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_68 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_335_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_69 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_69 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_336_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_70 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_70 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_337_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_71 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_71 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_338_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_72 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_72 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_339_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_73 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_73 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_340_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_74 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_74 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_341_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_75 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_75 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_342_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_76 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_76 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_343_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_77 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_77 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_344_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_78 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_78 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_345_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_79 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_79 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_346_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_80 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_80 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_347_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_81 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_81 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_348_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_82 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_82 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_349_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_83 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_83 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_350_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_84 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_84 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_351_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_85 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_85 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_352_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_86 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_86 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_353_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_87 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_87 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_354_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_88 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_88 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_355_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_89 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_89 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_356_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_90 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_90 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_357_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_91 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_91 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_358_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_92 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_92 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_359_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_93 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_93 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_360_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_94 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_94 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_361_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_95 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_95 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_362_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_96 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_96 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_363_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_97 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_97 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_364_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_98 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_98 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_365_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_99 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_99 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_366_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_100 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_100 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_367_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_101 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_101 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_368_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_102 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_102 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_369_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_103 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_103 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_370_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_104 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_104 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_371_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_105 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_105 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_372_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_106 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_106 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_373_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_107 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_107 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_374_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_108 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_108 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_375_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_109 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_109 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_376_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_110 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_110 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_377_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_111 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_111 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_378_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_112 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_112 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_379_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_113 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_113 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_380_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_114 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_114 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_381_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_115 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_115 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_382_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_116 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_116 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_383_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_117 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_117 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_384_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_118 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_118 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_385_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_119 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_119 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_386_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_120 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_120 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_387_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_121 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_121 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_388_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_122 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_122 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_389_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_123 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_123 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_390_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_124 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_124 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_391_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_125 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_125 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_392_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_126 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_126 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_393_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_127 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_127 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_394_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_128 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_128 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_395_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_129 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_129 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_396_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_130 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_130 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_397_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_131 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_131 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_398_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_132 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_132 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_399_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_133 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_133 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_400_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_134 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_134 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_401_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_135 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_135 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_402_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_136 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_136 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_403_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_137 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_137 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_404_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_138 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_138 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_405_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_139 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_139 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_406_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_140 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_140 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_407_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_141 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_141 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_408_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_142 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_142 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_409_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_143 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_143 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_410_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_144 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_144 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_411_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_145 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_145 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_412_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_146 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_146 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_413_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_147 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_147 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_414_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_148 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_148 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_415_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_149 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_149 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_416_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_150 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_150 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_417_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_151 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_151 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_418_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_152 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_152 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_419_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_153 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_153 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_420_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_154 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_154 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_421_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_155 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_155 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_422_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_156 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_156 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_423_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_157 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_157 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_424_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_158 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_158 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_425_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_159 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_159 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_426_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_160 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_160 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_427_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_161 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_161 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_428_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_162 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_162 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_429_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_163 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_163 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_430_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_164 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_164 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_431_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_165 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_165 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_432_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_166 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_166 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_433_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_167 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_167 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_434_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_168 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_168 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_435_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_169 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_169 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_436_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_170 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_170 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_437_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_171 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_171 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_438_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_172 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_172 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_439_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_173 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_173 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_440_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_174 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_174 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_441_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_175 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_175 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_442_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_176 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_176 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_443_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_177 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_177 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_444_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_178 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_178 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_445_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_179 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_179 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_446_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_180 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_180 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_447_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_181 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_181 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_448_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_182 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_182 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_449_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_183 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_183 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_450_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_184 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_184 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_451_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_185 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_185 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_452_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_186 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_186 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_453_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_187 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_187 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_454_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_188 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_188 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_455_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_189 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_189 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_456_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_190 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_190 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_457_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_191 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_191 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_458_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_192 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_192 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_459_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_193 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_193 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_460_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_194 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_194 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_461_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_195 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_195 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_462_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_196 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_196 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_463_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_197 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_197 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_464_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_198 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_198 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_465_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_199 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_199 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_466_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_200 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_200 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_467_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_201 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_201 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_468_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_202 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_202 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_469_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_203 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_203 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_470_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_204 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_204 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_471_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_205 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_205 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_472_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_206 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_206 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_473_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_207 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_207 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_474_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_208 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_208 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_475_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_209 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_209 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_476_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_210 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_210 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_477_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_211 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_211 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_478_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_212 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_212 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_479_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_213 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_213 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_480_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_214 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_214 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_481_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_215 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_215 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_482_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_216 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_216 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_483_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_217 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_217 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_484_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_218 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_218 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_485_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_219 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_219 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_486_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_220 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_220 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_487_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_221 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_221 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_488_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_222 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_222 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_489_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_223 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_223 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_490_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_224 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_224 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_491_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_225 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_225 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_492_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_226 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_226 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_493_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_227 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_227 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_494_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_228 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_228 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_495_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_229 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_229 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_496_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_230 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_230 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_497_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_231 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_231 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_498_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_232 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_232 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_499_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_233 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_233 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_500_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_234 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_234 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_501_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_235 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_235 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_502_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_236 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_236 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_503_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_237 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_237 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_504_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_238 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_238 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_505_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_239 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_239 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_506_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_240 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_240 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_507_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_241 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_241 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_508_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_242 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_242 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_509_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_243 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_243 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_510_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_244 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_244 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_511_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_245 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_245 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_512_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_246 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_246 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_513_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_247 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_247 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_514_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_248 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_248 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_515_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_249 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_249 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_516_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_250 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_250 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_517_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_251 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_251 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_518_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_252 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_252 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_519_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_253 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_253 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_520_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_254 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_254 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_521_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_255 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_255 <= {_T_538,_T_535};
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      fghr <= 8'h0;
    end else begin
      fghr <= _T_339 | _T_338;
    end
  end
  always @(posedge rvclkhdr_538_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_0 <= 2'h0;
    end else if (bht_bank_sel_1_0_0) begin
      if (_T_8870) begin
        bht_bank_rd_data_out_1_0 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_0 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_538_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_1 <= 2'h0;
    end else if (bht_bank_sel_1_0_1) begin
      if (_T_8879) begin
        bht_bank_rd_data_out_1_1 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_1 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_538_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_2 <= 2'h0;
    end else if (bht_bank_sel_1_0_2) begin
      if (_T_8888) begin
        bht_bank_rd_data_out_1_2 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_2 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_538_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_3 <= 2'h0;
    end else if (bht_bank_sel_1_0_3) begin
      if (_T_8897) begin
        bht_bank_rd_data_out_1_3 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_3 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_538_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_4 <= 2'h0;
    end else if (bht_bank_sel_1_0_4) begin
      if (_T_8906) begin
        bht_bank_rd_data_out_1_4 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_4 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_538_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_5 <= 2'h0;
    end else if (bht_bank_sel_1_0_5) begin
      if (_T_8915) begin
        bht_bank_rd_data_out_1_5 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_5 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_538_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_6 <= 2'h0;
    end else if (bht_bank_sel_1_0_6) begin
      if (_T_8924) begin
        bht_bank_rd_data_out_1_6 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_6 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_538_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_7 <= 2'h0;
    end else if (bht_bank_sel_1_0_7) begin
      if (_T_8933) begin
        bht_bank_rd_data_out_1_7 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_7 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_538_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_8 <= 2'h0;
    end else if (bht_bank_sel_1_0_8) begin
      if (_T_8942) begin
        bht_bank_rd_data_out_1_8 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_8 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_538_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_9 <= 2'h0;
    end else if (bht_bank_sel_1_0_9) begin
      if (_T_8951) begin
        bht_bank_rd_data_out_1_9 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_9 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_538_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_10 <= 2'h0;
    end else if (bht_bank_sel_1_0_10) begin
      if (_T_8960) begin
        bht_bank_rd_data_out_1_10 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_10 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_538_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_11 <= 2'h0;
    end else if (bht_bank_sel_1_0_11) begin
      if (_T_8969) begin
        bht_bank_rd_data_out_1_11 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_11 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_538_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_12 <= 2'h0;
    end else if (bht_bank_sel_1_0_12) begin
      if (_T_8978) begin
        bht_bank_rd_data_out_1_12 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_12 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_538_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_13 <= 2'h0;
    end else if (bht_bank_sel_1_0_13) begin
      if (_T_8987) begin
        bht_bank_rd_data_out_1_13 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_13 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_538_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_14 <= 2'h0;
    end else if (bht_bank_sel_1_0_14) begin
      if (_T_8996) begin
        bht_bank_rd_data_out_1_14 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_14 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_538_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_15 <= 2'h0;
    end else if (bht_bank_sel_1_0_15) begin
      if (_T_9005) begin
        bht_bank_rd_data_out_1_15 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_15 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_539_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_16 <= 2'h0;
    end else if (bht_bank_sel_1_1_0) begin
      if (_T_9014) begin
        bht_bank_rd_data_out_1_16 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_16 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_539_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_17 <= 2'h0;
    end else if (bht_bank_sel_1_1_1) begin
      if (_T_9023) begin
        bht_bank_rd_data_out_1_17 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_17 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_539_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_18 <= 2'h0;
    end else if (bht_bank_sel_1_1_2) begin
      if (_T_9032) begin
        bht_bank_rd_data_out_1_18 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_18 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_539_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_19 <= 2'h0;
    end else if (bht_bank_sel_1_1_3) begin
      if (_T_9041) begin
        bht_bank_rd_data_out_1_19 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_19 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_539_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_20 <= 2'h0;
    end else if (bht_bank_sel_1_1_4) begin
      if (_T_9050) begin
        bht_bank_rd_data_out_1_20 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_20 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_539_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_21 <= 2'h0;
    end else if (bht_bank_sel_1_1_5) begin
      if (_T_9059) begin
        bht_bank_rd_data_out_1_21 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_21 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_539_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_22 <= 2'h0;
    end else if (bht_bank_sel_1_1_6) begin
      if (_T_9068) begin
        bht_bank_rd_data_out_1_22 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_22 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_539_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_23 <= 2'h0;
    end else if (bht_bank_sel_1_1_7) begin
      if (_T_9077) begin
        bht_bank_rd_data_out_1_23 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_23 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_539_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_24 <= 2'h0;
    end else if (bht_bank_sel_1_1_8) begin
      if (_T_9086) begin
        bht_bank_rd_data_out_1_24 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_24 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_539_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_25 <= 2'h0;
    end else if (bht_bank_sel_1_1_9) begin
      if (_T_9095) begin
        bht_bank_rd_data_out_1_25 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_25 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_539_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_26 <= 2'h0;
    end else if (bht_bank_sel_1_1_10) begin
      if (_T_9104) begin
        bht_bank_rd_data_out_1_26 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_26 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_539_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_27 <= 2'h0;
    end else if (bht_bank_sel_1_1_11) begin
      if (_T_9113) begin
        bht_bank_rd_data_out_1_27 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_27 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_539_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_28 <= 2'h0;
    end else if (bht_bank_sel_1_1_12) begin
      if (_T_9122) begin
        bht_bank_rd_data_out_1_28 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_28 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_539_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_29 <= 2'h0;
    end else if (bht_bank_sel_1_1_13) begin
      if (_T_9131) begin
        bht_bank_rd_data_out_1_29 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_29 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_539_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_30 <= 2'h0;
    end else if (bht_bank_sel_1_1_14) begin
      if (_T_9140) begin
        bht_bank_rd_data_out_1_30 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_30 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_539_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_31 <= 2'h0;
    end else if (bht_bank_sel_1_1_15) begin
      if (_T_9149) begin
        bht_bank_rd_data_out_1_31 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_31 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_540_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_32 <= 2'h0;
    end else if (bht_bank_sel_1_2_0) begin
      if (_T_9158) begin
        bht_bank_rd_data_out_1_32 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_32 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_540_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_33 <= 2'h0;
    end else if (bht_bank_sel_1_2_1) begin
      if (_T_9167) begin
        bht_bank_rd_data_out_1_33 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_33 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_540_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_34 <= 2'h0;
    end else if (bht_bank_sel_1_2_2) begin
      if (_T_9176) begin
        bht_bank_rd_data_out_1_34 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_34 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_540_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_35 <= 2'h0;
    end else if (bht_bank_sel_1_2_3) begin
      if (_T_9185) begin
        bht_bank_rd_data_out_1_35 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_35 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_540_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_36 <= 2'h0;
    end else if (bht_bank_sel_1_2_4) begin
      if (_T_9194) begin
        bht_bank_rd_data_out_1_36 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_36 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_540_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_37 <= 2'h0;
    end else if (bht_bank_sel_1_2_5) begin
      if (_T_9203) begin
        bht_bank_rd_data_out_1_37 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_37 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_540_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_38 <= 2'h0;
    end else if (bht_bank_sel_1_2_6) begin
      if (_T_9212) begin
        bht_bank_rd_data_out_1_38 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_38 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_540_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_39 <= 2'h0;
    end else if (bht_bank_sel_1_2_7) begin
      if (_T_9221) begin
        bht_bank_rd_data_out_1_39 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_39 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_540_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_40 <= 2'h0;
    end else if (bht_bank_sel_1_2_8) begin
      if (_T_9230) begin
        bht_bank_rd_data_out_1_40 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_40 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_540_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_41 <= 2'h0;
    end else if (bht_bank_sel_1_2_9) begin
      if (_T_9239) begin
        bht_bank_rd_data_out_1_41 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_41 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_540_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_42 <= 2'h0;
    end else if (bht_bank_sel_1_2_10) begin
      if (_T_9248) begin
        bht_bank_rd_data_out_1_42 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_42 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_540_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_43 <= 2'h0;
    end else if (bht_bank_sel_1_2_11) begin
      if (_T_9257) begin
        bht_bank_rd_data_out_1_43 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_43 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_540_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_44 <= 2'h0;
    end else if (bht_bank_sel_1_2_12) begin
      if (_T_9266) begin
        bht_bank_rd_data_out_1_44 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_44 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_540_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_45 <= 2'h0;
    end else if (bht_bank_sel_1_2_13) begin
      if (_T_9275) begin
        bht_bank_rd_data_out_1_45 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_45 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_540_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_46 <= 2'h0;
    end else if (bht_bank_sel_1_2_14) begin
      if (_T_9284) begin
        bht_bank_rd_data_out_1_46 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_46 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_540_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_47 <= 2'h0;
    end else if (bht_bank_sel_1_2_15) begin
      if (_T_9293) begin
        bht_bank_rd_data_out_1_47 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_47 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_541_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_48 <= 2'h0;
    end else if (bht_bank_sel_1_3_0) begin
      if (_T_9302) begin
        bht_bank_rd_data_out_1_48 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_48 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_541_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_49 <= 2'h0;
    end else if (bht_bank_sel_1_3_1) begin
      if (_T_9311) begin
        bht_bank_rd_data_out_1_49 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_49 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_541_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_50 <= 2'h0;
    end else if (bht_bank_sel_1_3_2) begin
      if (_T_9320) begin
        bht_bank_rd_data_out_1_50 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_50 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_541_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_51 <= 2'h0;
    end else if (bht_bank_sel_1_3_3) begin
      if (_T_9329) begin
        bht_bank_rd_data_out_1_51 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_51 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_541_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_52 <= 2'h0;
    end else if (bht_bank_sel_1_3_4) begin
      if (_T_9338) begin
        bht_bank_rd_data_out_1_52 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_52 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_541_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_53 <= 2'h0;
    end else if (bht_bank_sel_1_3_5) begin
      if (_T_9347) begin
        bht_bank_rd_data_out_1_53 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_53 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_541_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_54 <= 2'h0;
    end else if (bht_bank_sel_1_3_6) begin
      if (_T_9356) begin
        bht_bank_rd_data_out_1_54 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_54 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_541_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_55 <= 2'h0;
    end else if (bht_bank_sel_1_3_7) begin
      if (_T_9365) begin
        bht_bank_rd_data_out_1_55 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_55 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_541_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_56 <= 2'h0;
    end else if (bht_bank_sel_1_3_8) begin
      if (_T_9374) begin
        bht_bank_rd_data_out_1_56 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_56 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_541_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_57 <= 2'h0;
    end else if (bht_bank_sel_1_3_9) begin
      if (_T_9383) begin
        bht_bank_rd_data_out_1_57 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_57 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_541_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_58 <= 2'h0;
    end else if (bht_bank_sel_1_3_10) begin
      if (_T_9392) begin
        bht_bank_rd_data_out_1_58 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_58 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_541_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_59 <= 2'h0;
    end else if (bht_bank_sel_1_3_11) begin
      if (_T_9401) begin
        bht_bank_rd_data_out_1_59 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_59 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_541_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_60 <= 2'h0;
    end else if (bht_bank_sel_1_3_12) begin
      if (_T_9410) begin
        bht_bank_rd_data_out_1_60 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_60 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_541_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_61 <= 2'h0;
    end else if (bht_bank_sel_1_3_13) begin
      if (_T_9419) begin
        bht_bank_rd_data_out_1_61 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_61 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_541_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_62 <= 2'h0;
    end else if (bht_bank_sel_1_3_14) begin
      if (_T_9428) begin
        bht_bank_rd_data_out_1_62 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_62 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_541_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_63 <= 2'h0;
    end else if (bht_bank_sel_1_3_15) begin
      if (_T_9437) begin
        bht_bank_rd_data_out_1_63 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_63 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_542_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_64 <= 2'h0;
    end else if (bht_bank_sel_1_4_0) begin
      if (_T_9446) begin
        bht_bank_rd_data_out_1_64 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_64 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_542_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_65 <= 2'h0;
    end else if (bht_bank_sel_1_4_1) begin
      if (_T_9455) begin
        bht_bank_rd_data_out_1_65 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_65 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_542_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_66 <= 2'h0;
    end else if (bht_bank_sel_1_4_2) begin
      if (_T_9464) begin
        bht_bank_rd_data_out_1_66 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_66 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_542_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_67 <= 2'h0;
    end else if (bht_bank_sel_1_4_3) begin
      if (_T_9473) begin
        bht_bank_rd_data_out_1_67 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_67 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_542_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_68 <= 2'h0;
    end else if (bht_bank_sel_1_4_4) begin
      if (_T_9482) begin
        bht_bank_rd_data_out_1_68 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_68 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_542_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_69 <= 2'h0;
    end else if (bht_bank_sel_1_4_5) begin
      if (_T_9491) begin
        bht_bank_rd_data_out_1_69 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_69 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_542_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_70 <= 2'h0;
    end else if (bht_bank_sel_1_4_6) begin
      if (_T_9500) begin
        bht_bank_rd_data_out_1_70 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_70 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_542_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_71 <= 2'h0;
    end else if (bht_bank_sel_1_4_7) begin
      if (_T_9509) begin
        bht_bank_rd_data_out_1_71 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_71 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_542_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_72 <= 2'h0;
    end else if (bht_bank_sel_1_4_8) begin
      if (_T_9518) begin
        bht_bank_rd_data_out_1_72 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_72 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_542_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_73 <= 2'h0;
    end else if (bht_bank_sel_1_4_9) begin
      if (_T_9527) begin
        bht_bank_rd_data_out_1_73 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_73 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_542_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_74 <= 2'h0;
    end else if (bht_bank_sel_1_4_10) begin
      if (_T_9536) begin
        bht_bank_rd_data_out_1_74 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_74 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_542_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_75 <= 2'h0;
    end else if (bht_bank_sel_1_4_11) begin
      if (_T_9545) begin
        bht_bank_rd_data_out_1_75 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_75 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_542_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_76 <= 2'h0;
    end else if (bht_bank_sel_1_4_12) begin
      if (_T_9554) begin
        bht_bank_rd_data_out_1_76 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_76 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_542_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_77 <= 2'h0;
    end else if (bht_bank_sel_1_4_13) begin
      if (_T_9563) begin
        bht_bank_rd_data_out_1_77 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_77 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_542_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_78 <= 2'h0;
    end else if (bht_bank_sel_1_4_14) begin
      if (_T_9572) begin
        bht_bank_rd_data_out_1_78 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_78 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_542_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_79 <= 2'h0;
    end else if (bht_bank_sel_1_4_15) begin
      if (_T_9581) begin
        bht_bank_rd_data_out_1_79 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_79 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_543_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_80 <= 2'h0;
    end else if (bht_bank_sel_1_5_0) begin
      if (_T_9590) begin
        bht_bank_rd_data_out_1_80 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_80 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_543_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_81 <= 2'h0;
    end else if (bht_bank_sel_1_5_1) begin
      if (_T_9599) begin
        bht_bank_rd_data_out_1_81 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_81 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_543_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_82 <= 2'h0;
    end else if (bht_bank_sel_1_5_2) begin
      if (_T_9608) begin
        bht_bank_rd_data_out_1_82 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_82 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_543_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_83 <= 2'h0;
    end else if (bht_bank_sel_1_5_3) begin
      if (_T_9617) begin
        bht_bank_rd_data_out_1_83 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_83 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_543_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_84 <= 2'h0;
    end else if (bht_bank_sel_1_5_4) begin
      if (_T_9626) begin
        bht_bank_rd_data_out_1_84 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_84 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_543_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_85 <= 2'h0;
    end else if (bht_bank_sel_1_5_5) begin
      if (_T_9635) begin
        bht_bank_rd_data_out_1_85 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_85 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_543_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_86 <= 2'h0;
    end else if (bht_bank_sel_1_5_6) begin
      if (_T_9644) begin
        bht_bank_rd_data_out_1_86 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_86 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_543_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_87 <= 2'h0;
    end else if (bht_bank_sel_1_5_7) begin
      if (_T_9653) begin
        bht_bank_rd_data_out_1_87 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_87 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_543_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_88 <= 2'h0;
    end else if (bht_bank_sel_1_5_8) begin
      if (_T_9662) begin
        bht_bank_rd_data_out_1_88 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_88 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_543_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_89 <= 2'h0;
    end else if (bht_bank_sel_1_5_9) begin
      if (_T_9671) begin
        bht_bank_rd_data_out_1_89 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_89 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_543_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_90 <= 2'h0;
    end else if (bht_bank_sel_1_5_10) begin
      if (_T_9680) begin
        bht_bank_rd_data_out_1_90 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_90 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_543_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_91 <= 2'h0;
    end else if (bht_bank_sel_1_5_11) begin
      if (_T_9689) begin
        bht_bank_rd_data_out_1_91 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_91 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_543_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_92 <= 2'h0;
    end else if (bht_bank_sel_1_5_12) begin
      if (_T_9698) begin
        bht_bank_rd_data_out_1_92 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_92 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_543_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_93 <= 2'h0;
    end else if (bht_bank_sel_1_5_13) begin
      if (_T_9707) begin
        bht_bank_rd_data_out_1_93 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_93 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_543_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_94 <= 2'h0;
    end else if (bht_bank_sel_1_5_14) begin
      if (_T_9716) begin
        bht_bank_rd_data_out_1_94 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_94 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_543_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_95 <= 2'h0;
    end else if (bht_bank_sel_1_5_15) begin
      if (_T_9725) begin
        bht_bank_rd_data_out_1_95 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_95 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_544_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_96 <= 2'h0;
    end else if (bht_bank_sel_1_6_0) begin
      if (_T_9734) begin
        bht_bank_rd_data_out_1_96 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_96 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_544_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_97 <= 2'h0;
    end else if (bht_bank_sel_1_6_1) begin
      if (_T_9743) begin
        bht_bank_rd_data_out_1_97 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_97 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_544_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_98 <= 2'h0;
    end else if (bht_bank_sel_1_6_2) begin
      if (_T_9752) begin
        bht_bank_rd_data_out_1_98 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_98 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_544_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_99 <= 2'h0;
    end else if (bht_bank_sel_1_6_3) begin
      if (_T_9761) begin
        bht_bank_rd_data_out_1_99 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_99 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_544_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_100 <= 2'h0;
    end else if (bht_bank_sel_1_6_4) begin
      if (_T_9770) begin
        bht_bank_rd_data_out_1_100 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_100 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_544_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_101 <= 2'h0;
    end else if (bht_bank_sel_1_6_5) begin
      if (_T_9779) begin
        bht_bank_rd_data_out_1_101 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_101 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_544_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_102 <= 2'h0;
    end else if (bht_bank_sel_1_6_6) begin
      if (_T_9788) begin
        bht_bank_rd_data_out_1_102 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_102 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_544_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_103 <= 2'h0;
    end else if (bht_bank_sel_1_6_7) begin
      if (_T_9797) begin
        bht_bank_rd_data_out_1_103 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_103 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_544_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_104 <= 2'h0;
    end else if (bht_bank_sel_1_6_8) begin
      if (_T_9806) begin
        bht_bank_rd_data_out_1_104 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_104 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_544_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_105 <= 2'h0;
    end else if (bht_bank_sel_1_6_9) begin
      if (_T_9815) begin
        bht_bank_rd_data_out_1_105 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_105 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_544_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_106 <= 2'h0;
    end else if (bht_bank_sel_1_6_10) begin
      if (_T_9824) begin
        bht_bank_rd_data_out_1_106 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_106 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_544_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_107 <= 2'h0;
    end else if (bht_bank_sel_1_6_11) begin
      if (_T_9833) begin
        bht_bank_rd_data_out_1_107 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_107 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_544_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_108 <= 2'h0;
    end else if (bht_bank_sel_1_6_12) begin
      if (_T_9842) begin
        bht_bank_rd_data_out_1_108 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_108 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_544_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_109 <= 2'h0;
    end else if (bht_bank_sel_1_6_13) begin
      if (_T_9851) begin
        bht_bank_rd_data_out_1_109 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_109 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_544_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_110 <= 2'h0;
    end else if (bht_bank_sel_1_6_14) begin
      if (_T_9860) begin
        bht_bank_rd_data_out_1_110 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_110 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_544_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_111 <= 2'h0;
    end else if (bht_bank_sel_1_6_15) begin
      if (_T_9869) begin
        bht_bank_rd_data_out_1_111 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_111 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_545_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_112 <= 2'h0;
    end else if (bht_bank_sel_1_7_0) begin
      if (_T_9878) begin
        bht_bank_rd_data_out_1_112 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_112 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_545_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_113 <= 2'h0;
    end else if (bht_bank_sel_1_7_1) begin
      if (_T_9887) begin
        bht_bank_rd_data_out_1_113 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_113 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_545_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_114 <= 2'h0;
    end else if (bht_bank_sel_1_7_2) begin
      if (_T_9896) begin
        bht_bank_rd_data_out_1_114 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_114 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_545_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_115 <= 2'h0;
    end else if (bht_bank_sel_1_7_3) begin
      if (_T_9905) begin
        bht_bank_rd_data_out_1_115 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_115 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_545_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_116 <= 2'h0;
    end else if (bht_bank_sel_1_7_4) begin
      if (_T_9914) begin
        bht_bank_rd_data_out_1_116 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_116 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_545_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_117 <= 2'h0;
    end else if (bht_bank_sel_1_7_5) begin
      if (_T_9923) begin
        bht_bank_rd_data_out_1_117 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_117 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_545_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_118 <= 2'h0;
    end else if (bht_bank_sel_1_7_6) begin
      if (_T_9932) begin
        bht_bank_rd_data_out_1_118 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_118 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_545_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_119 <= 2'h0;
    end else if (bht_bank_sel_1_7_7) begin
      if (_T_9941) begin
        bht_bank_rd_data_out_1_119 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_119 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_545_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_120 <= 2'h0;
    end else if (bht_bank_sel_1_7_8) begin
      if (_T_9950) begin
        bht_bank_rd_data_out_1_120 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_120 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_545_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_121 <= 2'h0;
    end else if (bht_bank_sel_1_7_9) begin
      if (_T_9959) begin
        bht_bank_rd_data_out_1_121 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_121 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_545_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_122 <= 2'h0;
    end else if (bht_bank_sel_1_7_10) begin
      if (_T_9968) begin
        bht_bank_rd_data_out_1_122 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_122 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_545_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_123 <= 2'h0;
    end else if (bht_bank_sel_1_7_11) begin
      if (_T_9977) begin
        bht_bank_rd_data_out_1_123 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_123 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_545_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_124 <= 2'h0;
    end else if (bht_bank_sel_1_7_12) begin
      if (_T_9986) begin
        bht_bank_rd_data_out_1_124 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_124 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_545_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_125 <= 2'h0;
    end else if (bht_bank_sel_1_7_13) begin
      if (_T_9995) begin
        bht_bank_rd_data_out_1_125 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_125 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_545_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_126 <= 2'h0;
    end else if (bht_bank_sel_1_7_14) begin
      if (_T_10004) begin
        bht_bank_rd_data_out_1_126 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_126 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_545_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_127 <= 2'h0;
    end else if (bht_bank_sel_1_7_15) begin
      if (_T_10013) begin
        bht_bank_rd_data_out_1_127 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_127 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_546_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_128 <= 2'h0;
    end else if (bht_bank_sel_1_8_0) begin
      if (_T_10022) begin
        bht_bank_rd_data_out_1_128 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_128 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_546_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_129 <= 2'h0;
    end else if (bht_bank_sel_1_8_1) begin
      if (_T_10031) begin
        bht_bank_rd_data_out_1_129 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_129 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_546_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_130 <= 2'h0;
    end else if (bht_bank_sel_1_8_2) begin
      if (_T_10040) begin
        bht_bank_rd_data_out_1_130 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_130 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_546_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_131 <= 2'h0;
    end else if (bht_bank_sel_1_8_3) begin
      if (_T_10049) begin
        bht_bank_rd_data_out_1_131 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_131 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_546_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_132 <= 2'h0;
    end else if (bht_bank_sel_1_8_4) begin
      if (_T_10058) begin
        bht_bank_rd_data_out_1_132 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_132 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_546_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_133 <= 2'h0;
    end else if (bht_bank_sel_1_8_5) begin
      if (_T_10067) begin
        bht_bank_rd_data_out_1_133 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_133 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_546_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_134 <= 2'h0;
    end else if (bht_bank_sel_1_8_6) begin
      if (_T_10076) begin
        bht_bank_rd_data_out_1_134 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_134 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_546_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_135 <= 2'h0;
    end else if (bht_bank_sel_1_8_7) begin
      if (_T_10085) begin
        bht_bank_rd_data_out_1_135 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_135 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_546_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_136 <= 2'h0;
    end else if (bht_bank_sel_1_8_8) begin
      if (_T_10094) begin
        bht_bank_rd_data_out_1_136 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_136 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_546_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_137 <= 2'h0;
    end else if (bht_bank_sel_1_8_9) begin
      if (_T_10103) begin
        bht_bank_rd_data_out_1_137 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_137 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_546_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_138 <= 2'h0;
    end else if (bht_bank_sel_1_8_10) begin
      if (_T_10112) begin
        bht_bank_rd_data_out_1_138 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_138 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_546_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_139 <= 2'h0;
    end else if (bht_bank_sel_1_8_11) begin
      if (_T_10121) begin
        bht_bank_rd_data_out_1_139 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_139 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_546_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_140 <= 2'h0;
    end else if (bht_bank_sel_1_8_12) begin
      if (_T_10130) begin
        bht_bank_rd_data_out_1_140 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_140 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_546_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_141 <= 2'h0;
    end else if (bht_bank_sel_1_8_13) begin
      if (_T_10139) begin
        bht_bank_rd_data_out_1_141 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_141 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_546_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_142 <= 2'h0;
    end else if (bht_bank_sel_1_8_14) begin
      if (_T_10148) begin
        bht_bank_rd_data_out_1_142 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_142 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_546_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_143 <= 2'h0;
    end else if (bht_bank_sel_1_8_15) begin
      if (_T_10157) begin
        bht_bank_rd_data_out_1_143 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_143 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_547_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_144 <= 2'h0;
    end else if (bht_bank_sel_1_9_0) begin
      if (_T_10166) begin
        bht_bank_rd_data_out_1_144 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_144 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_547_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_145 <= 2'h0;
    end else if (bht_bank_sel_1_9_1) begin
      if (_T_10175) begin
        bht_bank_rd_data_out_1_145 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_145 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_547_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_146 <= 2'h0;
    end else if (bht_bank_sel_1_9_2) begin
      if (_T_10184) begin
        bht_bank_rd_data_out_1_146 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_146 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_547_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_147 <= 2'h0;
    end else if (bht_bank_sel_1_9_3) begin
      if (_T_10193) begin
        bht_bank_rd_data_out_1_147 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_147 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_547_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_148 <= 2'h0;
    end else if (bht_bank_sel_1_9_4) begin
      if (_T_10202) begin
        bht_bank_rd_data_out_1_148 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_148 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_547_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_149 <= 2'h0;
    end else if (bht_bank_sel_1_9_5) begin
      if (_T_10211) begin
        bht_bank_rd_data_out_1_149 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_149 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_547_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_150 <= 2'h0;
    end else if (bht_bank_sel_1_9_6) begin
      if (_T_10220) begin
        bht_bank_rd_data_out_1_150 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_150 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_547_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_151 <= 2'h0;
    end else if (bht_bank_sel_1_9_7) begin
      if (_T_10229) begin
        bht_bank_rd_data_out_1_151 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_151 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_547_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_152 <= 2'h0;
    end else if (bht_bank_sel_1_9_8) begin
      if (_T_10238) begin
        bht_bank_rd_data_out_1_152 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_152 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_547_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_153 <= 2'h0;
    end else if (bht_bank_sel_1_9_9) begin
      if (_T_10247) begin
        bht_bank_rd_data_out_1_153 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_153 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_547_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_154 <= 2'h0;
    end else if (bht_bank_sel_1_9_10) begin
      if (_T_10256) begin
        bht_bank_rd_data_out_1_154 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_154 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_547_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_155 <= 2'h0;
    end else if (bht_bank_sel_1_9_11) begin
      if (_T_10265) begin
        bht_bank_rd_data_out_1_155 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_155 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_547_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_156 <= 2'h0;
    end else if (bht_bank_sel_1_9_12) begin
      if (_T_10274) begin
        bht_bank_rd_data_out_1_156 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_156 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_547_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_157 <= 2'h0;
    end else if (bht_bank_sel_1_9_13) begin
      if (_T_10283) begin
        bht_bank_rd_data_out_1_157 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_157 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_547_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_158 <= 2'h0;
    end else if (bht_bank_sel_1_9_14) begin
      if (_T_10292) begin
        bht_bank_rd_data_out_1_158 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_158 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_547_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_159 <= 2'h0;
    end else if (bht_bank_sel_1_9_15) begin
      if (_T_10301) begin
        bht_bank_rd_data_out_1_159 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_159 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_548_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_160 <= 2'h0;
    end else if (bht_bank_sel_1_10_0) begin
      if (_T_10310) begin
        bht_bank_rd_data_out_1_160 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_160 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_548_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_161 <= 2'h0;
    end else if (bht_bank_sel_1_10_1) begin
      if (_T_10319) begin
        bht_bank_rd_data_out_1_161 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_161 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_548_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_162 <= 2'h0;
    end else if (bht_bank_sel_1_10_2) begin
      if (_T_10328) begin
        bht_bank_rd_data_out_1_162 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_162 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_548_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_163 <= 2'h0;
    end else if (bht_bank_sel_1_10_3) begin
      if (_T_10337) begin
        bht_bank_rd_data_out_1_163 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_163 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_548_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_164 <= 2'h0;
    end else if (bht_bank_sel_1_10_4) begin
      if (_T_10346) begin
        bht_bank_rd_data_out_1_164 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_164 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_548_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_165 <= 2'h0;
    end else if (bht_bank_sel_1_10_5) begin
      if (_T_10355) begin
        bht_bank_rd_data_out_1_165 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_165 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_548_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_166 <= 2'h0;
    end else if (bht_bank_sel_1_10_6) begin
      if (_T_10364) begin
        bht_bank_rd_data_out_1_166 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_166 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_548_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_167 <= 2'h0;
    end else if (bht_bank_sel_1_10_7) begin
      if (_T_10373) begin
        bht_bank_rd_data_out_1_167 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_167 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_548_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_168 <= 2'h0;
    end else if (bht_bank_sel_1_10_8) begin
      if (_T_10382) begin
        bht_bank_rd_data_out_1_168 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_168 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_548_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_169 <= 2'h0;
    end else if (bht_bank_sel_1_10_9) begin
      if (_T_10391) begin
        bht_bank_rd_data_out_1_169 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_169 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_548_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_170 <= 2'h0;
    end else if (bht_bank_sel_1_10_10) begin
      if (_T_10400) begin
        bht_bank_rd_data_out_1_170 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_170 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_548_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_171 <= 2'h0;
    end else if (bht_bank_sel_1_10_11) begin
      if (_T_10409) begin
        bht_bank_rd_data_out_1_171 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_171 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_548_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_172 <= 2'h0;
    end else if (bht_bank_sel_1_10_12) begin
      if (_T_10418) begin
        bht_bank_rd_data_out_1_172 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_172 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_548_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_173 <= 2'h0;
    end else if (bht_bank_sel_1_10_13) begin
      if (_T_10427) begin
        bht_bank_rd_data_out_1_173 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_173 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_548_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_174 <= 2'h0;
    end else if (bht_bank_sel_1_10_14) begin
      if (_T_10436) begin
        bht_bank_rd_data_out_1_174 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_174 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_548_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_175 <= 2'h0;
    end else if (bht_bank_sel_1_10_15) begin
      if (_T_10445) begin
        bht_bank_rd_data_out_1_175 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_175 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_549_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_176 <= 2'h0;
    end else if (bht_bank_sel_1_11_0) begin
      if (_T_10454) begin
        bht_bank_rd_data_out_1_176 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_176 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_549_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_177 <= 2'h0;
    end else if (bht_bank_sel_1_11_1) begin
      if (_T_10463) begin
        bht_bank_rd_data_out_1_177 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_177 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_549_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_178 <= 2'h0;
    end else if (bht_bank_sel_1_11_2) begin
      if (_T_10472) begin
        bht_bank_rd_data_out_1_178 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_178 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_549_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_179 <= 2'h0;
    end else if (bht_bank_sel_1_11_3) begin
      if (_T_10481) begin
        bht_bank_rd_data_out_1_179 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_179 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_549_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_180 <= 2'h0;
    end else if (bht_bank_sel_1_11_4) begin
      if (_T_10490) begin
        bht_bank_rd_data_out_1_180 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_180 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_549_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_181 <= 2'h0;
    end else if (bht_bank_sel_1_11_5) begin
      if (_T_10499) begin
        bht_bank_rd_data_out_1_181 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_181 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_549_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_182 <= 2'h0;
    end else if (bht_bank_sel_1_11_6) begin
      if (_T_10508) begin
        bht_bank_rd_data_out_1_182 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_182 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_549_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_183 <= 2'h0;
    end else if (bht_bank_sel_1_11_7) begin
      if (_T_10517) begin
        bht_bank_rd_data_out_1_183 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_183 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_549_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_184 <= 2'h0;
    end else if (bht_bank_sel_1_11_8) begin
      if (_T_10526) begin
        bht_bank_rd_data_out_1_184 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_184 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_549_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_185 <= 2'h0;
    end else if (bht_bank_sel_1_11_9) begin
      if (_T_10535) begin
        bht_bank_rd_data_out_1_185 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_185 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_549_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_186 <= 2'h0;
    end else if (bht_bank_sel_1_11_10) begin
      if (_T_10544) begin
        bht_bank_rd_data_out_1_186 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_186 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_549_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_187 <= 2'h0;
    end else if (bht_bank_sel_1_11_11) begin
      if (_T_10553) begin
        bht_bank_rd_data_out_1_187 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_187 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_549_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_188 <= 2'h0;
    end else if (bht_bank_sel_1_11_12) begin
      if (_T_10562) begin
        bht_bank_rd_data_out_1_188 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_188 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_549_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_189 <= 2'h0;
    end else if (bht_bank_sel_1_11_13) begin
      if (_T_10571) begin
        bht_bank_rd_data_out_1_189 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_189 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_549_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_190 <= 2'h0;
    end else if (bht_bank_sel_1_11_14) begin
      if (_T_10580) begin
        bht_bank_rd_data_out_1_190 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_190 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_549_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_191 <= 2'h0;
    end else if (bht_bank_sel_1_11_15) begin
      if (_T_10589) begin
        bht_bank_rd_data_out_1_191 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_191 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_550_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_192 <= 2'h0;
    end else if (bht_bank_sel_1_12_0) begin
      if (_T_10598) begin
        bht_bank_rd_data_out_1_192 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_192 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_550_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_193 <= 2'h0;
    end else if (bht_bank_sel_1_12_1) begin
      if (_T_10607) begin
        bht_bank_rd_data_out_1_193 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_193 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_550_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_194 <= 2'h0;
    end else if (bht_bank_sel_1_12_2) begin
      if (_T_10616) begin
        bht_bank_rd_data_out_1_194 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_194 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_550_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_195 <= 2'h0;
    end else if (bht_bank_sel_1_12_3) begin
      if (_T_10625) begin
        bht_bank_rd_data_out_1_195 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_195 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_550_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_196 <= 2'h0;
    end else if (bht_bank_sel_1_12_4) begin
      if (_T_10634) begin
        bht_bank_rd_data_out_1_196 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_196 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_550_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_197 <= 2'h0;
    end else if (bht_bank_sel_1_12_5) begin
      if (_T_10643) begin
        bht_bank_rd_data_out_1_197 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_197 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_550_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_198 <= 2'h0;
    end else if (bht_bank_sel_1_12_6) begin
      if (_T_10652) begin
        bht_bank_rd_data_out_1_198 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_198 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_550_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_199 <= 2'h0;
    end else if (bht_bank_sel_1_12_7) begin
      if (_T_10661) begin
        bht_bank_rd_data_out_1_199 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_199 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_550_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_200 <= 2'h0;
    end else if (bht_bank_sel_1_12_8) begin
      if (_T_10670) begin
        bht_bank_rd_data_out_1_200 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_200 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_550_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_201 <= 2'h0;
    end else if (bht_bank_sel_1_12_9) begin
      if (_T_10679) begin
        bht_bank_rd_data_out_1_201 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_201 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_550_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_202 <= 2'h0;
    end else if (bht_bank_sel_1_12_10) begin
      if (_T_10688) begin
        bht_bank_rd_data_out_1_202 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_202 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_550_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_203 <= 2'h0;
    end else if (bht_bank_sel_1_12_11) begin
      if (_T_10697) begin
        bht_bank_rd_data_out_1_203 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_203 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_550_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_204 <= 2'h0;
    end else if (bht_bank_sel_1_12_12) begin
      if (_T_10706) begin
        bht_bank_rd_data_out_1_204 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_204 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_550_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_205 <= 2'h0;
    end else if (bht_bank_sel_1_12_13) begin
      if (_T_10715) begin
        bht_bank_rd_data_out_1_205 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_205 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_550_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_206 <= 2'h0;
    end else if (bht_bank_sel_1_12_14) begin
      if (_T_10724) begin
        bht_bank_rd_data_out_1_206 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_206 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_550_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_207 <= 2'h0;
    end else if (bht_bank_sel_1_12_15) begin
      if (_T_10733) begin
        bht_bank_rd_data_out_1_207 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_207 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_551_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_208 <= 2'h0;
    end else if (bht_bank_sel_1_13_0) begin
      if (_T_10742) begin
        bht_bank_rd_data_out_1_208 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_208 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_551_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_209 <= 2'h0;
    end else if (bht_bank_sel_1_13_1) begin
      if (_T_10751) begin
        bht_bank_rd_data_out_1_209 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_209 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_551_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_210 <= 2'h0;
    end else if (bht_bank_sel_1_13_2) begin
      if (_T_10760) begin
        bht_bank_rd_data_out_1_210 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_210 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_551_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_211 <= 2'h0;
    end else if (bht_bank_sel_1_13_3) begin
      if (_T_10769) begin
        bht_bank_rd_data_out_1_211 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_211 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_551_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_212 <= 2'h0;
    end else if (bht_bank_sel_1_13_4) begin
      if (_T_10778) begin
        bht_bank_rd_data_out_1_212 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_212 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_551_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_213 <= 2'h0;
    end else if (bht_bank_sel_1_13_5) begin
      if (_T_10787) begin
        bht_bank_rd_data_out_1_213 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_213 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_551_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_214 <= 2'h0;
    end else if (bht_bank_sel_1_13_6) begin
      if (_T_10796) begin
        bht_bank_rd_data_out_1_214 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_214 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_551_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_215 <= 2'h0;
    end else if (bht_bank_sel_1_13_7) begin
      if (_T_10805) begin
        bht_bank_rd_data_out_1_215 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_215 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_551_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_216 <= 2'h0;
    end else if (bht_bank_sel_1_13_8) begin
      if (_T_10814) begin
        bht_bank_rd_data_out_1_216 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_216 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_551_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_217 <= 2'h0;
    end else if (bht_bank_sel_1_13_9) begin
      if (_T_10823) begin
        bht_bank_rd_data_out_1_217 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_217 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_551_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_218 <= 2'h0;
    end else if (bht_bank_sel_1_13_10) begin
      if (_T_10832) begin
        bht_bank_rd_data_out_1_218 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_218 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_551_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_219 <= 2'h0;
    end else if (bht_bank_sel_1_13_11) begin
      if (_T_10841) begin
        bht_bank_rd_data_out_1_219 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_219 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_551_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_220 <= 2'h0;
    end else if (bht_bank_sel_1_13_12) begin
      if (_T_10850) begin
        bht_bank_rd_data_out_1_220 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_220 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_551_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_221 <= 2'h0;
    end else if (bht_bank_sel_1_13_13) begin
      if (_T_10859) begin
        bht_bank_rd_data_out_1_221 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_221 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_551_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_222 <= 2'h0;
    end else if (bht_bank_sel_1_13_14) begin
      if (_T_10868) begin
        bht_bank_rd_data_out_1_222 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_222 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_551_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_223 <= 2'h0;
    end else if (bht_bank_sel_1_13_15) begin
      if (_T_10877) begin
        bht_bank_rd_data_out_1_223 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_223 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_552_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_224 <= 2'h0;
    end else if (bht_bank_sel_1_14_0) begin
      if (_T_10886) begin
        bht_bank_rd_data_out_1_224 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_224 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_552_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_225 <= 2'h0;
    end else if (bht_bank_sel_1_14_1) begin
      if (_T_10895) begin
        bht_bank_rd_data_out_1_225 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_225 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_552_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_226 <= 2'h0;
    end else if (bht_bank_sel_1_14_2) begin
      if (_T_10904) begin
        bht_bank_rd_data_out_1_226 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_226 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_552_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_227 <= 2'h0;
    end else if (bht_bank_sel_1_14_3) begin
      if (_T_10913) begin
        bht_bank_rd_data_out_1_227 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_227 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_552_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_228 <= 2'h0;
    end else if (bht_bank_sel_1_14_4) begin
      if (_T_10922) begin
        bht_bank_rd_data_out_1_228 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_228 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_552_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_229 <= 2'h0;
    end else if (bht_bank_sel_1_14_5) begin
      if (_T_10931) begin
        bht_bank_rd_data_out_1_229 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_229 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_552_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_230 <= 2'h0;
    end else if (bht_bank_sel_1_14_6) begin
      if (_T_10940) begin
        bht_bank_rd_data_out_1_230 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_230 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_552_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_231 <= 2'h0;
    end else if (bht_bank_sel_1_14_7) begin
      if (_T_10949) begin
        bht_bank_rd_data_out_1_231 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_231 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_552_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_232 <= 2'h0;
    end else if (bht_bank_sel_1_14_8) begin
      if (_T_10958) begin
        bht_bank_rd_data_out_1_232 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_232 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_552_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_233 <= 2'h0;
    end else if (bht_bank_sel_1_14_9) begin
      if (_T_10967) begin
        bht_bank_rd_data_out_1_233 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_233 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_552_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_234 <= 2'h0;
    end else if (bht_bank_sel_1_14_10) begin
      if (_T_10976) begin
        bht_bank_rd_data_out_1_234 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_234 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_552_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_235 <= 2'h0;
    end else if (bht_bank_sel_1_14_11) begin
      if (_T_10985) begin
        bht_bank_rd_data_out_1_235 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_235 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_552_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_236 <= 2'h0;
    end else if (bht_bank_sel_1_14_12) begin
      if (_T_10994) begin
        bht_bank_rd_data_out_1_236 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_236 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_552_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_237 <= 2'h0;
    end else if (bht_bank_sel_1_14_13) begin
      if (_T_11003) begin
        bht_bank_rd_data_out_1_237 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_237 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_552_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_238 <= 2'h0;
    end else if (bht_bank_sel_1_14_14) begin
      if (_T_11012) begin
        bht_bank_rd_data_out_1_238 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_238 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_552_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_239 <= 2'h0;
    end else if (bht_bank_sel_1_14_15) begin
      if (_T_11021) begin
        bht_bank_rd_data_out_1_239 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_239 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_553_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_240 <= 2'h0;
    end else if (bht_bank_sel_1_15_0) begin
      if (_T_11030) begin
        bht_bank_rd_data_out_1_240 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_240 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_553_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_241 <= 2'h0;
    end else if (bht_bank_sel_1_15_1) begin
      if (_T_11039) begin
        bht_bank_rd_data_out_1_241 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_241 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_553_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_242 <= 2'h0;
    end else if (bht_bank_sel_1_15_2) begin
      if (_T_11048) begin
        bht_bank_rd_data_out_1_242 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_242 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_553_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_243 <= 2'h0;
    end else if (bht_bank_sel_1_15_3) begin
      if (_T_11057) begin
        bht_bank_rd_data_out_1_243 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_243 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_553_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_244 <= 2'h0;
    end else if (bht_bank_sel_1_15_4) begin
      if (_T_11066) begin
        bht_bank_rd_data_out_1_244 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_244 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_553_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_245 <= 2'h0;
    end else if (bht_bank_sel_1_15_5) begin
      if (_T_11075) begin
        bht_bank_rd_data_out_1_245 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_245 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_553_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_246 <= 2'h0;
    end else if (bht_bank_sel_1_15_6) begin
      if (_T_11084) begin
        bht_bank_rd_data_out_1_246 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_246 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_553_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_247 <= 2'h0;
    end else if (bht_bank_sel_1_15_7) begin
      if (_T_11093) begin
        bht_bank_rd_data_out_1_247 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_247 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_553_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_248 <= 2'h0;
    end else if (bht_bank_sel_1_15_8) begin
      if (_T_11102) begin
        bht_bank_rd_data_out_1_248 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_248 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_553_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_249 <= 2'h0;
    end else if (bht_bank_sel_1_15_9) begin
      if (_T_11111) begin
        bht_bank_rd_data_out_1_249 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_249 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_553_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_250 <= 2'h0;
    end else if (bht_bank_sel_1_15_10) begin
      if (_T_11120) begin
        bht_bank_rd_data_out_1_250 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_250 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_553_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_251 <= 2'h0;
    end else if (bht_bank_sel_1_15_11) begin
      if (_T_11129) begin
        bht_bank_rd_data_out_1_251 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_251 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_553_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_252 <= 2'h0;
    end else if (bht_bank_sel_1_15_12) begin
      if (_T_11138) begin
        bht_bank_rd_data_out_1_252 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_252 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_553_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_253 <= 2'h0;
    end else if (bht_bank_sel_1_15_13) begin
      if (_T_11147) begin
        bht_bank_rd_data_out_1_253 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_253 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_553_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_254 <= 2'h0;
    end else if (bht_bank_sel_1_15_14) begin
      if (_T_11156) begin
        bht_bank_rd_data_out_1_254 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_254 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_553_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_255 <= 2'h0;
    end else if (bht_bank_sel_1_15_15) begin
      if (_T_11165) begin
        bht_bank_rd_data_out_1_255 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_255 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_522_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_0 <= 2'h0;
    end else if (bht_bank_sel_0_0_0) begin
      if (_T_6566) begin
        bht_bank_rd_data_out_0_0 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_0 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_522_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_1 <= 2'h0;
    end else if (bht_bank_sel_0_0_1) begin
      if (_T_6575) begin
        bht_bank_rd_data_out_0_1 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_1 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_522_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_2 <= 2'h0;
    end else if (bht_bank_sel_0_0_2) begin
      if (_T_6584) begin
        bht_bank_rd_data_out_0_2 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_2 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_522_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_3 <= 2'h0;
    end else if (bht_bank_sel_0_0_3) begin
      if (_T_6593) begin
        bht_bank_rd_data_out_0_3 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_3 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_522_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_4 <= 2'h0;
    end else if (bht_bank_sel_0_0_4) begin
      if (_T_6602) begin
        bht_bank_rd_data_out_0_4 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_4 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_522_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_5 <= 2'h0;
    end else if (bht_bank_sel_0_0_5) begin
      if (_T_6611) begin
        bht_bank_rd_data_out_0_5 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_5 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_522_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_6 <= 2'h0;
    end else if (bht_bank_sel_0_0_6) begin
      if (_T_6620) begin
        bht_bank_rd_data_out_0_6 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_6 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_522_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_7 <= 2'h0;
    end else if (bht_bank_sel_0_0_7) begin
      if (_T_6629) begin
        bht_bank_rd_data_out_0_7 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_7 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_522_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_8 <= 2'h0;
    end else if (bht_bank_sel_0_0_8) begin
      if (_T_6638) begin
        bht_bank_rd_data_out_0_8 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_8 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_522_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_9 <= 2'h0;
    end else if (bht_bank_sel_0_0_9) begin
      if (_T_6647) begin
        bht_bank_rd_data_out_0_9 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_9 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_522_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_10 <= 2'h0;
    end else if (bht_bank_sel_0_0_10) begin
      if (_T_6656) begin
        bht_bank_rd_data_out_0_10 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_10 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_522_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_11 <= 2'h0;
    end else if (bht_bank_sel_0_0_11) begin
      if (_T_6665) begin
        bht_bank_rd_data_out_0_11 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_11 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_522_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_12 <= 2'h0;
    end else if (bht_bank_sel_0_0_12) begin
      if (_T_6674) begin
        bht_bank_rd_data_out_0_12 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_12 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_522_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_13 <= 2'h0;
    end else if (bht_bank_sel_0_0_13) begin
      if (_T_6683) begin
        bht_bank_rd_data_out_0_13 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_13 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_522_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_14 <= 2'h0;
    end else if (bht_bank_sel_0_0_14) begin
      if (_T_6692) begin
        bht_bank_rd_data_out_0_14 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_14 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_522_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_15 <= 2'h0;
    end else if (bht_bank_sel_0_0_15) begin
      if (_T_6701) begin
        bht_bank_rd_data_out_0_15 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_15 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_523_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_16 <= 2'h0;
    end else if (bht_bank_sel_0_1_0) begin
      if (_T_6710) begin
        bht_bank_rd_data_out_0_16 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_16 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_523_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_17 <= 2'h0;
    end else if (bht_bank_sel_0_1_1) begin
      if (_T_6719) begin
        bht_bank_rd_data_out_0_17 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_17 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_523_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_18 <= 2'h0;
    end else if (bht_bank_sel_0_1_2) begin
      if (_T_6728) begin
        bht_bank_rd_data_out_0_18 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_18 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_523_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_19 <= 2'h0;
    end else if (bht_bank_sel_0_1_3) begin
      if (_T_6737) begin
        bht_bank_rd_data_out_0_19 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_19 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_523_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_20 <= 2'h0;
    end else if (bht_bank_sel_0_1_4) begin
      if (_T_6746) begin
        bht_bank_rd_data_out_0_20 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_20 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_523_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_21 <= 2'h0;
    end else if (bht_bank_sel_0_1_5) begin
      if (_T_6755) begin
        bht_bank_rd_data_out_0_21 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_21 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_523_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_22 <= 2'h0;
    end else if (bht_bank_sel_0_1_6) begin
      if (_T_6764) begin
        bht_bank_rd_data_out_0_22 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_22 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_523_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_23 <= 2'h0;
    end else if (bht_bank_sel_0_1_7) begin
      if (_T_6773) begin
        bht_bank_rd_data_out_0_23 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_23 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_523_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_24 <= 2'h0;
    end else if (bht_bank_sel_0_1_8) begin
      if (_T_6782) begin
        bht_bank_rd_data_out_0_24 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_24 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_523_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_25 <= 2'h0;
    end else if (bht_bank_sel_0_1_9) begin
      if (_T_6791) begin
        bht_bank_rd_data_out_0_25 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_25 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_523_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_26 <= 2'h0;
    end else if (bht_bank_sel_0_1_10) begin
      if (_T_6800) begin
        bht_bank_rd_data_out_0_26 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_26 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_523_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_27 <= 2'h0;
    end else if (bht_bank_sel_0_1_11) begin
      if (_T_6809) begin
        bht_bank_rd_data_out_0_27 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_27 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_523_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_28 <= 2'h0;
    end else if (bht_bank_sel_0_1_12) begin
      if (_T_6818) begin
        bht_bank_rd_data_out_0_28 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_28 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_523_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_29 <= 2'h0;
    end else if (bht_bank_sel_0_1_13) begin
      if (_T_6827) begin
        bht_bank_rd_data_out_0_29 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_29 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_523_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_30 <= 2'h0;
    end else if (bht_bank_sel_0_1_14) begin
      if (_T_6836) begin
        bht_bank_rd_data_out_0_30 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_30 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_523_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_31 <= 2'h0;
    end else if (bht_bank_sel_0_1_15) begin
      if (_T_6845) begin
        bht_bank_rd_data_out_0_31 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_31 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_524_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_32 <= 2'h0;
    end else if (bht_bank_sel_0_2_0) begin
      if (_T_6854) begin
        bht_bank_rd_data_out_0_32 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_32 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_524_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_33 <= 2'h0;
    end else if (bht_bank_sel_0_2_1) begin
      if (_T_6863) begin
        bht_bank_rd_data_out_0_33 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_33 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_524_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_34 <= 2'h0;
    end else if (bht_bank_sel_0_2_2) begin
      if (_T_6872) begin
        bht_bank_rd_data_out_0_34 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_34 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_524_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_35 <= 2'h0;
    end else if (bht_bank_sel_0_2_3) begin
      if (_T_6881) begin
        bht_bank_rd_data_out_0_35 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_35 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_524_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_36 <= 2'h0;
    end else if (bht_bank_sel_0_2_4) begin
      if (_T_6890) begin
        bht_bank_rd_data_out_0_36 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_36 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_524_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_37 <= 2'h0;
    end else if (bht_bank_sel_0_2_5) begin
      if (_T_6899) begin
        bht_bank_rd_data_out_0_37 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_37 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_524_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_38 <= 2'h0;
    end else if (bht_bank_sel_0_2_6) begin
      if (_T_6908) begin
        bht_bank_rd_data_out_0_38 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_38 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_524_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_39 <= 2'h0;
    end else if (bht_bank_sel_0_2_7) begin
      if (_T_6917) begin
        bht_bank_rd_data_out_0_39 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_39 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_524_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_40 <= 2'h0;
    end else if (bht_bank_sel_0_2_8) begin
      if (_T_6926) begin
        bht_bank_rd_data_out_0_40 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_40 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_524_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_41 <= 2'h0;
    end else if (bht_bank_sel_0_2_9) begin
      if (_T_6935) begin
        bht_bank_rd_data_out_0_41 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_41 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_524_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_42 <= 2'h0;
    end else if (bht_bank_sel_0_2_10) begin
      if (_T_6944) begin
        bht_bank_rd_data_out_0_42 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_42 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_524_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_43 <= 2'h0;
    end else if (bht_bank_sel_0_2_11) begin
      if (_T_6953) begin
        bht_bank_rd_data_out_0_43 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_43 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_524_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_44 <= 2'h0;
    end else if (bht_bank_sel_0_2_12) begin
      if (_T_6962) begin
        bht_bank_rd_data_out_0_44 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_44 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_524_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_45 <= 2'h0;
    end else if (bht_bank_sel_0_2_13) begin
      if (_T_6971) begin
        bht_bank_rd_data_out_0_45 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_45 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_524_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_46 <= 2'h0;
    end else if (bht_bank_sel_0_2_14) begin
      if (_T_6980) begin
        bht_bank_rd_data_out_0_46 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_46 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_524_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_47 <= 2'h0;
    end else if (bht_bank_sel_0_2_15) begin
      if (_T_6989) begin
        bht_bank_rd_data_out_0_47 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_47 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_525_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_48 <= 2'h0;
    end else if (bht_bank_sel_0_3_0) begin
      if (_T_6998) begin
        bht_bank_rd_data_out_0_48 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_48 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_525_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_49 <= 2'h0;
    end else if (bht_bank_sel_0_3_1) begin
      if (_T_7007) begin
        bht_bank_rd_data_out_0_49 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_49 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_525_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_50 <= 2'h0;
    end else if (bht_bank_sel_0_3_2) begin
      if (_T_7016) begin
        bht_bank_rd_data_out_0_50 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_50 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_525_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_51 <= 2'h0;
    end else if (bht_bank_sel_0_3_3) begin
      if (_T_7025) begin
        bht_bank_rd_data_out_0_51 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_51 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_525_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_52 <= 2'h0;
    end else if (bht_bank_sel_0_3_4) begin
      if (_T_7034) begin
        bht_bank_rd_data_out_0_52 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_52 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_525_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_53 <= 2'h0;
    end else if (bht_bank_sel_0_3_5) begin
      if (_T_7043) begin
        bht_bank_rd_data_out_0_53 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_53 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_525_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_54 <= 2'h0;
    end else if (bht_bank_sel_0_3_6) begin
      if (_T_7052) begin
        bht_bank_rd_data_out_0_54 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_54 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_525_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_55 <= 2'h0;
    end else if (bht_bank_sel_0_3_7) begin
      if (_T_7061) begin
        bht_bank_rd_data_out_0_55 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_55 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_525_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_56 <= 2'h0;
    end else if (bht_bank_sel_0_3_8) begin
      if (_T_7070) begin
        bht_bank_rd_data_out_0_56 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_56 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_525_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_57 <= 2'h0;
    end else if (bht_bank_sel_0_3_9) begin
      if (_T_7079) begin
        bht_bank_rd_data_out_0_57 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_57 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_525_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_58 <= 2'h0;
    end else if (bht_bank_sel_0_3_10) begin
      if (_T_7088) begin
        bht_bank_rd_data_out_0_58 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_58 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_525_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_59 <= 2'h0;
    end else if (bht_bank_sel_0_3_11) begin
      if (_T_7097) begin
        bht_bank_rd_data_out_0_59 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_59 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_525_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_60 <= 2'h0;
    end else if (bht_bank_sel_0_3_12) begin
      if (_T_7106) begin
        bht_bank_rd_data_out_0_60 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_60 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_525_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_61 <= 2'h0;
    end else if (bht_bank_sel_0_3_13) begin
      if (_T_7115) begin
        bht_bank_rd_data_out_0_61 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_61 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_525_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_62 <= 2'h0;
    end else if (bht_bank_sel_0_3_14) begin
      if (_T_7124) begin
        bht_bank_rd_data_out_0_62 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_62 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_525_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_63 <= 2'h0;
    end else if (bht_bank_sel_0_3_15) begin
      if (_T_7133) begin
        bht_bank_rd_data_out_0_63 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_63 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_526_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_64 <= 2'h0;
    end else if (bht_bank_sel_0_4_0) begin
      if (_T_7142) begin
        bht_bank_rd_data_out_0_64 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_64 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_526_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_65 <= 2'h0;
    end else if (bht_bank_sel_0_4_1) begin
      if (_T_7151) begin
        bht_bank_rd_data_out_0_65 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_65 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_526_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_66 <= 2'h0;
    end else if (bht_bank_sel_0_4_2) begin
      if (_T_7160) begin
        bht_bank_rd_data_out_0_66 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_66 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_526_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_67 <= 2'h0;
    end else if (bht_bank_sel_0_4_3) begin
      if (_T_7169) begin
        bht_bank_rd_data_out_0_67 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_67 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_526_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_68 <= 2'h0;
    end else if (bht_bank_sel_0_4_4) begin
      if (_T_7178) begin
        bht_bank_rd_data_out_0_68 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_68 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_526_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_69 <= 2'h0;
    end else if (bht_bank_sel_0_4_5) begin
      if (_T_7187) begin
        bht_bank_rd_data_out_0_69 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_69 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_526_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_70 <= 2'h0;
    end else if (bht_bank_sel_0_4_6) begin
      if (_T_7196) begin
        bht_bank_rd_data_out_0_70 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_70 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_526_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_71 <= 2'h0;
    end else if (bht_bank_sel_0_4_7) begin
      if (_T_7205) begin
        bht_bank_rd_data_out_0_71 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_71 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_526_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_72 <= 2'h0;
    end else if (bht_bank_sel_0_4_8) begin
      if (_T_7214) begin
        bht_bank_rd_data_out_0_72 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_72 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_526_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_73 <= 2'h0;
    end else if (bht_bank_sel_0_4_9) begin
      if (_T_7223) begin
        bht_bank_rd_data_out_0_73 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_73 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_526_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_74 <= 2'h0;
    end else if (bht_bank_sel_0_4_10) begin
      if (_T_7232) begin
        bht_bank_rd_data_out_0_74 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_74 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_526_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_75 <= 2'h0;
    end else if (bht_bank_sel_0_4_11) begin
      if (_T_7241) begin
        bht_bank_rd_data_out_0_75 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_75 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_526_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_76 <= 2'h0;
    end else if (bht_bank_sel_0_4_12) begin
      if (_T_7250) begin
        bht_bank_rd_data_out_0_76 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_76 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_526_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_77 <= 2'h0;
    end else if (bht_bank_sel_0_4_13) begin
      if (_T_7259) begin
        bht_bank_rd_data_out_0_77 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_77 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_526_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_78 <= 2'h0;
    end else if (bht_bank_sel_0_4_14) begin
      if (_T_7268) begin
        bht_bank_rd_data_out_0_78 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_78 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_526_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_79 <= 2'h0;
    end else if (bht_bank_sel_0_4_15) begin
      if (_T_7277) begin
        bht_bank_rd_data_out_0_79 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_79 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_527_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_80 <= 2'h0;
    end else if (bht_bank_sel_0_5_0) begin
      if (_T_7286) begin
        bht_bank_rd_data_out_0_80 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_80 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_527_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_81 <= 2'h0;
    end else if (bht_bank_sel_0_5_1) begin
      if (_T_7295) begin
        bht_bank_rd_data_out_0_81 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_81 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_527_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_82 <= 2'h0;
    end else if (bht_bank_sel_0_5_2) begin
      if (_T_7304) begin
        bht_bank_rd_data_out_0_82 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_82 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_527_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_83 <= 2'h0;
    end else if (bht_bank_sel_0_5_3) begin
      if (_T_7313) begin
        bht_bank_rd_data_out_0_83 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_83 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_527_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_84 <= 2'h0;
    end else if (bht_bank_sel_0_5_4) begin
      if (_T_7322) begin
        bht_bank_rd_data_out_0_84 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_84 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_527_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_85 <= 2'h0;
    end else if (bht_bank_sel_0_5_5) begin
      if (_T_7331) begin
        bht_bank_rd_data_out_0_85 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_85 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_527_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_86 <= 2'h0;
    end else if (bht_bank_sel_0_5_6) begin
      if (_T_7340) begin
        bht_bank_rd_data_out_0_86 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_86 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_527_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_87 <= 2'h0;
    end else if (bht_bank_sel_0_5_7) begin
      if (_T_7349) begin
        bht_bank_rd_data_out_0_87 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_87 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_527_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_88 <= 2'h0;
    end else if (bht_bank_sel_0_5_8) begin
      if (_T_7358) begin
        bht_bank_rd_data_out_0_88 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_88 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_527_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_89 <= 2'h0;
    end else if (bht_bank_sel_0_5_9) begin
      if (_T_7367) begin
        bht_bank_rd_data_out_0_89 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_89 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_527_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_90 <= 2'h0;
    end else if (bht_bank_sel_0_5_10) begin
      if (_T_7376) begin
        bht_bank_rd_data_out_0_90 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_90 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_527_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_91 <= 2'h0;
    end else if (bht_bank_sel_0_5_11) begin
      if (_T_7385) begin
        bht_bank_rd_data_out_0_91 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_91 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_527_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_92 <= 2'h0;
    end else if (bht_bank_sel_0_5_12) begin
      if (_T_7394) begin
        bht_bank_rd_data_out_0_92 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_92 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_527_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_93 <= 2'h0;
    end else if (bht_bank_sel_0_5_13) begin
      if (_T_7403) begin
        bht_bank_rd_data_out_0_93 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_93 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_527_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_94 <= 2'h0;
    end else if (bht_bank_sel_0_5_14) begin
      if (_T_7412) begin
        bht_bank_rd_data_out_0_94 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_94 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_527_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_95 <= 2'h0;
    end else if (bht_bank_sel_0_5_15) begin
      if (_T_7421) begin
        bht_bank_rd_data_out_0_95 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_95 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_528_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_96 <= 2'h0;
    end else if (bht_bank_sel_0_6_0) begin
      if (_T_7430) begin
        bht_bank_rd_data_out_0_96 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_96 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_528_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_97 <= 2'h0;
    end else if (bht_bank_sel_0_6_1) begin
      if (_T_7439) begin
        bht_bank_rd_data_out_0_97 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_97 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_528_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_98 <= 2'h0;
    end else if (bht_bank_sel_0_6_2) begin
      if (_T_7448) begin
        bht_bank_rd_data_out_0_98 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_98 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_528_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_99 <= 2'h0;
    end else if (bht_bank_sel_0_6_3) begin
      if (_T_7457) begin
        bht_bank_rd_data_out_0_99 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_99 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_528_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_100 <= 2'h0;
    end else if (bht_bank_sel_0_6_4) begin
      if (_T_7466) begin
        bht_bank_rd_data_out_0_100 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_100 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_528_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_101 <= 2'h0;
    end else if (bht_bank_sel_0_6_5) begin
      if (_T_7475) begin
        bht_bank_rd_data_out_0_101 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_101 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_528_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_102 <= 2'h0;
    end else if (bht_bank_sel_0_6_6) begin
      if (_T_7484) begin
        bht_bank_rd_data_out_0_102 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_102 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_528_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_103 <= 2'h0;
    end else if (bht_bank_sel_0_6_7) begin
      if (_T_7493) begin
        bht_bank_rd_data_out_0_103 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_103 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_528_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_104 <= 2'h0;
    end else if (bht_bank_sel_0_6_8) begin
      if (_T_7502) begin
        bht_bank_rd_data_out_0_104 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_104 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_528_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_105 <= 2'h0;
    end else if (bht_bank_sel_0_6_9) begin
      if (_T_7511) begin
        bht_bank_rd_data_out_0_105 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_105 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_528_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_106 <= 2'h0;
    end else if (bht_bank_sel_0_6_10) begin
      if (_T_7520) begin
        bht_bank_rd_data_out_0_106 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_106 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_528_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_107 <= 2'h0;
    end else if (bht_bank_sel_0_6_11) begin
      if (_T_7529) begin
        bht_bank_rd_data_out_0_107 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_107 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_528_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_108 <= 2'h0;
    end else if (bht_bank_sel_0_6_12) begin
      if (_T_7538) begin
        bht_bank_rd_data_out_0_108 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_108 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_528_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_109 <= 2'h0;
    end else if (bht_bank_sel_0_6_13) begin
      if (_T_7547) begin
        bht_bank_rd_data_out_0_109 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_109 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_528_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_110 <= 2'h0;
    end else if (bht_bank_sel_0_6_14) begin
      if (_T_7556) begin
        bht_bank_rd_data_out_0_110 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_110 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_528_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_111 <= 2'h0;
    end else if (bht_bank_sel_0_6_15) begin
      if (_T_7565) begin
        bht_bank_rd_data_out_0_111 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_111 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_529_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_112 <= 2'h0;
    end else if (bht_bank_sel_0_7_0) begin
      if (_T_7574) begin
        bht_bank_rd_data_out_0_112 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_112 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_529_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_113 <= 2'h0;
    end else if (bht_bank_sel_0_7_1) begin
      if (_T_7583) begin
        bht_bank_rd_data_out_0_113 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_113 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_529_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_114 <= 2'h0;
    end else if (bht_bank_sel_0_7_2) begin
      if (_T_7592) begin
        bht_bank_rd_data_out_0_114 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_114 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_529_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_115 <= 2'h0;
    end else if (bht_bank_sel_0_7_3) begin
      if (_T_7601) begin
        bht_bank_rd_data_out_0_115 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_115 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_529_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_116 <= 2'h0;
    end else if (bht_bank_sel_0_7_4) begin
      if (_T_7610) begin
        bht_bank_rd_data_out_0_116 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_116 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_529_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_117 <= 2'h0;
    end else if (bht_bank_sel_0_7_5) begin
      if (_T_7619) begin
        bht_bank_rd_data_out_0_117 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_117 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_529_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_118 <= 2'h0;
    end else if (bht_bank_sel_0_7_6) begin
      if (_T_7628) begin
        bht_bank_rd_data_out_0_118 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_118 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_529_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_119 <= 2'h0;
    end else if (bht_bank_sel_0_7_7) begin
      if (_T_7637) begin
        bht_bank_rd_data_out_0_119 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_119 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_529_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_120 <= 2'h0;
    end else if (bht_bank_sel_0_7_8) begin
      if (_T_7646) begin
        bht_bank_rd_data_out_0_120 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_120 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_529_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_121 <= 2'h0;
    end else if (bht_bank_sel_0_7_9) begin
      if (_T_7655) begin
        bht_bank_rd_data_out_0_121 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_121 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_529_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_122 <= 2'h0;
    end else if (bht_bank_sel_0_7_10) begin
      if (_T_7664) begin
        bht_bank_rd_data_out_0_122 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_122 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_529_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_123 <= 2'h0;
    end else if (bht_bank_sel_0_7_11) begin
      if (_T_7673) begin
        bht_bank_rd_data_out_0_123 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_123 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_529_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_124 <= 2'h0;
    end else if (bht_bank_sel_0_7_12) begin
      if (_T_7682) begin
        bht_bank_rd_data_out_0_124 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_124 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_529_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_125 <= 2'h0;
    end else if (bht_bank_sel_0_7_13) begin
      if (_T_7691) begin
        bht_bank_rd_data_out_0_125 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_125 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_529_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_126 <= 2'h0;
    end else if (bht_bank_sel_0_7_14) begin
      if (_T_7700) begin
        bht_bank_rd_data_out_0_126 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_126 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_529_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_127 <= 2'h0;
    end else if (bht_bank_sel_0_7_15) begin
      if (_T_7709) begin
        bht_bank_rd_data_out_0_127 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_127 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_530_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_128 <= 2'h0;
    end else if (bht_bank_sel_0_8_0) begin
      if (_T_7718) begin
        bht_bank_rd_data_out_0_128 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_128 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_530_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_129 <= 2'h0;
    end else if (bht_bank_sel_0_8_1) begin
      if (_T_7727) begin
        bht_bank_rd_data_out_0_129 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_129 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_530_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_130 <= 2'h0;
    end else if (bht_bank_sel_0_8_2) begin
      if (_T_7736) begin
        bht_bank_rd_data_out_0_130 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_130 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_530_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_131 <= 2'h0;
    end else if (bht_bank_sel_0_8_3) begin
      if (_T_7745) begin
        bht_bank_rd_data_out_0_131 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_131 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_530_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_132 <= 2'h0;
    end else if (bht_bank_sel_0_8_4) begin
      if (_T_7754) begin
        bht_bank_rd_data_out_0_132 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_132 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_530_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_133 <= 2'h0;
    end else if (bht_bank_sel_0_8_5) begin
      if (_T_7763) begin
        bht_bank_rd_data_out_0_133 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_133 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_530_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_134 <= 2'h0;
    end else if (bht_bank_sel_0_8_6) begin
      if (_T_7772) begin
        bht_bank_rd_data_out_0_134 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_134 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_530_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_135 <= 2'h0;
    end else if (bht_bank_sel_0_8_7) begin
      if (_T_7781) begin
        bht_bank_rd_data_out_0_135 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_135 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_530_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_136 <= 2'h0;
    end else if (bht_bank_sel_0_8_8) begin
      if (_T_7790) begin
        bht_bank_rd_data_out_0_136 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_136 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_530_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_137 <= 2'h0;
    end else if (bht_bank_sel_0_8_9) begin
      if (_T_7799) begin
        bht_bank_rd_data_out_0_137 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_137 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_530_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_138 <= 2'h0;
    end else if (bht_bank_sel_0_8_10) begin
      if (_T_7808) begin
        bht_bank_rd_data_out_0_138 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_138 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_530_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_139 <= 2'h0;
    end else if (bht_bank_sel_0_8_11) begin
      if (_T_7817) begin
        bht_bank_rd_data_out_0_139 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_139 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_530_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_140 <= 2'h0;
    end else if (bht_bank_sel_0_8_12) begin
      if (_T_7826) begin
        bht_bank_rd_data_out_0_140 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_140 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_530_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_141 <= 2'h0;
    end else if (bht_bank_sel_0_8_13) begin
      if (_T_7835) begin
        bht_bank_rd_data_out_0_141 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_141 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_530_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_142 <= 2'h0;
    end else if (bht_bank_sel_0_8_14) begin
      if (_T_7844) begin
        bht_bank_rd_data_out_0_142 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_142 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_530_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_143 <= 2'h0;
    end else if (bht_bank_sel_0_8_15) begin
      if (_T_7853) begin
        bht_bank_rd_data_out_0_143 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_143 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_531_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_144 <= 2'h0;
    end else if (bht_bank_sel_0_9_0) begin
      if (_T_7862) begin
        bht_bank_rd_data_out_0_144 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_144 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_531_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_145 <= 2'h0;
    end else if (bht_bank_sel_0_9_1) begin
      if (_T_7871) begin
        bht_bank_rd_data_out_0_145 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_145 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_531_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_146 <= 2'h0;
    end else if (bht_bank_sel_0_9_2) begin
      if (_T_7880) begin
        bht_bank_rd_data_out_0_146 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_146 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_531_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_147 <= 2'h0;
    end else if (bht_bank_sel_0_9_3) begin
      if (_T_7889) begin
        bht_bank_rd_data_out_0_147 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_147 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_531_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_148 <= 2'h0;
    end else if (bht_bank_sel_0_9_4) begin
      if (_T_7898) begin
        bht_bank_rd_data_out_0_148 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_148 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_531_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_149 <= 2'h0;
    end else if (bht_bank_sel_0_9_5) begin
      if (_T_7907) begin
        bht_bank_rd_data_out_0_149 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_149 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_531_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_150 <= 2'h0;
    end else if (bht_bank_sel_0_9_6) begin
      if (_T_7916) begin
        bht_bank_rd_data_out_0_150 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_150 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_531_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_151 <= 2'h0;
    end else if (bht_bank_sel_0_9_7) begin
      if (_T_7925) begin
        bht_bank_rd_data_out_0_151 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_151 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_531_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_152 <= 2'h0;
    end else if (bht_bank_sel_0_9_8) begin
      if (_T_7934) begin
        bht_bank_rd_data_out_0_152 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_152 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_531_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_153 <= 2'h0;
    end else if (bht_bank_sel_0_9_9) begin
      if (_T_7943) begin
        bht_bank_rd_data_out_0_153 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_153 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_531_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_154 <= 2'h0;
    end else if (bht_bank_sel_0_9_10) begin
      if (_T_7952) begin
        bht_bank_rd_data_out_0_154 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_154 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_531_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_155 <= 2'h0;
    end else if (bht_bank_sel_0_9_11) begin
      if (_T_7961) begin
        bht_bank_rd_data_out_0_155 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_155 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_531_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_156 <= 2'h0;
    end else if (bht_bank_sel_0_9_12) begin
      if (_T_7970) begin
        bht_bank_rd_data_out_0_156 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_156 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_531_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_157 <= 2'h0;
    end else if (bht_bank_sel_0_9_13) begin
      if (_T_7979) begin
        bht_bank_rd_data_out_0_157 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_157 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_531_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_158 <= 2'h0;
    end else if (bht_bank_sel_0_9_14) begin
      if (_T_7988) begin
        bht_bank_rd_data_out_0_158 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_158 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_531_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_159 <= 2'h0;
    end else if (bht_bank_sel_0_9_15) begin
      if (_T_7997) begin
        bht_bank_rd_data_out_0_159 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_159 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_532_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_160 <= 2'h0;
    end else if (bht_bank_sel_0_10_0) begin
      if (_T_8006) begin
        bht_bank_rd_data_out_0_160 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_160 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_532_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_161 <= 2'h0;
    end else if (bht_bank_sel_0_10_1) begin
      if (_T_8015) begin
        bht_bank_rd_data_out_0_161 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_161 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_532_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_162 <= 2'h0;
    end else if (bht_bank_sel_0_10_2) begin
      if (_T_8024) begin
        bht_bank_rd_data_out_0_162 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_162 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_532_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_163 <= 2'h0;
    end else if (bht_bank_sel_0_10_3) begin
      if (_T_8033) begin
        bht_bank_rd_data_out_0_163 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_163 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_532_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_164 <= 2'h0;
    end else if (bht_bank_sel_0_10_4) begin
      if (_T_8042) begin
        bht_bank_rd_data_out_0_164 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_164 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_532_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_165 <= 2'h0;
    end else if (bht_bank_sel_0_10_5) begin
      if (_T_8051) begin
        bht_bank_rd_data_out_0_165 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_165 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_532_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_166 <= 2'h0;
    end else if (bht_bank_sel_0_10_6) begin
      if (_T_8060) begin
        bht_bank_rd_data_out_0_166 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_166 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_532_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_167 <= 2'h0;
    end else if (bht_bank_sel_0_10_7) begin
      if (_T_8069) begin
        bht_bank_rd_data_out_0_167 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_167 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_532_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_168 <= 2'h0;
    end else if (bht_bank_sel_0_10_8) begin
      if (_T_8078) begin
        bht_bank_rd_data_out_0_168 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_168 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_532_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_169 <= 2'h0;
    end else if (bht_bank_sel_0_10_9) begin
      if (_T_8087) begin
        bht_bank_rd_data_out_0_169 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_169 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_532_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_170 <= 2'h0;
    end else if (bht_bank_sel_0_10_10) begin
      if (_T_8096) begin
        bht_bank_rd_data_out_0_170 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_170 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_532_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_171 <= 2'h0;
    end else if (bht_bank_sel_0_10_11) begin
      if (_T_8105) begin
        bht_bank_rd_data_out_0_171 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_171 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_532_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_172 <= 2'h0;
    end else if (bht_bank_sel_0_10_12) begin
      if (_T_8114) begin
        bht_bank_rd_data_out_0_172 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_172 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_532_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_173 <= 2'h0;
    end else if (bht_bank_sel_0_10_13) begin
      if (_T_8123) begin
        bht_bank_rd_data_out_0_173 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_173 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_532_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_174 <= 2'h0;
    end else if (bht_bank_sel_0_10_14) begin
      if (_T_8132) begin
        bht_bank_rd_data_out_0_174 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_174 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_532_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_175 <= 2'h0;
    end else if (bht_bank_sel_0_10_15) begin
      if (_T_8141) begin
        bht_bank_rd_data_out_0_175 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_175 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_533_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_176 <= 2'h0;
    end else if (bht_bank_sel_0_11_0) begin
      if (_T_8150) begin
        bht_bank_rd_data_out_0_176 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_176 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_533_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_177 <= 2'h0;
    end else if (bht_bank_sel_0_11_1) begin
      if (_T_8159) begin
        bht_bank_rd_data_out_0_177 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_177 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_533_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_178 <= 2'h0;
    end else if (bht_bank_sel_0_11_2) begin
      if (_T_8168) begin
        bht_bank_rd_data_out_0_178 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_178 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_533_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_179 <= 2'h0;
    end else if (bht_bank_sel_0_11_3) begin
      if (_T_8177) begin
        bht_bank_rd_data_out_0_179 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_179 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_533_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_180 <= 2'h0;
    end else if (bht_bank_sel_0_11_4) begin
      if (_T_8186) begin
        bht_bank_rd_data_out_0_180 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_180 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_533_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_181 <= 2'h0;
    end else if (bht_bank_sel_0_11_5) begin
      if (_T_8195) begin
        bht_bank_rd_data_out_0_181 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_181 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_533_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_182 <= 2'h0;
    end else if (bht_bank_sel_0_11_6) begin
      if (_T_8204) begin
        bht_bank_rd_data_out_0_182 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_182 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_533_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_183 <= 2'h0;
    end else if (bht_bank_sel_0_11_7) begin
      if (_T_8213) begin
        bht_bank_rd_data_out_0_183 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_183 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_533_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_184 <= 2'h0;
    end else if (bht_bank_sel_0_11_8) begin
      if (_T_8222) begin
        bht_bank_rd_data_out_0_184 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_184 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_533_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_185 <= 2'h0;
    end else if (bht_bank_sel_0_11_9) begin
      if (_T_8231) begin
        bht_bank_rd_data_out_0_185 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_185 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_533_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_186 <= 2'h0;
    end else if (bht_bank_sel_0_11_10) begin
      if (_T_8240) begin
        bht_bank_rd_data_out_0_186 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_186 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_533_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_187 <= 2'h0;
    end else if (bht_bank_sel_0_11_11) begin
      if (_T_8249) begin
        bht_bank_rd_data_out_0_187 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_187 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_533_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_188 <= 2'h0;
    end else if (bht_bank_sel_0_11_12) begin
      if (_T_8258) begin
        bht_bank_rd_data_out_0_188 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_188 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_533_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_189 <= 2'h0;
    end else if (bht_bank_sel_0_11_13) begin
      if (_T_8267) begin
        bht_bank_rd_data_out_0_189 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_189 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_533_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_190 <= 2'h0;
    end else if (bht_bank_sel_0_11_14) begin
      if (_T_8276) begin
        bht_bank_rd_data_out_0_190 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_190 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_533_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_191 <= 2'h0;
    end else if (bht_bank_sel_0_11_15) begin
      if (_T_8285) begin
        bht_bank_rd_data_out_0_191 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_191 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_534_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_192 <= 2'h0;
    end else if (bht_bank_sel_0_12_0) begin
      if (_T_8294) begin
        bht_bank_rd_data_out_0_192 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_192 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_534_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_193 <= 2'h0;
    end else if (bht_bank_sel_0_12_1) begin
      if (_T_8303) begin
        bht_bank_rd_data_out_0_193 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_193 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_534_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_194 <= 2'h0;
    end else if (bht_bank_sel_0_12_2) begin
      if (_T_8312) begin
        bht_bank_rd_data_out_0_194 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_194 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_534_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_195 <= 2'h0;
    end else if (bht_bank_sel_0_12_3) begin
      if (_T_8321) begin
        bht_bank_rd_data_out_0_195 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_195 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_534_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_196 <= 2'h0;
    end else if (bht_bank_sel_0_12_4) begin
      if (_T_8330) begin
        bht_bank_rd_data_out_0_196 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_196 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_534_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_197 <= 2'h0;
    end else if (bht_bank_sel_0_12_5) begin
      if (_T_8339) begin
        bht_bank_rd_data_out_0_197 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_197 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_534_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_198 <= 2'h0;
    end else if (bht_bank_sel_0_12_6) begin
      if (_T_8348) begin
        bht_bank_rd_data_out_0_198 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_198 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_534_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_199 <= 2'h0;
    end else if (bht_bank_sel_0_12_7) begin
      if (_T_8357) begin
        bht_bank_rd_data_out_0_199 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_199 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_534_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_200 <= 2'h0;
    end else if (bht_bank_sel_0_12_8) begin
      if (_T_8366) begin
        bht_bank_rd_data_out_0_200 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_200 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_534_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_201 <= 2'h0;
    end else if (bht_bank_sel_0_12_9) begin
      if (_T_8375) begin
        bht_bank_rd_data_out_0_201 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_201 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_534_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_202 <= 2'h0;
    end else if (bht_bank_sel_0_12_10) begin
      if (_T_8384) begin
        bht_bank_rd_data_out_0_202 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_202 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_534_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_203 <= 2'h0;
    end else if (bht_bank_sel_0_12_11) begin
      if (_T_8393) begin
        bht_bank_rd_data_out_0_203 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_203 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_534_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_204 <= 2'h0;
    end else if (bht_bank_sel_0_12_12) begin
      if (_T_8402) begin
        bht_bank_rd_data_out_0_204 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_204 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_534_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_205 <= 2'h0;
    end else if (bht_bank_sel_0_12_13) begin
      if (_T_8411) begin
        bht_bank_rd_data_out_0_205 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_205 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_534_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_206 <= 2'h0;
    end else if (bht_bank_sel_0_12_14) begin
      if (_T_8420) begin
        bht_bank_rd_data_out_0_206 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_206 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_534_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_207 <= 2'h0;
    end else if (bht_bank_sel_0_12_15) begin
      if (_T_8429) begin
        bht_bank_rd_data_out_0_207 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_207 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_535_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_208 <= 2'h0;
    end else if (bht_bank_sel_0_13_0) begin
      if (_T_8438) begin
        bht_bank_rd_data_out_0_208 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_208 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_535_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_209 <= 2'h0;
    end else if (bht_bank_sel_0_13_1) begin
      if (_T_8447) begin
        bht_bank_rd_data_out_0_209 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_209 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_535_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_210 <= 2'h0;
    end else if (bht_bank_sel_0_13_2) begin
      if (_T_8456) begin
        bht_bank_rd_data_out_0_210 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_210 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_535_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_211 <= 2'h0;
    end else if (bht_bank_sel_0_13_3) begin
      if (_T_8465) begin
        bht_bank_rd_data_out_0_211 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_211 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_535_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_212 <= 2'h0;
    end else if (bht_bank_sel_0_13_4) begin
      if (_T_8474) begin
        bht_bank_rd_data_out_0_212 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_212 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_535_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_213 <= 2'h0;
    end else if (bht_bank_sel_0_13_5) begin
      if (_T_8483) begin
        bht_bank_rd_data_out_0_213 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_213 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_535_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_214 <= 2'h0;
    end else if (bht_bank_sel_0_13_6) begin
      if (_T_8492) begin
        bht_bank_rd_data_out_0_214 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_214 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_535_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_215 <= 2'h0;
    end else if (bht_bank_sel_0_13_7) begin
      if (_T_8501) begin
        bht_bank_rd_data_out_0_215 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_215 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_535_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_216 <= 2'h0;
    end else if (bht_bank_sel_0_13_8) begin
      if (_T_8510) begin
        bht_bank_rd_data_out_0_216 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_216 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_535_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_217 <= 2'h0;
    end else if (bht_bank_sel_0_13_9) begin
      if (_T_8519) begin
        bht_bank_rd_data_out_0_217 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_217 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_535_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_218 <= 2'h0;
    end else if (bht_bank_sel_0_13_10) begin
      if (_T_8528) begin
        bht_bank_rd_data_out_0_218 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_218 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_535_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_219 <= 2'h0;
    end else if (bht_bank_sel_0_13_11) begin
      if (_T_8537) begin
        bht_bank_rd_data_out_0_219 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_219 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_535_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_220 <= 2'h0;
    end else if (bht_bank_sel_0_13_12) begin
      if (_T_8546) begin
        bht_bank_rd_data_out_0_220 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_220 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_535_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_221 <= 2'h0;
    end else if (bht_bank_sel_0_13_13) begin
      if (_T_8555) begin
        bht_bank_rd_data_out_0_221 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_221 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_535_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_222 <= 2'h0;
    end else if (bht_bank_sel_0_13_14) begin
      if (_T_8564) begin
        bht_bank_rd_data_out_0_222 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_222 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_535_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_223 <= 2'h0;
    end else if (bht_bank_sel_0_13_15) begin
      if (_T_8573) begin
        bht_bank_rd_data_out_0_223 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_223 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_536_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_224 <= 2'h0;
    end else if (bht_bank_sel_0_14_0) begin
      if (_T_8582) begin
        bht_bank_rd_data_out_0_224 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_224 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_536_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_225 <= 2'h0;
    end else if (bht_bank_sel_0_14_1) begin
      if (_T_8591) begin
        bht_bank_rd_data_out_0_225 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_225 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_536_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_226 <= 2'h0;
    end else if (bht_bank_sel_0_14_2) begin
      if (_T_8600) begin
        bht_bank_rd_data_out_0_226 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_226 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_536_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_227 <= 2'h0;
    end else if (bht_bank_sel_0_14_3) begin
      if (_T_8609) begin
        bht_bank_rd_data_out_0_227 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_227 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_536_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_228 <= 2'h0;
    end else if (bht_bank_sel_0_14_4) begin
      if (_T_8618) begin
        bht_bank_rd_data_out_0_228 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_228 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_536_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_229 <= 2'h0;
    end else if (bht_bank_sel_0_14_5) begin
      if (_T_8627) begin
        bht_bank_rd_data_out_0_229 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_229 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_536_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_230 <= 2'h0;
    end else if (bht_bank_sel_0_14_6) begin
      if (_T_8636) begin
        bht_bank_rd_data_out_0_230 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_230 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_536_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_231 <= 2'h0;
    end else if (bht_bank_sel_0_14_7) begin
      if (_T_8645) begin
        bht_bank_rd_data_out_0_231 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_231 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_536_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_232 <= 2'h0;
    end else if (bht_bank_sel_0_14_8) begin
      if (_T_8654) begin
        bht_bank_rd_data_out_0_232 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_232 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_536_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_233 <= 2'h0;
    end else if (bht_bank_sel_0_14_9) begin
      if (_T_8663) begin
        bht_bank_rd_data_out_0_233 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_233 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_536_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_234 <= 2'h0;
    end else if (bht_bank_sel_0_14_10) begin
      if (_T_8672) begin
        bht_bank_rd_data_out_0_234 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_234 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_536_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_235 <= 2'h0;
    end else if (bht_bank_sel_0_14_11) begin
      if (_T_8681) begin
        bht_bank_rd_data_out_0_235 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_235 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_536_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_236 <= 2'h0;
    end else if (bht_bank_sel_0_14_12) begin
      if (_T_8690) begin
        bht_bank_rd_data_out_0_236 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_236 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_536_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_237 <= 2'h0;
    end else if (bht_bank_sel_0_14_13) begin
      if (_T_8699) begin
        bht_bank_rd_data_out_0_237 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_237 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_536_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_238 <= 2'h0;
    end else if (bht_bank_sel_0_14_14) begin
      if (_T_8708) begin
        bht_bank_rd_data_out_0_238 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_238 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_536_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_239 <= 2'h0;
    end else if (bht_bank_sel_0_14_15) begin
      if (_T_8717) begin
        bht_bank_rd_data_out_0_239 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_239 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_537_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_240 <= 2'h0;
    end else if (bht_bank_sel_0_15_0) begin
      if (_T_8726) begin
        bht_bank_rd_data_out_0_240 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_240 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_537_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_241 <= 2'h0;
    end else if (bht_bank_sel_0_15_1) begin
      if (_T_8735) begin
        bht_bank_rd_data_out_0_241 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_241 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_537_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_242 <= 2'h0;
    end else if (bht_bank_sel_0_15_2) begin
      if (_T_8744) begin
        bht_bank_rd_data_out_0_242 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_242 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_537_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_243 <= 2'h0;
    end else if (bht_bank_sel_0_15_3) begin
      if (_T_8753) begin
        bht_bank_rd_data_out_0_243 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_243 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_537_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_244 <= 2'h0;
    end else if (bht_bank_sel_0_15_4) begin
      if (_T_8762) begin
        bht_bank_rd_data_out_0_244 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_244 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_537_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_245 <= 2'h0;
    end else if (bht_bank_sel_0_15_5) begin
      if (_T_8771) begin
        bht_bank_rd_data_out_0_245 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_245 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_537_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_246 <= 2'h0;
    end else if (bht_bank_sel_0_15_6) begin
      if (_T_8780) begin
        bht_bank_rd_data_out_0_246 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_246 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_537_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_247 <= 2'h0;
    end else if (bht_bank_sel_0_15_7) begin
      if (_T_8789) begin
        bht_bank_rd_data_out_0_247 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_247 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_537_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_248 <= 2'h0;
    end else if (bht_bank_sel_0_15_8) begin
      if (_T_8798) begin
        bht_bank_rd_data_out_0_248 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_248 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_537_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_249 <= 2'h0;
    end else if (bht_bank_sel_0_15_9) begin
      if (_T_8807) begin
        bht_bank_rd_data_out_0_249 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_249 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_537_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_250 <= 2'h0;
    end else if (bht_bank_sel_0_15_10) begin
      if (_T_8816) begin
        bht_bank_rd_data_out_0_250 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_250 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_537_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_251 <= 2'h0;
    end else if (bht_bank_sel_0_15_11) begin
      if (_T_8825) begin
        bht_bank_rd_data_out_0_251 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_251 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_537_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_252 <= 2'h0;
    end else if (bht_bank_sel_0_15_12) begin
      if (_T_8834) begin
        bht_bank_rd_data_out_0_252 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_252 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_537_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_253 <= 2'h0;
    end else if (bht_bank_sel_0_15_13) begin
      if (_T_8843) begin
        bht_bank_rd_data_out_0_253 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_253 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_537_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_254 <= 2'h0;
    end else if (bht_bank_sel_0_15_14) begin
      if (_T_8852) begin
        bht_bank_rd_data_out_0_254 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_254 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_537_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_255 <= 2'h0;
    end else if (bht_bank_sel_0_15_15) begin
      if (_T_8861) begin
        bht_bank_rd_data_out_0_255 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_255 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      exu_mp_way_f <= 1'h0;
    end else begin
      exu_mp_way_f <= io_exu_bp_exu_mp_pkt_bits_way;
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      exu_flush_final_d1 <= 1'h0;
    end else begin
      exu_flush_final_d1 <= io_exu_flush_final;
    end
  end
  always @(posedge rvclkhdr_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_lru_b0_f <= 256'h0;
    end else begin
      btb_lru_b0_f <= _T_183 | _T_185;
    end
  end
  always @(posedge rvclkhdr_1_io_l1clk or posedge reset) begin
    if (reset) begin
      ifc_fetch_adder_prior <= 30'h0;
    end else begin
      ifc_fetch_adder_prior <= io_ifc_fetch_addr_f[30:1];
    end
  end
  always @(posedge rvclkhdr_2_io_l1clk or posedge reset) begin
    if (reset) begin
      rets_out_0 <= 32'h0;
    end else begin
      rets_out_0 <= _T_482 | _T_483;
    end
  end
  always @(posedge rvclkhdr_3_io_l1clk or posedge reset) begin
    if (reset) begin
      rets_out_1 <= 32'h0;
    end else begin
      rets_out_1 <= _T_487 | _T_488;
    end
  end
  always @(posedge rvclkhdr_4_io_l1clk or posedge reset) begin
    if (reset) begin
      rets_out_2 <= 32'h0;
    end else begin
      rets_out_2 <= _T_492 | _T_493;
    end
  end
  always @(posedge rvclkhdr_5_io_l1clk or posedge reset) begin
    if (reset) begin
      rets_out_3 <= 32'h0;
    end else begin
      rets_out_3 <= _T_497 | _T_498;
    end
  end
  always @(posedge rvclkhdr_6_io_l1clk or posedge reset) begin
    if (reset) begin
      rets_out_4 <= 32'h0;
    end else begin
      rets_out_4 <= _T_502 | _T_503;
    end
  end
  always @(posedge rvclkhdr_7_io_l1clk or posedge reset) begin
    if (reset) begin
      rets_out_5 <= 32'h0;
    end else begin
      rets_out_5 <= _T_507 | _T_508;
    end
  end
  always @(posedge rvclkhdr_8_io_l1clk or posedge reset) begin
    if (reset) begin
      rets_out_6 <= 32'h0;
    end else begin
      rets_out_6 <= _T_512 | _T_513;
    end
  end
  always @(posedge rvclkhdr_9_io_l1clk or posedge reset) begin
    if (reset) begin
      rets_out_7 <= 32'h0;
    end else begin
      rets_out_7 <= rets_out_6;
    end
  end
endmodule
module ifu_compress_ctl(
  input  [15:0] io_din,
  output [31:0] io_dout
);
  wire  _T_2 = ~io_din[14]; // @[ifu_compress_ctl.scala 12:83]
  wire  _T_4 = ~io_din[13]; // @[ifu_compress_ctl.scala 12:83]
  wire  _T_7 = ~io_din[6]; // @[ifu_compress_ctl.scala 12:83]
  wire  _T_9 = ~io_din[5]; // @[ifu_compress_ctl.scala 12:83]
  wire  _T_11 = io_din[15] & _T_2; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_12 = _T_11 & _T_4; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_13 = _T_12 & io_din[10]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_14 = _T_13 & _T_7; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_15 = _T_14 & _T_9; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_16 = _T_15 & io_din[0]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_23 = ~io_din[11]; // @[ifu_compress_ctl.scala 12:83]
  wire  _T_28 = _T_12 & _T_23; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_29 = _T_28 & io_din[10]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_30 = _T_29 & io_din[0]; // @[ifu_compress_ctl.scala 12:110]
  wire  out_30 = _T_16 | _T_30; // @[ifu_compress_ctl.scala 17:53]
  wire  _T_38 = ~io_din[10]; // @[ifu_compress_ctl.scala 12:83]
  wire  _T_40 = ~io_din[9]; // @[ifu_compress_ctl.scala 12:83]
  wire  _T_42 = ~io_din[8]; // @[ifu_compress_ctl.scala 12:83]
  wire  _T_44 = ~io_din[7]; // @[ifu_compress_ctl.scala 12:83]
  wire  _T_50 = ~io_din[4]; // @[ifu_compress_ctl.scala 12:83]
  wire  _T_52 = ~io_din[3]; // @[ifu_compress_ctl.scala 12:83]
  wire  _T_54 = ~io_din[2]; // @[ifu_compress_ctl.scala 12:83]
  wire  _T_56 = _T_2 & io_din[12]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_57 = _T_56 & _T_23; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_58 = _T_57 & _T_38; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_59 = _T_58 & _T_40; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_60 = _T_59 & _T_42; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_61 = _T_60 & _T_44; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_62 = _T_61 & _T_7; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_63 = _T_62 & _T_9; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_64 = _T_63 & _T_50; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_65 = _T_64 & _T_52; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_66 = _T_65 & _T_54; // @[ifu_compress_ctl.scala 12:110]
  wire  out_20 = _T_66 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_79 = _T_28 & io_din[0]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_90 = _T_12 & _T_38; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_91 = _T_90 & io_din[0]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_92 = _T_79 | _T_91; // @[ifu_compress_ctl.scala 21:46]
  wire  _T_102 = _T_12 & io_din[6]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_103 = _T_102 & io_din[0]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_104 = _T_92 | _T_103; // @[ifu_compress_ctl.scala 21:80]
  wire  _T_114 = _T_12 & io_din[5]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_115 = _T_114 & io_din[0]; // @[ifu_compress_ctl.scala 12:110]
  wire  out_14 = _T_104 | _T_115; // @[ifu_compress_ctl.scala 21:113]
  wire  _T_128 = _T_12 & io_din[11]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_129 = _T_128 & _T_38; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_130 = _T_129 & io_din[0]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_142 = _T_128 & io_din[6]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_143 = _T_142 & io_din[0]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_144 = _T_130 | _T_143; // @[ifu_compress_ctl.scala 23:50]
  wire  _T_147 = ~io_din[0]; // @[ifu_compress_ctl.scala 23:101]
  wire  _T_148 = io_din[14] & _T_147; // @[ifu_compress_ctl.scala 23:99]
  wire  out_13 = _T_144 | _T_148; // @[ifu_compress_ctl.scala 23:86]
  wire  _T_161 = _T_102 & io_din[5]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_162 = _T_161 & io_din[0]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_175 = _T_162 | _T_79; // @[ifu_compress_ctl.scala 25:47]
  wire  _T_188 = _T_175 | _T_91; // @[ifu_compress_ctl.scala 25:81]
  wire  _T_190 = ~io_din[15]; // @[ifu_compress_ctl.scala 12:83]
  wire  _T_194 = _T_190 & _T_2; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_195 = _T_194 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_196 = _T_188 | _T_195; // @[ifu_compress_ctl.scala 25:115]
  wire  _T_200 = io_din[15] & io_din[14]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_201 = _T_200 & io_din[13]; // @[ifu_compress_ctl.scala 12:110]
  wire  out_12 = _T_196 | _T_201; // @[ifu_compress_ctl.scala 26:26]
  wire  _T_217 = _T_11 & _T_7; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_218 = _T_217 & _T_9; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_219 = _T_218 & _T_50; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_220 = _T_219 & _T_52; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_221 = _T_220 & _T_54; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_224 = _T_221 & _T_147; // @[ifu_compress_ctl.scala 28:53]
  wire  _T_228 = _T_2 & io_din[13]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_229 = _T_224 | _T_228; // @[ifu_compress_ctl.scala 28:67]
  wire  _T_234 = _T_200 & io_din[0]; // @[ifu_compress_ctl.scala 12:110]
  wire  out_6 = _T_229 | _T_234; // @[ifu_compress_ctl.scala 28:88]
  wire  _T_239 = io_din[15] & _T_147; // @[ifu_compress_ctl.scala 30:24]
  wire  _T_243 = io_din[15] & io_din[11]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_244 = _T_243 & io_din[10]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_245 = _T_239 | _T_244; // @[ifu_compress_ctl.scala 30:39]
  wire  _T_249 = io_din[13] & _T_42; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_250 = _T_245 | _T_249; // @[ifu_compress_ctl.scala 30:63]
  wire  _T_253 = io_din[13] & io_din[7]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_254 = _T_250 | _T_253; // @[ifu_compress_ctl.scala 30:83]
  wire  _T_257 = io_din[13] & io_din[9]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_258 = _T_254 | _T_257; // @[ifu_compress_ctl.scala 30:102]
  wire  _T_261 = io_din[13] & io_din[10]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_262 = _T_258 | _T_261; // @[ifu_compress_ctl.scala 31:22]
  wire  _T_265 = io_din[13] & io_din[11]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_266 = _T_262 | _T_265; // @[ifu_compress_ctl.scala 31:42]
  wire  _T_271 = _T_266 | _T_228; // @[ifu_compress_ctl.scala 31:62]
  wire  out_5 = _T_271 | _T_200; // @[ifu_compress_ctl.scala 31:83]
  wire  _T_288 = _T_2 & _T_23; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_289 = _T_288 & _T_38; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_290 = _T_289 & _T_40; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_291 = _T_290 & _T_42; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_292 = _T_291 & _T_44; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_295 = _T_292 & _T_147; // @[ifu_compress_ctl.scala 33:50]
  wire  _T_303 = _T_194 & _T_147; // @[ifu_compress_ctl.scala 33:87]
  wire  _T_304 = _T_295 | _T_303; // @[ifu_compress_ctl.scala 33:65]
  wire  _T_308 = _T_2 & io_din[6]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_311 = _T_308 & _T_147; // @[ifu_compress_ctl.scala 34:23]
  wire  _T_312 = _T_304 | _T_311; // @[ifu_compress_ctl.scala 33:102]
  wire  _T_317 = _T_190 & io_din[14]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_318 = _T_317 & io_din[0]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_319 = _T_312 | _T_318; // @[ifu_compress_ctl.scala 34:38]
  wire  _T_323 = _T_2 & io_din[5]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_326 = _T_323 & _T_147; // @[ifu_compress_ctl.scala 34:82]
  wire  _T_327 = _T_319 | _T_326; // @[ifu_compress_ctl.scala 34:62]
  wire  _T_331 = _T_2 & io_din[4]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_334 = _T_331 & _T_147; // @[ifu_compress_ctl.scala 35:23]
  wire  _T_335 = _T_327 | _T_334; // @[ifu_compress_ctl.scala 34:97]
  wire  _T_339 = _T_2 & io_din[3]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_342 = _T_339 & _T_147; // @[ifu_compress_ctl.scala 35:58]
  wire  _T_343 = _T_335 | _T_342; // @[ifu_compress_ctl.scala 35:38]
  wire  _T_347 = _T_2 & io_din[2]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_350 = _T_347 & _T_147; // @[ifu_compress_ctl.scala 35:93]
  wire  _T_351 = _T_343 | _T_350; // @[ifu_compress_ctl.scala 35:73]
  wire  _T_357 = _T_2 & _T_4; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_358 = _T_357 & io_din[0]; // @[ifu_compress_ctl.scala 12:110]
  wire  out_4 = _T_351 | _T_358; // @[ifu_compress_ctl.scala 35:108]
  wire  _T_380 = _T_56 & io_din[11]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_381 = _T_380 & _T_7; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_382 = _T_381 & _T_9; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_383 = _T_382 & _T_50; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_384 = _T_383 & _T_52; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_385 = _T_384 & _T_54; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_386 = _T_385 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_403 = _T_56 & io_din[10]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_404 = _T_403 & _T_7; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_405 = _T_404 & _T_9; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_406 = _T_405 & _T_50; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_407 = _T_406 & _T_52; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_408 = _T_407 & _T_54; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_409 = _T_408 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_410 = _T_386 | _T_409; // @[ifu_compress_ctl.scala 40:59]
  wire  _T_427 = _T_56 & io_din[9]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_428 = _T_427 & _T_7; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_429 = _T_428 & _T_9; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_430 = _T_429 & _T_50; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_431 = _T_430 & _T_52; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_432 = _T_431 & _T_54; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_433 = _T_432 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_434 = _T_410 | _T_433; // @[ifu_compress_ctl.scala 40:107]
  wire  _T_451 = _T_56 & io_din[8]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_452 = _T_451 & _T_7; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_453 = _T_452 & _T_9; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_454 = _T_453 & _T_50; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_455 = _T_454 & _T_52; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_456 = _T_455 & _T_54; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_457 = _T_456 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_458 = _T_434 | _T_457; // @[ifu_compress_ctl.scala 41:50]
  wire  _T_475 = _T_56 & io_din[7]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_476 = _T_475 & _T_7; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_477 = _T_476 & _T_9; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_478 = _T_477 & _T_50; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_479 = _T_478 & _T_52; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_480 = _T_479 & _T_54; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_481 = _T_480 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_482 = _T_458 | _T_481; // @[ifu_compress_ctl.scala 41:94]
  wire  _T_487 = ~io_din[12]; // @[ifu_compress_ctl.scala 12:83]
  wire  _T_499 = _T_11 & _T_487; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_500 = _T_499 & _T_7; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_501 = _T_500 & _T_9; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_502 = _T_501 & _T_50; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_503 = _T_502 & _T_52; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_504 = _T_503 & _T_54; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_507 = _T_504 & _T_147; // @[ifu_compress_ctl.scala 42:94]
  wire  _T_508 = _T_482 | _T_507; // @[ifu_compress_ctl.scala 42:49]
  wire  _T_514 = _T_190 & io_din[13]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_515 = _T_514 & _T_42; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_516 = _T_508 | _T_515; // @[ifu_compress_ctl.scala 42:109]
  wire  _T_522 = _T_514 & io_din[7]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_523 = _T_516 | _T_522; // @[ifu_compress_ctl.scala 43:26]
  wire  _T_529 = _T_514 & io_din[9]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_530 = _T_523 | _T_529; // @[ifu_compress_ctl.scala 43:48]
  wire  _T_536 = _T_514 & io_din[10]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_537 = _T_530 | _T_536; // @[ifu_compress_ctl.scala 43:70]
  wire  _T_543 = _T_514 & io_din[11]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_544 = _T_537 | _T_543; // @[ifu_compress_ctl.scala 43:93]
  wire  out_2 = _T_544 | _T_228; // @[ifu_compress_ctl.scala 44:26]
  wire [4:0] rs2d = io_din[6:2]; // @[ifu_compress_ctl.scala 50:20]
  wire [4:0] rdd = io_din[11:7]; // @[ifu_compress_ctl.scala 51:19]
  wire [4:0] rdpd = {2'h1,io_din[9:7]}; // @[Cat.scala 29:58]
  wire [4:0] rs2pd = {2'h1,io_din[4:2]}; // @[Cat.scala 29:58]
  wire  _T_557 = _T_308 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_564 = _T_317 & io_din[11]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_565 = _T_564 & io_din[0]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_566 = _T_557 | _T_565; // @[ifu_compress_ctl.scala 55:33]
  wire  _T_572 = _T_323 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_573 = _T_566 | _T_572; // @[ifu_compress_ctl.scala 55:58]
  wire  _T_580 = _T_317 & io_din[10]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_581 = _T_580 & io_din[0]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_582 = _T_573 | _T_581; // @[ifu_compress_ctl.scala 55:79]
  wire  _T_588 = _T_331 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_589 = _T_582 | _T_588; // @[ifu_compress_ctl.scala 55:104]
  wire  _T_596 = _T_317 & io_din[9]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_597 = _T_596 & io_din[0]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_598 = _T_589 | _T_597; // @[ifu_compress_ctl.scala 56:24]
  wire  _T_604 = _T_339 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_605 = _T_598 | _T_604; // @[ifu_compress_ctl.scala 56:48]
  wire  _T_613 = _T_317 & _T_42; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_614 = _T_613 & io_din[0]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_615 = _T_605 | _T_614; // @[ifu_compress_ctl.scala 56:69]
  wire  _T_621 = _T_347 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_622 = _T_615 | _T_621; // @[ifu_compress_ctl.scala 56:94]
  wire  _T_629 = _T_317 & io_din[7]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_630 = _T_629 & io_din[0]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_631 = _T_622 | _T_630; // @[ifu_compress_ctl.scala 57:22]
  wire  _T_635 = _T_190 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_636 = _T_631 | _T_635; // @[ifu_compress_ctl.scala 57:46]
  wire  _T_642 = _T_190 & _T_4; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_643 = _T_642 & io_din[0]; // @[ifu_compress_ctl.scala 12:110]
  wire  rdrd = _T_636 | _T_643; // @[ifu_compress_ctl.scala 57:65]
  wire  _T_651 = _T_380 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_659 = _T_403 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_660 = _T_651 | _T_659; // @[ifu_compress_ctl.scala 59:38]
  wire  _T_668 = _T_427 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_669 = _T_660 | _T_668; // @[ifu_compress_ctl.scala 59:63]
  wire  _T_677 = _T_451 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_678 = _T_669 | _T_677; // @[ifu_compress_ctl.scala 59:87]
  wire  _T_686 = _T_475 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_687 = _T_678 | _T_686; // @[ifu_compress_ctl.scala 60:27]
  wire  _T_703 = _T_2 & _T_487; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_704 = _T_703 & _T_7; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_705 = _T_704 & _T_9; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_706 = _T_705 & _T_50; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_707 = _T_706 & _T_52; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_708 = _T_707 & _T_54; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_709 = _T_708 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_710 = _T_687 | _T_709; // @[ifu_compress_ctl.scala 60:51]
  wire  _T_717 = _T_56 & io_din[6]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_718 = _T_717 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_719 = _T_710 | _T_718; // @[ifu_compress_ctl.scala 60:89]
  wire  _T_726 = _T_56 & io_din[5]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_727 = _T_726 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_728 = _T_719 | _T_727; // @[ifu_compress_ctl.scala 61:27]
  wire  _T_735 = _T_56 & io_din[4]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_736 = _T_735 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_737 = _T_728 | _T_736; // @[ifu_compress_ctl.scala 61:51]
  wire  _T_744 = _T_56 & io_din[3]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_745 = _T_744 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_746 = _T_737 | _T_745; // @[ifu_compress_ctl.scala 61:75]
  wire  _T_753 = _T_56 & io_din[2]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_754 = _T_753 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_755 = _T_746 | _T_754; // @[ifu_compress_ctl.scala 61:99]
  wire  _T_764 = _T_194 & _T_4; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_765 = _T_764 & io_din[0]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_766 = _T_755 | _T_765; // @[ifu_compress_ctl.scala 62:27]
  wire  rdrs1 = _T_766 | _T_195; // @[ifu_compress_ctl.scala 62:54]
  wire  _T_777 = io_din[15] & io_din[6]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_778 = _T_777 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_782 = io_din[15] & io_din[5]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_783 = _T_782 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_784 = _T_778 | _T_783; // @[ifu_compress_ctl.scala 64:34]
  wire  _T_788 = io_din[15] & io_din[4]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_789 = _T_788 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_790 = _T_784 | _T_789; // @[ifu_compress_ctl.scala 64:54]
  wire  _T_794 = io_din[15] & io_din[3]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_795 = _T_794 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_796 = _T_790 | _T_795; // @[ifu_compress_ctl.scala 64:74]
  wire  _T_800 = io_din[15] & io_din[2]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_801 = _T_800 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_802 = _T_796 | _T_801; // @[ifu_compress_ctl.scala 64:94]
  wire  _T_807 = _T_200 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  rs2rs2 = _T_802 | _T_807; // @[ifu_compress_ctl.scala 64:114]
  wire  rdprd = _T_12 & io_din[0]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_820 = io_din[15] & _T_4; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_821 = _T_820 & io_din[0]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_827 = _T_821 | _T_234; // @[ifu_compress_ctl.scala 68:36]
  wire  _T_830 = ~io_din[1]; // @[ifu_compress_ctl.scala 12:83]
  wire  _T_831 = io_din[14] & _T_830; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_834 = _T_831 & _T_147; // @[ifu_compress_ctl.scala 68:76]
  wire  rdprs1 = _T_827 | _T_834; // @[ifu_compress_ctl.scala 68:57]
  wire  _T_846 = _T_128 & io_din[10]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_847 = _T_846 & io_din[0]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_851 = io_din[15] & _T_830; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_854 = _T_851 & _T_147; // @[ifu_compress_ctl.scala 70:66]
  wire  rs2prs2 = _T_847 | _T_854; // @[ifu_compress_ctl.scala 70:47]
  wire  _T_859 = _T_190 & _T_830; // @[ifu_compress_ctl.scala 12:110]
  wire  rs2prd = _T_859 & _T_147; // @[ifu_compress_ctl.scala 72:33]
  wire  _T_866 = _T_2 & _T_830; // @[ifu_compress_ctl.scala 12:110]
  wire  uimm9_2 = _T_866 & _T_147; // @[ifu_compress_ctl.scala 74:34]
  wire  _T_875 = _T_317 & _T_830; // @[ifu_compress_ctl.scala 12:110]
  wire  ulwimm6_2 = _T_875 & _T_147; // @[ifu_compress_ctl.scala 76:39]
  wire  ulwspimm7_2 = _T_317 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_897 = _T_317 & io_din[13]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_898 = _T_897 & _T_23; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_899 = _T_898 & _T_38; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_900 = _T_899 & _T_40; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_901 = _T_900 & io_din[8]; // @[ifu_compress_ctl.scala 12:110]
  wire  rdeq2 = _T_901 & _T_44; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1027 = _T_194 & io_din[13]; // @[ifu_compress_ctl.scala 12:110]
  wire  rdeq1 = _T_482 | _T_1027; // @[ifu_compress_ctl.scala 84:42]
  wire  _T_1050 = io_din[14] & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1051 = rdeq2 | _T_1050; // @[ifu_compress_ctl.scala 86:53]
  wire  rs1eq2 = _T_1051 | uimm9_2; // @[ifu_compress_ctl.scala 86:71]
  wire  _T_1092 = _T_357 & io_din[11]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1093 = _T_1092 & _T_38; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1094 = _T_1093 & io_din[0]; // @[ifu_compress_ctl.scala 12:110]
  wire  simm5_0 = _T_1094 | _T_643; // @[ifu_compress_ctl.scala 92:45]
  wire  _T_1112 = _T_897 & io_din[7]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1121 = _T_897 & _T_42; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1122 = _T_1112 | _T_1121; // @[ifu_compress_ctl.scala 96:44]
  wire  _T_1130 = _T_897 & io_din[9]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1131 = _T_1122 | _T_1130; // @[ifu_compress_ctl.scala 96:70]
  wire  _T_1139 = _T_897 & io_din[10]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1140 = _T_1131 | _T_1139; // @[ifu_compress_ctl.scala 96:95]
  wire  _T_1148 = _T_897 & io_din[11]; // @[ifu_compress_ctl.scala 12:110]
  wire  sluimm17_12 = _T_1140 | _T_1148; // @[ifu_compress_ctl.scala 96:121]
  wire  uimm5_0 = _T_79 | _T_195; // @[ifu_compress_ctl.scala 98:45]
  wire [6:0] l1_6 = {out_6,out_5,out_4,_T_228,out_2,1'h1,1'h1}; // @[Cat.scala 29:58]
  wire [4:0] _T_1192 = rdrd ? rdd : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_1193 = rdprd ? rdpd : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_1194 = rs2prd ? rs2pd : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_1195 = rdeq1 ? 5'h1 : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_1196 = rdeq2 ? 5'h2 : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_1197 = _T_1192 | _T_1193; // @[Mux.scala 27:72]
  wire [4:0] _T_1198 = _T_1197 | _T_1194; // @[Mux.scala 27:72]
  wire [4:0] _T_1199 = _T_1198 | _T_1195; // @[Mux.scala 27:72]
  wire [4:0] l1_11 = _T_1199 | _T_1196; // @[Mux.scala 27:72]
  wire [4:0] _T_1210 = rdrs1 ? rdd : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_1211 = rdprs1 ? rdpd : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_1212 = rs1eq2 ? 5'h2 : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_1213 = _T_1210 | _T_1211; // @[Mux.scala 27:72]
  wire [4:0] l1_19 = _T_1213 | _T_1212; // @[Mux.scala 27:72]
  wire [4:0] _T_1219 = {3'h0,1'h0,out_20}; // @[Cat.scala 29:58]
  wire [4:0] _T_1222 = rs2rs2 ? rs2d : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_1223 = rs2prs2 ? rs2pd : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_1224 = _T_1222 | _T_1223; // @[Mux.scala 27:72]
  wire [4:0] l1_24 = _T_1219 | _T_1224; // @[ifu_compress_ctl.scala 114:67]
  wire [14:0] _T_1232 = {out_14,out_13,out_12,l1_11,l1_6}; // @[Cat.scala 29:58]
  wire [31:0] l1 = {1'h0,out_30,2'h0,3'h0,l1_24,l1_19,_T_1232}; // @[Cat.scala 29:58]
  wire [5:0] simm5d = {io_din[12],rs2d}; // @[Cat.scala 29:58]
  wire [5:0] simm9d = {io_din[12],io_din[4:3],io_din[5],io_din[2],io_din[6]}; // @[Cat.scala 29:58]
  wire [10:0] sjald_1 = {io_din[12],io_din[8],io_din[10:9],io_din[6],io_din[7],io_din[2],io_din[11],io_din[5:4],io_din[3]}; // @[Cat.scala 29:58]
  wire [19:0] sjald = {io_din[12],io_din[12],io_din[12],io_din[12],io_din[12],io_din[12],io_din[12],io_din[12],io_din[12],sjald_1}; // @[Cat.scala 29:58]
  wire [9:0] _T_1296 = {io_din[12],io_din[12],io_din[12],io_din[12],io_din[12],io_din[12],io_din[12],io_din[12],io_din[12],io_din[12]}; // @[Cat.scala 29:58]
  wire [19:0] sluimmd = {_T_1296,io_din[12],io_din[12],io_din[12],io_din[12],io_din[12],rs2d}; // @[Cat.scala 29:58]
  wire [11:0] _T_1314 = {simm5d[5],simm5d[5],simm5d[5],simm5d[5],simm5d[5],simm5d[5],simm5d[5],simm5d[4:0]}; // @[Cat.scala 29:58]
  wire [11:0] _T_1317 = {2'h0,io_din[10:7],io_din[12:11],io_din[5],io_din[6],2'h0}; // @[Cat.scala 29:58]
  wire [11:0] _T_1325 = {simm9d[5],simm9d[5],simm9d[5],simm9d[4:0],4'h0}; // @[Cat.scala 29:58]
  wire [11:0] _T_1328 = {5'h0,io_din[5],io_din[12:10],io_din[6],2'h0}; // @[Cat.scala 29:58]
  wire [11:0] _T_1331 = {4'h0,io_din[3:2],io_din[12],io_din[6:4],2'h0}; // @[Cat.scala 29:58]
  wire [11:0] _T_1333 = {6'h0,io_din[12],rs2d}; // @[Cat.scala 29:58]
  wire [11:0] _T_1339 = {sjald[19],sjald[9:0],sjald[10]}; // @[Cat.scala 29:58]
  wire [11:0] _T_1342 = simm5_0 ? _T_1314 : 12'h0; // @[Mux.scala 27:72]
  wire [11:0] _T_1343 = uimm9_2 ? _T_1317 : 12'h0; // @[Mux.scala 27:72]
  wire [11:0] _T_1344 = rdeq2 ? _T_1325 : 12'h0; // @[Mux.scala 27:72]
  wire [11:0] _T_1345 = ulwimm6_2 ? _T_1328 : 12'h0; // @[Mux.scala 27:72]
  wire [11:0] _T_1346 = ulwspimm7_2 ? _T_1331 : 12'h0; // @[Mux.scala 27:72]
  wire [11:0] _T_1347 = uimm5_0 ? _T_1333 : 12'h0; // @[Mux.scala 27:72]
  wire [11:0] _T_1348 = _T_228 ? _T_1339 : 12'h0; // @[Mux.scala 27:72]
  wire [11:0] _T_1349 = sluimm17_12 ? sluimmd[19:8] : 12'h0; // @[Mux.scala 27:72]
  wire [11:0] _T_1350 = _T_1342 | _T_1343; // @[Mux.scala 27:72]
  wire [11:0] _T_1351 = _T_1350 | _T_1344; // @[Mux.scala 27:72]
  wire [11:0] _T_1352 = _T_1351 | _T_1345; // @[Mux.scala 27:72]
  wire [11:0] _T_1353 = _T_1352 | _T_1346; // @[Mux.scala 27:72]
  wire [11:0] _T_1354 = _T_1353 | _T_1347; // @[Mux.scala 27:72]
  wire [11:0] _T_1355 = _T_1354 | _T_1348; // @[Mux.scala 27:72]
  wire [11:0] _T_1356 = _T_1355 | _T_1349; // @[Mux.scala 27:72]
  wire [11:0] l2_31 = l1[31:20] | _T_1356; // @[ifu_compress_ctl.scala 133:25]
  wire [7:0] _T_1363 = _T_228 ? sjald[19:12] : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_1364 = sluimm17_12 ? sluimmd[7:0] : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_1365 = _T_1363 | _T_1364; // @[Mux.scala 27:72]
  wire [7:0] l2_19 = l1[19:12] | _T_1365; // @[ifu_compress_ctl.scala 143:25]
  wire [31:0] l2 = {l2_31,l2_19,l1[11:0]}; // @[Cat.scala 29:58]
  wire [8:0] sbr8d = {io_din[12],io_din[6],io_din[5],io_din[2],io_din[11],io_din[10],io_din[4],io_din[3],1'h0}; // @[Cat.scala 29:58]
  wire [6:0] uswimm6d = {io_din[5],io_din[12:10],io_din[6],2'h0}; // @[Cat.scala 29:58]
  wire [7:0] uswspimm7d = {io_din[8:7],io_din[12:9],2'h0}; // @[Cat.scala 29:58]
  wire [6:0] _T_1400 = {sbr8d[8],sbr8d[8],sbr8d[8],sbr8d[8],sbr8d[7:5]}; // @[Cat.scala 29:58]
  wire [6:0] _T_1403 = {5'h0,uswimm6d[6:5]}; // @[Cat.scala 29:58]
  wire [6:0] _T_1406 = {4'h0,uswspimm7d[7:5]}; // @[Cat.scala 29:58]
  wire [6:0] _T_1407 = _T_234 ? _T_1400 : 7'h0; // @[Mux.scala 27:72]
  wire [6:0] _T_1408 = _T_854 ? _T_1403 : 7'h0; // @[Mux.scala 27:72]
  wire [6:0] _T_1409 = _T_807 ? _T_1406 : 7'h0; // @[Mux.scala 27:72]
  wire [6:0] _T_1410 = _T_1407 | _T_1408; // @[Mux.scala 27:72]
  wire [6:0] _T_1411 = _T_1410 | _T_1409; // @[Mux.scala 27:72]
  wire [6:0] l3_31 = l2[31:25] | _T_1411; // @[ifu_compress_ctl.scala 151:25]
  wire [12:0] l3_24 = l2[24:12]; // @[ifu_compress_ctl.scala 154:17]
  wire [4:0] _T_1417 = {sbr8d[4:1],sbr8d[8]}; // @[Cat.scala 29:58]
  wire [4:0] _T_1422 = _T_234 ? _T_1417 : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_1423 = _T_854 ? uswimm6d[4:0] : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_1424 = _T_807 ? uswspimm7d[4:0] : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_1425 = _T_1422 | _T_1423; // @[Mux.scala 27:72]
  wire [4:0] _T_1426 = _T_1425 | _T_1424; // @[Mux.scala 27:72]
  wire [4:0] l3_11 = l2[11:7] | _T_1426; // @[ifu_compress_ctl.scala 156:24]
  wire [31:0] l3 = {l3_31,l3_24,l3_11,l2[6:0]}; // @[Cat.scala 29:58]
  wire  _T_1437 = _T_4 & _T_487; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1438 = _T_1437 & io_din[11]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1439 = _T_1438 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1442 = _T_1439 & _T_147; // @[ifu_compress_ctl.scala 162:39]
  wire  _T_1450 = _T_1437 & io_din[6]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1451 = _T_1450 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1454 = _T_1451 & _T_147; // @[ifu_compress_ctl.scala 162:79]
  wire  _T_1455 = _T_1442 | _T_1454; // @[ifu_compress_ctl.scala 162:54]
  wire  _T_1464 = _T_642 & io_din[11]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1465 = _T_1464 & _T_830; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1466 = _T_1455 | _T_1465; // @[ifu_compress_ctl.scala 162:94]
  wire  _T_1474 = _T_1437 & io_din[5]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1475 = _T_1474 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1478 = _T_1475 & _T_147; // @[ifu_compress_ctl.scala 163:55]
  wire  _T_1479 = _T_1466 | _T_1478; // @[ifu_compress_ctl.scala 163:30]
  wire  _T_1487 = _T_1437 & io_din[10]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1488 = _T_1487 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1491 = _T_1488 & _T_147; // @[ifu_compress_ctl.scala 163:96]
  wire  _T_1492 = _T_1479 | _T_1491; // @[ifu_compress_ctl.scala 163:70]
  wire  _T_1501 = _T_642 & io_din[6]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1502 = _T_1501 & _T_830; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1503 = _T_1492 | _T_1502; // @[ifu_compress_ctl.scala 163:111]
  wire  _T_1510 = io_din[15] & _T_487; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1511 = _T_1510 & _T_830; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1512 = _T_1511 & io_din[0]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1513 = _T_1503 | _T_1512; // @[ifu_compress_ctl.scala 164:29]
  wire  _T_1521 = _T_1437 & io_din[9]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1522 = _T_1521 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1525 = _T_1522 & _T_147; // @[ifu_compress_ctl.scala 164:79]
  wire  _T_1526 = _T_1513 | _T_1525; // @[ifu_compress_ctl.scala 164:54]
  wire  _T_1533 = _T_487 & io_din[6]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1534 = _T_1533 & _T_830; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1535 = _T_1534 & io_din[0]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1536 = _T_1526 | _T_1535; // @[ifu_compress_ctl.scala 164:94]
  wire  _T_1545 = _T_642 & io_din[5]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1546 = _T_1545 & _T_830; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1547 = _T_1536 | _T_1546; // @[ifu_compress_ctl.scala 164:118]
  wire  _T_1555 = _T_1437 & io_din[8]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1556 = _T_1555 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1559 = _T_1556 & _T_147; // @[ifu_compress_ctl.scala 165:28]
  wire  _T_1560 = _T_1547 | _T_1559; // @[ifu_compress_ctl.scala 164:144]
  wire  _T_1567 = _T_487 & io_din[5]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1568 = _T_1567 & _T_830; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1569 = _T_1568 & io_din[0]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1570 = _T_1560 | _T_1569; // @[ifu_compress_ctl.scala 165:43]
  wire  _T_1579 = _T_642 & io_din[10]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1580 = _T_1579 & _T_830; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1581 = _T_1570 | _T_1580; // @[ifu_compress_ctl.scala 165:67]
  wire  _T_1589 = _T_1437 & io_din[7]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1590 = _T_1589 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1593 = _T_1590 & _T_147; // @[ifu_compress_ctl.scala 166:28]
  wire  _T_1594 = _T_1581 | _T_1593; // @[ifu_compress_ctl.scala 165:94]
  wire  _T_1602 = io_din[12] & io_din[11]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1603 = _T_1602 & _T_38; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1604 = _T_1603 & _T_830; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1605 = _T_1604 & io_din[0]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1606 = _T_1594 | _T_1605; // @[ifu_compress_ctl.scala 166:43]
  wire  _T_1615 = _T_642 & io_din[9]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1616 = _T_1615 & _T_830; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1617 = _T_1606 | _T_1616; // @[ifu_compress_ctl.scala 166:71]
  wire  _T_1625 = _T_1437 & io_din[4]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1626 = _T_1625 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1629 = _T_1626 & _T_147; // @[ifu_compress_ctl.scala 167:28]
  wire  _T_1630 = _T_1617 | _T_1629; // @[ifu_compress_ctl.scala 166:97]
  wire  _T_1636 = io_din[13] & io_din[12]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1637 = _T_1636 & _T_830; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1638 = _T_1637 & io_din[0]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1639 = _T_1630 | _T_1638; // @[ifu_compress_ctl.scala 167:43]
  wire  _T_1648 = _T_642 & io_din[8]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1649 = _T_1648 & _T_830; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1650 = _T_1639 | _T_1649; // @[ifu_compress_ctl.scala 167:67]
  wire  _T_1658 = _T_1437 & io_din[3]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1659 = _T_1658 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1662 = _T_1659 & _T_147; // @[ifu_compress_ctl.scala 168:28]
  wire  _T_1663 = _T_1650 | _T_1662; // @[ifu_compress_ctl.scala 167:93]
  wire  _T_1669 = io_din[13] & io_din[4]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1670 = _T_1669 & _T_830; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1671 = _T_1670 & io_din[0]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1672 = _T_1663 | _T_1671; // @[ifu_compress_ctl.scala 168:43]
  wire  _T_1680 = _T_1437 & io_din[2]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1681 = _T_1680 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1684 = _T_1681 & _T_147; // @[ifu_compress_ctl.scala 168:91]
  wire  _T_1685 = _T_1672 | _T_1684; // @[ifu_compress_ctl.scala 168:66]
  wire  _T_1694 = _T_642 & io_din[7]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1695 = _T_1694 & _T_830; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1696 = _T_1685 | _T_1695; // @[ifu_compress_ctl.scala 168:106]
  wire  _T_1702 = io_din[13] & io_din[3]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1703 = _T_1702 & _T_830; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1704 = _T_1703 & io_din[0]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1705 = _T_1696 | _T_1704; // @[ifu_compress_ctl.scala 169:29]
  wire  _T_1711 = io_din[13] & io_din[2]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1712 = _T_1711 & _T_830; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1713 = _T_1712 & io_din[0]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1714 = _T_1705 | _T_1713; // @[ifu_compress_ctl.scala 169:52]
  wire  _T_1720 = io_din[14] & _T_4; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1721 = _T_1720 & _T_830; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1722 = _T_1714 | _T_1721; // @[ifu_compress_ctl.scala 169:75]
  wire  _T_1731 = _T_703 & _T_830; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1732 = _T_1731 & io_din[0]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1733 = _T_1722 | _T_1732; // @[ifu_compress_ctl.scala 169:98]
  wire  _T_1740 = _T_820 & io_din[12]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1741 = _T_1740 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1744 = _T_1741 & _T_147; // @[ifu_compress_ctl.scala 170:54]
  wire  _T_1745 = _T_1733 | _T_1744; // @[ifu_compress_ctl.scala 170:29]
  wire  _T_1754 = _T_642 & _T_487; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1755 = _T_1754 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1758 = _T_1755 & _T_147; // @[ifu_compress_ctl.scala 170:96]
  wire  _T_1759 = _T_1745 | _T_1758; // @[ifu_compress_ctl.scala 170:69]
  wire  _T_1768 = _T_642 & io_din[12]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1769 = _T_1768 & _T_830; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1770 = _T_1759 | _T_1769; // @[ifu_compress_ctl.scala 170:111]
  wire  _T_1777 = _T_1720 & _T_147; // @[ifu_compress_ctl.scala 171:50]
  wire  legal = _T_1770 | _T_1777; // @[ifu_compress_ctl.scala 171:30]
  wire [9:0] _T_1787 = {legal,legal,legal,legal,legal,legal,legal,legal,legal,legal}; // @[Cat.scala 29:58]
  wire [18:0] _T_1796 = {_T_1787,legal,legal,legal,legal,legal,legal,legal,legal,legal}; // @[Cat.scala 29:58]
  wire [27:0] _T_1805 = {_T_1796,legal,legal,legal,legal,legal,legal,legal,legal,legal}; // @[Cat.scala 29:58]
  wire [31:0] _T_1809 = {_T_1805,legal,legal,legal,legal}; // @[Cat.scala 29:58]
  assign io_dout = l3 & _T_1809; // @[ifu_compress_ctl.scala 173:10]
endmodule
module ifu_aln_ctl(
  input         clock,
  input         reset,
  input         io_scan_mode,
  input         io_active_clk,
  input         io_ifu_async_error_start,
  input         io_iccm_rd_ecc_double_err,
  input         io_ic_access_fault_f,
  input  [1:0]  io_ic_access_fault_type_f,
  input  [7:0]  io_ifu_bp_fghr_f,
  input  [30:0] io_ifu_bp_btb_target_f,
  input  [11:0] io_ifu_bp_poffset_f,
  input  [1:0]  io_ifu_bp_hist0_f,
  input  [1:0]  io_ifu_bp_hist1_f,
  input  [1:0]  io_ifu_bp_pc4_f,
  input  [1:0]  io_ifu_bp_way_f,
  input  [1:0]  io_ifu_bp_valid_f,
  input  [1:0]  io_ifu_bp_ret_f,
  input         io_exu_flush_final,
  input         io_dec_aln_aln_dec_dec_i0_decode_d,
  output [15:0] io_dec_aln_aln_dec_ifu_i0_cinst,
  output        io_dec_aln_aln_ib_ifu_i0_icaf,
  output [1:0]  io_dec_aln_aln_ib_ifu_i0_icaf_type,
  output        io_dec_aln_aln_ib_ifu_i0_icaf_f1,
  output        io_dec_aln_aln_ib_ifu_i0_dbecc,
  output [7:0]  io_dec_aln_aln_ib_ifu_i0_bp_index,
  output [7:0]  io_dec_aln_aln_ib_ifu_i0_bp_fghr,
  output [4:0]  io_dec_aln_aln_ib_ifu_i0_bp_btag,
  output        io_dec_aln_aln_ib_ifu_i0_valid,
  output [31:0] io_dec_aln_aln_ib_ifu_i0_instr,
  output [30:0] io_dec_aln_aln_ib_ifu_i0_pc,
  output        io_dec_aln_aln_ib_ifu_i0_pc4,
  output        io_dec_aln_aln_ib_i0_brp_valid,
  output [11:0] io_dec_aln_aln_ib_i0_brp_bits_toffset,
  output [1:0]  io_dec_aln_aln_ib_i0_brp_bits_hist,
  output        io_dec_aln_aln_ib_i0_brp_bits_br_error,
  output        io_dec_aln_aln_ib_i0_brp_bits_br_start_error,
  output [30:0] io_dec_aln_aln_ib_i0_brp_bits_prett,
  output        io_dec_aln_aln_ib_i0_brp_bits_way,
  output        io_dec_aln_aln_ib_i0_brp_bits_ret,
  output        io_dec_aln_ifu_pmu_instr_aligned,
  input  [31:0] io_ifu_fetch_data_f,
  input  [1:0]  io_ifu_fetch_val,
  input  [30:0] io_ifu_fetch_pc,
  output        io_ifu_fb_consume1,
  output        io_ifu_fb_consume2
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
`endif // RANDOMIZE_REG_INIT
  wire  rvclkhdr_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_1_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_1_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_1_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_1_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_2_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_2_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_2_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_2_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_3_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_3_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_3_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_3_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_4_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_4_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_4_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_4_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_5_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_5_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_5_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_5_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_6_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_6_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_6_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_6_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_7_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_7_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_7_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_7_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_8_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_8_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_8_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_8_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_9_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_9_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_9_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_9_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_10_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_10_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_10_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_10_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_11_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_11_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_11_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_11_io_scan_mode; // @[lib.scala 368:23]
  wire [15:0] decompressed_io_din; // @[ifu_aln_ctl.scala 352:28]
  wire [31:0] decompressed_io_dout; // @[ifu_aln_ctl.scala 352:28]
  reg  error_stall; // @[ifu_aln_ctl.scala 102:51]
  wire  _T = error_stall | io_ifu_async_error_start; // @[ifu_aln_ctl.scala 99:34]
  wire  _T_1 = ~io_exu_flush_final; // @[ifu_aln_ctl.scala 99:64]
  reg [1:0] wrptr; // @[ifu_aln_ctl.scala 104:48]
  reg [1:0] rdptr; // @[ifu_aln_ctl.scala 106:48]
  reg [1:0] f2val; // @[ifu_aln_ctl.scala 108:48]
  reg [1:0] f1val; // @[ifu_aln_ctl.scala 109:48]
  reg [1:0] f0val; // @[ifu_aln_ctl.scala 110:48]
  reg  q2off; // @[ifu_aln_ctl.scala 112:48]
  reg  q1off; // @[ifu_aln_ctl.scala 113:48]
  reg  q0off; // @[ifu_aln_ctl.scala 114:48]
  wire  _T_785 = ~error_stall; // @[ifu_aln_ctl.scala 395:55]
  wire  i0_shift = io_dec_aln_aln_dec_dec_i0_decode_d & _T_785; // @[ifu_aln_ctl.scala 395:53]
  wire  _T_186 = rdptr == 2'h0; // @[ifu_aln_ctl.scala 169:31]
  wire  _T_189 = _T_186 & q0off; // @[Mux.scala 27:72]
  wire  _T_187 = rdptr == 2'h1; // @[ifu_aln_ctl.scala 170:11]
  wire  _T_190 = _T_187 & q1off; // @[Mux.scala 27:72]
  wire  _T_192 = _T_189 | _T_190; // @[Mux.scala 27:72]
  wire  _T_188 = rdptr == 2'h2; // @[ifu_aln_ctl.scala 171:11]
  wire  _T_191 = _T_188 & q2off; // @[Mux.scala 27:72]
  wire  q0ptr = _T_192 | _T_191; // @[Mux.scala 27:72]
  wire  _T_202 = ~q0ptr; // @[ifu_aln_ctl.scala 175:26]
  wire [1:0] q0sel = {q0ptr,_T_202}; // @[Cat.scala 29:58]
  wire [2:0] qren = {_T_188,_T_187,_T_186}; // @[Cat.scala 29:58]
  reg [31:0] q1; // @[lib.scala 374:16]
  reg [31:0] q0; // @[lib.scala 374:16]
  wire [63:0] _T_479 = {q1,q0}; // @[Cat.scala 29:58]
  wire [63:0] _T_486 = qren[0] ? _T_479 : 64'h0; // @[Mux.scala 27:72]
  reg [31:0] q2; // @[lib.scala 374:16]
  wire [63:0] _T_482 = {q2,q1}; // @[Cat.scala 29:58]
  wire [63:0] _T_487 = qren[1] ? _T_482 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_489 = _T_486 | _T_487; // @[Mux.scala 27:72]
  wire [63:0] _T_485 = {q0,q2}; // @[Cat.scala 29:58]
  wire [63:0] _T_488 = qren[2] ? _T_485 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] qeff = _T_489 | _T_488; // @[Mux.scala 27:72]
  wire [31:0] q0eff = qeff[31:0]; // @[ifu_aln_ctl.scala 294:42]
  wire [31:0] _T_496 = q0sel[0] ? q0eff : 32'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_497 = q0sel[1] ? q0eff[31:16] : 16'h0; // @[Mux.scala 27:72]
  wire [31:0] _GEN_0 = {{16'd0}, _T_497}; // @[Mux.scala 27:72]
  wire [31:0] q0final = _T_496 | _GEN_0; // @[Mux.scala 27:72]
  wire [31:0] _T_520 = f0val[1] ? q0final : 32'h0; // @[Mux.scala 27:72]
  wire  _T_513 = ~f0val[1]; // @[ifu_aln_ctl.scala 301:58]
  wire  _T_515 = _T_513 & f0val[0]; // @[ifu_aln_ctl.scala 301:68]
  wire  _T_197 = _T_186 & q1off; // @[Mux.scala 27:72]
  wire  _T_198 = _T_187 & q2off; // @[Mux.scala 27:72]
  wire  _T_200 = _T_197 | _T_198; // @[Mux.scala 27:72]
  wire  _T_199 = _T_188 & q0off; // @[Mux.scala 27:72]
  wire  q1ptr = _T_200 | _T_199; // @[Mux.scala 27:72]
  wire  _T_203 = ~q1ptr; // @[ifu_aln_ctl.scala 177:26]
  wire [1:0] q1sel = {q1ptr,_T_203}; // @[Cat.scala 29:58]
  wire [31:0] q1eff = qeff[63:32]; // @[ifu_aln_ctl.scala 294:29]
  wire [15:0] _T_506 = q1sel[0] ? q1eff[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_507 = q1sel[1] ? q1eff[31:16] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] q1final = _T_506 | _T_507; // @[Mux.scala 27:72]
  wire [31:0] _T_519 = {q1final,q0final[15:0]}; // @[Cat.scala 29:58]
  wire [31:0] _T_521 = _T_515 ? _T_519 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] aligndata = _T_520 | _T_521; // @[Mux.scala 27:72]
  wire  first4B = aligndata[1:0] == 2'h3; // @[ifu_aln_ctl.scala 334:29]
  wire  first2B = ~first4B; // @[ifu_aln_ctl.scala 336:17]
  wire  shift_2B = i0_shift & first2B; // @[ifu_aln_ctl.scala 399:24]
  wire [1:0] _T_443 = {1'h0,f0val[1]}; // @[Cat.scala 29:58]
  wire [1:0] _T_448 = shift_2B ? _T_443 : 2'h0; // @[Mux.scala 27:72]
  wire  _T_444 = ~shift_2B; // @[ifu_aln_ctl.scala 284:18]
  wire  shift_4B = i0_shift & first4B; // @[ifu_aln_ctl.scala 400:24]
  wire  _T_445 = ~shift_4B; // @[ifu_aln_ctl.scala 284:30]
  wire  _T_446 = _T_444 & _T_445; // @[ifu_aln_ctl.scala 284:28]
  wire [1:0] _T_449 = _T_446 ? f0val : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] sf0val = _T_448 | _T_449; // @[Mux.scala 27:72]
  wire  sf0_valid = sf0val[0]; // @[ifu_aln_ctl.scala 235:22]
  wire  _T_351 = ~sf0_valid; // @[ifu_aln_ctl.scala 256:26]
  wire  _T_802 = f0val[0] & _T_513; // @[ifu_aln_ctl.scala 403:28]
  wire  f1_shift_2B = _T_802 & shift_4B; // @[ifu_aln_ctl.scala 403:40]
  wire  _T_417 = f1_shift_2B & f1val[1]; // @[Mux.scala 27:72]
  wire  _T_416 = ~f1_shift_2B; // @[ifu_aln_ctl.scala 277:53]
  wire [1:0] _T_418 = _T_416 ? f1val : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _GEN_1 = {{1'd0}, _T_417}; // @[Mux.scala 27:72]
  wire [1:0] sf1val = _GEN_1 | _T_418; // @[Mux.scala 27:72]
  wire  sf1_valid = sf1val[0]; // @[ifu_aln_ctl.scala 234:22]
  wire  _T_352 = _T_351 & sf1_valid; // @[ifu_aln_ctl.scala 256:37]
  wire  f2_valid = f2val[0]; // @[ifu_aln_ctl.scala 233:20]
  wire  _T_353 = _T_352 & f2_valid; // @[ifu_aln_ctl.scala 256:50]
  wire  ifvalid = io_ifu_fetch_val[0]; // @[ifu_aln_ctl.scala 244:30]
  wire  _T_354 = _T_353 & ifvalid; // @[ifu_aln_ctl.scala 256:62]
  wire  _T_355 = sf0_valid & sf1_valid; // @[ifu_aln_ctl.scala 257:37]
  wire  _T_356 = ~f2_valid; // @[ifu_aln_ctl.scala 257:52]
  wire  _T_357 = _T_355 & _T_356; // @[ifu_aln_ctl.scala 257:50]
  wire  _T_358 = _T_357 & ifvalid; // @[ifu_aln_ctl.scala 257:62]
  wire  fetch_to_f2 = _T_354 | _T_358; // @[ifu_aln_ctl.scala 256:74]
  reg [30:0] f2pc; // @[lib.scala 374:16]
  wire  _T_335 = ~sf1_valid; // @[ifu_aln_ctl.scala 252:39]
  wire  _T_336 = _T_351 & _T_335; // @[ifu_aln_ctl.scala 252:37]
  wire  _T_337 = _T_336 & f2_valid; // @[ifu_aln_ctl.scala 252:50]
  wire  _T_338 = _T_337 & ifvalid; // @[ifu_aln_ctl.scala 252:62]
  wire  _T_342 = _T_352 & _T_356; // @[ifu_aln_ctl.scala 253:50]
  wire  _T_343 = _T_342 & ifvalid; // @[ifu_aln_ctl.scala 253:62]
  wire  _T_344 = _T_338 | _T_343; // @[ifu_aln_ctl.scala 252:74]
  wire  _T_346 = sf0_valid & _T_335; // @[ifu_aln_ctl.scala 254:37]
  wire  _T_348 = _T_346 & _T_356; // @[ifu_aln_ctl.scala 254:50]
  wire  _T_349 = _T_348 & ifvalid; // @[ifu_aln_ctl.scala 254:62]
  wire  fetch_to_f1 = _T_344 | _T_349; // @[ifu_aln_ctl.scala 253:74]
  wire  _T_25 = fetch_to_f1 | _T_353; // @[ifu_aln_ctl.scala 134:33]
  reg [30:0] f1pc; // @[lib.scala 374:16]
  wire  _T_332 = _T_336 & _T_356; // @[ifu_aln_ctl.scala 251:50]
  wire  fetch_to_f0 = _T_332 & ifvalid; // @[ifu_aln_ctl.scala 251:62]
  wire  _T_27 = fetch_to_f0 | _T_337; // @[ifu_aln_ctl.scala 135:33]
  wire  _T_28 = _T_27 | _T_352; // @[ifu_aln_ctl.scala 135:47]
  wire  _T_29 = _T_28 | shift_2B; // @[ifu_aln_ctl.scala 135:61]
  reg [30:0] f0pc; // @[lib.scala 374:16]
  wire  _T_35 = wrptr == 2'h2; // @[ifu_aln_ctl.scala 139:21]
  wire  _T_36 = _T_35 & ifvalid; // @[ifu_aln_ctl.scala 139:29]
  wire  _T_37 = wrptr == 2'h1; // @[ifu_aln_ctl.scala 139:46]
  wire  _T_38 = _T_37 & ifvalid; // @[ifu_aln_ctl.scala 139:54]
  wire  _T_39 = wrptr == 2'h0; // @[ifu_aln_ctl.scala 139:71]
  wire  _T_40 = _T_39 & ifvalid; // @[ifu_aln_ctl.scala 139:79]
  wire [2:0] qwen = {_T_36,_T_38,_T_40}; // @[Cat.scala 29:58]
  reg [11:0] brdata2; // @[lib.scala 374:16]
  reg [11:0] brdata1; // @[lib.scala 374:16]
  reg [11:0] brdata0; // @[lib.scala 374:16]
  reg [54:0] misc2; // @[lib.scala 374:16]
  reg [54:0] misc1; // @[lib.scala 374:16]
  reg [54:0] misc0; // @[lib.scala 374:16]
  wire  _T_44 = qren[0] & io_ifu_fb_consume1; // @[ifu_aln_ctl.scala 143:34]
  wire  _T_46 = _T_44 & _T_1; // @[ifu_aln_ctl.scala 143:55]
  wire  _T_49 = qren[1] & io_ifu_fb_consume1; // @[ifu_aln_ctl.scala 144:14]
  wire  _T_51 = _T_49 & _T_1; // @[ifu_aln_ctl.scala 144:35]
  wire  _T_59 = qren[0] & io_ifu_fb_consume2; // @[ifu_aln_ctl.scala 146:14]
  wire  _T_61 = _T_59 & _T_1; // @[ifu_aln_ctl.scala 146:35]
  wire  _T_69 = qren[2] & io_ifu_fb_consume2; // @[ifu_aln_ctl.scala 148:14]
  wire  _T_71 = _T_69 & _T_1; // @[ifu_aln_ctl.scala 148:35]
  wire  _T_73 = ~io_ifu_fb_consume1; // @[ifu_aln_ctl.scala 149:6]
  wire  _T_74 = ~io_ifu_fb_consume2; // @[ifu_aln_ctl.scala 149:28]
  wire  _T_75 = _T_73 & _T_74; // @[ifu_aln_ctl.scala 149:26]
  wire  _T_77 = _T_75 & _T_1; // @[ifu_aln_ctl.scala 149:48]
  wire [1:0] _T_80 = _T_51 ? 2'h2 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_82 = _T_61 ? 2'h2 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_85 = _T_77 ? rdptr : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _GEN_2 = {{1'd0}, _T_46}; // @[Mux.scala 27:72]
  wire [1:0] _T_86 = _GEN_2 | _T_80; // @[Mux.scala 27:72]
  wire [1:0] _T_88 = _T_86 | _T_82; // @[Mux.scala 27:72]
  wire [1:0] _GEN_3 = {{1'd0}, _T_71}; // @[Mux.scala 27:72]
  wire [1:0] _T_90 = _T_88 | _GEN_3; // @[Mux.scala 27:72]
  wire  _T_95 = qwen[0] & _T_1; // @[ifu_aln_ctl.scala 152:34]
  wire  _T_99 = qwen[1] & _T_1; // @[ifu_aln_ctl.scala 153:14]
  wire  _T_105 = ~ifvalid; // @[ifu_aln_ctl.scala 155:6]
  wire  _T_107 = _T_105 & _T_1; // @[ifu_aln_ctl.scala 155:15]
  wire [1:0] _T_110 = _T_99 ? 2'h2 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_112 = _T_107 ? wrptr : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _GEN_4 = {{1'd0}, _T_95}; // @[Mux.scala 27:72]
  wire [1:0] _T_113 = _GEN_4 | _T_110; // @[Mux.scala 27:72]
  wire  _T_118 = ~qwen[2]; // @[ifu_aln_ctl.scala 157:26]
  wire  _T_120 = _T_118 & _T_188; // @[ifu_aln_ctl.scala 157:35]
  wire  _T_795 = shift_2B & f0val[0]; // @[Mux.scala 27:72]
  wire  _T_796 = shift_4B & _T_802; // @[Mux.scala 27:72]
  wire  f0_shift_2B = _T_795 | _T_796; // @[Mux.scala 27:72]
  wire  _T_122 = q2off | f0_shift_2B; // @[ifu_aln_ctl.scala 157:74]
  wire  _T_126 = _T_118 & _T_187; // @[ifu_aln_ctl.scala 158:15]
  wire  _T_128 = q2off | f1_shift_2B; // @[ifu_aln_ctl.scala 158:54]
  wire  _T_132 = _T_118 & _T_186; // @[ifu_aln_ctl.scala 159:15]
  wire  _T_134 = _T_120 & _T_122; // @[Mux.scala 27:72]
  wire  _T_135 = _T_126 & _T_128; // @[Mux.scala 27:72]
  wire  _T_136 = _T_132 & q2off; // @[Mux.scala 27:72]
  wire  _T_137 = _T_134 | _T_135; // @[Mux.scala 27:72]
  wire  _T_141 = ~qwen[1]; // @[ifu_aln_ctl.scala 161:26]
  wire  _T_143 = _T_141 & _T_187; // @[ifu_aln_ctl.scala 161:35]
  wire  _T_145 = q1off | f0_shift_2B; // @[ifu_aln_ctl.scala 161:74]
  wire  _T_149 = _T_141 & _T_186; // @[ifu_aln_ctl.scala 162:15]
  wire  _T_151 = q1off | f1_shift_2B; // @[ifu_aln_ctl.scala 162:54]
  wire  _T_155 = _T_141 & _T_188; // @[ifu_aln_ctl.scala 163:15]
  wire  _T_157 = _T_143 & _T_145; // @[Mux.scala 27:72]
  wire  _T_158 = _T_149 & _T_151; // @[Mux.scala 27:72]
  wire  _T_159 = _T_155 & q1off; // @[Mux.scala 27:72]
  wire  _T_160 = _T_157 | _T_158; // @[Mux.scala 27:72]
  wire  _T_164 = ~qwen[0]; // @[ifu_aln_ctl.scala 165:26]
  wire  _T_166 = _T_164 & _T_186; // @[ifu_aln_ctl.scala 165:35]
  wire  _T_168 = q0off | f0_shift_2B; // @[ifu_aln_ctl.scala 165:76]
  wire  _T_172 = _T_164 & _T_188; // @[ifu_aln_ctl.scala 166:35]
  wire  _T_174 = q0off | f1_shift_2B; // @[ifu_aln_ctl.scala 166:76]
  wire  _T_178 = _T_164 & _T_187; // @[ifu_aln_ctl.scala 167:35]
  wire  _T_180 = _T_166 & _T_168; // @[Mux.scala 27:72]
  wire  _T_181 = _T_172 & _T_174; // @[Mux.scala 27:72]
  wire  _T_182 = _T_178 & q0off; // @[Mux.scala 27:72]
  wire  _T_183 = _T_180 | _T_181; // @[Mux.scala 27:72]
  wire [50:0] _T_205 = {io_ifu_bp_btb_target_f,io_ifu_bp_poffset_f,io_ifu_bp_fghr_f}; // @[Cat.scala 29:58]
  wire [3:0] _T_207 = {io_iccm_rd_ecc_double_err,io_ic_access_fault_f,io_ic_access_fault_type_f}; // @[Cat.scala 29:58]
  wire [109:0] _T_211 = {misc1,misc0}; // @[Cat.scala 29:58]
  wire [109:0] _T_214 = {misc2,misc1}; // @[Cat.scala 29:58]
  wire [109:0] _T_217 = {misc0,misc2}; // @[Cat.scala 29:58]
  wire [109:0] _T_218 = qren[0] ? _T_211 : 110'h0; // @[Mux.scala 27:72]
  wire [109:0] _T_219 = qren[1] ? _T_214 : 110'h0; // @[Mux.scala 27:72]
  wire [109:0] _T_220 = qren[2] ? _T_217 : 110'h0; // @[Mux.scala 27:72]
  wire [109:0] _T_221 = _T_218 | _T_219; // @[Mux.scala 27:72]
  wire [109:0] misceff = _T_221 | _T_220; // @[Mux.scala 27:72]
  wire [54:0] misc1eff = misceff[109:55]; // @[ifu_aln_ctl.scala 186:25]
  wire [54:0] misc0eff = misceff[54:0]; // @[ifu_aln_ctl.scala 187:25]
  wire  f1dbecc = misc1eff[54]; // @[ifu_aln_ctl.scala 190:25]
  wire  f1icaf = misc1eff[53]; // @[ifu_aln_ctl.scala 191:21]
  wire [1:0] f1ictype = misc1eff[52:51]; // @[ifu_aln_ctl.scala 192:26]
  wire [30:0] f1prett = misc1eff[50:20]; // @[ifu_aln_ctl.scala 193:25]
  wire [11:0] f1poffset = misc1eff[19:8]; // @[ifu_aln_ctl.scala 194:27]
  wire [7:0] f1fghr = misc1eff[7:0]; // @[ifu_aln_ctl.scala 195:24]
  wire  f0dbecc = misc0eff[54]; // @[ifu_aln_ctl.scala 197:25]
  wire  f0icaf = misc0eff[53]; // @[ifu_aln_ctl.scala 198:21]
  wire [1:0] f0ictype = misc0eff[52:51]; // @[ifu_aln_ctl.scala 199:26]
  wire [30:0] f0prett = misc0eff[50:20]; // @[ifu_aln_ctl.scala 200:25]
  wire [11:0] f0poffset = misc0eff[19:8]; // @[ifu_aln_ctl.scala 201:27]
  wire [7:0] f0fghr = misc0eff[7:0]; // @[ifu_aln_ctl.scala 202:24]
  wire [5:0] _T_241 = {io_ifu_bp_hist1_f[0],io_ifu_bp_hist0_f[0],io_ifu_bp_pc4_f[0],io_ifu_bp_way_f[0],io_ifu_bp_valid_f[0],io_ifu_bp_ret_f[0]}; // @[Cat.scala 29:58]
  wire [5:0] _T_246 = {io_ifu_bp_hist1_f[1],io_ifu_bp_hist0_f[1],io_ifu_bp_pc4_f[1],io_ifu_bp_way_f[1],io_ifu_bp_valid_f[1],io_ifu_bp_ret_f[1]}; // @[Cat.scala 29:58]
  wire [23:0] _T_250 = {brdata1,brdata0}; // @[Cat.scala 29:58]
  wire [23:0] _T_253 = {brdata2,brdata1}; // @[Cat.scala 29:58]
  wire [23:0] _T_256 = {brdata0,brdata2}; // @[Cat.scala 29:58]
  wire [23:0] _T_257 = qren[0] ? _T_250 : 24'h0; // @[Mux.scala 27:72]
  wire [23:0] _T_258 = qren[1] ? _T_253 : 24'h0; // @[Mux.scala 27:72]
  wire [23:0] _T_259 = qren[2] ? _T_256 : 24'h0; // @[Mux.scala 27:72]
  wire [23:0] _T_260 = _T_257 | _T_258; // @[Mux.scala 27:72]
  wire [23:0] brdataeff = _T_260 | _T_259; // @[Mux.scala 27:72]
  wire [11:0] brdata0eff = brdataeff[11:0]; // @[ifu_aln_ctl.scala 213:43]
  wire [11:0] brdata1eff = brdataeff[23:12]; // @[ifu_aln_ctl.scala 213:61]
  wire [11:0] _T_267 = q0sel[0] ? brdata0eff : 12'h0; // @[Mux.scala 27:72]
  wire [5:0] _T_268 = q0sel[1] ? brdata0eff[11:6] : 6'h0; // @[Mux.scala 27:72]
  wire [11:0] _GEN_5 = {{6'd0}, _T_268}; // @[Mux.scala 27:72]
  wire [11:0] brdata0final = _T_267 | _GEN_5; // @[Mux.scala 27:72]
  wire [11:0] _T_275 = q1sel[0] ? brdata1eff : 12'h0; // @[Mux.scala 27:72]
  wire [5:0] _T_276 = q1sel[1] ? brdata1eff[11:6] : 6'h0; // @[Mux.scala 27:72]
  wire [11:0] _GEN_6 = {{6'd0}, _T_276}; // @[Mux.scala 27:72]
  wire [11:0] brdata1final = _T_275 | _GEN_6; // @[Mux.scala 27:72]
  wire [1:0] f0ret = {brdata0final[6],brdata0final[0]}; // @[Cat.scala 29:58]
  wire [1:0] f0brend = {brdata0final[7],brdata0final[1]}; // @[Cat.scala 29:58]
  wire [1:0] f0way = {brdata0final[8],brdata0final[2]}; // @[Cat.scala 29:58]
  wire [1:0] f0pc4 = {brdata0final[9],brdata0final[3]}; // @[Cat.scala 29:58]
  wire [1:0] f0hist0 = {brdata0final[10],brdata0final[4]}; // @[Cat.scala 29:58]
  wire [1:0] f0hist1 = {brdata0final[11],brdata0final[5]}; // @[Cat.scala 29:58]
  wire [1:0] f1ret = {brdata1final[6],brdata1final[0]}; // @[Cat.scala 29:58]
  wire [1:0] f1brend = {brdata1final[7],brdata1final[1]}; // @[Cat.scala 29:58]
  wire [1:0] f1way = {brdata1final[8],brdata1final[2]}; // @[Cat.scala 29:58]
  wire [1:0] f1pc4 = {brdata1final[9],brdata1final[3]}; // @[Cat.scala 29:58]
  wire [1:0] f1hist0 = {brdata1final[10],brdata1final[4]}; // @[Cat.scala 29:58]
  wire [1:0] f1hist1 = {brdata1final[11],brdata1final[5]}; // @[Cat.scala 29:58]
  wire  consume_fb0 = _T_351 & f0val[0]; // @[ifu_aln_ctl.scala 237:32]
  wire  consume_fb1 = _T_335 & f1val[0]; // @[ifu_aln_ctl.scala 238:32]
  wire  _T_311 = ~consume_fb1; // @[ifu_aln_ctl.scala 241:39]
  wire  _T_312 = consume_fb0 & _T_311; // @[ifu_aln_ctl.scala 241:37]
  wire  _T_315 = consume_fb0 & consume_fb1; // @[ifu_aln_ctl.scala 242:37]
  wire [30:0] f0pc_plus1 = f0pc + 31'h1; // @[ifu_aln_ctl.scala 259:25]
  wire [30:0] f1pc_plus1 = f1pc + 31'h1; // @[ifu_aln_ctl.scala 261:25]
  wire [30:0] _T_363 = f1_shift_2B ? 31'h7fffffff : 31'h0; // @[Bitwise.scala 72:12]
  wire [30:0] _T_364 = _T_363 & f1pc_plus1; // @[ifu_aln_ctl.scala 263:38]
  wire [30:0] _T_367 = _T_416 ? 31'h7fffffff : 31'h0; // @[Bitwise.scala 72:12]
  wire [30:0] _T_368 = _T_367 & f1pc; // @[ifu_aln_ctl.scala 263:78]
  wire [30:0] sf1pc = _T_364 | _T_368; // @[ifu_aln_ctl.scala 263:52]
  wire  _T_371 = ~fetch_to_f1; // @[ifu_aln_ctl.scala 267:6]
  wire  _T_372 = ~_T_353; // @[ifu_aln_ctl.scala 267:21]
  wire  _T_373 = _T_371 & _T_372; // @[ifu_aln_ctl.scala 267:19]
  wire [30:0] _T_375 = fetch_to_f1 ? io_ifu_fetch_pc : 31'h0; // @[Mux.scala 27:72]
  wire [30:0] _T_376 = _T_353 ? f2pc : 31'h0; // @[Mux.scala 27:72]
  wire [30:0] _T_377 = _T_373 ? sf1pc : 31'h0; // @[Mux.scala 27:72]
  wire [30:0] _T_378 = _T_375 | _T_376; // @[Mux.scala 27:72]
  wire  _T_384 = ~fetch_to_f0; // @[ifu_aln_ctl.scala 272:24]
  wire  _T_385 = ~_T_337; // @[ifu_aln_ctl.scala 272:39]
  wire  _T_386 = _T_384 & _T_385; // @[ifu_aln_ctl.scala 272:37]
  wire  _T_387 = ~_T_352; // @[ifu_aln_ctl.scala 272:54]
  wire  _T_388 = _T_386 & _T_387; // @[ifu_aln_ctl.scala 272:52]
  wire [30:0] _T_390 = fetch_to_f0 ? io_ifu_fetch_pc : 31'h0; // @[Mux.scala 27:72]
  wire [30:0] _T_391 = _T_337 ? f2pc : 31'h0; // @[Mux.scala 27:72]
  wire [30:0] _T_392 = _T_352 ? sf1pc : 31'h0; // @[Mux.scala 27:72]
  wire [30:0] _T_393 = _T_388 ? f0pc_plus1 : 31'h0; // @[Mux.scala 27:72]
  wire [30:0] _T_394 = _T_390 | _T_391; // @[Mux.scala 27:72]
  wire [30:0] _T_395 = _T_394 | _T_392; // @[Mux.scala 27:72]
  wire  _T_399 = fetch_to_f2 & _T_1; // @[ifu_aln_ctl.scala 274:38]
  wire  _T_401 = ~fetch_to_f2; // @[ifu_aln_ctl.scala 275:25]
  wire  _T_403 = _T_401 & _T_372; // @[ifu_aln_ctl.scala 275:38]
  wire  _T_405 = _T_403 & _T_385; // @[ifu_aln_ctl.scala 275:53]
  wire  _T_407 = _T_405 & _T_1; // @[ifu_aln_ctl.scala 275:68]
  wire [1:0] _T_409 = _T_399 ? io_ifu_fetch_val : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_410 = _T_407 ? f2val : 2'h0; // @[Mux.scala 27:72]
  wire  _T_422 = fetch_to_f1 & _T_1; // @[ifu_aln_ctl.scala 279:39]
  wire  _T_425 = _T_353 & _T_1; // @[ifu_aln_ctl.scala 280:54]
  wire  _T_431 = _T_373 & _T_387; // @[ifu_aln_ctl.scala 281:54]
  wire  _T_433 = _T_431 & _T_1; // @[ifu_aln_ctl.scala 281:69]
  wire [1:0] _T_435 = _T_422 ? io_ifu_fetch_val : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_436 = _T_425 ? f2val : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_437 = _T_433 ? sf1val : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_438 = _T_435 | _T_436; // @[Mux.scala 27:72]
  wire  _T_453 = fetch_to_f0 & _T_1; // @[ifu_aln_ctl.scala 286:38]
  wire  _T_456 = _T_337 & _T_1; // @[ifu_aln_ctl.scala 287:54]
  wire  _T_459 = _T_352 & _T_1; // @[ifu_aln_ctl.scala 288:69]
  wire  _T_467 = _T_388 & _T_1; // @[ifu_aln_ctl.scala 289:69]
  wire [1:0] _T_469 = _T_453 ? io_ifu_fetch_val : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_470 = _T_456 ? f2val : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_471 = _T_459 ? sf1val : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_472 = _T_467 ? sf0val : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_473 = _T_469 | _T_470; // @[Mux.scala 27:72]
  wire [1:0] _T_474 = _T_473 | _T_471; // @[Mux.scala 27:72]
  wire [1:0] _T_530 = {f1val[0],1'h1}; // @[Cat.scala 29:58]
  wire [1:0] _T_531 = f0val[1] ? 2'h3 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_532 = _T_515 ? _T_530 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] alignval = _T_531 | _T_532; // @[Mux.scala 27:72]
  wire [1:0] _T_542 = {f1icaf,f0icaf}; // @[Cat.scala 29:58]
  wire  _T_543 = f0val[1] & f0icaf; // @[Mux.scala 27:72]
  wire [1:0] _T_544 = _T_515 ? _T_542 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _GEN_7 = {{1'd0}, _T_543}; // @[Mux.scala 27:72]
  wire [1:0] alignicaf = _GEN_7 | _T_544; // @[Mux.scala 27:72]
  wire [1:0] _T_549 = f0dbecc ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [1:0] _T_555 = {f1dbecc,f0dbecc}; // @[Cat.scala 29:58]
  wire [1:0] _T_556 = f0val[1] ? _T_549 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_557 = _T_515 ? _T_555 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] aligndbecc = _T_556 | _T_557; // @[Mux.scala 27:72]
  wire [1:0] _T_568 = {f1brend[0],f0brend[0]}; // @[Cat.scala 29:58]
  wire [1:0] _T_569 = f0val[1] ? f0brend : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_570 = _T_515 ? _T_568 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] alignbrend = _T_569 | _T_570; // @[Mux.scala 27:72]
  wire [1:0] _T_581 = {f1pc4[0],f0pc4[0]}; // @[Cat.scala 29:58]
  wire [1:0] _T_582 = f0val[1] ? f0pc4 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_583 = _T_515 ? _T_581 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] alignpc4 = _T_582 | _T_583; // @[Mux.scala 27:72]
  wire [1:0] _T_594 = {f1ret[0],f0ret[0]}; // @[Cat.scala 29:58]
  wire [1:0] _T_595 = f0val[1] ? f0ret : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_596 = _T_515 ? _T_594 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] alignret = _T_595 | _T_596; // @[Mux.scala 27:72]
  wire [1:0] _T_607 = {f1way[0],f0way[0]}; // @[Cat.scala 29:58]
  wire [1:0] _T_608 = f0val[1] ? f0way : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_609 = _T_515 ? _T_607 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] alignway = _T_608 | _T_609; // @[Mux.scala 27:72]
  wire [1:0] _T_620 = {f1hist1[0],f0hist1[0]}; // @[Cat.scala 29:58]
  wire [1:0] _T_621 = f0val[1] ? f0hist1 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_622 = _T_515 ? _T_620 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] alignhist1 = _T_621 | _T_622; // @[Mux.scala 27:72]
  wire [1:0] _T_633 = {f1hist0[0],f0hist0[0]}; // @[Cat.scala 29:58]
  wire [1:0] _T_634 = f0val[1] ? f0hist0 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_635 = _T_515 ? _T_633 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] alignhist0 = _T_634 | _T_635; // @[Mux.scala 27:72]
  wire [30:0] _T_647 = f0val[1] ? f0pc_plus1 : 31'h0; // @[Mux.scala 27:72]
  wire [30:0] _T_648 = _T_515 ? f1pc : 31'h0; // @[Mux.scala 27:72]
  wire [30:0] secondpc = _T_647 | _T_648; // @[Mux.scala 27:72]
  wire  _T_657 = first4B & alignval[1]; // @[Mux.scala 27:72]
  wire  _T_658 = first2B & alignval[0]; // @[Mux.scala 27:72]
  wire  _T_662 = |alignicaf; // @[ifu_aln_ctl.scala 340:74]
  wire  _T_665 = first4B & _T_662; // @[Mux.scala 27:72]
  wire  _T_666 = first2B & alignicaf[0]; // @[Mux.scala 27:72]
  wire  _T_671 = first4B & _T_513; // @[ifu_aln_ctl.scala 342:54]
  wire  _T_673 = _T_671 & f0val[0]; // @[ifu_aln_ctl.scala 342:66]
  wire  _T_675 = ~alignicaf[0]; // @[ifu_aln_ctl.scala 342:79]
  wire  _T_676 = _T_673 & _T_675; // @[ifu_aln_ctl.scala 342:77]
  wire  _T_678 = ~aligndbecc[0]; // @[ifu_aln_ctl.scala 342:95]
  wire  _T_679 = _T_676 & _T_678; // @[ifu_aln_ctl.scala 342:93]
  wire  icaf_eff = alignicaf[1] | aligndbecc[1]; // @[ifu_aln_ctl.scala 344:31]
  wire  _T_684 = first4B & icaf_eff; // @[ifu_aln_ctl.scala 346:47]
  wire  _T_687 = |aligndbecc; // @[ifu_aln_ctl.scala 348:74]
  wire  _T_690 = first4B & _T_687; // @[Mux.scala 27:72]
  wire  _T_691 = first2B & aligndbecc[0]; // @[Mux.scala 27:72]
  wire [31:0] _T_696 = first4B ? aligndata : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_697 = first2B ? decompressed_io_dout : 32'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_702 = f0pc[8:1] ^ f0pc[16:9]; // @[lib.scala 51:47]
  wire [7:0] firstpc_hash = _T_702 ^ f0pc[24:17]; // @[lib.scala 51:85]
  wire [7:0] _T_706 = secondpc[8:1] ^ secondpc[16:9]; // @[lib.scala 51:47]
  wire [7:0] secondpc_hash = _T_706 ^ secondpc[24:17]; // @[lib.scala 51:85]
  wire [4:0] _T_712 = f0pc[13:9] ^ f0pc[18:14]; // @[lib.scala 42:111]
  wire [4:0] firstbrtag_hash = _T_712 ^ f0pc[23:19]; // @[lib.scala 42:111]
  wire [4:0] _T_717 = secondpc[13:9] ^ secondpc[18:14]; // @[lib.scala 42:111]
  wire [4:0] secondbrtag_hash = _T_717 ^ secondpc[23:19]; // @[lib.scala 42:111]
  wire  _T_719 = first2B & alignbrend[0]; // @[ifu_aln_ctl.scala 365:45]
  wire  _T_721 = first4B & alignbrend[1]; // @[ifu_aln_ctl.scala 365:73]
  wire  _T_722 = _T_719 | _T_721; // @[ifu_aln_ctl.scala 365:62]
  wire  _T_726 = _T_657 & alignbrend[0]; // @[ifu_aln_ctl.scala 365:115]
  wire  _T_729 = first2B & alignret[0]; // @[ifu_aln_ctl.scala 367:49]
  wire  _T_731 = first4B & alignret[1]; // @[ifu_aln_ctl.scala 367:75]
  wire  _T_734 = first2B & alignpc4[0]; // @[ifu_aln_ctl.scala 369:29]
  wire  _T_736 = first4B & alignpc4[1]; // @[ifu_aln_ctl.scala 369:55]
  wire  i0_brp_pc4 = _T_734 | _T_736; // @[ifu_aln_ctl.scala 369:44]
  wire  _T_738 = first2B | alignbrend[0]; // @[ifu_aln_ctl.scala 371:53]
  wire  _T_744 = first2B & alignhist1[0]; // @[ifu_aln_ctl.scala 373:54]
  wire  _T_746 = first4B & alignhist1[1]; // @[ifu_aln_ctl.scala 373:82]
  wire  _T_747 = _T_744 | _T_746; // @[ifu_aln_ctl.scala 373:71]
  wire  _T_749 = first2B & alignhist0[0]; // @[ifu_aln_ctl.scala 374:14]
  wire  _T_751 = first4B & alignhist0[1]; // @[ifu_aln_ctl.scala 374:42]
  wire  _T_752 = _T_749 | _T_751; // @[ifu_aln_ctl.scala 374:31]
  wire  i0_ends_f1 = first4B & _T_515; // @[ifu_aln_ctl.scala 376:28]
  wire  _T_768 = io_dec_aln_aln_ib_i0_brp_valid & i0_brp_pc4; // @[ifu_aln_ctl.scala 385:77]
  wire  _T_769 = _T_768 & first2B; // @[ifu_aln_ctl.scala 385:91]
  wire  _T_770 = ~i0_brp_pc4; // @[ifu_aln_ctl.scala 385:139]
  wire  _T_771 = io_dec_aln_aln_ib_i0_brp_valid & _T_770; // @[ifu_aln_ctl.scala 385:137]
  wire  _T_772 = _T_771 & first4B; // @[ifu_aln_ctl.scala 385:151]
  rvclkhdr rvclkhdr ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_io_l1clk),
    .io_clk(rvclkhdr_io_clk),
    .io_en(rvclkhdr_io_en),
    .io_scan_mode(rvclkhdr_io_scan_mode)
  );
  rvclkhdr rvclkhdr_1 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_1_io_l1clk),
    .io_clk(rvclkhdr_1_io_clk),
    .io_en(rvclkhdr_1_io_en),
    .io_scan_mode(rvclkhdr_1_io_scan_mode)
  );
  rvclkhdr rvclkhdr_2 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_2_io_l1clk),
    .io_clk(rvclkhdr_2_io_clk),
    .io_en(rvclkhdr_2_io_en),
    .io_scan_mode(rvclkhdr_2_io_scan_mode)
  );
  rvclkhdr rvclkhdr_3 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_3_io_l1clk),
    .io_clk(rvclkhdr_3_io_clk),
    .io_en(rvclkhdr_3_io_en),
    .io_scan_mode(rvclkhdr_3_io_scan_mode)
  );
  rvclkhdr rvclkhdr_4 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_4_io_l1clk),
    .io_clk(rvclkhdr_4_io_clk),
    .io_en(rvclkhdr_4_io_en),
    .io_scan_mode(rvclkhdr_4_io_scan_mode)
  );
  rvclkhdr rvclkhdr_5 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_5_io_l1clk),
    .io_clk(rvclkhdr_5_io_clk),
    .io_en(rvclkhdr_5_io_en),
    .io_scan_mode(rvclkhdr_5_io_scan_mode)
  );
  rvclkhdr rvclkhdr_6 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_6_io_l1clk),
    .io_clk(rvclkhdr_6_io_clk),
    .io_en(rvclkhdr_6_io_en),
    .io_scan_mode(rvclkhdr_6_io_scan_mode)
  );
  rvclkhdr rvclkhdr_7 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_7_io_l1clk),
    .io_clk(rvclkhdr_7_io_clk),
    .io_en(rvclkhdr_7_io_en),
    .io_scan_mode(rvclkhdr_7_io_scan_mode)
  );
  rvclkhdr rvclkhdr_8 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_8_io_l1clk),
    .io_clk(rvclkhdr_8_io_clk),
    .io_en(rvclkhdr_8_io_en),
    .io_scan_mode(rvclkhdr_8_io_scan_mode)
  );
  rvclkhdr rvclkhdr_9 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_9_io_l1clk),
    .io_clk(rvclkhdr_9_io_clk),
    .io_en(rvclkhdr_9_io_en),
    .io_scan_mode(rvclkhdr_9_io_scan_mode)
  );
  rvclkhdr rvclkhdr_10 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_10_io_l1clk),
    .io_clk(rvclkhdr_10_io_clk),
    .io_en(rvclkhdr_10_io_en),
    .io_scan_mode(rvclkhdr_10_io_scan_mode)
  );
  rvclkhdr rvclkhdr_11 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_11_io_l1clk),
    .io_clk(rvclkhdr_11_io_clk),
    .io_en(rvclkhdr_11_io_en),
    .io_scan_mode(rvclkhdr_11_io_scan_mode)
  );
  ifu_compress_ctl decompressed ( // @[ifu_aln_ctl.scala 352:28]
    .io_din(decompressed_io_din),
    .io_dout(decompressed_io_dout)
  );
  assign io_dec_aln_aln_dec_ifu_i0_cinst = aligndata[15:0]; // @[ifu_aln_ctl.scala 331:35]
  assign io_dec_aln_aln_ib_ifu_i0_icaf = _T_665 | _T_666; // @[ifu_aln_ctl.scala 340:33]
  assign io_dec_aln_aln_ib_ifu_i0_icaf_type = _T_679 ? f1ictype : f0ictype; // @[ifu_aln_ctl.scala 342:38]
  assign io_dec_aln_aln_ib_ifu_i0_icaf_f1 = _T_684 & _T_515; // @[ifu_aln_ctl.scala 346:36]
  assign io_dec_aln_aln_ib_ifu_i0_dbecc = _T_690 | _T_691; // @[ifu_aln_ctl.scala 348:34]
  assign io_dec_aln_aln_ib_ifu_i0_bp_index = _T_738 ? firstpc_hash : secondpc_hash; // @[ifu_aln_ctl.scala 387:37]
  assign io_dec_aln_aln_ib_ifu_i0_bp_fghr = i0_ends_f1 ? f1fghr : f0fghr; // @[ifu_aln_ctl.scala 389:36]
  assign io_dec_aln_aln_ib_ifu_i0_bp_btag = _T_738 ? firstbrtag_hash : secondbrtag_hash; // @[ifu_aln_ctl.scala 391:36]
  assign io_dec_aln_aln_ib_ifu_i0_valid = _T_657 | _T_658; // @[ifu_aln_ctl.scala 338:34]
  assign io_dec_aln_aln_ib_ifu_i0_instr = _T_696 | _T_697; // @[ifu_aln_ctl.scala 354:34]
  assign io_dec_aln_aln_ib_ifu_i0_pc = f0pc; // @[ifu_aln_ctl.scala 325:31]
  assign io_dec_aln_aln_ib_ifu_i0_pc4 = aligndata[1:0] == 2'h3; // @[ifu_aln_ctl.scala 329:32]
  assign io_dec_aln_aln_ib_i0_brp_valid = _T_722 | _T_726; // @[ifu_aln_ctl.scala 365:34]
  assign io_dec_aln_aln_ib_i0_brp_bits_toffset = i0_ends_f1 ? f1poffset : f0poffset; // @[ifu_aln_ctl.scala 377:41]
  assign io_dec_aln_aln_ib_i0_brp_bits_hist = {_T_747,_T_752}; // @[ifu_aln_ctl.scala 373:38]
  assign io_dec_aln_aln_ib_i0_brp_bits_br_error = _T_769 | _T_772; // @[ifu_aln_ctl.scala 385:42]
  assign io_dec_aln_aln_ib_i0_brp_bits_br_start_error = _T_657 & alignbrend[0]; // @[ifu_aln_ctl.scala 381:49]
  assign io_dec_aln_aln_ib_i0_brp_bits_prett = i0_ends_f1 ? f1prett : f0prett; // @[ifu_aln_ctl.scala 379:39]
  assign io_dec_aln_aln_ib_i0_brp_bits_way = _T_738 ? alignway[0] : alignway[1]; // @[ifu_aln_ctl.scala 371:37]
  assign io_dec_aln_aln_ib_i0_brp_bits_ret = _T_729 | _T_731; // @[ifu_aln_ctl.scala 367:37]
  assign io_dec_aln_ifu_pmu_instr_aligned = io_dec_aln_aln_dec_dec_i0_decode_d & _T_785; // @[ifu_aln_ctl.scala 397:36]
  assign io_ifu_fb_consume1 = _T_312 & _T_1; // @[ifu_aln_ctl.scala 241:22]
  assign io_ifu_fb_consume2 = _T_315 & _T_1; // @[ifu_aln_ctl.scala 242:22]
  assign rvclkhdr_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_io_en = _T_354 | _T_358; // @[lib.scala 371:17]
  assign rvclkhdr_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_1_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_1_io_en = _T_25 | f1_shift_2B; // @[lib.scala 371:17]
  assign rvclkhdr_1_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_2_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_2_io_en = _T_29 | shift_4B; // @[lib.scala 371:17]
  assign rvclkhdr_2_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_3_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_3_io_en = qwen[2]; // @[lib.scala 371:17]
  assign rvclkhdr_3_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_4_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_4_io_en = qwen[1]; // @[lib.scala 371:17]
  assign rvclkhdr_4_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_5_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_5_io_en = qwen[0]; // @[lib.scala 371:17]
  assign rvclkhdr_5_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_6_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_6_io_en = qwen[2]; // @[lib.scala 371:17]
  assign rvclkhdr_6_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_7_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_7_io_en = qwen[1]; // @[lib.scala 371:17]
  assign rvclkhdr_7_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_8_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_8_io_en = qwen[0]; // @[lib.scala 371:17]
  assign rvclkhdr_8_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_9_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_9_io_en = qwen[2]; // @[lib.scala 371:17]
  assign rvclkhdr_9_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_10_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_10_io_en = qwen[1]; // @[lib.scala 371:17]
  assign rvclkhdr_10_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_11_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_11_io_en = qwen[0]; // @[lib.scala 371:17]
  assign rvclkhdr_11_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign decompressed_io_din = aligndata[15:0]; // @[ifu_aln_ctl.scala 393:23]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  error_stall = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  wrptr = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  rdptr = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  f2val = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  f1val = _RAND_4[1:0];
  _RAND_5 = {1{`RANDOM}};
  f0val = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  q2off = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  q1off = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  q0off = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  q1 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  q0 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  q2 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  f2pc = _RAND_12[30:0];
  _RAND_13 = {1{`RANDOM}};
  f1pc = _RAND_13[30:0];
  _RAND_14 = {1{`RANDOM}};
  f0pc = _RAND_14[30:0];
  _RAND_15 = {1{`RANDOM}};
  brdata2 = _RAND_15[11:0];
  _RAND_16 = {1{`RANDOM}};
  brdata1 = _RAND_16[11:0];
  _RAND_17 = {1{`RANDOM}};
  brdata0 = _RAND_17[11:0];
  _RAND_18 = {2{`RANDOM}};
  misc2 = _RAND_18[54:0];
  _RAND_19 = {2{`RANDOM}};
  misc1 = _RAND_19[54:0];
  _RAND_20 = {2{`RANDOM}};
  misc0 = _RAND_20[54:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    error_stall = 1'h0;
  end
  if (reset) begin
    wrptr = 2'h0;
  end
  if (reset) begin
    rdptr = 2'h0;
  end
  if (reset) begin
    f2val = 2'h0;
  end
  if (reset) begin
    f1val = 2'h0;
  end
  if (reset) begin
    f0val = 2'h0;
  end
  if (reset) begin
    q2off = 1'h0;
  end
  if (reset) begin
    q1off = 1'h0;
  end
  if (reset) begin
    q0off = 1'h0;
  end
  if (reset) begin
    q1 = 32'h0;
  end
  if (reset) begin
    q0 = 32'h0;
  end
  if (reset) begin
    q2 = 32'h0;
  end
  if (reset) begin
    f2pc = 31'h0;
  end
  if (reset) begin
    f1pc = 31'h0;
  end
  if (reset) begin
    f0pc = 31'h0;
  end
  if (reset) begin
    brdata2 = 12'h0;
  end
  if (reset) begin
    brdata1 = 12'h0;
  end
  if (reset) begin
    brdata0 = 12'h0;
  end
  if (reset) begin
    misc2 = 55'h0;
  end
  if (reset) begin
    misc1 = 55'h0;
  end
  if (reset) begin
    misc0 = 55'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      error_stall <= 1'h0;
    end else begin
      error_stall <= _T & _T_1;
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      wrptr <= 2'h0;
    end else begin
      wrptr <= _T_113 | _T_112;
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      rdptr <= 2'h0;
    end else begin
      rdptr <= _T_90 | _T_85;
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      f2val <= 2'h0;
    end else begin
      f2val <= _T_409 | _T_410;
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      f1val <= 2'h0;
    end else begin
      f1val <= _T_438 | _T_437;
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      f0val <= 2'h0;
    end else begin
      f0val <= _T_474 | _T_472;
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      q2off <= 1'h0;
    end else begin
      q2off <= _T_137 | _T_136;
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      q1off <= 1'h0;
    end else begin
      q1off <= _T_160 | _T_159;
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      q0off <= 1'h0;
    end else begin
      q0off <= _T_183 | _T_182;
    end
  end
  always @(posedge rvclkhdr_10_io_l1clk or posedge reset) begin
    if (reset) begin
      q1 <= 32'h0;
    end else begin
      q1 <= io_ifu_fetch_data_f;
    end
  end
  always @(posedge rvclkhdr_11_io_l1clk or posedge reset) begin
    if (reset) begin
      q0 <= 32'h0;
    end else begin
      q0 <= io_ifu_fetch_data_f;
    end
  end
  always @(posedge rvclkhdr_9_io_l1clk or posedge reset) begin
    if (reset) begin
      q2 <= 32'h0;
    end else begin
      q2 <= io_ifu_fetch_data_f;
    end
  end
  always @(posedge rvclkhdr_io_l1clk or posedge reset) begin
    if (reset) begin
      f2pc <= 31'h0;
    end else begin
      f2pc <= io_ifu_fetch_pc;
    end
  end
  always @(posedge rvclkhdr_1_io_l1clk or posedge reset) begin
    if (reset) begin
      f1pc <= 31'h0;
    end else begin
      f1pc <= _T_378 | _T_377;
    end
  end
  always @(posedge rvclkhdr_2_io_l1clk or posedge reset) begin
    if (reset) begin
      f0pc <= 31'h0;
    end else begin
      f0pc <= _T_395 | _T_393;
    end
  end
  always @(posedge rvclkhdr_3_io_l1clk or posedge reset) begin
    if (reset) begin
      brdata2 <= 12'h0;
    end else begin
      brdata2 <= {_T_246,_T_241};
    end
  end
  always @(posedge rvclkhdr_4_io_l1clk or posedge reset) begin
    if (reset) begin
      brdata1 <= 12'h0;
    end else begin
      brdata1 <= {_T_246,_T_241};
    end
  end
  always @(posedge rvclkhdr_5_io_l1clk or posedge reset) begin
    if (reset) begin
      brdata0 <= 12'h0;
    end else begin
      brdata0 <= {_T_246,_T_241};
    end
  end
  always @(posedge rvclkhdr_6_io_l1clk or posedge reset) begin
    if (reset) begin
      misc2 <= 55'h0;
    end else begin
      misc2 <= {_T_207,_T_205};
    end
  end
  always @(posedge rvclkhdr_7_io_l1clk or posedge reset) begin
    if (reset) begin
      misc1 <= 55'h0;
    end else begin
      misc1 <= {_T_207,_T_205};
    end
  end
  always @(posedge rvclkhdr_8_io_l1clk or posedge reset) begin
    if (reset) begin
      misc0 <= 55'h0;
    end else begin
      misc0 <= {_T_207,_T_205};
    end
  end
endmodule
module ifu_ifc_ctl(
  input         clock,
  input         reset,
  input         io_exu_flush_final,
  input  [30:0] io_exu_flush_path_final,
  input         io_free_clk,
  input         io_active_clk,
  input         io_scan_mode,
  input         io_ic_hit_f,
  input         io_ifu_ic_mb_empty,
  input         io_ifu_fb_consume1,
  input         io_ifu_fb_consume2,
  input         io_ifu_bp_hit_taken_f,
  input  [30:0] io_ifu_bp_btb_target_f,
  input         io_ic_dma_active,
  input         io_dec_ifc_dec_tlu_flush_noredir_wb,
  input  [31:0] io_dec_ifc_dec_tlu_mrac_ff,
  output        io_dec_ifc_ifu_pmu_fetch_stall,
  input         io_dma_ifc_dma_iccm_stall_any,
  output [30:0] io_ifc_fetch_addr_f,
  output [30:0] io_ifc_fetch_addr_bf,
  output        io_ifc_fetch_req_f,
  output        io_ifc_fetch_uncacheable_bf,
  output        io_ifc_fetch_req_bf,
  output        io_ifc_fetch_req_bf_raw,
  output        io_ifc_iccm_access_bf,
  output        io_ifc_region_acc_fault_bf,
  output        io_ifc_dma_access_ok
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  wire  rvclkhdr_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_io_scan_mode; // @[lib.scala 368:23]
  reg  dma_iccm_stall_any_f; // @[ifu_ifc_ctl.scala 63:58]
  wire  dma_stall = io_ic_dma_active | dma_iccm_stall_any_f; // @[ifu_ifc_ctl.scala 62:36]
  reg  miss_a; // @[ifu_ifc_ctl.scala 65:44]
  wire  _T_2 = ~io_exu_flush_final; // @[ifu_ifc_ctl.scala 67:26]
  wire  _T_3 = ~io_ifc_fetch_req_f; // @[ifu_ifc_ctl.scala 67:49]
  wire  _T_4 = ~io_ic_hit_f; // @[ifu_ifc_ctl.scala 67:71]
  wire  _T_5 = _T_3 | _T_4; // @[ifu_ifc_ctl.scala 67:69]
  wire  sel_last_addr_bf = _T_2 & _T_5; // @[ifu_ifc_ctl.scala 67:46]
  wire  _T_7 = _T_2 & io_ifc_fetch_req_f; // @[ifu_ifc_ctl.scala 68:46]
  wire  _T_8 = _T_7 & io_ifu_bp_hit_taken_f; // @[ifu_ifc_ctl.scala 68:67]
  wire  sel_btb_addr_bf = _T_8 & io_ic_hit_f; // @[ifu_ifc_ctl.scala 68:92]
  wire  _T_11 = ~io_ifu_bp_hit_taken_f; // @[ifu_ifc_ctl.scala 69:69]
  wire  _T_12 = _T_7 & _T_11; // @[ifu_ifc_ctl.scala 69:67]
  wire  sel_next_addr_bf = _T_12 & io_ic_hit_f; // @[ifu_ifc_ctl.scala 69:92]
  wire [30:0] _T_17 = io_exu_flush_final ? io_exu_flush_path_final : 31'h0; // @[Mux.scala 27:72]
  wire [30:0] _T_18 = sel_last_addr_bf ? io_ifc_fetch_addr_f : 31'h0; // @[Mux.scala 27:72]
  wire [30:0] _T_19 = sel_btb_addr_bf ? io_ifu_bp_btb_target_f : 31'h0; // @[Mux.scala 27:72]
  wire [29:0] address_upper = io_ifc_fetch_addr_f[30:1] + 30'h1; // @[ifu_ifc_ctl.scala 78:48]
  wire  _T_29 = address_upper[4] ^ io_ifc_fetch_addr_f[5]; // @[ifu_ifc_ctl.scala 79:63]
  wire  _T_30 = ~_T_29; // @[ifu_ifc_ctl.scala 79:24]
  wire  fetch_addr_next_0 = _T_30 & io_ifc_fetch_addr_f[0]; // @[ifu_ifc_ctl.scala 79:109]
  wire [30:0] fetch_addr_next = {address_upper,fetch_addr_next_0}; // @[Cat.scala 29:58]
  wire [30:0] _T_20 = sel_next_addr_bf ? fetch_addr_next : 31'h0; // @[Mux.scala 27:72]
  wire [30:0] _T_21 = _T_17 | _T_18; // @[Mux.scala 27:72]
  wire [30:0] _T_22 = _T_21 | _T_19; // @[Mux.scala 27:72]
  reg [1:0] state; // @[ifu_ifc_ctl.scala 104:45]
  wire  idle = state == 2'h0; // @[ifu_ifc_ctl.scala 123:17]
  wire  _T_35 = io_ifu_fb_consume2 | io_ifu_fb_consume1; // @[ifu_ifc_ctl.scala 86:91]
  wire  _T_36 = ~_T_35; // @[ifu_ifc_ctl.scala 86:70]
  wire [3:0] _T_121 = io_exu_flush_final ? 4'h1 : 4'h0; // @[Mux.scala 27:72]
  wire  _T_81 = ~io_ifu_fb_consume2; // @[ifu_ifc_ctl.scala 109:38]
  wire  _T_82 = io_ifu_fb_consume1 & _T_81; // @[ifu_ifc_ctl.scala 109:36]
  wire  _T_48 = io_ifc_fetch_req_f & _T_4; // @[ifu_ifc_ctl.scala 91:32]
  wire  miss_f = _T_48 & _T_2; // @[ifu_ifc_ctl.scala 91:47]
  wire  _T_84 = _T_3 | miss_f; // @[ifu_ifc_ctl.scala 109:81]
  wire  _T_85 = _T_82 & _T_84; // @[ifu_ifc_ctl.scala 109:58]
  wire  _T_86 = io_ifu_fb_consume2 & io_ifc_fetch_req_f; // @[ifu_ifc_ctl.scala 110:25]
  wire  fb_right = _T_85 | _T_86; // @[ifu_ifc_ctl.scala 109:92]
  wire  _T_98 = _T_2 & fb_right; // @[ifu_ifc_ctl.scala 117:16]
  reg [3:0] fb_write_f; // @[ifu_ifc_ctl.scala 128:50]
  wire [3:0] _T_101 = {1'h0,fb_write_f[3:1]}; // @[Cat.scala 29:58]
  wire [3:0] _T_122 = _T_98 ? _T_101 : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_126 = _T_121 | _T_122; // @[Mux.scala 27:72]
  wire  fb_right2 = io_ifu_fb_consume2 & _T_84; // @[ifu_ifc_ctl.scala 112:36]
  wire  _T_103 = _T_2 & fb_right2; // @[ifu_ifc_ctl.scala 118:16]
  wire [3:0] _T_106 = {2'h0,fb_write_f[3:2]}; // @[Cat.scala 29:58]
  wire [3:0] _T_123 = _T_103 ? _T_106 : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_127 = _T_126 | _T_123; // @[Mux.scala 27:72]
  wire  _T_91 = io_ifu_fb_consume1 | io_ifu_fb_consume2; // @[ifu_ifc_ctl.scala 113:56]
  wire  _T_92 = ~_T_91; // @[ifu_ifc_ctl.scala 113:35]
  wire  _T_93 = io_ifc_fetch_req_f & _T_92; // @[ifu_ifc_ctl.scala 113:33]
  wire  _T_94 = ~miss_f; // @[ifu_ifc_ctl.scala 113:80]
  wire  fb_left = _T_93 & _T_94; // @[ifu_ifc_ctl.scala 113:78]
  wire  _T_108 = _T_2 & fb_left; // @[ifu_ifc_ctl.scala 119:16]
  wire [3:0] _T_111 = {fb_write_f[2:0],1'h0}; // @[Cat.scala 29:58]
  wire [3:0] _T_124 = _T_108 ? _T_111 : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_128 = _T_127 | _T_124; // @[Mux.scala 27:72]
  wire  _T_113 = ~fb_right; // @[ifu_ifc_ctl.scala 120:18]
  wire  _T_114 = _T_2 & _T_113; // @[ifu_ifc_ctl.scala 120:16]
  wire  _T_115 = ~fb_right2; // @[ifu_ifc_ctl.scala 120:30]
  wire  _T_116 = _T_114 & _T_115; // @[ifu_ifc_ctl.scala 120:28]
  wire  _T_117 = ~fb_left; // @[ifu_ifc_ctl.scala 120:43]
  wire  _T_118 = _T_116 & _T_117; // @[ifu_ifc_ctl.scala 120:41]
  wire [3:0] _T_125 = _T_118 ? fb_write_f : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] fb_write_ns = _T_128 | _T_125; // @[Mux.scala 27:72]
  wire  fb_full_f_ns = fb_write_ns[3]; // @[ifu_ifc_ctl.scala 126:30]
  wire  _T_37 = fb_full_f_ns & _T_36; // @[ifu_ifc_ctl.scala 86:68]
  wire  _T_38 = ~_T_37; // @[ifu_ifc_ctl.scala 86:53]
  wire  _T_39 = io_ifc_fetch_req_bf_raw & _T_38; // @[ifu_ifc_ctl.scala 86:51]
  wire  _T_40 = ~dma_stall; // @[ifu_ifc_ctl.scala 87:5]
  wire  _T_41 = _T_39 & _T_40; // @[ifu_ifc_ctl.scala 86:114]
  wire  _T_44 = ~io_dec_ifc_dec_tlu_flush_noredir_wb; // @[ifu_ifc_ctl.scala 87:39]
  wire  _T_51 = io_ifu_ic_mb_empty | io_exu_flush_final; // @[ifu_ifc_ctl.scala 93:39]
  wire  _T_53 = _T_51 & _T_40; // @[ifu_ifc_ctl.scala 93:61]
  wire  _T_55 = _T_53 & _T_94; // @[ifu_ifc_ctl.scala 93:74]
  wire  _T_56 = ~miss_a; // @[ifu_ifc_ctl.scala 93:86]
  wire  mb_empty_mod = _T_55 & _T_56; // @[ifu_ifc_ctl.scala 93:84]
  wire  goto_idle = io_exu_flush_final & io_dec_ifc_dec_tlu_flush_noredir_wb; // @[ifu_ifc_ctl.scala 95:35]
  wire  _T_60 = io_exu_flush_final & _T_44; // @[ifu_ifc_ctl.scala 97:36]
  wire  leave_idle = _T_60 & idle; // @[ifu_ifc_ctl.scala 97:75]
  wire  _T_63 = ~state[1]; // @[ifu_ifc_ctl.scala 99:23]
  wire  _T_65 = _T_63 & state[0]; // @[ifu_ifc_ctl.scala 99:33]
  wire  _T_66 = _T_65 & miss_f; // @[ifu_ifc_ctl.scala 99:44]
  wire  _T_67 = ~goto_idle; // @[ifu_ifc_ctl.scala 99:55]
  wire  _T_68 = _T_66 & _T_67; // @[ifu_ifc_ctl.scala 99:53]
  wire  _T_70 = ~mb_empty_mod; // @[ifu_ifc_ctl.scala 100:17]
  wire  _T_71 = state[1] & _T_70; // @[ifu_ifc_ctl.scala 100:15]
  wire  _T_73 = _T_71 & _T_67; // @[ifu_ifc_ctl.scala 100:31]
  wire  next_state_1 = _T_68 | _T_73; // @[ifu_ifc_ctl.scala 99:67]
  wire  _T_75 = _T_67 & leave_idle; // @[ifu_ifc_ctl.scala 102:34]
  wire  _T_78 = state[0] & _T_67; // @[ifu_ifc_ctl.scala 102:60]
  wire  next_state_0 = _T_75 | _T_78; // @[ifu_ifc_ctl.scala 102:48]
  wire  wfm = state == 2'h3; // @[ifu_ifc_ctl.scala 124:16]
  reg  fb_full_f; // @[ifu_ifc_ctl.scala 127:52]
  wire  _T_136 = _T_35 | io_exu_flush_final; // @[ifu_ifc_ctl.scala 131:61]
  wire  _T_137 = ~_T_136; // @[ifu_ifc_ctl.scala 131:19]
  wire  _T_138 = fb_full_f & _T_137; // @[ifu_ifc_ctl.scala 131:17]
  wire  _T_139 = _T_138 | dma_stall; // @[ifu_ifc_ctl.scala 131:84]
  wire  _T_140 = io_ifc_fetch_req_bf_raw & _T_139; // @[ifu_ifc_ctl.scala 130:68]
  wire [31:0] _T_142 = {io_ifc_fetch_addr_bf,1'h0}; // @[Cat.scala 29:58]
  wire  iccm_acc_in_region_bf = _T_142[31:28] == 4'he; // @[lib.scala 84:47]
  wire  iccm_acc_in_range_bf = _T_142[31:16] == 16'hee00; // @[lib.scala 87:29]
  wire  _T_145 = ~io_ifc_iccm_access_bf; // @[ifu_ifc_ctl.scala 138:30]
  wire  _T_148 = fb_full_f & _T_36; // @[ifu_ifc_ctl.scala 139:16]
  wire  _T_149 = _T_145 | _T_148; // @[ifu_ifc_ctl.scala 138:53]
  wire  _T_150 = ~io_ifc_fetch_req_bf; // @[ifu_ifc_ctl.scala 140:13]
  wire  _T_151 = wfm & _T_150; // @[ifu_ifc_ctl.scala 140:11]
  wire  _T_152 = _T_149 | _T_151; // @[ifu_ifc_ctl.scala 139:62]
  wire  _T_153 = _T_152 | idle; // @[ifu_ifc_ctl.scala 140:35]
  wire  _T_155 = _T_153 & _T_2; // @[ifu_ifc_ctl.scala 140:44]
  wire  _T_157 = ~iccm_acc_in_range_bf; // @[ifu_ifc_ctl.scala 142:33]
  wire [4:0] _T_160 = {io_ifc_fetch_addr_bf[30:27],1'h0}; // @[Cat.scala 29:58]
  wire [31:0] _T_161 = io_dec_ifc_dec_tlu_mrac_ff >> _T_160; // @[ifu_ifc_ctl.scala 143:61]
  reg  _T_164; // @[ifu_ifc_ctl.scala 145:57]
  reg [30:0] _T_166; // @[lib.scala 374:16]
  rvclkhdr rvclkhdr ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_io_l1clk),
    .io_clk(rvclkhdr_io_clk),
    .io_en(rvclkhdr_io_en),
    .io_scan_mode(rvclkhdr_io_scan_mode)
  );
  assign io_dec_ifc_ifu_pmu_fetch_stall = wfm | _T_140; // @[ifu_ifc_ctl.scala 130:34]
  assign io_ifc_fetch_addr_f = _T_166; // @[ifu_ifc_ctl.scala 147:23]
  assign io_ifc_fetch_addr_bf = _T_22 | _T_20; // @[ifu_ifc_ctl.scala 73:24]
  assign io_ifc_fetch_req_f = _T_164; // @[ifu_ifc_ctl.scala 145:22]
  assign io_ifc_fetch_uncacheable_bf = ~_T_161[0]; // @[ifu_ifc_ctl.scala 143:31]
  assign io_ifc_fetch_req_bf = _T_41 & _T_44; // @[ifu_ifc_ctl.scala 86:23]
  assign io_ifc_fetch_req_bf_raw = ~idle; // @[ifu_ifc_ctl.scala 84:27]
  assign io_ifc_iccm_access_bf = _T_142[31:16] == 16'hee00; // @[ifu_ifc_ctl.scala 137:25]
  assign io_ifc_region_acc_fault_bf = _T_157 & iccm_acc_in_region_bf; // @[ifu_ifc_ctl.scala 142:30]
  assign io_ifc_dma_access_ok = _T_155 | dma_iccm_stall_any_f; // @[ifu_ifc_ctl.scala 138:24]
  assign rvclkhdr_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_io_en = io_exu_flush_final | io_ifc_fetch_req_f; // @[lib.scala 371:17]
  assign rvclkhdr_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  dma_iccm_stall_any_f = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  miss_a = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  state = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  fb_write_f = _RAND_3[3:0];
  _RAND_4 = {1{`RANDOM}};
  fb_full_f = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  _T_164 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  _T_166 = _RAND_6[30:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    dma_iccm_stall_any_f = 1'h0;
  end
  if (reset) begin
    miss_a = 1'h0;
  end
  if (reset) begin
    state = 2'h0;
  end
  if (reset) begin
    fb_write_f = 4'h0;
  end
  if (reset) begin
    fb_full_f = 1'h0;
  end
  if (reset) begin
    _T_164 = 1'h0;
  end
  if (reset) begin
    _T_166 = 31'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      dma_iccm_stall_any_f <= 1'h0;
    end else begin
      dma_iccm_stall_any_f <= io_dma_ifc_dma_iccm_stall_any;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      miss_a <= 1'h0;
    end else begin
      miss_a <= _T_48 & _T_2;
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      state <= 2'h0;
    end else begin
      state <= {next_state_1,next_state_0};
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      fb_write_f <= 4'h0;
    end else begin
      fb_write_f <= _T_128 | _T_125;
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      fb_full_f <= 1'h0;
    end else begin
      fb_full_f <= fb_write_ns[3];
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      _T_164 <= 1'h0;
    end else begin
      _T_164 <= io_ifc_fetch_req_bf;
    end
  end
  always @(posedge rvclkhdr_io_l1clk or posedge reset) begin
    if (reset) begin
      _T_166 <= 31'h0;
    end else begin
      _T_166 <= io_ifc_fetch_addr_bf;
    end
  end
endmodule
module ifu(
  input         clock,
  input         reset,
  input         io_exu_flush_final,
  input  [30:0] io_exu_flush_path_final,
  input         io_free_clk,
  input         io_active_clk,
  input         io_ifu_dec_dec_aln_aln_dec_dec_i0_decode_d,
  output [15:0] io_ifu_dec_dec_aln_aln_dec_ifu_i0_cinst,
  output        io_ifu_dec_dec_aln_aln_ib_ifu_i0_icaf,
  output [1:0]  io_ifu_dec_dec_aln_aln_ib_ifu_i0_icaf_type,
  output        io_ifu_dec_dec_aln_aln_ib_ifu_i0_icaf_f1,
  output        io_ifu_dec_dec_aln_aln_ib_ifu_i0_dbecc,
  output [7:0]  io_ifu_dec_dec_aln_aln_ib_ifu_i0_bp_index,
  output [7:0]  io_ifu_dec_dec_aln_aln_ib_ifu_i0_bp_fghr,
  output [4:0]  io_ifu_dec_dec_aln_aln_ib_ifu_i0_bp_btag,
  output        io_ifu_dec_dec_aln_aln_ib_ifu_i0_valid,
  output [31:0] io_ifu_dec_dec_aln_aln_ib_ifu_i0_instr,
  output [30:0] io_ifu_dec_dec_aln_aln_ib_ifu_i0_pc,
  output        io_ifu_dec_dec_aln_aln_ib_ifu_i0_pc4,
  output        io_ifu_dec_dec_aln_aln_ib_i0_brp_valid,
  output [11:0] io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_toffset,
  output [1:0]  io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_hist,
  output        io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_br_error,
  output        io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_br_start_error,
  output [30:0] io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_prett,
  output        io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_way,
  output        io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_ret,
  output        io_ifu_dec_dec_aln_ifu_pmu_instr_aligned,
  input         io_ifu_dec_dec_mem_ctrl_dec_tlu_flush_err_wb,
  input         io_ifu_dec_dec_mem_ctrl_dec_tlu_i0_commit_cmt,
  input         io_ifu_dec_dec_mem_ctrl_dec_tlu_force_halt,
  input         io_ifu_dec_dec_mem_ctrl_dec_tlu_fence_i_wb,
  input  [70:0] io_ifu_dec_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_wrdata,
  input  [16:0] io_ifu_dec_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_dicawics,
  input         io_ifu_dec_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_rd_valid,
  input         io_ifu_dec_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_wr_valid,
  input         io_ifu_dec_dec_mem_ctrl_dec_tlu_core_ecc_disable,
  output        io_ifu_dec_dec_mem_ctrl_ifu_pmu_ic_miss,
  output        io_ifu_dec_dec_mem_ctrl_ifu_pmu_ic_hit,
  output        io_ifu_dec_dec_mem_ctrl_ifu_pmu_bus_error,
  output        io_ifu_dec_dec_mem_ctrl_ifu_pmu_bus_busy,
  output        io_ifu_dec_dec_mem_ctrl_ifu_ic_error_start,
  output        io_ifu_dec_dec_mem_ctrl_ifu_iccm_rd_ecc_single_err,
  output [70:0] io_ifu_dec_dec_mem_ctrl_ifu_ic_debug_rd_data,
  output        io_ifu_dec_dec_mem_ctrl_ifu_ic_debug_rd_data_valid,
  output        io_ifu_dec_dec_mem_ctrl_ifu_miss_state_idle,
  input         io_ifu_dec_dec_ifc_dec_tlu_flush_noredir_wb,
  input  [31:0] io_ifu_dec_dec_ifc_dec_tlu_mrac_ff,
  output        io_ifu_dec_dec_ifc_ifu_pmu_fetch_stall,
  input         io_ifu_dec_dec_bp_dec_tlu_br0_r_pkt_valid,
  input  [1:0]  io_ifu_dec_dec_bp_dec_tlu_br0_r_pkt_bits_hist,
  input         io_ifu_dec_dec_bp_dec_tlu_br0_r_pkt_bits_br_error,
  input         io_ifu_dec_dec_bp_dec_tlu_br0_r_pkt_bits_br_start_error,
  input         io_ifu_dec_dec_bp_dec_tlu_br0_r_pkt_bits_way,
  input         io_ifu_dec_dec_bp_dec_tlu_br0_r_pkt_bits_middle,
  input         io_ifu_dec_dec_bp_dec_tlu_flush_leak_one_wb,
  input         io_ifu_dec_dec_bp_dec_tlu_bpred_disable,
  input  [7:0]  io_exu_ifu_exu_bp_exu_i0_br_index_r,
  input  [7:0]  io_exu_ifu_exu_bp_exu_i0_br_fghr_r,
  input         io_exu_ifu_exu_bp_exu_mp_pkt_bits_misp,
  input         io_exu_ifu_exu_bp_exu_mp_pkt_bits_ataken,
  input         io_exu_ifu_exu_bp_exu_mp_pkt_bits_boffset,
  input         io_exu_ifu_exu_bp_exu_mp_pkt_bits_pc4,
  input  [1:0]  io_exu_ifu_exu_bp_exu_mp_pkt_bits_hist,
  input  [11:0] io_exu_ifu_exu_bp_exu_mp_pkt_bits_toffset,
  input         io_exu_ifu_exu_bp_exu_mp_pkt_bits_pcall,
  input         io_exu_ifu_exu_bp_exu_mp_pkt_bits_pret,
  input         io_exu_ifu_exu_bp_exu_mp_pkt_bits_pja,
  input         io_exu_ifu_exu_bp_exu_mp_pkt_bits_way,
  input  [7:0]  io_exu_ifu_exu_bp_exu_mp_eghr,
  input  [7:0]  io_exu_ifu_exu_bp_exu_mp_fghr,
  input  [7:0]  io_exu_ifu_exu_bp_exu_mp_index,
  input  [4:0]  io_exu_ifu_exu_bp_exu_mp_btag,
  output [14:0] io_iccm_rw_addr,
  output        io_iccm_buf_correct_ecc,
  output        io_iccm_correction_state,
  output        io_iccm_wren,
  output        io_iccm_rden,
  output [2:0]  io_iccm_wr_size,
  output [77:0] io_iccm_wr_data,
  input  [63:0] io_iccm_rd_data,
  input  [77:0] io_iccm_rd_data_ecc,
  output [30:0] io_ic_rw_addr,
  output [1:0]  io_ic_tag_valid,
  output        io_ic_rd_en,
  output [70:0] io_ic_debug_wr_data,
  output [9:0]  io_ic_debug_addr,
  input  [63:0] io_ic_rd_data,
  input  [70:0] io_ic_debug_rd_data,
  input  [25:0] io_ic_tag_debug_rd_data,
  input  [1:0]  io_ic_eccerr,
  input  [1:0]  io_ic_rd_hit,
  input         io_ic_tag_perr,
  output        io_ic_debug_rd_en,
  output        io_ic_debug_wr_en,
  output        io_ic_debug_tag_array,
  output [1:0]  io_ic_debug_way,
  output [63:0] io_ic_premux_data,
  output        io_ic_sel_premux_data,
  output        io_ifu_ar_valid,
  output [31:0] io_ifu_ar_bits_addr,
  input         io_ifu_bus_clk_en,
  input         io_ifu_dma_dma_ifc_dma_iccm_stall_any,
  input         io_ifu_dma_dma_mem_ctl_dma_iccm_req,
  input  [31:0] io_ifu_dma_dma_mem_ctl_dma_mem_addr,
  input  [2:0]  io_ifu_dma_dma_mem_ctl_dma_mem_sz,
  input         io_ifu_dma_dma_mem_ctl_dma_mem_write,
  input  [63:0] io_ifu_dma_dma_mem_ctl_dma_mem_wdata,
  input  [2:0]  io_ifu_dma_dma_mem_ctl_dma_mem_tag,
  output        io_iccm_dma_ecc_error,
  output        io_iccm_dma_rvalid,
  output [63:0] io_iccm_dma_rdata,
  output [2:0]  io_iccm_dma_rtag,
  output        io_iccm_ready,
  output        io_iccm_dma_sb_error,
  input         io_dec_tlu_flush_lower_wb,
  input         io_scan_mode
);
  wire  mem_ctl_clock; // @[ifu.scala 34:23]
  wire  mem_ctl_reset; // @[ifu.scala 34:23]
  wire  mem_ctl_io_free_clk; // @[ifu.scala 34:23]
  wire  mem_ctl_io_active_clk; // @[ifu.scala 34:23]
  wire  mem_ctl_io_exu_flush_final; // @[ifu.scala 34:23]
  wire  mem_ctl_io_dec_mem_ctrl_dec_tlu_flush_err_wb; // @[ifu.scala 34:23]
  wire  mem_ctl_io_dec_mem_ctrl_dec_tlu_i0_commit_cmt; // @[ifu.scala 34:23]
  wire  mem_ctl_io_dec_mem_ctrl_dec_tlu_force_halt; // @[ifu.scala 34:23]
  wire  mem_ctl_io_dec_mem_ctrl_dec_tlu_fence_i_wb; // @[ifu.scala 34:23]
  wire [70:0] mem_ctl_io_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_wrdata; // @[ifu.scala 34:23]
  wire [16:0] mem_ctl_io_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_dicawics; // @[ifu.scala 34:23]
  wire  mem_ctl_io_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_rd_valid; // @[ifu.scala 34:23]
  wire  mem_ctl_io_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_wr_valid; // @[ifu.scala 34:23]
  wire  mem_ctl_io_dec_mem_ctrl_dec_tlu_core_ecc_disable; // @[ifu.scala 34:23]
  wire  mem_ctl_io_dec_mem_ctrl_ifu_pmu_ic_miss; // @[ifu.scala 34:23]
  wire  mem_ctl_io_dec_mem_ctrl_ifu_pmu_ic_hit; // @[ifu.scala 34:23]
  wire  mem_ctl_io_dec_mem_ctrl_ifu_pmu_bus_error; // @[ifu.scala 34:23]
  wire  mem_ctl_io_dec_mem_ctrl_ifu_pmu_bus_busy; // @[ifu.scala 34:23]
  wire  mem_ctl_io_dec_mem_ctrl_ifu_ic_error_start; // @[ifu.scala 34:23]
  wire  mem_ctl_io_dec_mem_ctrl_ifu_iccm_rd_ecc_single_err; // @[ifu.scala 34:23]
  wire [70:0] mem_ctl_io_dec_mem_ctrl_ifu_ic_debug_rd_data; // @[ifu.scala 34:23]
  wire  mem_ctl_io_dec_mem_ctrl_ifu_ic_debug_rd_data_valid; // @[ifu.scala 34:23]
  wire  mem_ctl_io_dec_mem_ctrl_ifu_miss_state_idle; // @[ifu.scala 34:23]
  wire [30:0] mem_ctl_io_ifc_fetch_addr_bf; // @[ifu.scala 34:23]
  wire  mem_ctl_io_ifc_fetch_uncacheable_bf; // @[ifu.scala 34:23]
  wire  mem_ctl_io_ifc_fetch_req_bf; // @[ifu.scala 34:23]
  wire  mem_ctl_io_ifc_fetch_req_bf_raw; // @[ifu.scala 34:23]
  wire  mem_ctl_io_ifc_iccm_access_bf; // @[ifu.scala 34:23]
  wire  mem_ctl_io_ifc_region_acc_fault_bf; // @[ifu.scala 34:23]
  wire  mem_ctl_io_ifc_dma_access_ok; // @[ifu.scala 34:23]
  wire  mem_ctl_io_ifu_bp_hit_taken_f; // @[ifu.scala 34:23]
  wire  mem_ctl_io_ifu_bp_inst_mask_f; // @[ifu.scala 34:23]
  wire  mem_ctl_io_ifu_axi_ar_valid; // @[ifu.scala 34:23]
  wire [31:0] mem_ctl_io_ifu_axi_ar_bits_addr; // @[ifu.scala 34:23]
  wire  mem_ctl_io_ifu_bus_clk_en; // @[ifu.scala 34:23]
  wire  mem_ctl_io_dma_mem_ctl_dma_iccm_req; // @[ifu.scala 34:23]
  wire [31:0] mem_ctl_io_dma_mem_ctl_dma_mem_addr; // @[ifu.scala 34:23]
  wire [2:0] mem_ctl_io_dma_mem_ctl_dma_mem_sz; // @[ifu.scala 34:23]
  wire  mem_ctl_io_dma_mem_ctl_dma_mem_write; // @[ifu.scala 34:23]
  wire [63:0] mem_ctl_io_dma_mem_ctl_dma_mem_wdata; // @[ifu.scala 34:23]
  wire [2:0] mem_ctl_io_dma_mem_ctl_dma_mem_tag; // @[ifu.scala 34:23]
  wire [14:0] mem_ctl_io_iccm_rw_addr; // @[ifu.scala 34:23]
  wire  mem_ctl_io_iccm_buf_correct_ecc; // @[ifu.scala 34:23]
  wire  mem_ctl_io_iccm_correction_state; // @[ifu.scala 34:23]
  wire  mem_ctl_io_iccm_wren; // @[ifu.scala 34:23]
  wire  mem_ctl_io_iccm_rden; // @[ifu.scala 34:23]
  wire [2:0] mem_ctl_io_iccm_wr_size; // @[ifu.scala 34:23]
  wire [77:0] mem_ctl_io_iccm_wr_data; // @[ifu.scala 34:23]
  wire [63:0] mem_ctl_io_iccm_rd_data; // @[ifu.scala 34:23]
  wire [77:0] mem_ctl_io_iccm_rd_data_ecc; // @[ifu.scala 34:23]
  wire [30:0] mem_ctl_io_ic_rw_addr; // @[ifu.scala 34:23]
  wire [1:0] mem_ctl_io_ic_tag_valid; // @[ifu.scala 34:23]
  wire  mem_ctl_io_ic_rd_en; // @[ifu.scala 34:23]
  wire [70:0] mem_ctl_io_ic_debug_wr_data; // @[ifu.scala 34:23]
  wire [9:0] mem_ctl_io_ic_debug_addr; // @[ifu.scala 34:23]
  wire [63:0] mem_ctl_io_ic_rd_data; // @[ifu.scala 34:23]
  wire [70:0] mem_ctl_io_ic_debug_rd_data; // @[ifu.scala 34:23]
  wire [25:0] mem_ctl_io_ic_tag_debug_rd_data; // @[ifu.scala 34:23]
  wire [1:0] mem_ctl_io_ic_eccerr; // @[ifu.scala 34:23]
  wire [1:0] mem_ctl_io_ic_rd_hit; // @[ifu.scala 34:23]
  wire  mem_ctl_io_ic_tag_perr; // @[ifu.scala 34:23]
  wire  mem_ctl_io_ic_debug_rd_en; // @[ifu.scala 34:23]
  wire  mem_ctl_io_ic_debug_wr_en; // @[ifu.scala 34:23]
  wire  mem_ctl_io_ic_debug_tag_array; // @[ifu.scala 34:23]
  wire [1:0] mem_ctl_io_ic_debug_way; // @[ifu.scala 34:23]
  wire [63:0] mem_ctl_io_ic_premux_data; // @[ifu.scala 34:23]
  wire  mem_ctl_io_ic_sel_premux_data; // @[ifu.scala 34:23]
  wire [1:0] mem_ctl_io_ifu_fetch_val; // @[ifu.scala 34:23]
  wire  mem_ctl_io_ifu_ic_mb_empty; // @[ifu.scala 34:23]
  wire  mem_ctl_io_ic_dma_active; // @[ifu.scala 34:23]
  wire  mem_ctl_io_iccm_dma_ecc_error; // @[ifu.scala 34:23]
  wire  mem_ctl_io_iccm_dma_rvalid; // @[ifu.scala 34:23]
  wire [63:0] mem_ctl_io_iccm_dma_rdata; // @[ifu.scala 34:23]
  wire [2:0] mem_ctl_io_iccm_dma_rtag; // @[ifu.scala 34:23]
  wire  mem_ctl_io_iccm_ready; // @[ifu.scala 34:23]
  wire  mem_ctl_io_dec_tlu_flush_lower_wb; // @[ifu.scala 34:23]
  wire  mem_ctl_io_iccm_rd_ecc_double_err; // @[ifu.scala 34:23]
  wire  mem_ctl_io_iccm_dma_sb_error; // @[ifu.scala 34:23]
  wire  mem_ctl_io_ic_hit_f; // @[ifu.scala 34:23]
  wire  mem_ctl_io_ic_access_fault_f; // @[ifu.scala 34:23]
  wire [1:0] mem_ctl_io_ic_access_fault_type_f; // @[ifu.scala 34:23]
  wire  mem_ctl_io_ifu_async_error_start; // @[ifu.scala 34:23]
  wire [1:0] mem_ctl_io_ic_fetch_val_f; // @[ifu.scala 34:23]
  wire [31:0] mem_ctl_io_ic_data_f; // @[ifu.scala 34:23]
  wire  mem_ctl_io_scan_mode; // @[ifu.scala 34:23]
  wire  bp_ctl_clock; // @[ifu.scala 35:22]
  wire  bp_ctl_reset; // @[ifu.scala 35:22]
  wire  bp_ctl_io_active_clk; // @[ifu.scala 35:22]
  wire  bp_ctl_io_ic_hit_f; // @[ifu.scala 35:22]
  wire  bp_ctl_io_exu_flush_final; // @[ifu.scala 35:22]
  wire [30:0] bp_ctl_io_ifc_fetch_addr_f; // @[ifu.scala 35:22]
  wire  bp_ctl_io_ifc_fetch_req_f; // @[ifu.scala 35:22]
  wire  bp_ctl_io_dec_bp_dec_tlu_br0_r_pkt_valid; // @[ifu.scala 35:22]
  wire [1:0] bp_ctl_io_dec_bp_dec_tlu_br0_r_pkt_bits_hist; // @[ifu.scala 35:22]
  wire  bp_ctl_io_dec_bp_dec_tlu_br0_r_pkt_bits_br_error; // @[ifu.scala 35:22]
  wire  bp_ctl_io_dec_bp_dec_tlu_br0_r_pkt_bits_br_start_error; // @[ifu.scala 35:22]
  wire  bp_ctl_io_dec_bp_dec_tlu_br0_r_pkt_bits_way; // @[ifu.scala 35:22]
  wire  bp_ctl_io_dec_bp_dec_tlu_br0_r_pkt_bits_middle; // @[ifu.scala 35:22]
  wire  bp_ctl_io_dec_bp_dec_tlu_flush_leak_one_wb; // @[ifu.scala 35:22]
  wire  bp_ctl_io_dec_bp_dec_tlu_bpred_disable; // @[ifu.scala 35:22]
  wire  bp_ctl_io_dec_tlu_flush_lower_wb; // @[ifu.scala 35:22]
  wire [7:0] bp_ctl_io_exu_bp_exu_i0_br_index_r; // @[ifu.scala 35:22]
  wire [7:0] bp_ctl_io_exu_bp_exu_i0_br_fghr_r; // @[ifu.scala 35:22]
  wire  bp_ctl_io_exu_bp_exu_mp_pkt_bits_misp; // @[ifu.scala 35:22]
  wire  bp_ctl_io_exu_bp_exu_mp_pkt_bits_ataken; // @[ifu.scala 35:22]
  wire  bp_ctl_io_exu_bp_exu_mp_pkt_bits_boffset; // @[ifu.scala 35:22]
  wire  bp_ctl_io_exu_bp_exu_mp_pkt_bits_pc4; // @[ifu.scala 35:22]
  wire [1:0] bp_ctl_io_exu_bp_exu_mp_pkt_bits_hist; // @[ifu.scala 35:22]
  wire [11:0] bp_ctl_io_exu_bp_exu_mp_pkt_bits_toffset; // @[ifu.scala 35:22]
  wire  bp_ctl_io_exu_bp_exu_mp_pkt_bits_pcall; // @[ifu.scala 35:22]
  wire  bp_ctl_io_exu_bp_exu_mp_pkt_bits_pret; // @[ifu.scala 35:22]
  wire  bp_ctl_io_exu_bp_exu_mp_pkt_bits_pja; // @[ifu.scala 35:22]
  wire  bp_ctl_io_exu_bp_exu_mp_pkt_bits_way; // @[ifu.scala 35:22]
  wire [7:0] bp_ctl_io_exu_bp_exu_mp_eghr; // @[ifu.scala 35:22]
  wire [7:0] bp_ctl_io_exu_bp_exu_mp_fghr; // @[ifu.scala 35:22]
  wire [7:0] bp_ctl_io_exu_bp_exu_mp_index; // @[ifu.scala 35:22]
  wire [4:0] bp_ctl_io_exu_bp_exu_mp_btag; // @[ifu.scala 35:22]
  wire  bp_ctl_io_ifu_bp_hit_taken_f; // @[ifu.scala 35:22]
  wire [30:0] bp_ctl_io_ifu_bp_btb_target_f; // @[ifu.scala 35:22]
  wire  bp_ctl_io_ifu_bp_inst_mask_f; // @[ifu.scala 35:22]
  wire [7:0] bp_ctl_io_ifu_bp_fghr_f; // @[ifu.scala 35:22]
  wire [1:0] bp_ctl_io_ifu_bp_way_f; // @[ifu.scala 35:22]
  wire [1:0] bp_ctl_io_ifu_bp_ret_f; // @[ifu.scala 35:22]
  wire [1:0] bp_ctl_io_ifu_bp_hist1_f; // @[ifu.scala 35:22]
  wire [1:0] bp_ctl_io_ifu_bp_hist0_f; // @[ifu.scala 35:22]
  wire [1:0] bp_ctl_io_ifu_bp_pc4_f; // @[ifu.scala 35:22]
  wire [1:0] bp_ctl_io_ifu_bp_valid_f; // @[ifu.scala 35:22]
  wire [11:0] bp_ctl_io_ifu_bp_poffset_f; // @[ifu.scala 35:22]
  wire  bp_ctl_io_scan_mode; // @[ifu.scala 35:22]
  wire  aln_ctl_clock; // @[ifu.scala 36:23]
  wire  aln_ctl_reset; // @[ifu.scala 36:23]
  wire  aln_ctl_io_scan_mode; // @[ifu.scala 36:23]
  wire  aln_ctl_io_active_clk; // @[ifu.scala 36:23]
  wire  aln_ctl_io_ifu_async_error_start; // @[ifu.scala 36:23]
  wire  aln_ctl_io_iccm_rd_ecc_double_err; // @[ifu.scala 36:23]
  wire  aln_ctl_io_ic_access_fault_f; // @[ifu.scala 36:23]
  wire [1:0] aln_ctl_io_ic_access_fault_type_f; // @[ifu.scala 36:23]
  wire [7:0] aln_ctl_io_ifu_bp_fghr_f; // @[ifu.scala 36:23]
  wire [30:0] aln_ctl_io_ifu_bp_btb_target_f; // @[ifu.scala 36:23]
  wire [11:0] aln_ctl_io_ifu_bp_poffset_f; // @[ifu.scala 36:23]
  wire [1:0] aln_ctl_io_ifu_bp_hist0_f; // @[ifu.scala 36:23]
  wire [1:0] aln_ctl_io_ifu_bp_hist1_f; // @[ifu.scala 36:23]
  wire [1:0] aln_ctl_io_ifu_bp_pc4_f; // @[ifu.scala 36:23]
  wire [1:0] aln_ctl_io_ifu_bp_way_f; // @[ifu.scala 36:23]
  wire [1:0] aln_ctl_io_ifu_bp_valid_f; // @[ifu.scala 36:23]
  wire [1:0] aln_ctl_io_ifu_bp_ret_f; // @[ifu.scala 36:23]
  wire  aln_ctl_io_exu_flush_final; // @[ifu.scala 36:23]
  wire  aln_ctl_io_dec_aln_aln_dec_dec_i0_decode_d; // @[ifu.scala 36:23]
  wire [15:0] aln_ctl_io_dec_aln_aln_dec_ifu_i0_cinst; // @[ifu.scala 36:23]
  wire  aln_ctl_io_dec_aln_aln_ib_ifu_i0_icaf; // @[ifu.scala 36:23]
  wire [1:0] aln_ctl_io_dec_aln_aln_ib_ifu_i0_icaf_type; // @[ifu.scala 36:23]
  wire  aln_ctl_io_dec_aln_aln_ib_ifu_i0_icaf_f1; // @[ifu.scala 36:23]
  wire  aln_ctl_io_dec_aln_aln_ib_ifu_i0_dbecc; // @[ifu.scala 36:23]
  wire [7:0] aln_ctl_io_dec_aln_aln_ib_ifu_i0_bp_index; // @[ifu.scala 36:23]
  wire [7:0] aln_ctl_io_dec_aln_aln_ib_ifu_i0_bp_fghr; // @[ifu.scala 36:23]
  wire [4:0] aln_ctl_io_dec_aln_aln_ib_ifu_i0_bp_btag; // @[ifu.scala 36:23]
  wire  aln_ctl_io_dec_aln_aln_ib_ifu_i0_valid; // @[ifu.scala 36:23]
  wire [31:0] aln_ctl_io_dec_aln_aln_ib_ifu_i0_instr; // @[ifu.scala 36:23]
  wire [30:0] aln_ctl_io_dec_aln_aln_ib_ifu_i0_pc; // @[ifu.scala 36:23]
  wire  aln_ctl_io_dec_aln_aln_ib_ifu_i0_pc4; // @[ifu.scala 36:23]
  wire  aln_ctl_io_dec_aln_aln_ib_i0_brp_valid; // @[ifu.scala 36:23]
  wire [11:0] aln_ctl_io_dec_aln_aln_ib_i0_brp_bits_toffset; // @[ifu.scala 36:23]
  wire [1:0] aln_ctl_io_dec_aln_aln_ib_i0_brp_bits_hist; // @[ifu.scala 36:23]
  wire  aln_ctl_io_dec_aln_aln_ib_i0_brp_bits_br_error; // @[ifu.scala 36:23]
  wire  aln_ctl_io_dec_aln_aln_ib_i0_brp_bits_br_start_error; // @[ifu.scala 36:23]
  wire [30:0] aln_ctl_io_dec_aln_aln_ib_i0_brp_bits_prett; // @[ifu.scala 36:23]
  wire  aln_ctl_io_dec_aln_aln_ib_i0_brp_bits_way; // @[ifu.scala 36:23]
  wire  aln_ctl_io_dec_aln_aln_ib_i0_brp_bits_ret; // @[ifu.scala 36:23]
  wire  aln_ctl_io_dec_aln_ifu_pmu_instr_aligned; // @[ifu.scala 36:23]
  wire [31:0] aln_ctl_io_ifu_fetch_data_f; // @[ifu.scala 36:23]
  wire [1:0] aln_ctl_io_ifu_fetch_val; // @[ifu.scala 36:23]
  wire [30:0] aln_ctl_io_ifu_fetch_pc; // @[ifu.scala 36:23]
  wire  aln_ctl_io_ifu_fb_consume1; // @[ifu.scala 36:23]
  wire  aln_ctl_io_ifu_fb_consume2; // @[ifu.scala 36:23]
  wire  ifc_ctl_clock; // @[ifu.scala 37:23]
  wire  ifc_ctl_reset; // @[ifu.scala 37:23]
  wire  ifc_ctl_io_exu_flush_final; // @[ifu.scala 37:23]
  wire [30:0] ifc_ctl_io_exu_flush_path_final; // @[ifu.scala 37:23]
  wire  ifc_ctl_io_free_clk; // @[ifu.scala 37:23]
  wire  ifc_ctl_io_active_clk; // @[ifu.scala 37:23]
  wire  ifc_ctl_io_scan_mode; // @[ifu.scala 37:23]
  wire  ifc_ctl_io_ic_hit_f; // @[ifu.scala 37:23]
  wire  ifc_ctl_io_ifu_ic_mb_empty; // @[ifu.scala 37:23]
  wire  ifc_ctl_io_ifu_fb_consume1; // @[ifu.scala 37:23]
  wire  ifc_ctl_io_ifu_fb_consume2; // @[ifu.scala 37:23]
  wire  ifc_ctl_io_ifu_bp_hit_taken_f; // @[ifu.scala 37:23]
  wire [30:0] ifc_ctl_io_ifu_bp_btb_target_f; // @[ifu.scala 37:23]
  wire  ifc_ctl_io_ic_dma_active; // @[ifu.scala 37:23]
  wire  ifc_ctl_io_dec_ifc_dec_tlu_flush_noredir_wb; // @[ifu.scala 37:23]
  wire [31:0] ifc_ctl_io_dec_ifc_dec_tlu_mrac_ff; // @[ifu.scala 37:23]
  wire  ifc_ctl_io_dec_ifc_ifu_pmu_fetch_stall; // @[ifu.scala 37:23]
  wire  ifc_ctl_io_dma_ifc_dma_iccm_stall_any; // @[ifu.scala 37:23]
  wire [30:0] ifc_ctl_io_ifc_fetch_addr_f; // @[ifu.scala 37:23]
  wire [30:0] ifc_ctl_io_ifc_fetch_addr_bf; // @[ifu.scala 37:23]
  wire  ifc_ctl_io_ifc_fetch_req_f; // @[ifu.scala 37:23]
  wire  ifc_ctl_io_ifc_fetch_uncacheable_bf; // @[ifu.scala 37:23]
  wire  ifc_ctl_io_ifc_fetch_req_bf; // @[ifu.scala 37:23]
  wire  ifc_ctl_io_ifc_fetch_req_bf_raw; // @[ifu.scala 37:23]
  wire  ifc_ctl_io_ifc_iccm_access_bf; // @[ifu.scala 37:23]
  wire  ifc_ctl_io_ifc_region_acc_fault_bf; // @[ifu.scala 37:23]
  wire  ifc_ctl_io_ifc_dma_access_ok; // @[ifu.scala 37:23]
  ifu_mem_ctl mem_ctl ( // @[ifu.scala 34:23]
    .clock(mem_ctl_clock),
    .reset(mem_ctl_reset),
    .io_free_clk(mem_ctl_io_free_clk),
    .io_active_clk(mem_ctl_io_active_clk),
    .io_exu_flush_final(mem_ctl_io_exu_flush_final),
    .io_dec_mem_ctrl_dec_tlu_flush_err_wb(mem_ctl_io_dec_mem_ctrl_dec_tlu_flush_err_wb),
    .io_dec_mem_ctrl_dec_tlu_i0_commit_cmt(mem_ctl_io_dec_mem_ctrl_dec_tlu_i0_commit_cmt),
    .io_dec_mem_ctrl_dec_tlu_force_halt(mem_ctl_io_dec_mem_ctrl_dec_tlu_force_halt),
    .io_dec_mem_ctrl_dec_tlu_fence_i_wb(mem_ctl_io_dec_mem_ctrl_dec_tlu_fence_i_wb),
    .io_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_wrdata(mem_ctl_io_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_wrdata),
    .io_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_dicawics(mem_ctl_io_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_dicawics),
    .io_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_rd_valid(mem_ctl_io_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_rd_valid),
    .io_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_wr_valid(mem_ctl_io_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_wr_valid),
    .io_dec_mem_ctrl_dec_tlu_core_ecc_disable(mem_ctl_io_dec_mem_ctrl_dec_tlu_core_ecc_disable),
    .io_dec_mem_ctrl_ifu_pmu_ic_miss(mem_ctl_io_dec_mem_ctrl_ifu_pmu_ic_miss),
    .io_dec_mem_ctrl_ifu_pmu_ic_hit(mem_ctl_io_dec_mem_ctrl_ifu_pmu_ic_hit),
    .io_dec_mem_ctrl_ifu_pmu_bus_error(mem_ctl_io_dec_mem_ctrl_ifu_pmu_bus_error),
    .io_dec_mem_ctrl_ifu_pmu_bus_busy(mem_ctl_io_dec_mem_ctrl_ifu_pmu_bus_busy),
    .io_dec_mem_ctrl_ifu_ic_error_start(mem_ctl_io_dec_mem_ctrl_ifu_ic_error_start),
    .io_dec_mem_ctrl_ifu_iccm_rd_ecc_single_err(mem_ctl_io_dec_mem_ctrl_ifu_iccm_rd_ecc_single_err),
    .io_dec_mem_ctrl_ifu_ic_debug_rd_data(mem_ctl_io_dec_mem_ctrl_ifu_ic_debug_rd_data),
    .io_dec_mem_ctrl_ifu_ic_debug_rd_data_valid(mem_ctl_io_dec_mem_ctrl_ifu_ic_debug_rd_data_valid),
    .io_dec_mem_ctrl_ifu_miss_state_idle(mem_ctl_io_dec_mem_ctrl_ifu_miss_state_idle),
    .io_ifc_fetch_addr_bf(mem_ctl_io_ifc_fetch_addr_bf),
    .io_ifc_fetch_uncacheable_bf(mem_ctl_io_ifc_fetch_uncacheable_bf),
    .io_ifc_fetch_req_bf(mem_ctl_io_ifc_fetch_req_bf),
    .io_ifc_fetch_req_bf_raw(mem_ctl_io_ifc_fetch_req_bf_raw),
    .io_ifc_iccm_access_bf(mem_ctl_io_ifc_iccm_access_bf),
    .io_ifc_region_acc_fault_bf(mem_ctl_io_ifc_region_acc_fault_bf),
    .io_ifc_dma_access_ok(mem_ctl_io_ifc_dma_access_ok),
    .io_ifu_bp_hit_taken_f(mem_ctl_io_ifu_bp_hit_taken_f),
    .io_ifu_bp_inst_mask_f(mem_ctl_io_ifu_bp_inst_mask_f),
    .io_ifu_axi_ar_valid(mem_ctl_io_ifu_axi_ar_valid),
    .io_ifu_axi_ar_bits_addr(mem_ctl_io_ifu_axi_ar_bits_addr),
    .io_ifu_bus_clk_en(mem_ctl_io_ifu_bus_clk_en),
    .io_dma_mem_ctl_dma_iccm_req(mem_ctl_io_dma_mem_ctl_dma_iccm_req),
    .io_dma_mem_ctl_dma_mem_addr(mem_ctl_io_dma_mem_ctl_dma_mem_addr),
    .io_dma_mem_ctl_dma_mem_sz(mem_ctl_io_dma_mem_ctl_dma_mem_sz),
    .io_dma_mem_ctl_dma_mem_write(mem_ctl_io_dma_mem_ctl_dma_mem_write),
    .io_dma_mem_ctl_dma_mem_wdata(mem_ctl_io_dma_mem_ctl_dma_mem_wdata),
    .io_dma_mem_ctl_dma_mem_tag(mem_ctl_io_dma_mem_ctl_dma_mem_tag),
    .io_iccm_rw_addr(mem_ctl_io_iccm_rw_addr),
    .io_iccm_buf_correct_ecc(mem_ctl_io_iccm_buf_correct_ecc),
    .io_iccm_correction_state(mem_ctl_io_iccm_correction_state),
    .io_iccm_wren(mem_ctl_io_iccm_wren),
    .io_iccm_rden(mem_ctl_io_iccm_rden),
    .io_iccm_wr_size(mem_ctl_io_iccm_wr_size),
    .io_iccm_wr_data(mem_ctl_io_iccm_wr_data),
    .io_iccm_rd_data(mem_ctl_io_iccm_rd_data),
    .io_iccm_rd_data_ecc(mem_ctl_io_iccm_rd_data_ecc),
    .io_ic_rw_addr(mem_ctl_io_ic_rw_addr),
    .io_ic_tag_valid(mem_ctl_io_ic_tag_valid),
    .io_ic_rd_en(mem_ctl_io_ic_rd_en),
    .io_ic_debug_wr_data(mem_ctl_io_ic_debug_wr_data),
    .io_ic_debug_addr(mem_ctl_io_ic_debug_addr),
    .io_ic_rd_data(mem_ctl_io_ic_rd_data),
    .io_ic_debug_rd_data(mem_ctl_io_ic_debug_rd_data),
    .io_ic_tag_debug_rd_data(mem_ctl_io_ic_tag_debug_rd_data),
    .io_ic_eccerr(mem_ctl_io_ic_eccerr),
    .io_ic_rd_hit(mem_ctl_io_ic_rd_hit),
    .io_ic_tag_perr(mem_ctl_io_ic_tag_perr),
    .io_ic_debug_rd_en(mem_ctl_io_ic_debug_rd_en),
    .io_ic_debug_wr_en(mem_ctl_io_ic_debug_wr_en),
    .io_ic_debug_tag_array(mem_ctl_io_ic_debug_tag_array),
    .io_ic_debug_way(mem_ctl_io_ic_debug_way),
    .io_ic_premux_data(mem_ctl_io_ic_premux_data),
    .io_ic_sel_premux_data(mem_ctl_io_ic_sel_premux_data),
    .io_ifu_fetch_val(mem_ctl_io_ifu_fetch_val),
    .io_ifu_ic_mb_empty(mem_ctl_io_ifu_ic_mb_empty),
    .io_ic_dma_active(mem_ctl_io_ic_dma_active),
    .io_iccm_dma_ecc_error(mem_ctl_io_iccm_dma_ecc_error),
    .io_iccm_dma_rvalid(mem_ctl_io_iccm_dma_rvalid),
    .io_iccm_dma_rdata(mem_ctl_io_iccm_dma_rdata),
    .io_iccm_dma_rtag(mem_ctl_io_iccm_dma_rtag),
    .io_iccm_ready(mem_ctl_io_iccm_ready),
    .io_dec_tlu_flush_lower_wb(mem_ctl_io_dec_tlu_flush_lower_wb),
    .io_iccm_rd_ecc_double_err(mem_ctl_io_iccm_rd_ecc_double_err),
    .io_iccm_dma_sb_error(mem_ctl_io_iccm_dma_sb_error),
    .io_ic_hit_f(mem_ctl_io_ic_hit_f),
    .io_ic_access_fault_f(mem_ctl_io_ic_access_fault_f),
    .io_ic_access_fault_type_f(mem_ctl_io_ic_access_fault_type_f),
    .io_ifu_async_error_start(mem_ctl_io_ifu_async_error_start),
    .io_ic_fetch_val_f(mem_ctl_io_ic_fetch_val_f),
    .io_ic_data_f(mem_ctl_io_ic_data_f),
    .io_scan_mode(mem_ctl_io_scan_mode)
  );
  ifu_bp_ctl bp_ctl ( // @[ifu.scala 35:22]
    .clock(bp_ctl_clock),
    .reset(bp_ctl_reset),
    .io_active_clk(bp_ctl_io_active_clk),
    .io_ic_hit_f(bp_ctl_io_ic_hit_f),
    .io_exu_flush_final(bp_ctl_io_exu_flush_final),
    .io_ifc_fetch_addr_f(bp_ctl_io_ifc_fetch_addr_f),
    .io_ifc_fetch_req_f(bp_ctl_io_ifc_fetch_req_f),
    .io_dec_bp_dec_tlu_br0_r_pkt_valid(bp_ctl_io_dec_bp_dec_tlu_br0_r_pkt_valid),
    .io_dec_bp_dec_tlu_br0_r_pkt_bits_hist(bp_ctl_io_dec_bp_dec_tlu_br0_r_pkt_bits_hist),
    .io_dec_bp_dec_tlu_br0_r_pkt_bits_br_error(bp_ctl_io_dec_bp_dec_tlu_br0_r_pkt_bits_br_error),
    .io_dec_bp_dec_tlu_br0_r_pkt_bits_br_start_error(bp_ctl_io_dec_bp_dec_tlu_br0_r_pkt_bits_br_start_error),
    .io_dec_bp_dec_tlu_br0_r_pkt_bits_way(bp_ctl_io_dec_bp_dec_tlu_br0_r_pkt_bits_way),
    .io_dec_bp_dec_tlu_br0_r_pkt_bits_middle(bp_ctl_io_dec_bp_dec_tlu_br0_r_pkt_bits_middle),
    .io_dec_bp_dec_tlu_flush_leak_one_wb(bp_ctl_io_dec_bp_dec_tlu_flush_leak_one_wb),
    .io_dec_bp_dec_tlu_bpred_disable(bp_ctl_io_dec_bp_dec_tlu_bpred_disable),
    .io_dec_tlu_flush_lower_wb(bp_ctl_io_dec_tlu_flush_lower_wb),
    .io_exu_bp_exu_i0_br_index_r(bp_ctl_io_exu_bp_exu_i0_br_index_r),
    .io_exu_bp_exu_i0_br_fghr_r(bp_ctl_io_exu_bp_exu_i0_br_fghr_r),
    .io_exu_bp_exu_mp_pkt_bits_misp(bp_ctl_io_exu_bp_exu_mp_pkt_bits_misp),
    .io_exu_bp_exu_mp_pkt_bits_ataken(bp_ctl_io_exu_bp_exu_mp_pkt_bits_ataken),
    .io_exu_bp_exu_mp_pkt_bits_boffset(bp_ctl_io_exu_bp_exu_mp_pkt_bits_boffset),
    .io_exu_bp_exu_mp_pkt_bits_pc4(bp_ctl_io_exu_bp_exu_mp_pkt_bits_pc4),
    .io_exu_bp_exu_mp_pkt_bits_hist(bp_ctl_io_exu_bp_exu_mp_pkt_bits_hist),
    .io_exu_bp_exu_mp_pkt_bits_toffset(bp_ctl_io_exu_bp_exu_mp_pkt_bits_toffset),
    .io_exu_bp_exu_mp_pkt_bits_pcall(bp_ctl_io_exu_bp_exu_mp_pkt_bits_pcall),
    .io_exu_bp_exu_mp_pkt_bits_pret(bp_ctl_io_exu_bp_exu_mp_pkt_bits_pret),
    .io_exu_bp_exu_mp_pkt_bits_pja(bp_ctl_io_exu_bp_exu_mp_pkt_bits_pja),
    .io_exu_bp_exu_mp_pkt_bits_way(bp_ctl_io_exu_bp_exu_mp_pkt_bits_way),
    .io_exu_bp_exu_mp_eghr(bp_ctl_io_exu_bp_exu_mp_eghr),
    .io_exu_bp_exu_mp_fghr(bp_ctl_io_exu_bp_exu_mp_fghr),
    .io_exu_bp_exu_mp_index(bp_ctl_io_exu_bp_exu_mp_index),
    .io_exu_bp_exu_mp_btag(bp_ctl_io_exu_bp_exu_mp_btag),
    .io_ifu_bp_hit_taken_f(bp_ctl_io_ifu_bp_hit_taken_f),
    .io_ifu_bp_btb_target_f(bp_ctl_io_ifu_bp_btb_target_f),
    .io_ifu_bp_inst_mask_f(bp_ctl_io_ifu_bp_inst_mask_f),
    .io_ifu_bp_fghr_f(bp_ctl_io_ifu_bp_fghr_f),
    .io_ifu_bp_way_f(bp_ctl_io_ifu_bp_way_f),
    .io_ifu_bp_ret_f(bp_ctl_io_ifu_bp_ret_f),
    .io_ifu_bp_hist1_f(bp_ctl_io_ifu_bp_hist1_f),
    .io_ifu_bp_hist0_f(bp_ctl_io_ifu_bp_hist0_f),
    .io_ifu_bp_pc4_f(bp_ctl_io_ifu_bp_pc4_f),
    .io_ifu_bp_valid_f(bp_ctl_io_ifu_bp_valid_f),
    .io_ifu_bp_poffset_f(bp_ctl_io_ifu_bp_poffset_f),
    .io_scan_mode(bp_ctl_io_scan_mode)
  );
  ifu_aln_ctl aln_ctl ( // @[ifu.scala 36:23]
    .clock(aln_ctl_clock),
    .reset(aln_ctl_reset),
    .io_scan_mode(aln_ctl_io_scan_mode),
    .io_active_clk(aln_ctl_io_active_clk),
    .io_ifu_async_error_start(aln_ctl_io_ifu_async_error_start),
    .io_iccm_rd_ecc_double_err(aln_ctl_io_iccm_rd_ecc_double_err),
    .io_ic_access_fault_f(aln_ctl_io_ic_access_fault_f),
    .io_ic_access_fault_type_f(aln_ctl_io_ic_access_fault_type_f),
    .io_ifu_bp_fghr_f(aln_ctl_io_ifu_bp_fghr_f),
    .io_ifu_bp_btb_target_f(aln_ctl_io_ifu_bp_btb_target_f),
    .io_ifu_bp_poffset_f(aln_ctl_io_ifu_bp_poffset_f),
    .io_ifu_bp_hist0_f(aln_ctl_io_ifu_bp_hist0_f),
    .io_ifu_bp_hist1_f(aln_ctl_io_ifu_bp_hist1_f),
    .io_ifu_bp_pc4_f(aln_ctl_io_ifu_bp_pc4_f),
    .io_ifu_bp_way_f(aln_ctl_io_ifu_bp_way_f),
    .io_ifu_bp_valid_f(aln_ctl_io_ifu_bp_valid_f),
    .io_ifu_bp_ret_f(aln_ctl_io_ifu_bp_ret_f),
    .io_exu_flush_final(aln_ctl_io_exu_flush_final),
    .io_dec_aln_aln_dec_dec_i0_decode_d(aln_ctl_io_dec_aln_aln_dec_dec_i0_decode_d),
    .io_dec_aln_aln_dec_ifu_i0_cinst(aln_ctl_io_dec_aln_aln_dec_ifu_i0_cinst),
    .io_dec_aln_aln_ib_ifu_i0_icaf(aln_ctl_io_dec_aln_aln_ib_ifu_i0_icaf),
    .io_dec_aln_aln_ib_ifu_i0_icaf_type(aln_ctl_io_dec_aln_aln_ib_ifu_i0_icaf_type),
    .io_dec_aln_aln_ib_ifu_i0_icaf_f1(aln_ctl_io_dec_aln_aln_ib_ifu_i0_icaf_f1),
    .io_dec_aln_aln_ib_ifu_i0_dbecc(aln_ctl_io_dec_aln_aln_ib_ifu_i0_dbecc),
    .io_dec_aln_aln_ib_ifu_i0_bp_index(aln_ctl_io_dec_aln_aln_ib_ifu_i0_bp_index),
    .io_dec_aln_aln_ib_ifu_i0_bp_fghr(aln_ctl_io_dec_aln_aln_ib_ifu_i0_bp_fghr),
    .io_dec_aln_aln_ib_ifu_i0_bp_btag(aln_ctl_io_dec_aln_aln_ib_ifu_i0_bp_btag),
    .io_dec_aln_aln_ib_ifu_i0_valid(aln_ctl_io_dec_aln_aln_ib_ifu_i0_valid),
    .io_dec_aln_aln_ib_ifu_i0_instr(aln_ctl_io_dec_aln_aln_ib_ifu_i0_instr),
    .io_dec_aln_aln_ib_ifu_i0_pc(aln_ctl_io_dec_aln_aln_ib_ifu_i0_pc),
    .io_dec_aln_aln_ib_ifu_i0_pc4(aln_ctl_io_dec_aln_aln_ib_ifu_i0_pc4),
    .io_dec_aln_aln_ib_i0_brp_valid(aln_ctl_io_dec_aln_aln_ib_i0_brp_valid),
    .io_dec_aln_aln_ib_i0_brp_bits_toffset(aln_ctl_io_dec_aln_aln_ib_i0_brp_bits_toffset),
    .io_dec_aln_aln_ib_i0_brp_bits_hist(aln_ctl_io_dec_aln_aln_ib_i0_brp_bits_hist),
    .io_dec_aln_aln_ib_i0_brp_bits_br_error(aln_ctl_io_dec_aln_aln_ib_i0_brp_bits_br_error),
    .io_dec_aln_aln_ib_i0_brp_bits_br_start_error(aln_ctl_io_dec_aln_aln_ib_i0_brp_bits_br_start_error),
    .io_dec_aln_aln_ib_i0_brp_bits_prett(aln_ctl_io_dec_aln_aln_ib_i0_brp_bits_prett),
    .io_dec_aln_aln_ib_i0_brp_bits_way(aln_ctl_io_dec_aln_aln_ib_i0_brp_bits_way),
    .io_dec_aln_aln_ib_i0_brp_bits_ret(aln_ctl_io_dec_aln_aln_ib_i0_brp_bits_ret),
    .io_dec_aln_ifu_pmu_instr_aligned(aln_ctl_io_dec_aln_ifu_pmu_instr_aligned),
    .io_ifu_fetch_data_f(aln_ctl_io_ifu_fetch_data_f),
    .io_ifu_fetch_val(aln_ctl_io_ifu_fetch_val),
    .io_ifu_fetch_pc(aln_ctl_io_ifu_fetch_pc),
    .io_ifu_fb_consume1(aln_ctl_io_ifu_fb_consume1),
    .io_ifu_fb_consume2(aln_ctl_io_ifu_fb_consume2)
  );
  ifu_ifc_ctl ifc_ctl ( // @[ifu.scala 37:23]
    .clock(ifc_ctl_clock),
    .reset(ifc_ctl_reset),
    .io_exu_flush_final(ifc_ctl_io_exu_flush_final),
    .io_exu_flush_path_final(ifc_ctl_io_exu_flush_path_final),
    .io_free_clk(ifc_ctl_io_free_clk),
    .io_active_clk(ifc_ctl_io_active_clk),
    .io_scan_mode(ifc_ctl_io_scan_mode),
    .io_ic_hit_f(ifc_ctl_io_ic_hit_f),
    .io_ifu_ic_mb_empty(ifc_ctl_io_ifu_ic_mb_empty),
    .io_ifu_fb_consume1(ifc_ctl_io_ifu_fb_consume1),
    .io_ifu_fb_consume2(ifc_ctl_io_ifu_fb_consume2),
    .io_ifu_bp_hit_taken_f(ifc_ctl_io_ifu_bp_hit_taken_f),
    .io_ifu_bp_btb_target_f(ifc_ctl_io_ifu_bp_btb_target_f),
    .io_ic_dma_active(ifc_ctl_io_ic_dma_active),
    .io_dec_ifc_dec_tlu_flush_noredir_wb(ifc_ctl_io_dec_ifc_dec_tlu_flush_noredir_wb),
    .io_dec_ifc_dec_tlu_mrac_ff(ifc_ctl_io_dec_ifc_dec_tlu_mrac_ff),
    .io_dec_ifc_ifu_pmu_fetch_stall(ifc_ctl_io_dec_ifc_ifu_pmu_fetch_stall),
    .io_dma_ifc_dma_iccm_stall_any(ifc_ctl_io_dma_ifc_dma_iccm_stall_any),
    .io_ifc_fetch_addr_f(ifc_ctl_io_ifc_fetch_addr_f),
    .io_ifc_fetch_addr_bf(ifc_ctl_io_ifc_fetch_addr_bf),
    .io_ifc_fetch_req_f(ifc_ctl_io_ifc_fetch_req_f),
    .io_ifc_fetch_uncacheable_bf(ifc_ctl_io_ifc_fetch_uncacheable_bf),
    .io_ifc_fetch_req_bf(ifc_ctl_io_ifc_fetch_req_bf),
    .io_ifc_fetch_req_bf_raw(ifc_ctl_io_ifc_fetch_req_bf_raw),
    .io_ifc_iccm_access_bf(ifc_ctl_io_ifc_iccm_access_bf),
    .io_ifc_region_acc_fault_bf(ifc_ctl_io_ifc_region_acc_fault_bf),
    .io_ifc_dma_access_ok(ifc_ctl_io_ifc_dma_access_ok)
  );
  assign io_ifu_dec_dec_aln_aln_dec_ifu_i0_cinst = aln_ctl_io_dec_aln_aln_dec_ifu_i0_cinst; // @[ifu.scala 73:22]
  assign io_ifu_dec_dec_aln_aln_ib_ifu_i0_icaf = aln_ctl_io_dec_aln_aln_ib_ifu_i0_icaf; // @[ifu.scala 73:22]
  assign io_ifu_dec_dec_aln_aln_ib_ifu_i0_icaf_type = aln_ctl_io_dec_aln_aln_ib_ifu_i0_icaf_type; // @[ifu.scala 73:22]
  assign io_ifu_dec_dec_aln_aln_ib_ifu_i0_icaf_f1 = aln_ctl_io_dec_aln_aln_ib_ifu_i0_icaf_f1; // @[ifu.scala 73:22]
  assign io_ifu_dec_dec_aln_aln_ib_ifu_i0_dbecc = aln_ctl_io_dec_aln_aln_ib_ifu_i0_dbecc; // @[ifu.scala 73:22]
  assign io_ifu_dec_dec_aln_aln_ib_ifu_i0_bp_index = aln_ctl_io_dec_aln_aln_ib_ifu_i0_bp_index; // @[ifu.scala 73:22]
  assign io_ifu_dec_dec_aln_aln_ib_ifu_i0_bp_fghr = aln_ctl_io_dec_aln_aln_ib_ifu_i0_bp_fghr; // @[ifu.scala 73:22]
  assign io_ifu_dec_dec_aln_aln_ib_ifu_i0_bp_btag = aln_ctl_io_dec_aln_aln_ib_ifu_i0_bp_btag; // @[ifu.scala 73:22]
  assign io_ifu_dec_dec_aln_aln_ib_ifu_i0_valid = aln_ctl_io_dec_aln_aln_ib_ifu_i0_valid; // @[ifu.scala 73:22]
  assign io_ifu_dec_dec_aln_aln_ib_ifu_i0_instr = aln_ctl_io_dec_aln_aln_ib_ifu_i0_instr; // @[ifu.scala 73:22]
  assign io_ifu_dec_dec_aln_aln_ib_ifu_i0_pc = aln_ctl_io_dec_aln_aln_ib_ifu_i0_pc; // @[ifu.scala 73:22]
  assign io_ifu_dec_dec_aln_aln_ib_ifu_i0_pc4 = aln_ctl_io_dec_aln_aln_ib_ifu_i0_pc4; // @[ifu.scala 73:22]
  assign io_ifu_dec_dec_aln_aln_ib_i0_brp_valid = aln_ctl_io_dec_aln_aln_ib_i0_brp_valid; // @[ifu.scala 73:22]
  assign io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_toffset = aln_ctl_io_dec_aln_aln_ib_i0_brp_bits_toffset; // @[ifu.scala 73:22]
  assign io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_hist = aln_ctl_io_dec_aln_aln_ib_i0_brp_bits_hist; // @[ifu.scala 73:22]
  assign io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_br_error = aln_ctl_io_dec_aln_aln_ib_i0_brp_bits_br_error; // @[ifu.scala 73:22]
  assign io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_br_start_error = aln_ctl_io_dec_aln_aln_ib_i0_brp_bits_br_start_error; // @[ifu.scala 73:22]
  assign io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_prett = aln_ctl_io_dec_aln_aln_ib_i0_brp_bits_prett; // @[ifu.scala 73:22]
  assign io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_way = aln_ctl_io_dec_aln_aln_ib_i0_brp_bits_way; // @[ifu.scala 73:22]
  assign io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_ret = aln_ctl_io_dec_aln_aln_ib_i0_brp_bits_ret; // @[ifu.scala 73:22]
  assign io_ifu_dec_dec_aln_ifu_pmu_instr_aligned = aln_ctl_io_dec_aln_ifu_pmu_instr_aligned; // @[ifu.scala 73:22]
  assign io_ifu_dec_dec_mem_ctrl_ifu_pmu_ic_miss = mem_ctl_io_dec_mem_ctrl_ifu_pmu_ic_miss; // @[ifu.scala 93:27]
  assign io_ifu_dec_dec_mem_ctrl_ifu_pmu_ic_hit = mem_ctl_io_dec_mem_ctrl_ifu_pmu_ic_hit; // @[ifu.scala 93:27]
  assign io_ifu_dec_dec_mem_ctrl_ifu_pmu_bus_error = mem_ctl_io_dec_mem_ctrl_ifu_pmu_bus_error; // @[ifu.scala 93:27]
  assign io_ifu_dec_dec_mem_ctrl_ifu_pmu_bus_busy = mem_ctl_io_dec_mem_ctrl_ifu_pmu_bus_busy; // @[ifu.scala 93:27]
  assign io_ifu_dec_dec_mem_ctrl_ifu_ic_error_start = mem_ctl_io_dec_mem_ctrl_ifu_ic_error_start; // @[ifu.scala 93:27]
  assign io_ifu_dec_dec_mem_ctrl_ifu_iccm_rd_ecc_single_err = mem_ctl_io_dec_mem_ctrl_ifu_iccm_rd_ecc_single_err; // @[ifu.scala 93:27]
  assign io_ifu_dec_dec_mem_ctrl_ifu_ic_debug_rd_data = mem_ctl_io_dec_mem_ctrl_ifu_ic_debug_rd_data; // @[ifu.scala 93:27]
  assign io_ifu_dec_dec_mem_ctrl_ifu_ic_debug_rd_data_valid = mem_ctl_io_dec_mem_ctrl_ifu_ic_debug_rd_data_valid; // @[ifu.scala 93:27]
  assign io_ifu_dec_dec_mem_ctrl_ifu_miss_state_idle = mem_ctl_io_dec_mem_ctrl_ifu_miss_state_idle; // @[ifu.scala 93:27]
  assign io_ifu_dec_dec_ifc_ifu_pmu_fetch_stall = ifc_ctl_io_dec_ifc_ifu_pmu_fetch_stall; // @[ifu.scala 46:22]
  assign io_iccm_rw_addr = mem_ctl_io_iccm_rw_addr; // @[ifu.scala 107:19]
  assign io_iccm_buf_correct_ecc = mem_ctl_io_iccm_buf_correct_ecc; // @[ifu.scala 107:19]
  assign io_iccm_correction_state = mem_ctl_io_iccm_correction_state; // @[ifu.scala 107:19]
  assign io_iccm_wren = mem_ctl_io_iccm_wren; // @[ifu.scala 107:19]
  assign io_iccm_rden = mem_ctl_io_iccm_rden; // @[ifu.scala 107:19]
  assign io_iccm_wr_size = mem_ctl_io_iccm_wr_size; // @[ifu.scala 107:19]
  assign io_iccm_wr_data = mem_ctl_io_iccm_wr_data; // @[ifu.scala 107:19]
  assign io_ic_rw_addr = mem_ctl_io_ic_rw_addr; // @[ifu.scala 106:17]
  assign io_ic_tag_valid = mem_ctl_io_ic_tag_valid; // @[ifu.scala 106:17]
  assign io_ic_rd_en = mem_ctl_io_ic_rd_en; // @[ifu.scala 106:17]
  assign io_ic_debug_wr_data = mem_ctl_io_ic_debug_wr_data; // @[ifu.scala 106:17]
  assign io_ic_debug_addr = mem_ctl_io_ic_debug_addr; // @[ifu.scala 106:17]
  assign io_ic_debug_rd_en = mem_ctl_io_ic_debug_rd_en; // @[ifu.scala 106:17]
  assign io_ic_debug_wr_en = mem_ctl_io_ic_debug_wr_en; // @[ifu.scala 106:17]
  assign io_ic_debug_tag_array = mem_ctl_io_ic_debug_tag_array; // @[ifu.scala 106:17]
  assign io_ic_debug_way = mem_ctl_io_ic_debug_way; // @[ifu.scala 106:17]
  assign io_ic_premux_data = mem_ctl_io_ic_premux_data; // @[ifu.scala 106:17]
  assign io_ic_sel_premux_data = mem_ctl_io_ic_sel_premux_data; // @[ifu.scala 106:17]
  assign io_ifu_ar_valid = mem_ctl_io_ifu_axi_ar_valid; // @[ifu.scala 103:22]
  assign io_ifu_ar_bits_addr = mem_ctl_io_ifu_axi_ar_bits_addr; // @[ifu.scala 103:22]
  assign io_iccm_dma_ecc_error = mem_ctl_io_iccm_dma_ecc_error; // @[ifu.scala 113:25]
  assign io_iccm_dma_rvalid = mem_ctl_io_iccm_dma_rvalid; // @[ifu.scala 114:22]
  assign io_iccm_dma_rdata = mem_ctl_io_iccm_dma_rdata; // @[ifu.scala 115:21]
  assign io_iccm_dma_rtag = mem_ctl_io_iccm_dma_rtag; // @[ifu.scala 116:20]
  assign io_iccm_ready = mem_ctl_io_iccm_ready; // @[ifu.scala 117:17]
  assign io_iccm_dma_sb_error = mem_ctl_io_iccm_dma_sb_error; // @[ifu.scala 118:24]
  assign mem_ctl_clock = clock;
  assign mem_ctl_reset = reset;
  assign mem_ctl_io_free_clk = io_free_clk; // @[ifu.scala 90:23]
  assign mem_ctl_io_active_clk = io_active_clk; // @[ifu.scala 91:25]
  assign mem_ctl_io_exu_flush_final = io_exu_flush_final; // @[ifu.scala 92:30]
  assign mem_ctl_io_dec_mem_ctrl_dec_tlu_flush_err_wb = io_ifu_dec_dec_mem_ctrl_dec_tlu_flush_err_wb; // @[ifu.scala 93:27]
  assign mem_ctl_io_dec_mem_ctrl_dec_tlu_i0_commit_cmt = io_ifu_dec_dec_mem_ctrl_dec_tlu_i0_commit_cmt; // @[ifu.scala 93:27]
  assign mem_ctl_io_dec_mem_ctrl_dec_tlu_force_halt = io_ifu_dec_dec_mem_ctrl_dec_tlu_force_halt; // @[ifu.scala 93:27]
  assign mem_ctl_io_dec_mem_ctrl_dec_tlu_fence_i_wb = io_ifu_dec_dec_mem_ctrl_dec_tlu_fence_i_wb; // @[ifu.scala 93:27]
  assign mem_ctl_io_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_wrdata = io_ifu_dec_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_wrdata; // @[ifu.scala 93:27]
  assign mem_ctl_io_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_dicawics = io_ifu_dec_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_dicawics; // @[ifu.scala 93:27]
  assign mem_ctl_io_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_rd_valid = io_ifu_dec_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_rd_valid; // @[ifu.scala 93:27]
  assign mem_ctl_io_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_wr_valid = io_ifu_dec_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_wr_valid; // @[ifu.scala 93:27]
  assign mem_ctl_io_dec_mem_ctrl_dec_tlu_core_ecc_disable = io_ifu_dec_dec_mem_ctrl_dec_tlu_core_ecc_disable; // @[ifu.scala 93:27]
  assign mem_ctl_io_ifc_fetch_addr_bf = ifc_ctl_io_ifc_fetch_addr_bf; // @[ifu.scala 94:32]
  assign mem_ctl_io_ifc_fetch_uncacheable_bf = ifc_ctl_io_ifc_fetch_uncacheable_bf; // @[ifu.scala 95:39]
  assign mem_ctl_io_ifc_fetch_req_bf = ifc_ctl_io_ifc_fetch_req_bf; // @[ifu.scala 96:31]
  assign mem_ctl_io_ifc_fetch_req_bf_raw = ifc_ctl_io_ifc_fetch_req_bf_raw; // @[ifu.scala 97:35]
  assign mem_ctl_io_ifc_iccm_access_bf = ifc_ctl_io_ifc_iccm_access_bf; // @[ifu.scala 98:33]
  assign mem_ctl_io_ifc_region_acc_fault_bf = ifc_ctl_io_ifc_region_acc_fault_bf; // @[ifu.scala 99:38]
  assign mem_ctl_io_ifc_dma_access_ok = ifc_ctl_io_ifc_dma_access_ok; // @[ifu.scala 100:32]
  assign mem_ctl_io_ifu_bp_hit_taken_f = bp_ctl_io_ifu_bp_hit_taken_f; // @[ifu.scala 101:33]
  assign mem_ctl_io_ifu_bp_inst_mask_f = bp_ctl_io_ifu_bp_inst_mask_f; // @[ifu.scala 102:33]
  assign mem_ctl_io_ifu_bus_clk_en = io_ifu_bus_clk_en; // @[ifu.scala 104:29]
  assign mem_ctl_io_dma_mem_ctl_dma_iccm_req = io_ifu_dma_dma_mem_ctl_dma_iccm_req; // @[ifu.scala 105:26]
  assign mem_ctl_io_dma_mem_ctl_dma_mem_addr = io_ifu_dma_dma_mem_ctl_dma_mem_addr; // @[ifu.scala 105:26]
  assign mem_ctl_io_dma_mem_ctl_dma_mem_sz = io_ifu_dma_dma_mem_ctl_dma_mem_sz; // @[ifu.scala 105:26]
  assign mem_ctl_io_dma_mem_ctl_dma_mem_write = io_ifu_dma_dma_mem_ctl_dma_mem_write; // @[ifu.scala 105:26]
  assign mem_ctl_io_dma_mem_ctl_dma_mem_wdata = io_ifu_dma_dma_mem_ctl_dma_mem_wdata; // @[ifu.scala 105:26]
  assign mem_ctl_io_dma_mem_ctl_dma_mem_tag = io_ifu_dma_dma_mem_ctl_dma_mem_tag; // @[ifu.scala 105:26]
  assign mem_ctl_io_iccm_rd_data = io_iccm_rd_data; // @[ifu.scala 107:19]
  assign mem_ctl_io_iccm_rd_data_ecc = io_iccm_rd_data_ecc; // @[ifu.scala 107:19]
  assign mem_ctl_io_ic_rd_data = io_ic_rd_data; // @[ifu.scala 106:17]
  assign mem_ctl_io_ic_debug_rd_data = io_ic_debug_rd_data; // @[ifu.scala 106:17]
  assign mem_ctl_io_ic_tag_debug_rd_data = io_ic_tag_debug_rd_data; // @[ifu.scala 106:17]
  assign mem_ctl_io_ic_eccerr = io_ic_eccerr; // @[ifu.scala 106:17]
  assign mem_ctl_io_ic_rd_hit = io_ic_rd_hit; // @[ifu.scala 106:17]
  assign mem_ctl_io_ic_tag_perr = io_ic_tag_perr; // @[ifu.scala 106:17]
  assign mem_ctl_io_ifu_fetch_val = mem_ctl_io_ic_fetch_val_f; // @[ifu.scala 108:28]
  assign mem_ctl_io_dec_tlu_flush_lower_wb = io_dec_tlu_flush_lower_wb; // @[ifu.scala 109:37]
  assign mem_ctl_io_scan_mode = io_scan_mode; // @[ifu.scala 110:24]
  assign bp_ctl_clock = clock;
  assign bp_ctl_reset = reset;
  assign bp_ctl_io_active_clk = io_active_clk; // @[ifu.scala 80:24]
  assign bp_ctl_io_ic_hit_f = mem_ctl_io_ic_hit_f; // @[ifu.scala 81:22]
  assign bp_ctl_io_exu_flush_final = io_exu_flush_final; // @[ifu.scala 86:29]
  assign bp_ctl_io_ifc_fetch_addr_f = ifc_ctl_io_ifc_fetch_addr_f; // @[ifu.scala 82:30]
  assign bp_ctl_io_ifc_fetch_req_f = ifc_ctl_io_ifc_fetch_req_f; // @[ifu.scala 83:29]
  assign bp_ctl_io_dec_bp_dec_tlu_br0_r_pkt_valid = io_ifu_dec_dec_bp_dec_tlu_br0_r_pkt_valid; // @[ifu.scala 84:20]
  assign bp_ctl_io_dec_bp_dec_tlu_br0_r_pkt_bits_hist = io_ifu_dec_dec_bp_dec_tlu_br0_r_pkt_bits_hist; // @[ifu.scala 84:20]
  assign bp_ctl_io_dec_bp_dec_tlu_br0_r_pkt_bits_br_error = io_ifu_dec_dec_bp_dec_tlu_br0_r_pkt_bits_br_error; // @[ifu.scala 84:20]
  assign bp_ctl_io_dec_bp_dec_tlu_br0_r_pkt_bits_br_start_error = io_ifu_dec_dec_bp_dec_tlu_br0_r_pkt_bits_br_start_error; // @[ifu.scala 84:20]
  assign bp_ctl_io_dec_bp_dec_tlu_br0_r_pkt_bits_way = io_ifu_dec_dec_bp_dec_tlu_br0_r_pkt_bits_way; // @[ifu.scala 84:20]
  assign bp_ctl_io_dec_bp_dec_tlu_br0_r_pkt_bits_middle = io_ifu_dec_dec_bp_dec_tlu_br0_r_pkt_bits_middle; // @[ifu.scala 84:20]
  assign bp_ctl_io_dec_bp_dec_tlu_flush_leak_one_wb = io_ifu_dec_dec_bp_dec_tlu_flush_leak_one_wb; // @[ifu.scala 84:20]
  assign bp_ctl_io_dec_bp_dec_tlu_bpred_disable = io_ifu_dec_dec_bp_dec_tlu_bpred_disable; // @[ifu.scala 84:20]
  assign bp_ctl_io_dec_tlu_flush_lower_wb = io_dec_tlu_flush_lower_wb; // @[ifu.scala 87:36]
  assign bp_ctl_io_exu_bp_exu_i0_br_index_r = io_exu_ifu_exu_bp_exu_i0_br_index_r; // @[ifu.scala 85:20]
  assign bp_ctl_io_exu_bp_exu_i0_br_fghr_r = io_exu_ifu_exu_bp_exu_i0_br_fghr_r; // @[ifu.scala 85:20]
  assign bp_ctl_io_exu_bp_exu_mp_pkt_bits_misp = io_exu_ifu_exu_bp_exu_mp_pkt_bits_misp; // @[ifu.scala 85:20]
  assign bp_ctl_io_exu_bp_exu_mp_pkt_bits_ataken = io_exu_ifu_exu_bp_exu_mp_pkt_bits_ataken; // @[ifu.scala 85:20]
  assign bp_ctl_io_exu_bp_exu_mp_pkt_bits_boffset = io_exu_ifu_exu_bp_exu_mp_pkt_bits_boffset; // @[ifu.scala 85:20]
  assign bp_ctl_io_exu_bp_exu_mp_pkt_bits_pc4 = io_exu_ifu_exu_bp_exu_mp_pkt_bits_pc4; // @[ifu.scala 85:20]
  assign bp_ctl_io_exu_bp_exu_mp_pkt_bits_hist = io_exu_ifu_exu_bp_exu_mp_pkt_bits_hist; // @[ifu.scala 85:20]
  assign bp_ctl_io_exu_bp_exu_mp_pkt_bits_toffset = io_exu_ifu_exu_bp_exu_mp_pkt_bits_toffset; // @[ifu.scala 85:20]
  assign bp_ctl_io_exu_bp_exu_mp_pkt_bits_pcall = io_exu_ifu_exu_bp_exu_mp_pkt_bits_pcall; // @[ifu.scala 85:20]
  assign bp_ctl_io_exu_bp_exu_mp_pkt_bits_pret = io_exu_ifu_exu_bp_exu_mp_pkt_bits_pret; // @[ifu.scala 85:20]
  assign bp_ctl_io_exu_bp_exu_mp_pkt_bits_pja = io_exu_ifu_exu_bp_exu_mp_pkt_bits_pja; // @[ifu.scala 85:20]
  assign bp_ctl_io_exu_bp_exu_mp_pkt_bits_way = io_exu_ifu_exu_bp_exu_mp_pkt_bits_way; // @[ifu.scala 85:20]
  assign bp_ctl_io_exu_bp_exu_mp_eghr = io_exu_ifu_exu_bp_exu_mp_eghr; // @[ifu.scala 85:20]
  assign bp_ctl_io_exu_bp_exu_mp_fghr = io_exu_ifu_exu_bp_exu_mp_fghr; // @[ifu.scala 85:20]
  assign bp_ctl_io_exu_bp_exu_mp_index = io_exu_ifu_exu_bp_exu_mp_index; // @[ifu.scala 85:20]
  assign bp_ctl_io_exu_bp_exu_mp_btag = io_exu_ifu_exu_bp_exu_mp_btag; // @[ifu.scala 85:20]
  assign bp_ctl_io_scan_mode = io_scan_mode; // @[ifu.scala 79:23]
  assign aln_ctl_clock = clock;
  assign aln_ctl_reset = reset;
  assign aln_ctl_io_scan_mode = io_scan_mode; // @[ifu.scala 57:24]
  assign aln_ctl_io_active_clk = io_active_clk; // @[ifu.scala 58:25]
  assign aln_ctl_io_ifu_async_error_start = mem_ctl_io_ifu_async_error_start; // @[ifu.scala 59:36]
  assign aln_ctl_io_iccm_rd_ecc_double_err = mem_ctl_io_iccm_rd_ecc_double_err; // @[ifu.scala 60:37]
  assign aln_ctl_io_ic_access_fault_f = mem_ctl_io_ic_access_fault_f; // @[ifu.scala 61:32]
  assign aln_ctl_io_ic_access_fault_type_f = mem_ctl_io_ic_access_fault_type_f; // @[ifu.scala 62:37]
  assign aln_ctl_io_ifu_bp_fghr_f = bp_ctl_io_ifu_bp_fghr_f; // @[ifu.scala 63:28]
  assign aln_ctl_io_ifu_bp_btb_target_f = bp_ctl_io_ifu_bp_btb_target_f; // @[ifu.scala 64:34]
  assign aln_ctl_io_ifu_bp_poffset_f = bp_ctl_io_ifu_bp_poffset_f; // @[ifu.scala 65:31]
  assign aln_ctl_io_ifu_bp_hist0_f = bp_ctl_io_ifu_bp_hist0_f; // @[ifu.scala 66:29]
  assign aln_ctl_io_ifu_bp_hist1_f = bp_ctl_io_ifu_bp_hist1_f; // @[ifu.scala 67:29]
  assign aln_ctl_io_ifu_bp_pc4_f = bp_ctl_io_ifu_bp_pc4_f; // @[ifu.scala 68:27]
  assign aln_ctl_io_ifu_bp_way_f = bp_ctl_io_ifu_bp_way_f; // @[ifu.scala 69:27]
  assign aln_ctl_io_ifu_bp_valid_f = bp_ctl_io_ifu_bp_valid_f; // @[ifu.scala 70:29]
  assign aln_ctl_io_ifu_bp_ret_f = bp_ctl_io_ifu_bp_ret_f; // @[ifu.scala 71:27]
  assign aln_ctl_io_exu_flush_final = io_exu_flush_final; // @[ifu.scala 72:30]
  assign aln_ctl_io_dec_aln_aln_dec_dec_i0_decode_d = io_ifu_dec_dec_aln_aln_dec_dec_i0_decode_d; // @[ifu.scala 73:22]
  assign aln_ctl_io_ifu_fetch_data_f = mem_ctl_io_ic_data_f; // @[ifu.scala 74:31]
  assign aln_ctl_io_ifu_fetch_val = mem_ctl_io_ifu_fetch_val; // @[ifu.scala 75:28]
  assign aln_ctl_io_ifu_fetch_pc = ifc_ctl_io_ifc_fetch_addr_f; // @[ifu.scala 76:27]
  assign ifc_ctl_clock = clock;
  assign ifc_ctl_reset = reset;
  assign ifc_ctl_io_exu_flush_final = io_exu_flush_final; // @[ifu.scala 47:30]
  assign ifc_ctl_io_exu_flush_path_final = io_exu_flush_path_final; // @[ifu.scala 54:35]
  assign ifc_ctl_io_free_clk = io_free_clk; // @[ifu.scala 41:23]
  assign ifc_ctl_io_active_clk = io_active_clk; // @[ifu.scala 40:25]
  assign ifc_ctl_io_scan_mode = io_scan_mode; // @[ifu.scala 42:24]
  assign ifc_ctl_io_ic_hit_f = mem_ctl_io_ic_hit_f; // @[ifu.scala 43:23]
  assign ifc_ctl_io_ifu_ic_mb_empty = mem_ctl_io_ifu_ic_mb_empty; // @[ifu.scala 53:30]
  assign ifc_ctl_io_ifu_fb_consume1 = aln_ctl_io_ifu_fb_consume1; // @[ifu.scala 44:30]
  assign ifc_ctl_io_ifu_fb_consume2 = aln_ctl_io_ifu_fb_consume2; // @[ifu.scala 45:30]
  assign ifc_ctl_io_ifu_bp_hit_taken_f = bp_ctl_io_ifu_bp_hit_taken_f; // @[ifu.scala 48:33]
  assign ifc_ctl_io_ifu_bp_btb_target_f = bp_ctl_io_ifu_bp_btb_target_f; // @[ifu.scala 49:34]
  assign ifc_ctl_io_ic_dma_active = mem_ctl_io_ic_dma_active; // @[ifu.scala 50:28]
  assign ifc_ctl_io_dec_ifc_dec_tlu_flush_noredir_wb = io_ifu_dec_dec_ifc_dec_tlu_flush_noredir_wb; // @[ifu.scala 46:22]
  assign ifc_ctl_io_dec_ifc_dec_tlu_mrac_ff = io_ifu_dec_dec_ifc_dec_tlu_mrac_ff; // @[ifu.scala 46:22]
  assign ifc_ctl_io_dma_ifc_dma_iccm_stall_any = io_ifu_dma_dma_ifc_dma_iccm_stall_any; // @[ifu.scala 52:22]
endmodule
module dec_ib_ctl(
  input         io_ifu_ib_ifu_i0_icaf,
  input  [1:0]  io_ifu_ib_ifu_i0_icaf_type,
  input         io_ifu_ib_ifu_i0_icaf_f1,
  input         io_ifu_ib_ifu_i0_dbecc,
  input  [7:0]  io_ifu_ib_ifu_i0_bp_index,
  input  [7:0]  io_ifu_ib_ifu_i0_bp_fghr,
  input  [4:0]  io_ifu_ib_ifu_i0_bp_btag,
  input         io_ifu_ib_ifu_i0_valid,
  input  [31:0] io_ifu_ib_ifu_i0_instr,
  input  [30:0] io_ifu_ib_ifu_i0_pc,
  input         io_ifu_ib_ifu_i0_pc4,
  input         io_ifu_ib_i0_brp_valid,
  input  [11:0] io_ifu_ib_i0_brp_bits_toffset,
  input  [1:0]  io_ifu_ib_i0_brp_bits_hist,
  input         io_ifu_ib_i0_brp_bits_br_error,
  input         io_ifu_ib_i0_brp_bits_br_start_error,
  input  [30:0] io_ifu_ib_i0_brp_bits_prett,
  input         io_ifu_ib_i0_brp_bits_way,
  input         io_ifu_ib_i0_brp_bits_ret,
  output [30:0] io_ib_exu_dec_i0_pc_d,
  output        io_ib_exu_dec_debug_wdata_rs1_d,
  input         io_dbg_ib_dbg_cmd_valid,
  input         io_dbg_ib_dbg_cmd_write,
  input  [1:0]  io_dbg_ib_dbg_cmd_type,
  input  [31:0] io_dbg_ib_dbg_cmd_addr,
  output        io_dec_ib0_valid_d,
  output [1:0]  io_dec_i0_icaf_type_d,
  output [31:0] io_dec_i0_instr_d,
  output        io_dec_i0_pc4_d,
  output        io_dec_i0_brp_valid,
  output [11:0] io_dec_i0_brp_bits_toffset,
  output [1:0]  io_dec_i0_brp_bits_hist,
  output        io_dec_i0_brp_bits_br_error,
  output        io_dec_i0_brp_bits_br_start_error,
  output [30:0] io_dec_i0_brp_bits_prett,
  output        io_dec_i0_brp_bits_way,
  output        io_dec_i0_brp_bits_ret,
  output [7:0]  io_dec_i0_bp_index,
  output [7:0]  io_dec_i0_bp_fghr,
  output [4:0]  io_dec_i0_bp_btag,
  output        io_dec_i0_icaf_d,
  output        io_dec_i0_icaf_f1_d,
  output        io_dec_i0_dbecc_d,
  output        io_dec_debug_fence_d
);
  wire  _T = io_dbg_ib_dbg_cmd_type != 2'h2; // @[dec_ib_ctl.scala 52:74]
  wire  debug_valid = io_dbg_ib_dbg_cmd_valid & _T; // @[dec_ib_ctl.scala 52:48]
  wire  _T_1 = ~io_dbg_ib_dbg_cmd_write; // @[dec_ib_ctl.scala 53:38]
  wire  debug_read = debug_valid & _T_1; // @[dec_ib_ctl.scala 53:36]
  wire  debug_write = debug_valid & io_dbg_ib_dbg_cmd_write; // @[dec_ib_ctl.scala 54:36]
  wire  _T_2 = io_dbg_ib_dbg_cmd_type == 2'h0; // @[dec_ib_ctl.scala 56:62]
  wire  debug_read_gpr = debug_read & _T_2; // @[dec_ib_ctl.scala 56:37]
  wire  debug_write_gpr = debug_write & _T_2; // @[dec_ib_ctl.scala 57:37]
  wire  _T_4 = io_dbg_ib_dbg_cmd_type == 2'h1; // @[dec_ib_ctl.scala 58:62]
  wire  debug_read_csr = debug_read & _T_4; // @[dec_ib_ctl.scala 58:37]
  wire  debug_write_csr = debug_write & _T_4; // @[dec_ib_ctl.scala 59:37]
  wire [4:0] dreg = io_dbg_ib_dbg_cmd_addr[4:0]; // @[dec_ib_ctl.scala 61:47]
  wire [11:0] dcsr = io_dbg_ib_dbg_cmd_addr[11:0]; // @[dec_ib_ctl.scala 62:47]
  wire [31:0] _T_9 = {12'h0,dreg,15'h6033}; // @[Cat.scala 29:58]
  wire [31:0] _T_12 = {20'h6,dreg,7'h33}; // @[Cat.scala 29:58]
  wire [31:0] _T_14 = {dcsr,20'h2073}; // @[Cat.scala 29:58]
  wire [31:0] _T_16 = {dcsr,20'h1073}; // @[Cat.scala 29:58]
  wire [31:0] _T_17 = debug_read_gpr ? _T_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_18 = debug_write_gpr ? _T_12 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_19 = debug_read_csr ? _T_14 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_20 = debug_write_csr ? _T_16 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_21 = _T_17 | _T_18; // @[Mux.scala 27:72]
  wire [31:0] _T_22 = _T_21 | _T_19; // @[Mux.scala 27:72]
  wire [31:0] ib0_debug_in = _T_22 | _T_20; // @[Mux.scala 27:72]
  wire  _T_25 = dcsr == 12'h7c4; // @[dec_ib_ctl.scala 75:51]
  assign io_ib_exu_dec_i0_pc_d = io_ifu_ib_ifu_i0_pc; // @[dec_ib_ctl.scala 32:31]
  assign io_ib_exu_dec_debug_wdata_rs1_d = debug_write_gpr | debug_write_csr; // @[dec_ib_ctl.scala 72:35]
  assign io_dec_ib0_valid_d = io_ifu_ib_ifu_i0_valid | debug_valid; // @[dec_ib_ctl.scala 77:22]
  assign io_dec_i0_icaf_type_d = io_ifu_ib_ifu_i0_icaf_type; // @[dec_ib_ctl.scala 34:31]
  assign io_dec_i0_instr_d = debug_valid ? ib0_debug_in : io_ifu_ib_ifu_i0_instr; // @[dec_ib_ctl.scala 78:22]
  assign io_dec_i0_pc4_d = io_ifu_ib_ifu_i0_pc4; // @[dec_ib_ctl.scala 33:31]
  assign io_dec_i0_brp_valid = io_ifu_ib_i0_brp_valid; // @[dec_ib_ctl.scala 35:31]
  assign io_dec_i0_brp_bits_toffset = io_ifu_ib_i0_brp_bits_toffset; // @[dec_ib_ctl.scala 35:31]
  assign io_dec_i0_brp_bits_hist = io_ifu_ib_i0_brp_bits_hist; // @[dec_ib_ctl.scala 35:31]
  assign io_dec_i0_brp_bits_br_error = io_ifu_ib_i0_brp_bits_br_error; // @[dec_ib_ctl.scala 35:31]
  assign io_dec_i0_brp_bits_br_start_error = io_ifu_ib_i0_brp_bits_br_start_error; // @[dec_ib_ctl.scala 35:31]
  assign io_dec_i0_brp_bits_prett = io_ifu_ib_i0_brp_bits_prett; // @[dec_ib_ctl.scala 35:31]
  assign io_dec_i0_brp_bits_way = io_ifu_ib_i0_brp_bits_way; // @[dec_ib_ctl.scala 35:31]
  assign io_dec_i0_brp_bits_ret = io_ifu_ib_i0_brp_bits_ret; // @[dec_ib_ctl.scala 35:31]
  assign io_dec_i0_bp_index = io_ifu_ib_ifu_i0_bp_index; // @[dec_ib_ctl.scala 36:31]
  assign io_dec_i0_bp_fghr = io_ifu_ib_ifu_i0_bp_fghr; // @[dec_ib_ctl.scala 37:31]
  assign io_dec_i0_bp_btag = io_ifu_ib_ifu_i0_bp_btag; // @[dec_ib_ctl.scala 38:31]
  assign io_dec_i0_icaf_d = io_ifu_ib_ifu_i0_icaf; // @[dec_ib_ctl.scala 31:31]
  assign io_dec_i0_icaf_f1_d = io_ifu_ib_ifu_i0_icaf_f1; // @[dec_ib_ctl.scala 29:31]
  assign io_dec_i0_dbecc_d = io_ifu_ib_ifu_i0_dbecc; // @[dec_ib_ctl.scala 30:31]
  assign io_dec_debug_fence_d = debug_write_csr & _T_25; // @[dec_ib_ctl.scala 75:24]
endmodule
module dec_dec_ctl(
  input  [31:0] io_ins,
  output        io_out_alu,
  output        io_out_rs1,
  output        io_out_rs2,
  output        io_out_imm12,
  output        io_out_rd,
  output        io_out_shimm5,
  output        io_out_imm20,
  output        io_out_pc,
  output        io_out_load,
  output        io_out_store,
  output        io_out_lsu,
  output        io_out_add,
  output        io_out_sub,
  output        io_out_land,
  output        io_out_lor,
  output        io_out_lxor,
  output        io_out_sll,
  output        io_out_sra,
  output        io_out_srl,
  output        io_out_slt,
  output        io_out_unsign,
  output        io_out_condbr,
  output        io_out_beq,
  output        io_out_bne,
  output        io_out_bge,
  output        io_out_blt,
  output        io_out_jal,
  output        io_out_by,
  output        io_out_half,
  output        io_out_word,
  output        io_out_csr_read,
  output        io_out_csr_clr,
  output        io_out_csr_set,
  output        io_out_csr_write,
  output        io_out_csr_imm,
  output        io_out_presync,
  output        io_out_postsync,
  output        io_out_ebreak,
  output        io_out_ecall,
  output        io_out_mret,
  output        io_out_mul,
  output        io_out_rs1_sign,
  output        io_out_rs2_sign,
  output        io_out_low,
  output        io_out_div,
  output        io_out_rem,
  output        io_out_fence,
  output        io_out_fence_i,
  output        io_out_pm_alu,
  output        io_out_legal
);
  wire  _T_2 = io_ins[2] | io_ins[6]; // @[dec_dec_ctl.scala 20:27]
  wire  _T_4 = ~io_ins[25]; // @[dec_dec_ctl.scala 20:42]
  wire  _T_6 = _T_4 & io_ins[4]; // @[dec_dec_ctl.scala 20:53]
  wire  _T_7 = _T_2 | _T_6; // @[dec_dec_ctl.scala 20:39]
  wire  _T_9 = ~io_ins[5]; // @[dec_dec_ctl.scala 20:68]
  wire  _T_11 = _T_9 & io_ins[4]; // @[dec_dec_ctl.scala 20:78]
  wire  _T_14 = ~io_ins[14]; // @[dec_dec_ctl.scala 15:46]
  wire  _T_16 = ~io_ins[13]; // @[dec_dec_ctl.scala 15:46]
  wire  _T_18 = ~io_ins[2]; // @[dec_dec_ctl.scala 15:46]
  wire  _T_19 = _T_14 & _T_16; // @[dec_dec_ctl.scala 17:17]
  wire  _T_20 = _T_19 & _T_18; // @[dec_dec_ctl.scala 17:17]
  wire  _T_26 = _T_16 & io_ins[11]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_27 = _T_26 & _T_18; // @[dec_dec_ctl.scala 17:17]
  wire  _T_28 = _T_20 | _T_27; // @[dec_dec_ctl.scala 21:43]
  wire  _T_33 = io_ins[19] & io_ins[13]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_34 = _T_33 & _T_18; // @[dec_dec_ctl.scala 17:17]
  wire  _T_35 = _T_28 | _T_34; // @[dec_dec_ctl.scala 21:70]
  wire  _T_41 = _T_16 & io_ins[10]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_42 = _T_41 & _T_18; // @[dec_dec_ctl.scala 17:17]
  wire  _T_43 = _T_35 | _T_42; // @[dec_dec_ctl.scala 22:29]
  wire  _T_48 = io_ins[18] & io_ins[13]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_49 = _T_48 & _T_18; // @[dec_dec_ctl.scala 17:17]
  wire  _T_50 = _T_43 | _T_49; // @[dec_dec_ctl.scala 22:56]
  wire  _T_56 = _T_16 & io_ins[9]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_57 = _T_56 & _T_18; // @[dec_dec_ctl.scala 17:17]
  wire  _T_58 = _T_50 | _T_57; // @[dec_dec_ctl.scala 23:29]
  wire  _T_63 = io_ins[17] & io_ins[13]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_64 = _T_63 & _T_18; // @[dec_dec_ctl.scala 17:17]
  wire  _T_65 = _T_58 | _T_64; // @[dec_dec_ctl.scala 23:55]
  wire  _T_71 = _T_16 & io_ins[8]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_72 = _T_71 & _T_18; // @[dec_dec_ctl.scala 17:17]
  wire  _T_73 = _T_65 | _T_72; // @[dec_dec_ctl.scala 24:29]
  wire  _T_78 = io_ins[16] & io_ins[13]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_79 = _T_78 & _T_18; // @[dec_dec_ctl.scala 17:17]
  wire  _T_80 = _T_73 | _T_79; // @[dec_dec_ctl.scala 24:55]
  wire  _T_86 = _T_16 & io_ins[7]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_87 = _T_86 & _T_18; // @[dec_dec_ctl.scala 17:17]
  wire  _T_88 = _T_80 | _T_87; // @[dec_dec_ctl.scala 25:29]
  wire  _T_93 = io_ins[15] & io_ins[13]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_94 = _T_93 & _T_18; // @[dec_dec_ctl.scala 17:17]
  wire  _T_95 = _T_88 | _T_94; // @[dec_dec_ctl.scala 25:55]
  wire  _T_97 = ~io_ins[4]; // @[dec_dec_ctl.scala 15:46]
  wire  _T_99 = ~io_ins[3]; // @[dec_dec_ctl.scala 15:46]
  wire  _T_100 = _T_97 & _T_99; // @[dec_dec_ctl.scala 17:17]
  wire  _T_101 = _T_95 | _T_100; // @[dec_dec_ctl.scala 26:29]
  wire  _T_103 = ~io_ins[6]; // @[dec_dec_ctl.scala 15:46]
  wire  _T_106 = _T_103 & _T_18; // @[dec_dec_ctl.scala 17:17]
  wire  _T_113 = io_ins[5] & _T_97; // @[dec_dec_ctl.scala 17:17]
  wire  _T_114 = _T_113 & _T_18; // @[dec_dec_ctl.scala 17:17]
  wire  _T_120 = _T_103 & io_ins[5]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_121 = _T_120 & _T_18; // @[dec_dec_ctl.scala 17:17]
  wire  _T_129 = _T_100 & io_ins[2]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_136 = io_ins[13] & _T_9; // @[dec_dec_ctl.scala 17:17]
  wire  _T_137 = _T_136 & io_ins[4]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_138 = _T_137 & _T_18; // @[dec_dec_ctl.scala 17:17]
  wire  _T_139 = _T_129 | _T_138; // @[dec_dec_ctl.scala 28:42]
  wire  _T_143 = ~io_ins[12]; // @[dec_dec_ctl.scala 15:46]
  wire  _T_146 = _T_16 & _T_143; // @[dec_dec_ctl.scala 17:17]
  wire  _T_147 = _T_146 & io_ins[6]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_148 = _T_147 & io_ins[4]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_149 = _T_139 | _T_148; // @[dec_dec_ctl.scala 28:70]
  wire  _T_157 = _T_143 & _T_9; // @[dec_dec_ctl.scala 17:17]
  wire  _T_158 = _T_157 & io_ins[4]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_159 = _T_158 & _T_18; // @[dec_dec_ctl.scala 17:17]
  wire  _T_165 = _T_9 & _T_18; // @[dec_dec_ctl.scala 30:28]
  wire  _T_168 = io_ins[5] & io_ins[2]; // @[dec_dec_ctl.scala 30:55]
  wire  _T_169 = _T_165 | _T_168; // @[dec_dec_ctl.scala 30:42]
  wire  _T_180 = _T_16 & io_ins[12]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_181 = _T_180 & _T_9; // @[dec_dec_ctl.scala 17:17]
  wire  _T_182 = _T_181 & io_ins[4]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_186 = io_ins[5] & io_ins[3]; // @[dec_dec_ctl.scala 32:29]
  wire  _T_189 = io_ins[4] & io_ins[2]; // @[dec_dec_ctl.scala 32:53]
  wire  _T_195 = _T_9 & _T_99; // @[dec_dec_ctl.scala 33:28]
  wire  _T_197 = _T_195 & io_ins[2]; // @[dec_dec_ctl.scala 33:41]
  wire  _T_208 = _T_9 & _T_97; // @[dec_dec_ctl.scala 17:17]
  wire  _T_223 = _T_103 & _T_97; // @[dec_dec_ctl.scala 17:17]
  wire  _T_235 = _T_19 & _T_143; // @[dec_dec_ctl.scala 17:17]
  wire  _T_236 = _T_235 & _T_9; // @[dec_dec_ctl.scala 17:17]
  wire  _T_237 = _T_236 & io_ins[4]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_245 = _T_237 | _T_197; // @[dec_dec_ctl.scala 37:49]
  wire  _T_247 = ~io_ins[30]; // @[dec_dec_ctl.scala 15:46]
  wire  _T_261 = _T_247 & _T_4; // @[dec_dec_ctl.scala 17:17]
  wire  _T_262 = _T_261 & _T_14; // @[dec_dec_ctl.scala 17:17]
  wire  _T_263 = _T_262 & _T_16; // @[dec_dec_ctl.scala 17:17]
  wire  _T_264 = _T_263 & _T_143; // @[dec_dec_ctl.scala 17:17]
  wire  _T_265 = _T_264 & _T_103; // @[dec_dec_ctl.scala 17:17]
  wire  _T_266 = _T_265 & io_ins[4]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_267 = _T_266 & _T_18; // @[dec_dec_ctl.scala 17:17]
  wire  _T_278 = io_ins[30] & _T_143; // @[dec_dec_ctl.scala 17:17]
  wire  _T_279 = _T_278 & _T_103; // @[dec_dec_ctl.scala 17:17]
  wire  _T_280 = _T_279 & io_ins[5]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_281 = _T_280 & io_ins[4]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_282 = _T_281 & _T_18; // @[dec_dec_ctl.scala 17:17]
  wire  _T_293 = _T_4 & _T_14; // @[dec_dec_ctl.scala 17:17]
  wire  _T_294 = _T_293 & io_ins[13]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_295 = _T_294 & _T_103; // @[dec_dec_ctl.scala 17:17]
  wire  _T_296 = _T_295 & io_ins[4]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_297 = _T_296 & _T_18; // @[dec_dec_ctl.scala 17:17]
  wire  _T_298 = _T_282 | _T_297; // @[dec_dec_ctl.scala 39:49]
  wire  _T_307 = _T_14 & io_ins[13]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_308 = _T_307 & _T_9; // @[dec_dec_ctl.scala 17:17]
  wire  _T_309 = _T_308 & io_ins[4]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_310 = _T_309 & _T_18; // @[dec_dec_ctl.scala 17:17]
  wire  _T_311 = _T_298 | _T_310; // @[dec_dec_ctl.scala 39:85]
  wire  _T_317 = io_ins[6] & _T_97; // @[dec_dec_ctl.scala 17:17]
  wire  _T_318 = _T_317 & _T_18; // @[dec_dec_ctl.scala 17:17]
  wire  _T_327 = io_ins[14] & io_ins[13]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_328 = _T_327 & io_ins[12]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_329 = _T_328 & _T_9; // @[dec_dec_ctl.scala 17:17]
  wire  _T_330 = _T_329 & _T_18; // @[dec_dec_ctl.scala 17:17]
  wire  _T_340 = _T_4 & io_ins[14]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_341 = _T_340 & io_ins[13]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_342 = _T_341 & io_ins[12]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_343 = _T_342 & _T_103; // @[dec_dec_ctl.scala 17:17]
  wire  _T_344 = _T_343 & _T_18; // @[dec_dec_ctl.scala 17:17]
  wire  _T_349 = _T_103 & io_ins[3]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_362 = _T_341 & _T_143; // @[dec_dec_ctl.scala 17:17]
  wire  _T_363 = _T_362 & _T_103; // @[dec_dec_ctl.scala 17:17]
  wire  _T_364 = _T_363 & _T_18; // @[dec_dec_ctl.scala 17:17]
  wire  _T_365 = _T_349 | _T_364; // @[dec_dec_ctl.scala 42:37]
  wire  _T_369 = io_ins[5] & io_ins[4]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_370 = _T_369 & io_ins[2]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_371 = _T_365 | _T_370; // @[dec_dec_ctl.scala 42:74]
  wire  _T_381 = _T_371 | _T_148; // @[dec_dec_ctl.scala 43:26]
  wire  _T_391 = _T_327 & _T_143; // @[dec_dec_ctl.scala 17:17]
  wire  _T_392 = _T_391 & _T_9; // @[dec_dec_ctl.scala 17:17]
  wire  _T_393 = _T_392 & _T_18; // @[dec_dec_ctl.scala 17:17]
  wire  _T_406 = _T_340 & _T_16; // @[dec_dec_ctl.scala 17:17]
  wire  _T_407 = _T_406 & _T_143; // @[dec_dec_ctl.scala 17:17]
  wire  _T_408 = _T_407 & io_ins[4]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_409 = _T_408 & _T_18; // @[dec_dec_ctl.scala 17:17]
  wire  _T_420 = io_ins[14] & _T_16; // @[dec_dec_ctl.scala 17:17]
  wire  _T_421 = _T_420 & _T_143; // @[dec_dec_ctl.scala 17:17]
  wire  _T_422 = _T_421 & _T_9; // @[dec_dec_ctl.scala 17:17]
  wire  _T_423 = _T_422 & io_ins[4]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_424 = _T_423 & _T_18; // @[dec_dec_ctl.scala 17:17]
  wire  _T_439 = _T_293 & _T_16; // @[dec_dec_ctl.scala 17:17]
  wire  _T_440 = _T_439 & io_ins[12]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_441 = _T_440 & _T_103; // @[dec_dec_ctl.scala 17:17]
  wire  _T_442 = _T_441 & io_ins[4]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_453 = io_ins[30] & _T_16; // @[dec_dec_ctl.scala 17:17]
  wire  _T_454 = _T_453 & io_ins[12]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_455 = _T_454 & _T_103; // @[dec_dec_ctl.scala 17:17]
  wire  _T_456 = _T_455 & io_ins[4]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_472 = _T_261 & io_ins[14]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_473 = _T_472 & _T_16; // @[dec_dec_ctl.scala 17:17]
  wire  _T_474 = _T_473 & io_ins[12]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_475 = _T_474 & _T_103; // @[dec_dec_ctl.scala 17:17]
  wire  _T_476 = _T_475 & io_ins[4]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_515 = _T_307 & io_ins[12]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_516 = _T_515 & _T_9; // @[dec_dec_ctl.scala 17:17]
  wire  _T_517 = _T_516 & _T_18; // @[dec_dec_ctl.scala 17:17]
  wire  _T_524 = io_ins[13] & io_ins[6]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_525 = _T_524 & _T_97; // @[dec_dec_ctl.scala 17:17]
  wire  _T_526 = _T_525 & _T_18; // @[dec_dec_ctl.scala 17:17]
  wire  _T_527 = _T_517 | _T_526; // @[dec_dec_ctl.scala 50:51]
  wire  _T_533 = io_ins[14] & _T_9; // @[dec_dec_ctl.scala 17:17]
  wire  _T_534 = _T_533 & _T_97; // @[dec_dec_ctl.scala 17:17]
  wire  _T_535 = _T_527 | _T_534; // @[dec_dec_ctl.scala 50:79]
  wire  _T_548 = _T_294 & io_ins[12]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_549 = _T_548 & _T_103; // @[dec_dec_ctl.scala 17:17]
  wire  _T_550 = _T_549 & _T_18; // @[dec_dec_ctl.scala 17:17]
  wire  _T_551 = _T_535 | _T_550; // @[dec_dec_ctl.scala 51:29]
  wire  _T_560 = io_ins[25] & io_ins[14]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_561 = _T_560 & io_ins[12]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_562 = _T_561 & _T_103; // @[dec_dec_ctl.scala 17:17]
  wire  _T_563 = _T_562 & io_ins[5]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_564 = _T_563 & _T_18; // @[dec_dec_ctl.scala 17:17]
  wire  _T_582 = _T_14 & _T_143; // @[dec_dec_ctl.scala 17:17]
  wire  _T_583 = _T_582 & io_ins[6]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_584 = _T_583 & _T_97; // @[dec_dec_ctl.scala 17:17]
  wire  _T_594 = _T_14 & io_ins[12]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_595 = _T_594 & io_ins[6]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_596 = _T_595 & _T_97; // @[dec_dec_ctl.scala 17:17]
  wire  _T_605 = io_ins[14] & io_ins[12]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_606 = _T_605 & io_ins[5]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_607 = _T_606 & _T_97; // @[dec_dec_ctl.scala 17:17]
  wire  _T_617 = io_ins[14] & _T_143; // @[dec_dec_ctl.scala 17:17]
  wire  _T_618 = _T_617 & io_ins[5]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_619 = _T_618 & _T_97; // @[dec_dec_ctl.scala 17:17]
  wire  _T_635 = _T_146 & _T_103; // @[dec_dec_ctl.scala 17:17]
  wire  _T_636 = _T_635 & _T_97; // @[dec_dec_ctl.scala 17:17]
  wire  _T_645 = io_ins[12] & _T_103; // @[dec_dec_ctl.scala 17:17]
  wire  _T_646 = _T_645 & _T_97; // @[dec_dec_ctl.scala 17:17]
  wire  _T_653 = io_ins[13] & _T_103; // @[dec_dec_ctl.scala 17:17]
  wire  _T_659 = _T_524 & io_ins[4]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_663 = io_ins[7] & io_ins[6]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_664 = _T_663 & io_ins[4]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_665 = _T_659 | _T_664; // @[dec_dec_ctl.scala 62:44]
  wire  _T_669 = io_ins[8] & io_ins[6]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_670 = _T_669 & io_ins[4]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_671 = _T_665 | _T_670; // @[dec_dec_ctl.scala 62:67]
  wire  _T_675 = io_ins[9] & io_ins[6]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_676 = _T_675 & io_ins[4]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_677 = _T_671 | _T_676; // @[dec_dec_ctl.scala 63:26]
  wire  _T_681 = io_ins[10] & io_ins[6]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_682 = _T_681 & io_ins[4]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_683 = _T_677 | _T_682; // @[dec_dec_ctl.scala 63:49]
  wire  _T_687 = io_ins[11] & io_ins[6]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_688 = _T_687 & io_ins[4]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_696 = _T_93 & io_ins[12]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_697 = _T_696 & io_ins[6]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_698 = _T_697 & io_ins[4]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_705 = _T_78 & io_ins[12]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_706 = _T_705 & io_ins[6]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_707 = _T_706 & io_ins[4]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_708 = _T_698 | _T_707; // @[dec_dec_ctl.scala 65:49]
  wire  _T_715 = _T_63 & io_ins[12]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_716 = _T_715 & io_ins[6]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_717 = _T_716 & io_ins[4]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_718 = _T_708 | _T_717; // @[dec_dec_ctl.scala 65:79]
  wire  _T_725 = _T_48 & io_ins[12]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_726 = _T_725 & io_ins[6]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_727 = _T_726 & io_ins[4]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_728 = _T_718 | _T_727; // @[dec_dec_ctl.scala 66:33]
  wire  _T_735 = _T_33 & io_ins[12]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_736 = _T_735 & io_ins[6]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_737 = _T_736 & io_ins[4]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_745 = _T_180 & io_ins[6]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_753 = _T_420 & io_ins[6]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_754 = _T_753 & io_ins[4]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_759 = io_ins[15] & io_ins[14]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_760 = _T_759 & io_ins[6]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_761 = _T_760 & io_ins[4]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_762 = _T_754 | _T_761; // @[dec_dec_ctl.scala 69:47]
  wire  _T_767 = io_ins[16] & io_ins[14]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_768 = _T_767 & io_ins[6]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_769 = _T_768 & io_ins[4]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_770 = _T_762 | _T_769; // @[dec_dec_ctl.scala 69:74]
  wire  _T_775 = io_ins[17] & io_ins[14]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_776 = _T_775 & io_ins[6]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_777 = _T_776 & io_ins[4]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_778 = _T_770 | _T_777; // @[dec_dec_ctl.scala 70:30]
  wire  _T_783 = io_ins[18] & io_ins[14]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_784 = _T_783 & io_ins[6]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_785 = _T_784 & io_ins[4]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_786 = _T_778 | _T_785; // @[dec_dec_ctl.scala 70:57]
  wire  _T_791 = io_ins[19] & io_ins[14]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_792 = _T_791 & io_ins[6]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_793 = _T_792 & io_ins[4]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_800 = io_ins[15] & _T_143; // @[dec_dec_ctl.scala 17:17]
  wire  _T_801 = _T_800 & io_ins[6]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_802 = _T_801 & io_ins[4]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_808 = io_ins[16] & _T_143; // @[dec_dec_ctl.scala 17:17]
  wire  _T_809 = _T_808 & io_ins[6]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_810 = _T_809 & io_ins[4]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_811 = _T_802 | _T_810; // @[dec_dec_ctl.scala 72:47]
  wire  _T_817 = io_ins[17] & _T_143; // @[dec_dec_ctl.scala 17:17]
  wire  _T_818 = _T_817 & io_ins[6]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_819 = _T_818 & io_ins[4]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_820 = _T_811 | _T_819; // @[dec_dec_ctl.scala 72:75]
  wire  _T_826 = io_ins[18] & _T_143; // @[dec_dec_ctl.scala 17:17]
  wire  _T_827 = _T_826 & io_ins[6]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_828 = _T_827 & io_ins[4]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_829 = _T_820 | _T_828; // @[dec_dec_ctl.scala 73:31]
  wire  _T_835 = io_ins[19] & _T_143; // @[dec_dec_ctl.scala 17:17]
  wire  _T_836 = _T_835 & io_ins[6]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_837 = _T_836 & io_ins[4]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_840 = ~io_ins[22]; // @[dec_dec_ctl.scala 15:46]
  wire  _T_848 = _T_840 & io_ins[20]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_849 = _T_848 & _T_16; // @[dec_dec_ctl.scala 17:17]
  wire  _T_850 = _T_849 & _T_143; // @[dec_dec_ctl.scala 17:17]
  wire  _T_851 = _T_850 & io_ins[6]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_854 = ~io_ins[21]; // @[dec_dec_ctl.scala 15:46]
  wire  _T_856 = ~io_ins[20]; // @[dec_dec_ctl.scala 15:46]
  wire  _T_863 = _T_854 & _T_856; // @[dec_dec_ctl.scala 17:17]
  wire  _T_864 = _T_863 & _T_16; // @[dec_dec_ctl.scala 17:17]
  wire  _T_865 = _T_864 & _T_143; // @[dec_dec_ctl.scala 17:17]
  wire  _T_866 = _T_865 & io_ins[6]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_875 = io_ins[29] & _T_16; // @[dec_dec_ctl.scala 17:17]
  wire  _T_876 = _T_875 & _T_143; // @[dec_dec_ctl.scala 17:17]
  wire  _T_877 = _T_876 & io_ins[6]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_888 = io_ins[25] & _T_14; // @[dec_dec_ctl.scala 17:17]
  wire  _T_889 = _T_888 & _T_103; // @[dec_dec_ctl.scala 17:17]
  wire  _T_890 = _T_889 & io_ins[5]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_891 = _T_890 & io_ins[4]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_906 = _T_888 & io_ins[13]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_907 = _T_906 & _T_143; // @[dec_dec_ctl.scala 17:17]
  wire  _T_908 = _T_907 & _T_103; // @[dec_dec_ctl.scala 17:17]
  wire  _T_909 = _T_908 & io_ins[5]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_910 = _T_909 & io_ins[4]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_911 = _T_910 & _T_18; // @[dec_dec_ctl.scala 17:17]
  wire  _T_924 = _T_888 & _T_16; // @[dec_dec_ctl.scala 17:17]
  wire  _T_925 = _T_924 & io_ins[12]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_926 = _T_925 & _T_103; // @[dec_dec_ctl.scala 17:17]
  wire  _T_927 = _T_926 & io_ins[4]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_928 = _T_927 & _T_18; // @[dec_dec_ctl.scala 17:17]
  wire  _T_960 = _T_924 & _T_143; // @[dec_dec_ctl.scala 17:17]
  wire  _T_961 = _T_960 & io_ins[5]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_962 = _T_961 & io_ins[4]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_972 = _T_560 & _T_103; // @[dec_dec_ctl.scala 17:17]
  wire  _T_973 = _T_972 & io_ins[5]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_984 = _T_560 & io_ins[13]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_985 = _T_984 & _T_103; // @[dec_dec_ctl.scala 17:17]
  wire  _T_986 = _T_985 & io_ins[5]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_991 = _T_9 & io_ins[3]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_996 = io_ins[12] & _T_9; // @[dec_dec_ctl.scala 17:17]
  wire  _T_997 = _T_996 & io_ins[3]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1005 = io_ins[28] & io_ins[22]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1006 = _T_1005 & _T_16; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1007 = _T_1006 & _T_143; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1008 = _T_1007 & io_ins[4]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1012 = _T_1008 | _T_189; // @[dec_dec_ctl.scala 87:51]
  wire  _T_1018 = _T_4 & _T_103; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1019 = _T_1018 & io_ins[4]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1020 = _T_1012 | _T_1019; // @[dec_dec_ctl.scala 87:72]
  wire  _T_1036 = _T_86 & io_ins[6]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1037 = _T_1036 & io_ins[4]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1038 = _T_991 | _T_1037; // @[dec_dec_ctl.scala 89:41]
  wire  _T_1045 = _T_71 & io_ins[6]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1046 = _T_1045 & io_ins[4]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1047 = _T_1038 | _T_1046; // @[dec_dec_ctl.scala 89:68]
  wire  _T_1054 = _T_56 & io_ins[6]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1055 = _T_1054 & io_ins[4]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1056 = _T_1047 | _T_1055; // @[dec_dec_ctl.scala 90:30]
  wire  _T_1063 = _T_41 & io_ins[6]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1064 = _T_1063 & io_ins[4]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1065 = _T_1056 | _T_1064; // @[dec_dec_ctl.scala 90:57]
  wire  _T_1072 = _T_26 & io_ins[6]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1073 = _T_1072 & io_ins[4]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1074 = _T_1065 | _T_1073; // @[dec_dec_ctl.scala 91:31]
  wire  _T_1080 = _T_93 & io_ins[6]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1081 = _T_1080 & io_ins[4]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1082 = _T_1074 | _T_1081; // @[dec_dec_ctl.scala 91:59]
  wire  _T_1088 = _T_78 & io_ins[6]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1089 = _T_1088 & io_ins[4]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1090 = _T_1082 | _T_1089; // @[dec_dec_ctl.scala 92:30]
  wire  _T_1096 = _T_63 & io_ins[6]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1097 = _T_1096 & io_ins[4]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1098 = _T_1090 | _T_1097; // @[dec_dec_ctl.scala 92:57]
  wire  _T_1104 = _T_48 & io_ins[6]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1105 = _T_1104 & io_ins[4]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1106 = _T_1098 | _T_1105; // @[dec_dec_ctl.scala 93:30]
  wire  _T_1112 = _T_33 & io_ins[6]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1113 = _T_1112 & io_ins[4]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1129 = _T_840 & _T_16; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1130 = _T_1129 & _T_143; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1131 = _T_1130 & io_ins[6]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1132 = _T_1131 & io_ins[4]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1133 = _T_997 | _T_1132; // @[dec_dec_ctl.scala 95:45]
  wire  _T_1142 = _T_1133 | _T_1037; // @[dec_dec_ctl.scala 95:78]
  wire  _T_1151 = _T_1142 | _T_1046; // @[dec_dec_ctl.scala 96:30]
  wire  _T_1160 = _T_1151 | _T_1055; // @[dec_dec_ctl.scala 96:57]
  wire  _T_1169 = _T_1160 | _T_1064; // @[dec_dec_ctl.scala 97:30]
  wire  _T_1178 = _T_1169 | _T_1073; // @[dec_dec_ctl.scala 97:58]
  wire  _T_1186 = _T_1178 | _T_1081; // @[dec_dec_ctl.scala 98:31]
  wire  _T_1194 = _T_1186 | _T_1089; // @[dec_dec_ctl.scala 98:58]
  wire  _T_1202 = _T_1194 | _T_1097; // @[dec_dec_ctl.scala 99:30]
  wire  _T_1210 = _T_1202 | _T_1105; // @[dec_dec_ctl.scala 99:57]
  wire  _T_1220 = ~io_ins[31]; // @[dec_dec_ctl.scala 15:46]
  wire  _T_1226 = ~io_ins[27]; // @[dec_dec_ctl.scala 15:46]
  wire  _T_1228 = ~io_ins[26]; // @[dec_dec_ctl.scala 15:46]
  wire  _T_1232 = ~io_ins[24]; // @[dec_dec_ctl.scala 15:46]
  wire  _T_1234 = ~io_ins[23]; // @[dec_dec_ctl.scala 15:46]
  wire  _T_1241 = ~io_ins[19]; // @[dec_dec_ctl.scala 15:46]
  wire  _T_1243 = ~io_ins[18]; // @[dec_dec_ctl.scala 15:46]
  wire  _T_1245 = ~io_ins[17]; // @[dec_dec_ctl.scala 15:46]
  wire  _T_1247 = ~io_ins[16]; // @[dec_dec_ctl.scala 15:46]
  wire  _T_1249 = ~io_ins[15]; // @[dec_dec_ctl.scala 15:46]
  wire  _T_1253 = ~io_ins[11]; // @[dec_dec_ctl.scala 15:46]
  wire  _T_1255 = ~io_ins[10]; // @[dec_dec_ctl.scala 15:46]
  wire  _T_1257 = ~io_ins[9]; // @[dec_dec_ctl.scala 15:46]
  wire  _T_1259 = ~io_ins[8]; // @[dec_dec_ctl.scala 15:46]
  wire  _T_1261 = ~io_ins[7]; // @[dec_dec_ctl.scala 15:46]
  wire  _T_1271 = _T_1220 & _T_247; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1272 = _T_1271 & io_ins[29]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1273 = _T_1272 & io_ins[28]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1274 = _T_1273 & _T_1226; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1275 = _T_1274 & _T_1228; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1276 = _T_1275 & _T_4; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1277 = _T_1276 & _T_1232; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1278 = _T_1277 & _T_1234; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1279 = _T_1278 & _T_840; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1280 = _T_1279 & io_ins[21]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1281 = _T_1280 & _T_856; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1282 = _T_1281 & _T_1241; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1283 = _T_1282 & _T_1243; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1284 = _T_1283 & _T_1245; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1285 = _T_1284 & _T_1247; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1286 = _T_1285 & _T_1249; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1287 = _T_1286 & _T_14; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1288 = _T_1287 & _T_1253; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1289 = _T_1288 & _T_1255; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1290 = _T_1289 & _T_1257; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1291 = _T_1290 & _T_1259; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1292 = _T_1291 & _T_1261; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1293 = _T_1292 & io_ins[6]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1294 = _T_1293 & io_ins[5]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1295 = _T_1294 & io_ins[4]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1296 = _T_1295 & _T_99; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1297 = _T_1296 & _T_18; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1298 = _T_1297 & io_ins[1]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1299 = _T_1298 & io_ins[0]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1305 = ~io_ins[29]; // @[dec_dec_ctl.scala 15:46]
  wire  _T_1353 = _T_1271 & _T_1305; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1354 = _T_1353 & io_ins[28]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1355 = _T_1354 & _T_1226; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1356 = _T_1355 & _T_1228; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1357 = _T_1356 & _T_4; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1358 = _T_1357 & _T_1232; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1359 = _T_1358 & _T_1234; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1360 = _T_1359 & io_ins[22]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1361 = _T_1360 & _T_854; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1362 = _T_1361 & io_ins[20]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1363 = _T_1362 & _T_1241; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1364 = _T_1363 & _T_1243; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1365 = _T_1364 & _T_1245; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1366 = _T_1365 & _T_1247; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1367 = _T_1366 & _T_1249; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1368 = _T_1367 & _T_14; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1369 = _T_1368 & _T_1253; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1370 = _T_1369 & _T_1255; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1371 = _T_1370 & _T_1257; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1372 = _T_1371 & _T_1259; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1373 = _T_1372 & _T_1261; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1374 = _T_1373 & io_ins[6]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1375 = _T_1374 & io_ins[5]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1376 = _T_1375 & io_ins[4]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1377 = _T_1376 & _T_99; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1378 = _T_1377 & _T_18; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1379 = _T_1378 & io_ins[1]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1380 = _T_1379 & io_ins[0]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1381 = _T_1299 | _T_1380; // @[dec_dec_ctl.scala 101:136]
  wire  _T_1389 = ~io_ins[28]; // @[dec_dec_ctl.scala 15:46]
  wire  _T_1436 = _T_1353 & _T_1389; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1437 = _T_1436 & _T_1226; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1438 = _T_1437 & _T_1228; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1439 = _T_1438 & _T_4; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1440 = _T_1439 & _T_1232; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1441 = _T_1440 & _T_1234; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1442 = _T_1441 & _T_840; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1443 = _T_1442 & _T_854; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1444 = _T_1443 & _T_1241; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1445 = _T_1444 & _T_1243; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1446 = _T_1445 & _T_1245; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1447 = _T_1446 & _T_1247; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1448 = _T_1447 & _T_1249; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1449 = _T_1448 & _T_14; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1450 = _T_1449 & _T_1253; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1451 = _T_1450 & _T_1255; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1452 = _T_1451 & _T_1257; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1453 = _T_1452 & _T_1259; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1454 = _T_1453 & _T_1261; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1455 = _T_1454 & io_ins[5]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1456 = _T_1455 & io_ins[4]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1457 = _T_1456 & _T_99; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1458 = _T_1457 & _T_18; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1459 = _T_1458 & io_ins[1]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1460 = _T_1459 & io_ins[0]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1461 = _T_1381 | _T_1460; // @[dec_dec_ctl.scala 102:122]
  wire  _T_1489 = _T_1439 & _T_103; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1490 = _T_1489 & io_ins[4]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1491 = _T_1490 & _T_99; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1492 = _T_1491 & io_ins[1]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1493 = _T_1492 & io_ins[0]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1494 = _T_1461 | _T_1493; // @[dec_dec_ctl.scala 103:119]
  wire  _T_1521 = _T_1220 & _T_1305; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1522 = _T_1521 & _T_1389; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1523 = _T_1522 & _T_1226; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1524 = _T_1523 & _T_1228; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1525 = _T_1524 & _T_4; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1526 = _T_1525 & _T_14; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1527 = _T_1526 & _T_16; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1528 = _T_1527 & _T_143; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1529 = _T_1528 & _T_103; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1530 = _T_1529 & _T_99; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1531 = _T_1530 & _T_18; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1532 = _T_1531 & io_ins[1]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1533 = _T_1532 & io_ins[0]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1534 = _T_1494 | _T_1533; // @[dec_dec_ctl.scala 104:60]
  wire  _T_1563 = _T_1525 & io_ins[14]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1564 = _T_1563 & _T_16; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1565 = _T_1564 & io_ins[12]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1566 = _T_1565 & _T_103; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1567 = _T_1566 & io_ins[4]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1568 = _T_1567 & _T_99; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1569 = _T_1568 & io_ins[1]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1570 = _T_1569 & io_ins[0]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1571 = _T_1534 | _T_1570; // @[dec_dec_ctl.scala 105:69]
  wire  _T_1597 = _T_1438 & _T_103; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1598 = _T_1597 & io_ins[5]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1599 = _T_1598 & io_ins[4]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1600 = _T_1599 & _T_99; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1601 = _T_1600 & io_ins[1]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1602 = _T_1601 & io_ins[0]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1603 = _T_1571 | _T_1602; // @[dec_dec_ctl.scala 106:66]
  wire  _T_1620 = _T_235 & io_ins[6]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1621 = _T_1620 & io_ins[5]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1622 = _T_1621 & _T_97; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1623 = _T_1622 & _T_99; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1624 = _T_1623 & io_ins[1]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1625 = _T_1624 & io_ins[0]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1626 = _T_1603 | _T_1625; // @[dec_dec_ctl.scala 107:58]
  wire  _T_1638 = io_ins[14] & io_ins[6]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1639 = _T_1638 & io_ins[5]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1640 = _T_1639 & _T_97; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1641 = _T_1640 & _T_99; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1642 = _T_1641 & _T_18; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1643 = _T_1642 & io_ins[1]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1644 = _T_1643 & io_ins[0]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1645 = _T_1626 | _T_1644; // @[dec_dec_ctl.scala 108:46]
  wire  _T_1657 = _T_143 & _T_103; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1658 = _T_1657 & _T_9; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1659 = _T_1658 & io_ins[4]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1660 = _T_1659 & _T_99; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1661 = _T_1660 & io_ins[1]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1662 = _T_1661 & io_ins[0]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1663 = _T_1645 | _T_1662; // @[dec_dec_ctl.scala 109:40]
  wire  _T_1678 = _T_19 & io_ins[5]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1679 = _T_1678 & _T_97; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1680 = _T_1679 & _T_99; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1681 = _T_1680 & _T_18; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1682 = _T_1681 & io_ins[1]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1683 = _T_1682 & io_ins[0]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1684 = _T_1663 | _T_1683; // @[dec_dec_ctl.scala 110:39]
  wire  _T_1695 = io_ins[12] & io_ins[6]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1696 = _T_1695 & io_ins[5]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1697 = _T_1696 & io_ins[4]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1698 = _T_1697 & _T_99; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1699 = _T_1698 & _T_18; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1700 = _T_1699 & io_ins[1]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1701 = _T_1700 & io_ins[0]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1702 = _T_1684 | _T_1701; // @[dec_dec_ctl.scala 111:43]
  wire  _T_1771 = _T_1443 & _T_856; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1772 = _T_1771 & _T_1241; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1773 = _T_1772 & _T_1243; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1774 = _T_1773 & _T_1245; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1775 = _T_1774 & _T_1247; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1776 = _T_1775 & _T_1249; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1777 = _T_1776 & _T_14; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1778 = _T_1777 & _T_16; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1779 = _T_1778 & _T_1253; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1780 = _T_1779 & _T_1255; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1781 = _T_1780 & _T_1257; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1782 = _T_1781 & _T_1259; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1783 = _T_1782 & _T_1261; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1784 = _T_1783 & _T_103; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1785 = _T_1784 & _T_9; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1786 = _T_1785 & _T_97; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1787 = _T_1786 & io_ins[3]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1788 = _T_1787 & io_ins[2]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1789 = _T_1788 & io_ins[1]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1790 = _T_1789 & io_ins[0]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1791 = _T_1702 | _T_1790; // @[dec_dec_ctl.scala 112:39]
  wire  _T_1839 = _T_1436 & _T_1241; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1840 = _T_1839 & _T_1243; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1841 = _T_1840 & _T_1245; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1842 = _T_1841 & _T_1247; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1843 = _T_1842 & _T_1249; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1844 = _T_1843 & _T_14; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1845 = _T_1844 & _T_16; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1846 = _T_1845 & _T_143; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1847 = _T_1846 & _T_1253; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1848 = _T_1847 & _T_1255; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1849 = _T_1848 & _T_1257; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1850 = _T_1849 & _T_1259; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1851 = _T_1850 & _T_1261; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1852 = _T_1851 & _T_103; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1853 = _T_1852 & _T_9; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1854 = _T_1853 & _T_97; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1855 = _T_1854 & io_ins[3]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1856 = _T_1855 & io_ins[2]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1857 = _T_1856 & io_ins[1]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1858 = _T_1857 & io_ins[0]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1859 = _T_1791 | _T_1858; // @[dec_dec_ctl.scala 113:130]
  wire  _T_1871 = _T_524 & io_ins[5]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1872 = _T_1871 & io_ins[4]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1873 = _T_1872 & _T_99; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1874 = _T_1873 & _T_18; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1875 = _T_1874 & io_ins[1]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1876 = _T_1875 & io_ins[0]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1877 = _T_1859 | _T_1876; // @[dec_dec_ctl.scala 114:102]
  wire  _T_1892 = _T_16 & _T_103; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1893 = _T_1892 & _T_9; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1894 = _T_1893 & _T_97; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1895 = _T_1894 & _T_99; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1896 = _T_1895 & _T_18; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1897 = _T_1896 & io_ins[1]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1898 = _T_1897 & io_ins[0]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1899 = _T_1877 | _T_1898; // @[dec_dec_ctl.scala 115:39]
  wire  _T_1908 = io_ins[6] & io_ins[5]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1909 = _T_1908 & _T_97; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1910 = _T_1909 & io_ins[3]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1911 = _T_1910 & io_ins[2]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1912 = _T_1911 & io_ins[1]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1913 = _T_1912 & io_ins[0]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1914 = _T_1899 | _T_1913; // @[dec_dec_ctl.scala 116:43]
  wire  _T_1926 = _T_653 & _T_9; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1927 = _T_1926 & io_ins[4]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1928 = _T_1927 & _T_99; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1929 = _T_1928 & io_ins[1]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1930 = _T_1929 & io_ins[0]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1931 = _T_1914 | _T_1930; // @[dec_dec_ctl.scala 117:35]
  wire  _T_1947 = _T_582 & _T_103; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1948 = _T_1947 & _T_97; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1949 = _T_1948 & _T_99; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1950 = _T_1949 & _T_18; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1951 = _T_1950 & io_ins[1]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1952 = _T_1951 & io_ins[0]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1953 = _T_1931 | _T_1952; // @[dec_dec_ctl.scala 118:38]
  wire  _T_1962 = _T_103 & io_ins[4]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1963 = _T_1962 & _T_99; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1964 = _T_1963 & io_ins[2]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1965 = _T_1964 & io_ins[1]; // @[dec_dec_ctl.scala 17:17]
  wire  _T_1966 = _T_1965 & io_ins[0]; // @[dec_dec_ctl.scala 17:17]
  assign io_out_alu = _T_7 | _T_11; // @[dec_dec_ctl.scala 20:14]
  assign io_out_rs1 = _T_101 | _T_106; // @[dec_dec_ctl.scala 21:14]
  assign io_out_rs2 = _T_114 | _T_121; // @[dec_dec_ctl.scala 27:14]
  assign io_out_imm12 = _T_149 | _T_159; // @[dec_dec_ctl.scala 28:16]
  assign io_out_rd = _T_169 | io_ins[4]; // @[dec_dec_ctl.scala 30:13]
  assign io_out_shimm5 = _T_182 & _T_18; // @[dec_dec_ctl.scala 31:17]
  assign io_out_imm20 = _T_186 | _T_189; // @[dec_dec_ctl.scala 32:16]
  assign io_out_pc = _T_197 | _T_186; // @[dec_dec_ctl.scala 33:13]
  assign io_out_load = _T_208 & _T_18; // @[dec_dec_ctl.scala 34:15]
  assign io_out_store = _T_120 & _T_97; // @[dec_dec_ctl.scala 35:16]
  assign io_out_lsu = _T_223 & _T_18; // @[dec_dec_ctl.scala 36:14]
  assign io_out_add = _T_245 | _T_267; // @[dec_dec_ctl.scala 37:14]
  assign io_out_sub = _T_311 | _T_318; // @[dec_dec_ctl.scala 39:14]
  assign io_out_land = _T_330 | _T_344; // @[dec_dec_ctl.scala 41:15]
  assign io_out_lor = _T_381 | _T_393; // @[dec_dec_ctl.scala 42:14]
  assign io_out_lxor = _T_409 | _T_424; // @[dec_dec_ctl.scala 45:15]
  assign io_out_sll = _T_442 & _T_18; // @[dec_dec_ctl.scala 46:14]
  assign io_out_sra = _T_456 & _T_18; // @[dec_dec_ctl.scala 47:14]
  assign io_out_srl = _T_476 & _T_18; // @[dec_dec_ctl.scala 48:14]
  assign io_out_slt = _T_297 | _T_310; // @[dec_dec_ctl.scala 49:14]
  assign io_out_unsign = _T_551 | _T_564; // @[dec_dec_ctl.scala 50:17]
  assign io_out_condbr = _T_317 & _T_18; // @[dec_dec_ctl.scala 53:17]
  assign io_out_beq = _T_584 & _T_18; // @[dec_dec_ctl.scala 54:14]
  assign io_out_bne = _T_596 & _T_18; // @[dec_dec_ctl.scala 55:14]
  assign io_out_bge = _T_607 & _T_18; // @[dec_dec_ctl.scala 56:14]
  assign io_out_blt = _T_619 & _T_18; // @[dec_dec_ctl.scala 57:14]
  assign io_out_jal = io_ins[6] & io_ins[2]; // @[dec_dec_ctl.scala 58:14]
  assign io_out_by = _T_636 & _T_18; // @[dec_dec_ctl.scala 59:13]
  assign io_out_half = _T_646 & _T_18; // @[dec_dec_ctl.scala 60:15]
  assign io_out_word = _T_653 & _T_97; // @[dec_dec_ctl.scala 61:15]
  assign io_out_csr_read = _T_683 | _T_688; // @[dec_dec_ctl.scala 62:19]
  assign io_out_csr_clr = _T_728 | _T_737; // @[dec_dec_ctl.scala 65:18]
  assign io_out_csr_set = _T_829 | _T_837; // @[dec_dec_ctl.scala 72:18]
  assign io_out_csr_write = _T_745 & io_ins[4]; // @[dec_dec_ctl.scala 68:20]
  assign io_out_csr_imm = _T_786 | _T_793; // @[dec_dec_ctl.scala 69:18]
  assign io_out_presync = _T_1106 | _T_1113; // @[dec_dec_ctl.scala 89:18]
  assign io_out_postsync = _T_1210 | _T_1113; // @[dec_dec_ctl.scala 95:19]
  assign io_out_ebreak = _T_851 & io_ins[4]; // @[dec_dec_ctl.scala 75:17]
  assign io_out_ecall = _T_866 & io_ins[4]; // @[dec_dec_ctl.scala 76:16]
  assign io_out_mret = _T_877 & io_ins[4]; // @[dec_dec_ctl.scala 77:15]
  assign io_out_mul = _T_891 & _T_18; // @[dec_dec_ctl.scala 78:14]
  assign io_out_rs1_sign = _T_911 | _T_928; // @[dec_dec_ctl.scala 79:19]
  assign io_out_rs2_sign = _T_927 & _T_18; // @[dec_dec_ctl.scala 81:19]
  assign io_out_low = _T_962 & _T_18; // @[dec_dec_ctl.scala 82:14]
  assign io_out_div = _T_973 & _T_18; // @[dec_dec_ctl.scala 83:14]
  assign io_out_rem = _T_986 & _T_18; // @[dec_dec_ctl.scala 84:14]
  assign io_out_fence = _T_9 & io_ins[3]; // @[dec_dec_ctl.scala 85:16]
  assign io_out_fence_i = _T_996 & io_ins[3]; // @[dec_dec_ctl.scala 86:18]
  assign io_out_pm_alu = _T_1020 | _T_11; // @[dec_dec_ctl.scala 87:17]
  assign io_out_legal = _T_1953 | _T_1966; // @[dec_dec_ctl.scala 101:16]
endmodule
module dec_decode_ctl(
  input         clock,
  input         reset,
  output [1:0]  io_decode_exu_dec_data_en,
  output [1:0]  io_decode_exu_dec_ctl_en,
  output        io_decode_exu_i0_ap_land,
  output        io_decode_exu_i0_ap_lor,
  output        io_decode_exu_i0_ap_lxor,
  output        io_decode_exu_i0_ap_sll,
  output        io_decode_exu_i0_ap_srl,
  output        io_decode_exu_i0_ap_sra,
  output        io_decode_exu_i0_ap_beq,
  output        io_decode_exu_i0_ap_bne,
  output        io_decode_exu_i0_ap_blt,
  output        io_decode_exu_i0_ap_bge,
  output        io_decode_exu_i0_ap_add,
  output        io_decode_exu_i0_ap_sub,
  output        io_decode_exu_i0_ap_slt,
  output        io_decode_exu_i0_ap_unsign,
  output        io_decode_exu_i0_ap_jal,
  output        io_decode_exu_i0_ap_predict_t,
  output        io_decode_exu_i0_ap_predict_nt,
  output        io_decode_exu_i0_ap_csr_write,
  output        io_decode_exu_i0_ap_csr_imm,
  output        io_decode_exu_dec_i0_predict_p_d_valid,
  output        io_decode_exu_dec_i0_predict_p_d_bits_pc4,
  output [1:0]  io_decode_exu_dec_i0_predict_p_d_bits_hist,
  output [11:0] io_decode_exu_dec_i0_predict_p_d_bits_toffset,
  output        io_decode_exu_dec_i0_predict_p_d_bits_br_error,
  output        io_decode_exu_dec_i0_predict_p_d_bits_br_start_error,
  output [30:0] io_decode_exu_dec_i0_predict_p_d_bits_prett,
  output        io_decode_exu_dec_i0_predict_p_d_bits_pcall,
  output        io_decode_exu_dec_i0_predict_p_d_bits_pret,
  output        io_decode_exu_dec_i0_predict_p_d_bits_pja,
  output        io_decode_exu_dec_i0_predict_p_d_bits_way,
  output [7:0]  io_decode_exu_i0_predict_fghr_d,
  output [7:0]  io_decode_exu_i0_predict_index_d,
  output [4:0]  io_decode_exu_i0_predict_btag_d,
  output        io_decode_exu_dec_i0_rs1_en_d,
  output        io_decode_exu_dec_i0_rs2_en_d,
  output [31:0] io_decode_exu_dec_i0_immed_d,
  output [31:0] io_decode_exu_dec_i0_rs1_bypass_data_d,
  output [31:0] io_decode_exu_dec_i0_rs2_bypass_data_d,
  output        io_decode_exu_dec_i0_select_pc_d,
  output [1:0]  io_decode_exu_dec_i0_rs1_bypass_en_d,
  output [1:0]  io_decode_exu_dec_i0_rs2_bypass_en_d,
  output        io_decode_exu_mul_p_valid,
  output        io_decode_exu_mul_p_bits_rs1_sign,
  output        io_decode_exu_mul_p_bits_rs2_sign,
  output        io_decode_exu_mul_p_bits_low,
  output [30:0] io_decode_exu_pred_correct_npc_x,
  output        io_decode_exu_dec_extint_stall,
  input  [31:0] io_decode_exu_exu_i0_result_x,
  input  [31:0] io_decode_exu_exu_csr_rs1_x,
  output        io_dec_alu_dec_i0_alu_decode_d,
  output        io_dec_alu_dec_csr_ren_d,
  output [11:0] io_dec_alu_dec_i0_br_immed_d,
  input  [30:0] io_dec_alu_exu_i0_pc_x,
  output        io_dec_div_div_p_valid,
  output        io_dec_div_div_p_bits_unsign,
  output        io_dec_div_div_p_bits_rem,
  output        io_dec_div_dec_div_cancel,
  input         io_dctl_busbuff_lsu_nonblock_load_valid_m,
  input  [1:0]  io_dctl_busbuff_lsu_nonblock_load_tag_m,
  input         io_dctl_busbuff_lsu_nonblock_load_inv_r,
  input  [1:0]  io_dctl_busbuff_lsu_nonblock_load_inv_tag_r,
  input         io_dctl_busbuff_lsu_nonblock_load_data_valid,
  input         io_dctl_busbuff_lsu_nonblock_load_data_error,
  input  [1:0]  io_dctl_busbuff_lsu_nonblock_load_data_tag,
  input  [31:0] io_dctl_busbuff_lsu_nonblock_load_data,
  input         io_dctl_dma_dma_dccm_stall_any,
  output        io_dec_aln_dec_i0_decode_d,
  input  [15:0] io_dec_aln_ifu_i0_cinst,
  input  [31:0] io_dbg_dctl_dbg_cmd_wrdata,
  input         io_dec_tlu_flush_extint,
  input         io_dec_tlu_force_halt,
  output [31:0] io_dec_i0_inst_wb1,
  output [30:0] io_dec_i0_pc_wb1,
  input  [3:0]  io_dec_i0_trigger_match_d,
  input         io_dec_tlu_wr_pause_r,
  input         io_dec_tlu_pipelining_disable,
  input  [3:0]  io_lsu_trigger_match_m,
  input         io_lsu_pmu_misaligned_m,
  input         io_dec_tlu_debug_stall,
  input         io_dec_tlu_flush_leak_one_r,
  input         io_dec_debug_fence_d,
  input         io_dec_i0_icaf_d,
  input         io_dec_i0_icaf_f1_d,
  input  [1:0]  io_dec_i0_icaf_type_d,
  input         io_dec_i0_dbecc_d,
  input         io_dec_i0_brp_valid,
  input  [11:0] io_dec_i0_brp_bits_toffset,
  input  [1:0]  io_dec_i0_brp_bits_hist,
  input         io_dec_i0_brp_bits_br_error,
  input         io_dec_i0_brp_bits_br_start_error,
  input  [30:0] io_dec_i0_brp_bits_prett,
  input         io_dec_i0_brp_bits_way,
  input         io_dec_i0_brp_bits_ret,
  input  [7:0]  io_dec_i0_bp_index,
  input  [7:0]  io_dec_i0_bp_fghr,
  input  [4:0]  io_dec_i0_bp_btag,
  input         io_lsu_idle_any,
  input         io_lsu_load_stall_any,
  input         io_lsu_store_stall_any,
  input         io_exu_div_wren,
  input         io_dec_tlu_i0_kill_writeb_wb,
  input         io_dec_tlu_flush_lower_wb,
  input         io_dec_tlu_i0_kill_writeb_r,
  input         io_dec_tlu_flush_lower_r,
  input         io_dec_tlu_flush_pause_r,
  input         io_dec_tlu_presync_d,
  input         io_dec_tlu_postsync_d,
  input         io_dec_i0_pc4_d,
  input  [31:0] io_dec_csr_rddata_d,
  input         io_dec_csr_legal_d,
  input  [31:0] io_lsu_result_m,
  input  [31:0] io_lsu_result_corr_r,
  input         io_exu_flush_final,
  input  [31:0] io_dec_i0_instr_d,
  input         io_dec_ib0_valid_d,
  input         io_free_clk,
  input         io_active_clk,
  input         io_clk_override,
  output [4:0]  io_dec_i0_rs1_d,
  output [4:0]  io_dec_i0_rs2_d,
  output [4:0]  io_dec_i0_waddr_r,
  output        io_dec_i0_wen_r,
  output [31:0] io_dec_i0_wdata_r,
  output        io_lsu_p_valid,
  output        io_lsu_p_bits_fast_int,
  output        io_lsu_p_bits_by,
  output        io_lsu_p_bits_half,
  output        io_lsu_p_bits_word,
  output        io_lsu_p_bits_load,
  output        io_lsu_p_bits_store,
  output        io_lsu_p_bits_unsign,
  output        io_lsu_p_bits_store_data_bypass_d,
  output        io_lsu_p_bits_load_ldst_bypass_d,
  output [4:0]  io_div_waddr_wb,
  output        io_dec_lsu_valid_raw_d,
  output [11:0] io_dec_lsu_offset_d,
  output        io_dec_csr_wen_unq_d,
  output        io_dec_csr_any_unq_d,
  output [11:0] io_dec_csr_rdaddr_d,
  output        io_dec_csr_wen_r,
  output [11:0] io_dec_csr_wraddr_r,
  output [31:0] io_dec_csr_wrdata_r,
  output        io_dec_csr_stall_int_ff,
  output        io_dec_tlu_i0_valid_r,
  output        io_dec_tlu_packet_r_legal,
  output        io_dec_tlu_packet_r_icaf,
  output        io_dec_tlu_packet_r_icaf_f1,
  output [1:0]  io_dec_tlu_packet_r_icaf_type,
  output        io_dec_tlu_packet_r_fence_i,
  output [3:0]  io_dec_tlu_packet_r_i0trigger,
  output [3:0]  io_dec_tlu_packet_r_pmu_i0_itype,
  output        io_dec_tlu_packet_r_pmu_i0_br_unpred,
  output        io_dec_tlu_packet_r_pmu_divide,
  output        io_dec_tlu_packet_r_pmu_lsu_misaligned,
  output [30:0] io_dec_tlu_i0_pc_r,
  output [31:0] io_dec_illegal_inst,
  output        io_dec_pmu_instr_decoded,
  output        io_dec_pmu_decode_stall,
  output        io_dec_pmu_presync_stall,
  output        io_dec_pmu_postsync_stall,
  output        io_dec_nonblock_load_wen,
  output [4:0]  io_dec_nonblock_load_waddr,
  output        io_dec_pause_state,
  output        io_dec_pause_state_cg,
  output        io_dec_div_active,
  input         io_scan_mode
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
`endif // RANDOMIZE_REG_INIT
  wire  rvclkhdr_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_io_scan_mode; // @[lib.scala 343:22]
  wire [31:0] i0_dec_io_ins; // @[dec_decode_ctl.scala 356:22]
  wire  i0_dec_io_out_alu; // @[dec_decode_ctl.scala 356:22]
  wire  i0_dec_io_out_rs1; // @[dec_decode_ctl.scala 356:22]
  wire  i0_dec_io_out_rs2; // @[dec_decode_ctl.scala 356:22]
  wire  i0_dec_io_out_imm12; // @[dec_decode_ctl.scala 356:22]
  wire  i0_dec_io_out_rd; // @[dec_decode_ctl.scala 356:22]
  wire  i0_dec_io_out_shimm5; // @[dec_decode_ctl.scala 356:22]
  wire  i0_dec_io_out_imm20; // @[dec_decode_ctl.scala 356:22]
  wire  i0_dec_io_out_pc; // @[dec_decode_ctl.scala 356:22]
  wire  i0_dec_io_out_load; // @[dec_decode_ctl.scala 356:22]
  wire  i0_dec_io_out_store; // @[dec_decode_ctl.scala 356:22]
  wire  i0_dec_io_out_lsu; // @[dec_decode_ctl.scala 356:22]
  wire  i0_dec_io_out_add; // @[dec_decode_ctl.scala 356:22]
  wire  i0_dec_io_out_sub; // @[dec_decode_ctl.scala 356:22]
  wire  i0_dec_io_out_land; // @[dec_decode_ctl.scala 356:22]
  wire  i0_dec_io_out_lor; // @[dec_decode_ctl.scala 356:22]
  wire  i0_dec_io_out_lxor; // @[dec_decode_ctl.scala 356:22]
  wire  i0_dec_io_out_sll; // @[dec_decode_ctl.scala 356:22]
  wire  i0_dec_io_out_sra; // @[dec_decode_ctl.scala 356:22]
  wire  i0_dec_io_out_srl; // @[dec_decode_ctl.scala 356:22]
  wire  i0_dec_io_out_slt; // @[dec_decode_ctl.scala 356:22]
  wire  i0_dec_io_out_unsign; // @[dec_decode_ctl.scala 356:22]
  wire  i0_dec_io_out_condbr; // @[dec_decode_ctl.scala 356:22]
  wire  i0_dec_io_out_beq; // @[dec_decode_ctl.scala 356:22]
  wire  i0_dec_io_out_bne; // @[dec_decode_ctl.scala 356:22]
  wire  i0_dec_io_out_bge; // @[dec_decode_ctl.scala 356:22]
  wire  i0_dec_io_out_blt; // @[dec_decode_ctl.scala 356:22]
  wire  i0_dec_io_out_jal; // @[dec_decode_ctl.scala 356:22]
  wire  i0_dec_io_out_by; // @[dec_decode_ctl.scala 356:22]
  wire  i0_dec_io_out_half; // @[dec_decode_ctl.scala 356:22]
  wire  i0_dec_io_out_word; // @[dec_decode_ctl.scala 356:22]
  wire  i0_dec_io_out_csr_read; // @[dec_decode_ctl.scala 356:22]
  wire  i0_dec_io_out_csr_clr; // @[dec_decode_ctl.scala 356:22]
  wire  i0_dec_io_out_csr_set; // @[dec_decode_ctl.scala 356:22]
  wire  i0_dec_io_out_csr_write; // @[dec_decode_ctl.scala 356:22]
  wire  i0_dec_io_out_csr_imm; // @[dec_decode_ctl.scala 356:22]
  wire  i0_dec_io_out_presync; // @[dec_decode_ctl.scala 356:22]
  wire  i0_dec_io_out_postsync; // @[dec_decode_ctl.scala 356:22]
  wire  i0_dec_io_out_ebreak; // @[dec_decode_ctl.scala 356:22]
  wire  i0_dec_io_out_ecall; // @[dec_decode_ctl.scala 356:22]
  wire  i0_dec_io_out_mret; // @[dec_decode_ctl.scala 356:22]
  wire  i0_dec_io_out_mul; // @[dec_decode_ctl.scala 356:22]
  wire  i0_dec_io_out_rs1_sign; // @[dec_decode_ctl.scala 356:22]
  wire  i0_dec_io_out_rs2_sign; // @[dec_decode_ctl.scala 356:22]
  wire  i0_dec_io_out_low; // @[dec_decode_ctl.scala 356:22]
  wire  i0_dec_io_out_div; // @[dec_decode_ctl.scala 356:22]
  wire  i0_dec_io_out_rem; // @[dec_decode_ctl.scala 356:22]
  wire  i0_dec_io_out_fence; // @[dec_decode_ctl.scala 356:22]
  wire  i0_dec_io_out_fence_i; // @[dec_decode_ctl.scala 356:22]
  wire  i0_dec_io_out_pm_alu; // @[dec_decode_ctl.scala 356:22]
  wire  i0_dec_io_out_legal; // @[dec_decode_ctl.scala 356:22]
  wire  rvclkhdr_1_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_1_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_1_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_1_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_2_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_2_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_2_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_2_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_3_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_3_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_3_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_3_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_4_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_4_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_4_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_4_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_5_io_l1clk; // @[lib.scala 378:23]
  wire  rvclkhdr_5_io_clk; // @[lib.scala 378:23]
  wire  rvclkhdr_5_io_en; // @[lib.scala 378:23]
  wire  rvclkhdr_5_io_scan_mode; // @[lib.scala 378:23]
  wire  rvclkhdr_6_io_l1clk; // @[lib.scala 378:23]
  wire  rvclkhdr_6_io_clk; // @[lib.scala 378:23]
  wire  rvclkhdr_6_io_en; // @[lib.scala 378:23]
  wire  rvclkhdr_6_io_scan_mode; // @[lib.scala 378:23]
  wire  rvclkhdr_7_io_l1clk; // @[lib.scala 378:23]
  wire  rvclkhdr_7_io_clk; // @[lib.scala 378:23]
  wire  rvclkhdr_7_io_en; // @[lib.scala 378:23]
  wire  rvclkhdr_7_io_scan_mode; // @[lib.scala 378:23]
  wire  rvclkhdr_8_io_l1clk; // @[lib.scala 378:23]
  wire  rvclkhdr_8_io_clk; // @[lib.scala 378:23]
  wire  rvclkhdr_8_io_en; // @[lib.scala 378:23]
  wire  rvclkhdr_8_io_scan_mode; // @[lib.scala 378:23]
  wire  rvclkhdr_9_io_l1clk; // @[lib.scala 378:23]
  wire  rvclkhdr_9_io_clk; // @[lib.scala 378:23]
  wire  rvclkhdr_9_io_en; // @[lib.scala 378:23]
  wire  rvclkhdr_9_io_scan_mode; // @[lib.scala 378:23]
  wire  rvclkhdr_10_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_10_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_10_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_10_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_11_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_11_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_11_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_11_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_12_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_12_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_12_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_12_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_13_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_13_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_13_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_13_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_14_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_14_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_14_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_14_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_15_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_15_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_15_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_15_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_16_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_16_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_16_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_16_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_17_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_17_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_17_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_17_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_18_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_18_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_18_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_18_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_19_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_19_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_19_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_19_io_scan_mode; // @[lib.scala 368:23]
  reg  tlu_wr_pause_r1; // @[dec_decode_ctl.scala 463:55]
  wire  _T_1 = io_dec_tlu_wr_pause_r ^ tlu_wr_pause_r1; // @[dec_decode_ctl.scala 178:54]
  reg  tlu_wr_pause_r2; // @[dec_decode_ctl.scala 464:55]
  wire  _T_2 = tlu_wr_pause_r1 ^ tlu_wr_pause_r2; // @[dec_decode_ctl.scala 179:54]
  wire  _T_3 = _T_1 | _T_2; // @[dec_decode_ctl.scala 178:89]
  wire  _T_4 = io_dec_tlu_flush_extint ^ io_decode_exu_dec_extint_stall; // @[dec_decode_ctl.scala 180:54]
  wire  _T_5 = _T_3 | _T_4; // @[dec_decode_ctl.scala 179:89]
  reg  leak1_i1_stall; // @[dec_decode_ctl.scala 364:56]
  wire  _T_280 = ~io_dec_tlu_flush_lower_r; // @[dec_decode_ctl.scala 363:73]
  wire  _T_281 = leak1_i1_stall & _T_280; // @[dec_decode_ctl.scala 363:71]
  wire  leak1_i1_stall_in = io_dec_tlu_flush_leak_one_r | _T_281; // @[dec_decode_ctl.scala 363:53]
  wire  _T_6 = leak1_i1_stall_in ^ leak1_i1_stall; // @[dec_decode_ctl.scala 181:54]
  wire  _T_7 = _T_5 | _T_6; // @[dec_decode_ctl.scala 180:89]
  wire  _T_284 = io_dec_aln_dec_i0_decode_d & leak1_i1_stall; // @[dec_decode_ctl.scala 366:53]
  reg  leak1_i0_stall; // @[dec_decode_ctl.scala 367:56]
  wire  _T_286 = leak1_i0_stall & _T_280; // @[dec_decode_ctl.scala 366:89]
  wire  leak1_i0_stall_in = _T_284 | _T_286; // @[dec_decode_ctl.scala 366:71]
  wire  _T_8 = leak1_i0_stall_in ^ leak1_i0_stall; // @[dec_decode_ctl.scala 182:54]
  wire  _T_9 = _T_7 | _T_8; // @[dec_decode_ctl.scala 181:89]
  reg  pause_stall; // @[dec_decode_ctl.scala 461:50]
  wire  _T_415 = io_dec_tlu_wr_pause_r | pause_stall; // @[dec_decode_ctl.scala 460:44]
  wire  _T_408 = ~io_dec_tlu_flush_pause_r; // @[dec_decode_ctl.scala 459:49]
  wire  _T_409 = io_dec_tlu_flush_lower_r & _T_408; // @[dec_decode_ctl.scala 459:47]
  reg [31:0] write_csr_data; // @[lib.scala 374:16]
  wire [31:0] _T_412 = {31'h0,write_csr_data[0]}; // @[Cat.scala 29:58]
  wire  _T_413 = write_csr_data == _T_412; // @[dec_decode_ctl.scala 459:109]
  wire  _T_414 = pause_stall & _T_413; // @[dec_decode_ctl.scala 459:91]
  wire  clear_pause = _T_409 | _T_414; // @[dec_decode_ctl.scala 459:76]
  wire  _T_416 = ~clear_pause; // @[dec_decode_ctl.scala 460:61]
  wire  pause_state_in = _T_415 & _T_416; // @[dec_decode_ctl.scala 460:59]
  wire  _T_10 = pause_state_in ^ pause_stall; // @[dec_decode_ctl.scala 183:54]
  wire  _T_11 = _T_9 | _T_10; // @[dec_decode_ctl.scala 182:89]
  wire  _T_18 = ~leak1_i1_stall; // @[dec_decode_ctl.scala 192:80]
  wire  i0_brp_valid = io_dec_i0_brp_valid & _T_18; // @[dec_decode_ctl.scala 192:78]
  wire  i0_dp_raw_condbr = i0_dec_io_out_condbr; // @[dec_decode_ctl.scala 124:37 dec_decode_ctl.scala 358:12]
  wire  i0_dp_raw_jal = i0_dec_io_out_jal; // @[dec_decode_ctl.scala 124:37 dec_decode_ctl.scala 358:12]
  wire [19:0] i0_pcall_imm = {io_dec_i0_instr_d[31],io_dec_i0_instr_d[19:12],io_dec_i0_instr_d[20],io_dec_i0_instr_d[30:21]}; // @[Cat.scala 29:58]
  wire  _T_298 = i0_pcall_imm[19:12] == 8'hff; // @[dec_decode_ctl.scala 372:79]
  wire  _T_300 = i0_pcall_imm[19:12] == 8'h0; // @[dec_decode_ctl.scala 372:112]
  wire  i0_pcall_12b_offset = i0_pcall_imm[11] ? _T_298 : _T_300; // @[dec_decode_ctl.scala 372:33]
  wire  i0_dp_raw_imm20 = i0_dec_io_out_imm20; // @[dec_decode_ctl.scala 124:37 dec_decode_ctl.scala 358:12]
  wire  _T_301 = i0_pcall_12b_offset & i0_dp_raw_imm20; // @[dec_decode_ctl.scala 373:47]
  wire [4:0] i0r_rd = io_dec_i0_instr_d[11:7]; // @[dec_decode_ctl.scala 586:16]
  wire  _T_302 = i0r_rd == 5'h1; // @[dec_decode_ctl.scala 373:76]
  wire  _T_303 = i0r_rd == 5'h5; // @[dec_decode_ctl.scala 373:98]
  wire  _T_304 = _T_302 | _T_303; // @[dec_decode_ctl.scala 373:89]
  wire  i0_pcall_case = _T_301 & _T_304; // @[dec_decode_ctl.scala 373:65]
  wire  i0_pcall_raw = i0_dp_raw_jal & i0_pcall_case; // @[dec_decode_ctl.scala 375:38]
  wire  _T_20 = i0_dp_raw_condbr | i0_pcall_raw; // @[dec_decode_ctl.scala 203:92]
  wire  _T_309 = ~_T_304; // @[dec_decode_ctl.scala 374:67]
  wire  i0_pja_case = _T_301 & _T_309; // @[dec_decode_ctl.scala 374:65]
  wire  i0_pja_raw = i0_dp_raw_jal & i0_pja_case; // @[dec_decode_ctl.scala 377:38]
  wire  _T_21 = _T_20 | i0_pja_raw; // @[dec_decode_ctl.scala 203:107]
  wire  i0_dp_raw_imm12 = i0_dec_io_out_imm12; // @[dec_decode_ctl.scala 124:37 dec_decode_ctl.scala 358:12]
  wire  _T_325 = i0_dp_raw_jal & i0_dp_raw_imm12; // @[dec_decode_ctl.scala 381:37]
  wire  _T_326 = i0r_rd == 5'h0; // @[dec_decode_ctl.scala 381:65]
  wire  _T_327 = _T_325 & _T_326; // @[dec_decode_ctl.scala 381:55]
  wire [4:0] i0r_rs1 = io_dec_i0_instr_d[19:15]; // @[dec_decode_ctl.scala 584:16]
  wire  _T_328 = i0r_rs1 == 5'h1; // @[dec_decode_ctl.scala 381:89]
  wire  _T_329 = i0r_rs1 == 5'h5; // @[dec_decode_ctl.scala 381:111]
  wire  _T_330 = _T_328 | _T_329; // @[dec_decode_ctl.scala 381:101]
  wire  i0_pret_case = _T_327 & _T_330; // @[dec_decode_ctl.scala 381:79]
  wire  i0_pret_raw = i0_dp_raw_jal & i0_pret_case; // @[dec_decode_ctl.scala 382:32]
  wire  _T_22 = _T_21 | i0_pret_raw; // @[dec_decode_ctl.scala 203:120]
  wire  _T_23 = ~_T_22; // @[dec_decode_ctl.scala 203:73]
  wire  i0_notbr_error = i0_brp_valid & _T_23; // @[dec_decode_ctl.scala 203:71]
  wire  _T_31 = io_dec_i0_brp_bits_br_error | i0_notbr_error; // @[dec_decode_ctl.scala 208:87]
  wire  _T_25 = i0_brp_valid & io_dec_i0_brp_bits_hist[1]; // @[dec_decode_ctl.scala 206:72]
  wire  _T_314 = i0_pcall_raw | i0_pja_raw; // @[dec_decode_ctl.scala 379:41]
  wire [11:0] _T_323 = {io_dec_i0_instr_d[31],io_dec_i0_instr_d[7],io_dec_i0_instr_d[30:25],io_dec_i0_instr_d[11:8]}; // @[Cat.scala 29:58]
  wire [11:0] i0_br_offset = _T_314 ? i0_pcall_imm[11:0] : _T_323; // @[dec_decode_ctl.scala 379:26]
  wire  _T_26 = io_dec_i0_brp_bits_toffset != i0_br_offset; // @[dec_decode_ctl.scala 206:131]
  wire  _T_27 = _T_25 & _T_26; // @[dec_decode_ctl.scala 206:101]
  wire  _T_28 = ~i0_pret_raw; // @[dec_decode_ctl.scala 206:151]
  wire  i0_br_toffset_error = _T_27 & _T_28; // @[dec_decode_ctl.scala 206:149]
  wire  _T_32 = _T_31 | i0_br_toffset_error; // @[dec_decode_ctl.scala 208:104]
  wire  _T_29 = i0_brp_valid & io_dec_i0_brp_bits_ret; // @[dec_decode_ctl.scala 207:72]
  wire  i0_ret_error = _T_29 & _T_28; // @[dec_decode_ctl.scala 207:97]
  wire  i0_br_error = _T_32 | i0_ret_error; // @[dec_decode_ctl.scala 208:126]
  wire  _T_39 = i0_br_error | io_dec_i0_brp_bits_br_start_error; // @[dec_decode_ctl.scala 213:72]
  wire  i0_br_error_all = _T_39 & _T_18; // @[dec_decode_ctl.scala 213:109]
  wire  i0_icaf_d = io_dec_i0_icaf_d | io_dec_i0_dbecc_d; // @[dec_decode_ctl.scala 222:43]
  wire  _T_41 = i0_br_error_all | i0_icaf_d; // @[dec_decode_ctl.scala 225:25]
  wire  i0_dp_raw_postsync = i0_dec_io_out_postsync; // @[dec_decode_ctl.scala 124:37 dec_decode_ctl.scala 358:12]
  wire  i0_dp_postsync = _T_41 | i0_dp_raw_postsync; // @[dec_decode_ctl.scala 225:50]
  wire  _T_442 = i0_dp_postsync | io_dec_tlu_postsync_d; // @[dec_decode_ctl.scala 490:36]
  wire  debug_fence_i = io_dec_debug_fence_d & io_dbg_dctl_dbg_cmd_wrdata[0]; // @[dec_decode_ctl.scala 482:48]
  wire  _T_443 = _T_442 | debug_fence_i; // @[dec_decode_ctl.scala 490:60]
  wire  i0_dp_raw_csr_write = i0_dec_io_out_csr_write; // @[dec_decode_ctl.scala 124:37 dec_decode_ctl.scala 358:12]
  wire  i0_dp_csr_write = _T_41 ? 1'h0 : i0_dp_raw_csr_write; // @[dec_decode_ctl.scala 225:50]
  wire  _T_343 = ~io_dec_debug_fence_d; // @[dec_decode_ctl.scala 421:42]
  wire  i0_csr_write = i0_dp_csr_write & _T_343; // @[dec_decode_ctl.scala 421:40]
  wire  i0_dp_raw_csr_read = i0_dec_io_out_csr_read; // @[dec_decode_ctl.scala 124:37 dec_decode_ctl.scala 358:12]
  wire  i0_dp_csr_read = _T_41 ? 1'h0 : i0_dp_raw_csr_read; // @[dec_decode_ctl.scala 225:50]
  wire  _T_347 = ~i0_dp_csr_read; // @[dec_decode_ctl.scala 426:41]
  wire  i0_csr_write_only_d = i0_csr_write & _T_347; // @[dec_decode_ctl.scala 426:39]
  wire  _T_445 = io_dec_i0_instr_d[31:20] == 12'h7c2; // @[dec_decode_ctl.scala 490:112]
  wire  _T_446 = i0_csr_write_only_d & _T_445; // @[dec_decode_ctl.scala 490:99]
  wire  i0_postsync = _T_443 | _T_446; // @[dec_decode_ctl.scala 490:76]
  wire  i0_dp_raw_legal = i0_dec_io_out_legal; // @[dec_decode_ctl.scala 124:37 dec_decode_ctl.scala 358:12]
  wire  i0_dp_legal = _T_41 | i0_dp_raw_legal; // @[dec_decode_ctl.scala 225:50]
  wire  any_csr_d = i0_dp_csr_read | i0_csr_write; // @[dec_decode_ctl.scala 492:34]
  wire  _T_447 = ~any_csr_d; // @[dec_decode_ctl.scala 494:40]
  wire  _T_448 = _T_447 | io_dec_csr_legal_d; // @[dec_decode_ctl.scala 494:51]
  wire  i0_legal = i0_dp_legal & _T_448; // @[dec_decode_ctl.scala 494:37]
  wire  _T_507 = ~i0_legal; // @[dec_decode_ctl.scala 534:64]
  wire  _T_508 = i0_postsync | _T_507; // @[dec_decode_ctl.scala 534:62]
  wire  _T_509 = io_dec_aln_dec_i0_decode_d & _T_508; // @[dec_decode_ctl.scala 534:47]
  reg  postsync_stall; // @[dec_decode_ctl.scala 532:53]
  reg  x_d_valid; // @[lib.scala 384:16]
  wire  _T_510 = postsync_stall & x_d_valid; // @[dec_decode_ctl.scala 534:96]
  wire  ps_stall_in = _T_509 | _T_510; // @[dec_decode_ctl.scala 534:77]
  wire  _T_12 = ps_stall_in ^ postsync_stall; // @[dec_decode_ctl.scala 184:54]
  wire  _T_13 = _T_11 | _T_12; // @[dec_decode_ctl.scala 183:89]
  reg  flush_final_r; // @[dec_decode_ctl.scala 580:52]
  wire  _T_14 = io_exu_flush_final ^ flush_final_r; // @[dec_decode_ctl.scala 185:54]
  wire  _T_15 = _T_13 | _T_14; // @[dec_decode_ctl.scala 184:89]
  wire  shift_illegal = io_dec_aln_dec_i0_decode_d & _T_507; // @[dec_decode_ctl.scala 498:55]
  reg  illegal_lockout; // @[dec_decode_ctl.scala 502:54]
  wire  _T_469 = shift_illegal | illegal_lockout; // @[dec_decode_ctl.scala 501:40]
  wire  _T_470 = ~flush_final_r; // @[dec_decode_ctl.scala 501:61]
  wire  illegal_lockout_in = _T_469 & _T_470; // @[dec_decode_ctl.scala 501:59]
  wire  _T_16 = illegal_lockout_in ^ illegal_lockout; // @[dec_decode_ctl.scala 186:54]
  wire  i0_legal_decode_d = io_dec_aln_dec_i0_decode_d & i0_legal; // @[dec_decode_ctl.scala 608:54]
  wire  _T_33 = i0_br_error & i0_legal_decode_d; // @[dec_decode_ctl.scala 209:72]
  wire  _T_36 = io_dec_i0_brp_bits_br_start_error & i0_legal_decode_d; // @[dec_decode_ctl.scala 210:94]
  wire  i0_dp_raw_pm_alu = i0_dec_io_out_pm_alu; // @[dec_decode_ctl.scala 124:37 dec_decode_ctl.scala 358:12]
  wire  i0_dp_pm_alu = _T_41 ? 1'h0 : i0_dp_raw_pm_alu; // @[dec_decode_ctl.scala 225:50]
  wire  i0_dp_raw_fence_i = i0_dec_io_out_fence_i; // @[dec_decode_ctl.scala 124:37 dec_decode_ctl.scala 358:12]
  wire  i0_dp_fence_i = _T_41 ? 1'h0 : i0_dp_raw_fence_i; // @[dec_decode_ctl.scala 225:50]
  wire  i0_dp_raw_fence = i0_dec_io_out_fence; // @[dec_decode_ctl.scala 124:37 dec_decode_ctl.scala 358:12]
  wire  i0_dp_fence = _T_41 ? 1'h0 : i0_dp_raw_fence; // @[dec_decode_ctl.scala 225:50]
  wire  i0_dp_raw_rem = i0_dec_io_out_rem; // @[dec_decode_ctl.scala 124:37 dec_decode_ctl.scala 358:12]
  wire  i0_dp_raw_div = i0_dec_io_out_div; // @[dec_decode_ctl.scala 124:37 dec_decode_ctl.scala 358:12]
  wire  i0_dp_div = _T_41 ? 1'h0 : i0_dp_raw_div; // @[dec_decode_ctl.scala 225:50]
  wire  i0_dp_raw_low = i0_dec_io_out_low; // @[dec_decode_ctl.scala 124:37 dec_decode_ctl.scala 358:12]
  wire  i0_dp_raw_rs2_sign = i0_dec_io_out_rs2_sign; // @[dec_decode_ctl.scala 124:37 dec_decode_ctl.scala 358:12]
  wire  i0_dp_raw_rs1_sign = i0_dec_io_out_rs1_sign; // @[dec_decode_ctl.scala 124:37 dec_decode_ctl.scala 358:12]
  wire  i0_dp_raw_mul = i0_dec_io_out_mul; // @[dec_decode_ctl.scala 124:37 dec_decode_ctl.scala 358:12]
  wire  i0_dp_mul = _T_41 ? 1'h0 : i0_dp_raw_mul; // @[dec_decode_ctl.scala 225:50]
  wire  i0_dp_raw_mret = i0_dec_io_out_mret; // @[dec_decode_ctl.scala 124:37 dec_decode_ctl.scala 358:12]
  wire  i0_dp_mret = _T_41 ? 1'h0 : i0_dp_raw_mret; // @[dec_decode_ctl.scala 225:50]
  wire  i0_dp_raw_ecall = i0_dec_io_out_ecall; // @[dec_decode_ctl.scala 124:37 dec_decode_ctl.scala 358:12]
  wire  i0_dp_ecall = _T_41 ? 1'h0 : i0_dp_raw_ecall; // @[dec_decode_ctl.scala 225:50]
  wire  i0_dp_raw_ebreak = i0_dec_io_out_ebreak; // @[dec_decode_ctl.scala 124:37 dec_decode_ctl.scala 358:12]
  wire  i0_dp_ebreak = _T_41 ? 1'h0 : i0_dp_raw_ebreak; // @[dec_decode_ctl.scala 225:50]
  wire  i0_dp_raw_presync = i0_dec_io_out_presync; // @[dec_decode_ctl.scala 124:37 dec_decode_ctl.scala 358:12]
  wire  i0_dp_presync = _T_41 ? 1'h0 : i0_dp_raw_presync; // @[dec_decode_ctl.scala 225:50]
  wire  i0_dp_raw_csr_imm = i0_dec_io_out_csr_imm; // @[dec_decode_ctl.scala 124:37 dec_decode_ctl.scala 358:12]
  wire  i0_dp_csr_imm = _T_41 ? 1'h0 : i0_dp_raw_csr_imm; // @[dec_decode_ctl.scala 225:50]
  wire  i0_dp_raw_csr_set = i0_dec_io_out_csr_set; // @[dec_decode_ctl.scala 124:37 dec_decode_ctl.scala 358:12]
  wire  i0_dp_csr_set = _T_41 ? 1'h0 : i0_dp_raw_csr_set; // @[dec_decode_ctl.scala 225:50]
  wire  i0_dp_raw_csr_clr = i0_dec_io_out_csr_clr; // @[dec_decode_ctl.scala 124:37 dec_decode_ctl.scala 358:12]
  wire  i0_dp_csr_clr = _T_41 ? 1'h0 : i0_dp_raw_csr_clr; // @[dec_decode_ctl.scala 225:50]
  wire  i0_dp_raw_word = i0_dec_io_out_word; // @[dec_decode_ctl.scala 124:37 dec_decode_ctl.scala 358:12]
  wire  i0_dp_word = _T_41 ? 1'h0 : i0_dp_raw_word; // @[dec_decode_ctl.scala 225:50]
  wire  i0_dp_raw_half = i0_dec_io_out_half; // @[dec_decode_ctl.scala 124:37 dec_decode_ctl.scala 358:12]
  wire  i0_dp_half = _T_41 ? 1'h0 : i0_dp_raw_half; // @[dec_decode_ctl.scala 225:50]
  wire  i0_dp_raw_by = i0_dec_io_out_by; // @[dec_decode_ctl.scala 124:37 dec_decode_ctl.scala 358:12]
  wire  i0_dp_by = _T_41 ? 1'h0 : i0_dp_raw_by; // @[dec_decode_ctl.scala 225:50]
  wire  i0_dp_jal = _T_41 ? 1'h0 : i0_dp_raw_jal; // @[dec_decode_ctl.scala 225:50]
  wire  i0_dp_raw_blt = i0_dec_io_out_blt; // @[dec_decode_ctl.scala 124:37 dec_decode_ctl.scala 358:12]
  wire  i0_dp_raw_bge = i0_dec_io_out_bge; // @[dec_decode_ctl.scala 124:37 dec_decode_ctl.scala 358:12]
  wire  i0_dp_raw_bne = i0_dec_io_out_bne; // @[dec_decode_ctl.scala 124:37 dec_decode_ctl.scala 358:12]
  wire  i0_dp_raw_beq = i0_dec_io_out_beq; // @[dec_decode_ctl.scala 124:37 dec_decode_ctl.scala 358:12]
  wire  i0_dp_condbr = _T_41 ? 1'h0 : i0_dp_raw_condbr; // @[dec_decode_ctl.scala 225:50]
  wire  i0_dp_raw_unsign = i0_dec_io_out_unsign; // @[dec_decode_ctl.scala 124:37 dec_decode_ctl.scala 358:12]
  wire  i0_dp_unsign = _T_41 ? 1'h0 : i0_dp_raw_unsign; // @[dec_decode_ctl.scala 225:50]
  wire  i0_dp_raw_slt = i0_dec_io_out_slt; // @[dec_decode_ctl.scala 124:37 dec_decode_ctl.scala 358:12]
  wire  i0_dp_raw_srl = i0_dec_io_out_srl; // @[dec_decode_ctl.scala 124:37 dec_decode_ctl.scala 358:12]
  wire  i0_dp_raw_sra = i0_dec_io_out_sra; // @[dec_decode_ctl.scala 124:37 dec_decode_ctl.scala 358:12]
  wire  i0_dp_raw_sll = i0_dec_io_out_sll; // @[dec_decode_ctl.scala 124:37 dec_decode_ctl.scala 358:12]
  wire  i0_dp_raw_lxor = i0_dec_io_out_lxor; // @[dec_decode_ctl.scala 124:37 dec_decode_ctl.scala 358:12]
  wire  i0_dp_raw_lor = i0_dec_io_out_lor; // @[dec_decode_ctl.scala 124:37 dec_decode_ctl.scala 358:12]
  wire  i0_dp_raw_land = i0_dec_io_out_land; // @[dec_decode_ctl.scala 124:37 dec_decode_ctl.scala 358:12]
  wire  i0_dp_raw_sub = i0_dec_io_out_sub; // @[dec_decode_ctl.scala 124:37 dec_decode_ctl.scala 358:12]
  wire  i0_dp_raw_add = i0_dec_io_out_add; // @[dec_decode_ctl.scala 124:37 dec_decode_ctl.scala 358:12]
  wire  i0_dp_raw_lsu = i0_dec_io_out_lsu; // @[dec_decode_ctl.scala 124:37 dec_decode_ctl.scala 358:12]
  wire  i0_dp_lsu = _T_41 ? 1'h0 : i0_dp_raw_lsu; // @[dec_decode_ctl.scala 225:50]
  wire  i0_dp_raw_store = i0_dec_io_out_store; // @[dec_decode_ctl.scala 124:37 dec_decode_ctl.scala 358:12]
  wire  i0_dp_store = _T_41 ? 1'h0 : i0_dp_raw_store; // @[dec_decode_ctl.scala 225:50]
  wire  i0_dp_raw_load = i0_dec_io_out_load; // @[dec_decode_ctl.scala 124:37 dec_decode_ctl.scala 358:12]
  wire  i0_dp_load = _T_41 ? 1'h0 : i0_dp_raw_load; // @[dec_decode_ctl.scala 225:50]
  wire  i0_dp_raw_pc = i0_dec_io_out_pc; // @[dec_decode_ctl.scala 124:37 dec_decode_ctl.scala 358:12]
  wire  i0_dp_imm20 = _T_41 ? 1'h0 : i0_dp_raw_imm20; // @[dec_decode_ctl.scala 225:50]
  wire  i0_dp_raw_shimm5 = i0_dec_io_out_shimm5; // @[dec_decode_ctl.scala 124:37 dec_decode_ctl.scala 358:12]
  wire  i0_dp_shimm5 = _T_41 ? 1'h0 : i0_dp_raw_shimm5; // @[dec_decode_ctl.scala 225:50]
  wire  i0_dp_raw_rd = i0_dec_io_out_rd; // @[dec_decode_ctl.scala 124:37 dec_decode_ctl.scala 358:12]
  wire  i0_dp_rd = _T_41 ? 1'h0 : i0_dp_raw_rd; // @[dec_decode_ctl.scala 225:50]
  wire  i0_dp_imm12 = _T_41 ? 1'h0 : i0_dp_raw_imm12; // @[dec_decode_ctl.scala 225:50]
  wire  i0_dp_raw_rs2 = i0_dec_io_out_rs2; // @[dec_decode_ctl.scala 124:37 dec_decode_ctl.scala 358:12]
  wire  i0_dp_rs2 = _T_41 | i0_dp_raw_rs2; // @[dec_decode_ctl.scala 225:50]
  wire  i0_dp_raw_rs1 = i0_dec_io_out_rs1; // @[dec_decode_ctl.scala 124:37 dec_decode_ctl.scala 358:12]
  wire  i0_dp_rs1 = _T_41 | i0_dp_raw_rs1; // @[dec_decode_ctl.scala 225:50]
  wire  i0_dp_raw_alu = i0_dec_io_out_alu; // @[dec_decode_ctl.scala 124:37 dec_decode_ctl.scala 358:12]
  wire  i0_dp_alu = _T_41 | i0_dp_raw_alu; // @[dec_decode_ctl.scala 225:50]
  wire  i0_pcall = i0_dp_jal & i0_pcall_case; // @[dec_decode_ctl.scala 376:38]
  wire  _T_44 = i0_dp_condbr | i0_pcall; // @[dec_decode_ctl.scala 239:54]
  wire  i0_pja = i0_dp_jal & i0_pja_case; // @[dec_decode_ctl.scala 378:38]
  wire  _T_45 = _T_44 | i0_pja; // @[dec_decode_ctl.scala 239:65]
  wire  i0_pret = i0_dp_jal & i0_pret_case; // @[dec_decode_ctl.scala 383:32]
  wire  i0_predict_br = _T_45 | i0_pret; // @[dec_decode_ctl.scala 239:74]
  wire  _T_47 = io_dec_i0_brp_bits_hist[1] & i0_brp_valid; // @[dec_decode_ctl.scala 240:69]
  wire  _T_48 = ~_T_47; // @[dec_decode_ctl.scala 240:40]
  wire  i0_ap_pc2 = ~io_dec_i0_pc4_d; // @[dec_decode_ctl.scala 242:40]
  wire  cam_data_reset = io_dctl_busbuff_lsu_nonblock_load_data_valid | io_dctl_busbuff_lsu_nonblock_load_data_error; // @[dec_decode_ctl.scala 275:76]
  reg [2:0] cam_raw_0_bits_tag; // @[dec_decode_ctl.scala 311:47]
  wire [2:0] _GEN_123 = {{1'd0}, io_dctl_busbuff_lsu_nonblock_load_data_tag}; // @[dec_decode_ctl.scala 286:67]
  wire  _T_94 = _GEN_123 == cam_raw_0_bits_tag; // @[dec_decode_ctl.scala 286:67]
  wire  _T_95 = cam_data_reset & _T_94; // @[dec_decode_ctl.scala 286:45]
  reg  cam_raw_0_valid; // @[dec_decode_ctl.scala 311:47]
  wire  cam_data_reset_val_0 = _T_95 & cam_raw_0_valid; // @[dec_decode_ctl.scala 286:88]
  wire  cam_0_valid = cam_data_reset_val_0 ? 1'h0 : cam_raw_0_valid; // @[dec_decode_ctl.scala 290:39]
  wire  _T_51 = ~cam_0_valid; // @[dec_decode_ctl.scala 267:78]
  reg [2:0] cam_raw_1_bits_tag; // @[dec_decode_ctl.scala 311:47]
  wire  _T_120 = _GEN_123 == cam_raw_1_bits_tag; // @[dec_decode_ctl.scala 286:67]
  wire  _T_121 = cam_data_reset & _T_120; // @[dec_decode_ctl.scala 286:45]
  reg  cam_raw_1_valid; // @[dec_decode_ctl.scala 311:47]
  wire  cam_data_reset_val_1 = _T_121 & cam_raw_1_valid; // @[dec_decode_ctl.scala 286:88]
  wire  cam_1_valid = cam_data_reset_val_1 ? 1'h0 : cam_raw_1_valid; // @[dec_decode_ctl.scala 290:39]
  wire  _T_54 = ~cam_1_valid; // @[dec_decode_ctl.scala 267:78]
  wire  _T_57 = cam_0_valid & _T_54; // @[dec_decode_ctl.scala 267:126]
  wire [1:0] _T_59 = {io_dctl_busbuff_lsu_nonblock_load_valid_m, 1'h0}; // @[dec_decode_ctl.scala 267:158]
  reg [2:0] cam_raw_2_bits_tag; // @[dec_decode_ctl.scala 311:47]
  wire  _T_146 = _GEN_123 == cam_raw_2_bits_tag; // @[dec_decode_ctl.scala 286:67]
  wire  _T_147 = cam_data_reset & _T_146; // @[dec_decode_ctl.scala 286:45]
  reg  cam_raw_2_valid; // @[dec_decode_ctl.scala 311:47]
  wire  cam_data_reset_val_2 = _T_147 & cam_raw_2_valid; // @[dec_decode_ctl.scala 286:88]
  wire  cam_2_valid = cam_data_reset_val_2 ? 1'h0 : cam_raw_2_valid; // @[dec_decode_ctl.scala 290:39]
  wire  _T_60 = ~cam_2_valid; // @[dec_decode_ctl.scala 267:78]
  wire  _T_63 = cam_0_valid & cam_1_valid; // @[dec_decode_ctl.scala 267:126]
  wire  _T_66 = _T_63 & _T_60; // @[dec_decode_ctl.scala 267:126]
  wire [2:0] _T_68 = {io_dctl_busbuff_lsu_nonblock_load_valid_m, 2'h0}; // @[dec_decode_ctl.scala 267:158]
  reg [2:0] cam_raw_3_bits_tag; // @[dec_decode_ctl.scala 311:47]
  wire  _T_172 = _GEN_123 == cam_raw_3_bits_tag; // @[dec_decode_ctl.scala 286:67]
  wire  _T_173 = cam_data_reset & _T_172; // @[dec_decode_ctl.scala 286:45]
  reg  cam_raw_3_valid; // @[dec_decode_ctl.scala 311:47]
  wire  cam_data_reset_val_3 = _T_173 & cam_raw_3_valid; // @[dec_decode_ctl.scala 286:88]
  wire  cam_3_valid = cam_data_reset_val_3 ? 1'h0 : cam_raw_3_valid; // @[dec_decode_ctl.scala 290:39]
  wire  _T_69 = ~cam_3_valid; // @[dec_decode_ctl.scala 267:78]
  wire  _T_75 = _T_63 & cam_2_valid; // @[dec_decode_ctl.scala 267:126]
  wire  _T_78 = _T_75 & _T_69; // @[dec_decode_ctl.scala 267:126]
  wire [3:0] _T_80 = {io_dctl_busbuff_lsu_nonblock_load_valid_m, 3'h0}; // @[dec_decode_ctl.scala 267:158]
  wire  _T_81 = _T_51 & io_dctl_busbuff_lsu_nonblock_load_valid_m; // @[Mux.scala 27:72]
  wire [1:0] _T_82 = _T_57 ? _T_59 : 2'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_83 = _T_66 ? _T_68 : 3'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_84 = _T_78 ? _T_80 : 4'h0; // @[Mux.scala 27:72]
  wire [1:0] _GEN_127 = {{1'd0}, _T_81}; // @[Mux.scala 27:72]
  wire [1:0] _T_85 = _GEN_127 | _T_82; // @[Mux.scala 27:72]
  wire [2:0] _GEN_128 = {{1'd0}, _T_85}; // @[Mux.scala 27:72]
  wire [2:0] _T_86 = _GEN_128 | _T_83; // @[Mux.scala 27:72]
  wire [3:0] _GEN_129 = {{1'd0}, _T_86}; // @[Mux.scala 27:72]
  wire [3:0] cam_wen = _GEN_129 | _T_84; // @[Mux.scala 27:72]
  reg  x_d_bits_i0load; // @[lib.scala 384:16]
  reg [4:0] x_d_bits_i0rd; // @[lib.scala 384:16]
  wire [4:0] nonblock_load_rd = x_d_bits_i0load ? x_d_bits_i0rd : 5'h0; // @[dec_decode_ctl.scala 278:31]
  reg [2:0] _T_706; // @[dec_decode_ctl.scala 616:80]
  wire [3:0] i0_pipe_en = {io_dec_aln_dec_i0_decode_d,_T_706}; // @[Cat.scala 29:58]
  wire  _T_712 = |i0_pipe_en[2:1]; // @[dec_decode_ctl.scala 619:49]
  wire  i0_r_ctl_en = _T_712 | io_clk_override; // @[dec_decode_ctl.scala 619:53]
  reg  nonblock_load_valid_m_delay; // @[Reg.scala 27:20]
  reg  r_d_bits_i0load; // @[lib.scala 384:16]
  wire  i0_load_kill_wen_r = nonblock_load_valid_m_delay & r_d_bits_i0load; // @[dec_decode_ctl.scala 283:56]
  wire [2:0] _GEN_130 = {{1'd0}, io_dctl_busbuff_lsu_nonblock_load_inv_tag_r}; // @[dec_decode_ctl.scala 285:66]
  wire  _T_91 = _GEN_130 == cam_raw_0_bits_tag; // @[dec_decode_ctl.scala 285:66]
  wire  _T_92 = io_dctl_busbuff_lsu_nonblock_load_inv_r & _T_91; // @[dec_decode_ctl.scala 285:45]
  wire  cam_inv_reset_val_0 = _T_92 & cam_0_valid; // @[dec_decode_ctl.scala 285:87]
  reg  r_d_bits_i0v; // @[lib.scala 384:16]
  wire  _T_748 = ~io_dec_tlu_flush_lower_wb; // @[dec_decode_ctl.scala 651:51]
  wire  r_d_in_bits_i0v = r_d_bits_i0v & _T_748; // @[dec_decode_ctl.scala 651:49]
  wire  _T_759 = ~io_dec_tlu_i0_kill_writeb_r; // @[dec_decode_ctl.scala 659:47]
  wire  i0_wen_r = r_d_in_bits_i0v & _T_759; // @[dec_decode_ctl.scala 659:45]
  reg [4:0] r_d_bits_i0rd; // @[lib.scala 384:16]
  reg [4:0] cam_raw_0_bits_rd; // @[dec_decode_ctl.scala 311:47]
  wire  _T_103 = r_d_bits_i0rd == cam_raw_0_bits_rd; // @[dec_decode_ctl.scala 298:85]
  wire  _T_104 = i0_wen_r & _T_103; // @[dec_decode_ctl.scala 298:64]
  reg  cam_raw_0_bits_wb; // @[dec_decode_ctl.scala 311:47]
  wire  _T_106 = _T_104 & cam_raw_0_bits_wb; // @[dec_decode_ctl.scala 298:105]
  wire  _T_107 = cam_inv_reset_val_0 | _T_106; // @[dec_decode_ctl.scala 298:44]
  wire  _GEN_52 = _T_107 ? 1'h0 : cam_0_valid; // @[dec_decode_ctl.scala 298:131]
  wire  _GEN_55 = _T_107 ? 1'h0 : cam_raw_0_bits_wb; // @[dec_decode_ctl.scala 298:131]
  wire  _GEN_56 = cam_wen[0] | _GEN_52; // @[dec_decode_ctl.scala 293:28]
  wire  _GEN_57 = cam_wen[0] ? 1'h0 : _GEN_55; // @[dec_decode_ctl.scala 293:28]
  wire  _T_110 = nonblock_load_valid_m_delay & _T_91; // @[dec_decode_ctl.scala 303:44]
  wire  _T_112 = _T_110 & cam_0_valid; // @[dec_decode_ctl.scala 303:113]
  wire  nonblock_load_write_0 = _T_94 & cam_raw_0_valid; // @[dec_decode_ctl.scala 312:71]
  wire  _T_117 = _GEN_130 == cam_raw_1_bits_tag; // @[dec_decode_ctl.scala 285:66]
  wire  _T_118 = io_dctl_busbuff_lsu_nonblock_load_inv_r & _T_117; // @[dec_decode_ctl.scala 285:45]
  wire  cam_inv_reset_val_1 = _T_118 & cam_1_valid; // @[dec_decode_ctl.scala 285:87]
  reg [4:0] cam_raw_1_bits_rd; // @[dec_decode_ctl.scala 311:47]
  wire  _T_129 = r_d_bits_i0rd == cam_raw_1_bits_rd; // @[dec_decode_ctl.scala 298:85]
  wire  _T_130 = i0_wen_r & _T_129; // @[dec_decode_ctl.scala 298:64]
  reg  cam_raw_1_bits_wb; // @[dec_decode_ctl.scala 311:47]
  wire  _T_132 = _T_130 & cam_raw_1_bits_wb; // @[dec_decode_ctl.scala 298:105]
  wire  _T_133 = cam_inv_reset_val_1 | _T_132; // @[dec_decode_ctl.scala 298:44]
  wire  _GEN_63 = _T_133 ? 1'h0 : cam_1_valid; // @[dec_decode_ctl.scala 298:131]
  wire  _GEN_66 = _T_133 ? 1'h0 : cam_raw_1_bits_wb; // @[dec_decode_ctl.scala 298:131]
  wire  _GEN_67 = cam_wen[1] | _GEN_63; // @[dec_decode_ctl.scala 293:28]
  wire  _GEN_68 = cam_wen[1] ? 1'h0 : _GEN_66; // @[dec_decode_ctl.scala 293:28]
  wire  _T_136 = nonblock_load_valid_m_delay & _T_117; // @[dec_decode_ctl.scala 303:44]
  wire  _T_138 = _T_136 & cam_1_valid; // @[dec_decode_ctl.scala 303:113]
  wire  nonblock_load_write_1 = _T_120 & cam_raw_1_valid; // @[dec_decode_ctl.scala 312:71]
  wire  _T_143 = _GEN_130 == cam_raw_2_bits_tag; // @[dec_decode_ctl.scala 285:66]
  wire  _T_144 = io_dctl_busbuff_lsu_nonblock_load_inv_r & _T_143; // @[dec_decode_ctl.scala 285:45]
  wire  cam_inv_reset_val_2 = _T_144 & cam_2_valid; // @[dec_decode_ctl.scala 285:87]
  reg [4:0] cam_raw_2_bits_rd; // @[dec_decode_ctl.scala 311:47]
  wire  _T_155 = r_d_bits_i0rd == cam_raw_2_bits_rd; // @[dec_decode_ctl.scala 298:85]
  wire  _T_156 = i0_wen_r & _T_155; // @[dec_decode_ctl.scala 298:64]
  reg  cam_raw_2_bits_wb; // @[dec_decode_ctl.scala 311:47]
  wire  _T_158 = _T_156 & cam_raw_2_bits_wb; // @[dec_decode_ctl.scala 298:105]
  wire  _T_159 = cam_inv_reset_val_2 | _T_158; // @[dec_decode_ctl.scala 298:44]
  wire  _GEN_74 = _T_159 ? 1'h0 : cam_2_valid; // @[dec_decode_ctl.scala 298:131]
  wire  _GEN_77 = _T_159 ? 1'h0 : cam_raw_2_bits_wb; // @[dec_decode_ctl.scala 298:131]
  wire  _GEN_78 = cam_wen[2] | _GEN_74; // @[dec_decode_ctl.scala 293:28]
  wire  _GEN_79 = cam_wen[2] ? 1'h0 : _GEN_77; // @[dec_decode_ctl.scala 293:28]
  wire  _T_162 = nonblock_load_valid_m_delay & _T_143; // @[dec_decode_ctl.scala 303:44]
  wire  _T_164 = _T_162 & cam_2_valid; // @[dec_decode_ctl.scala 303:113]
  wire  nonblock_load_write_2 = _T_146 & cam_raw_2_valid; // @[dec_decode_ctl.scala 312:71]
  wire  _T_169 = _GEN_130 == cam_raw_3_bits_tag; // @[dec_decode_ctl.scala 285:66]
  wire  _T_170 = io_dctl_busbuff_lsu_nonblock_load_inv_r & _T_169; // @[dec_decode_ctl.scala 285:45]
  wire  cam_inv_reset_val_3 = _T_170 & cam_3_valid; // @[dec_decode_ctl.scala 285:87]
  reg [4:0] cam_raw_3_bits_rd; // @[dec_decode_ctl.scala 311:47]
  wire  _T_181 = r_d_bits_i0rd == cam_raw_3_bits_rd; // @[dec_decode_ctl.scala 298:85]
  wire  _T_182 = i0_wen_r & _T_181; // @[dec_decode_ctl.scala 298:64]
  reg  cam_raw_3_bits_wb; // @[dec_decode_ctl.scala 311:47]
  wire  _T_184 = _T_182 & cam_raw_3_bits_wb; // @[dec_decode_ctl.scala 298:105]
  wire  _T_185 = cam_inv_reset_val_3 | _T_184; // @[dec_decode_ctl.scala 298:44]
  wire  _GEN_85 = _T_185 ? 1'h0 : cam_3_valid; // @[dec_decode_ctl.scala 298:131]
  wire  _GEN_88 = _T_185 ? 1'h0 : cam_raw_3_bits_wb; // @[dec_decode_ctl.scala 298:131]
  wire  _GEN_89 = cam_wen[3] | _GEN_85; // @[dec_decode_ctl.scala 293:28]
  wire  _GEN_90 = cam_wen[3] ? 1'h0 : _GEN_88; // @[dec_decode_ctl.scala 293:28]
  wire  _T_188 = nonblock_load_valid_m_delay & _T_169; // @[dec_decode_ctl.scala 303:44]
  wire  _T_190 = _T_188 & cam_3_valid; // @[dec_decode_ctl.scala 303:113]
  wire  nonblock_load_write_3 = _T_172 & cam_raw_3_valid; // @[dec_decode_ctl.scala 312:71]
  wire  _T_195 = r_d_bits_i0rd == io_dec_nonblock_load_waddr; // @[dec_decode_ctl.scala 317:49]
  wire  nonblock_load_cancel = _T_195 & i0_wen_r; // @[dec_decode_ctl.scala 317:81]
  wire  _T_196 = nonblock_load_write_0 | nonblock_load_write_1; // @[dec_decode_ctl.scala 318:108]
  wire  _T_197 = _T_196 | nonblock_load_write_2; // @[dec_decode_ctl.scala 318:108]
  wire  _T_198 = _T_197 | nonblock_load_write_3; // @[dec_decode_ctl.scala 318:108]
  wire  _T_200 = io_dctl_busbuff_lsu_nonblock_load_data_valid & _T_198; // @[dec_decode_ctl.scala 318:77]
  wire  _T_201 = ~nonblock_load_cancel; // @[dec_decode_ctl.scala 318:122]
  wire  _T_203 = nonblock_load_rd == i0r_rs1; // @[dec_decode_ctl.scala 319:54]
  wire  _T_204 = _T_203 & io_dctl_busbuff_lsu_nonblock_load_valid_m; // @[dec_decode_ctl.scala 319:66]
  wire  _T_205 = _T_204 & io_decode_exu_dec_i0_rs1_en_d; // @[dec_decode_ctl.scala 319:110]
  wire [4:0] i0r_rs2 = io_dec_i0_instr_d[24:20]; // @[dec_decode_ctl.scala 585:16]
  wire  _T_206 = nonblock_load_rd == i0r_rs2; // @[dec_decode_ctl.scala 319:161]
  wire  _T_207 = _T_206 & io_dctl_busbuff_lsu_nonblock_load_valid_m; // @[dec_decode_ctl.scala 319:173]
  wire  _T_208 = _T_207 & io_decode_exu_dec_i0_rs2_en_d; // @[dec_decode_ctl.scala 319:217]
  wire  i0_nonblock_boundary_stall = _T_205 | _T_208; // @[dec_decode_ctl.scala 319:142]
  wire [4:0] _T_210 = nonblock_load_write_0 ? 5'h1f : 5'h0; // @[Bitwise.scala 72:12]
  wire [4:0] _T_211 = _T_210 & cam_raw_0_bits_rd; // @[dec_decode_ctl.scala 323:88]
  wire  _T_212 = io_decode_exu_dec_i0_rs1_en_d & cam_0_valid; // @[dec_decode_ctl.scala 323:137]
  wire  _T_213 = cam_raw_0_bits_rd == i0r_rs1; // @[dec_decode_ctl.scala 323:170]
  wire  _T_214 = _T_212 & _T_213; // @[dec_decode_ctl.scala 323:152]
  wire  _T_215 = io_decode_exu_dec_i0_rs2_en_d & cam_0_valid; // @[dec_decode_ctl.scala 323:214]
  wire  _T_216 = cam_raw_0_bits_rd == i0r_rs2; // @[dec_decode_ctl.scala 323:247]
  wire  _T_217 = _T_215 & _T_216; // @[dec_decode_ctl.scala 323:229]
  wire [4:0] _T_219 = nonblock_load_write_1 ? 5'h1f : 5'h0; // @[Bitwise.scala 72:12]
  wire [4:0] _T_220 = _T_219 & cam_raw_1_bits_rd; // @[dec_decode_ctl.scala 323:88]
  wire  _T_221 = io_decode_exu_dec_i0_rs1_en_d & cam_1_valid; // @[dec_decode_ctl.scala 323:137]
  wire  _T_222 = cam_raw_1_bits_rd == i0r_rs1; // @[dec_decode_ctl.scala 323:170]
  wire  _T_223 = _T_221 & _T_222; // @[dec_decode_ctl.scala 323:152]
  wire  _T_224 = io_decode_exu_dec_i0_rs2_en_d & cam_1_valid; // @[dec_decode_ctl.scala 323:214]
  wire  _T_225 = cam_raw_1_bits_rd == i0r_rs2; // @[dec_decode_ctl.scala 323:247]
  wire  _T_226 = _T_224 & _T_225; // @[dec_decode_ctl.scala 323:229]
  wire [4:0] _T_228 = nonblock_load_write_2 ? 5'h1f : 5'h0; // @[Bitwise.scala 72:12]
  wire [4:0] _T_229 = _T_228 & cam_raw_2_bits_rd; // @[dec_decode_ctl.scala 323:88]
  wire  _T_230 = io_decode_exu_dec_i0_rs1_en_d & cam_2_valid; // @[dec_decode_ctl.scala 323:137]
  wire  _T_231 = cam_raw_2_bits_rd == i0r_rs1; // @[dec_decode_ctl.scala 323:170]
  wire  _T_232 = _T_230 & _T_231; // @[dec_decode_ctl.scala 323:152]
  wire  _T_233 = io_decode_exu_dec_i0_rs2_en_d & cam_2_valid; // @[dec_decode_ctl.scala 323:214]
  wire  _T_234 = cam_raw_2_bits_rd == i0r_rs2; // @[dec_decode_ctl.scala 323:247]
  wire  _T_235 = _T_233 & _T_234; // @[dec_decode_ctl.scala 323:229]
  wire [4:0] _T_237 = nonblock_load_write_3 ? 5'h1f : 5'h0; // @[Bitwise.scala 72:12]
  wire [4:0] _T_238 = _T_237 & cam_raw_3_bits_rd; // @[dec_decode_ctl.scala 323:88]
  wire  _T_239 = io_decode_exu_dec_i0_rs1_en_d & cam_3_valid; // @[dec_decode_ctl.scala 323:137]
  wire  _T_240 = cam_raw_3_bits_rd == i0r_rs1; // @[dec_decode_ctl.scala 323:170]
  wire  _T_241 = _T_239 & _T_240; // @[dec_decode_ctl.scala 323:152]
  wire  _T_242 = io_decode_exu_dec_i0_rs2_en_d & cam_3_valid; // @[dec_decode_ctl.scala 323:214]
  wire  _T_243 = cam_raw_3_bits_rd == i0r_rs2; // @[dec_decode_ctl.scala 323:247]
  wire  _T_244 = _T_242 & _T_243; // @[dec_decode_ctl.scala 323:229]
  wire [4:0] _T_245 = _T_211 | _T_220; // @[dec_decode_ctl.scala 324:69]
  wire [4:0] _T_246 = _T_245 | _T_229; // @[dec_decode_ctl.scala 324:69]
  wire  _T_247 = _T_214 | _T_223; // @[dec_decode_ctl.scala 324:102]
  wire  _T_248 = _T_247 | _T_232; // @[dec_decode_ctl.scala 324:102]
  wire  ld_stall_1 = _T_248 | _T_241; // @[dec_decode_ctl.scala 324:102]
  wire  _T_249 = _T_217 | _T_226; // @[dec_decode_ctl.scala 324:134]
  wire  _T_250 = _T_249 | _T_235; // @[dec_decode_ctl.scala 324:134]
  wire  ld_stall_2 = _T_250 | _T_244; // @[dec_decode_ctl.scala 324:134]
  wire  _T_251 = ld_stall_1 | ld_stall_2; // @[dec_decode_ctl.scala 326:38]
  wire  i0_nonblock_load_stall = _T_251 | i0_nonblock_boundary_stall; // @[dec_decode_ctl.scala 326:51]
  wire  _T_253 = ~i0_predict_br; // @[dec_decode_ctl.scala 335:34]
  wire [3:0] _T_255 = i0_legal_decode_d ? 4'hf : 4'h0; // @[Bitwise.scala 72:12]
  wire  csr_read = i0_dp_csr_read & i0_legal_decode_d; // @[dec_decode_ctl.scala 419:36]
  wire  _T_256 = csr_read & io_dec_csr_wen_unq_d; // @[dec_decode_ctl.scala 347:16]
  wire  _T_258 = ~csr_read; // @[dec_decode_ctl.scala 348:6]
  wire  _T_259 = _T_258 & io_dec_csr_wen_unq_d; // @[dec_decode_ctl.scala 348:16]
  wire  _T_261 = ~io_dec_csr_wen_unq_d; // @[dec_decode_ctl.scala 349:18]
  wire  _T_262 = csr_read & _T_261; // @[dec_decode_ctl.scala 349:16]
  wire [3:0] _T_264 = i0_dp_mul ? 4'h1 : 4'h0; // @[Mux.scala 98:16]
  wire [3:0] _T_265 = i0_dp_load ? 4'h2 : _T_264; // @[Mux.scala 98:16]
  wire [3:0] _T_266 = i0_dp_store ? 4'h3 : _T_265; // @[Mux.scala 98:16]
  wire [3:0] _T_267 = i0_dp_pm_alu ? 4'h4 : _T_266; // @[Mux.scala 98:16]
  wire [3:0] _T_268 = _T_262 ? 4'h5 : _T_267; // @[Mux.scala 98:16]
  wire [3:0] _T_269 = _T_259 ? 4'h6 : _T_268; // @[Mux.scala 98:16]
  wire [3:0] _T_270 = _T_256 ? 4'h7 : _T_269; // @[Mux.scala 98:16]
  wire [3:0] _T_271 = i0_dp_ebreak ? 4'h8 : _T_270; // @[Mux.scala 98:16]
  wire [3:0] _T_272 = i0_dp_ecall ? 4'h9 : _T_271; // @[Mux.scala 98:16]
  wire [3:0] _T_273 = i0_dp_fence ? 4'ha : _T_272; // @[Mux.scala 98:16]
  wire [3:0] _T_274 = i0_dp_fence_i ? 4'hb : _T_273; // @[Mux.scala 98:16]
  wire [3:0] _T_275 = i0_dp_mret ? 4'hc : _T_274; // @[Mux.scala 98:16]
  wire [3:0] _T_276 = i0_dp_condbr ? 4'hd : _T_275; // @[Mux.scala 98:16]
  wire [3:0] _T_277 = i0_dp_jal ? 4'he : _T_276; // @[Mux.scala 98:16]
  reg  lsu_idle; // @[dec_decode_ctl.scala 360:45]
  wire  _T_333 = ~i0_pcall_case; // @[dec_decode_ctl.scala 384:35]
  wire  _T_334 = i0_dp_jal & _T_333; // @[dec_decode_ctl.scala 384:32]
  wire  _T_335 = ~i0_pja_case; // @[dec_decode_ctl.scala 384:52]
  wire  _T_336 = _T_334 & _T_335; // @[dec_decode_ctl.scala 384:50]
  wire  _T_337 = ~i0_pret_case; // @[dec_decode_ctl.scala 384:67]
  reg  _T_339; // @[dec_decode_ctl.scala 396:69]
  wire  lsu_decode_d = i0_legal_decode_d & i0_dp_lsu; // @[dec_decode_ctl.scala 538:40]
  wire  _T_907 = i0_dp_load | i0_dp_store; // @[dec_decode_ctl.scala 752:43]
  reg  x_d_bits_i0v; // @[lib.scala 384:16]
  wire  _T_881 = io_decode_exu_dec_i0_rs1_en_d & x_d_bits_i0v; // @[dec_decode_ctl.scala 732:59]
  wire  _T_882 = x_d_bits_i0rd == i0r_rs1; // @[dec_decode_ctl.scala 732:91]
  wire  i0_rs1_depend_i0_x = _T_881 & _T_882; // @[dec_decode_ctl.scala 732:74]
  wire  _T_883 = io_decode_exu_dec_i0_rs1_en_d & r_d_bits_i0v; // @[dec_decode_ctl.scala 733:59]
  wire  _T_884 = r_d_bits_i0rd == i0r_rs1; // @[dec_decode_ctl.scala 733:91]
  wire  i0_rs1_depend_i0_r = _T_883 & _T_884; // @[dec_decode_ctl.scala 733:74]
  wire [1:0] _T_896 = i0_rs1_depend_i0_r ? 2'h2 : 2'h0; // @[dec_decode_ctl.scala 739:63]
  wire [1:0] i0_rs1_depth_d = i0_rs1_depend_i0_x ? 2'h1 : _T_896; // @[dec_decode_ctl.scala 739:24]
  wire  _T_909 = _T_907 & i0_rs1_depth_d[0]; // @[dec_decode_ctl.scala 752:58]
  reg  i0_x_c_load; // @[Reg.scala 27:20]
  reg  i0_r_c_load; // @[Reg.scala 27:20]
  wire  _T_892_load = i0_rs1_depend_i0_r & i0_r_c_load; // @[dec_decode_ctl.scala 738:61]
  wire  i0_rs1_class_d_load = i0_rs1_depend_i0_x ? i0_x_c_load : _T_892_load; // @[dec_decode_ctl.scala 738:24]
  wire  load_ldst_bypass_d = _T_909 & i0_rs1_class_d_load; // @[dec_decode_ctl.scala 752:78]
  wire  _T_885 = io_decode_exu_dec_i0_rs2_en_d & x_d_bits_i0v; // @[dec_decode_ctl.scala 735:59]
  wire  _T_886 = x_d_bits_i0rd == i0r_rs2; // @[dec_decode_ctl.scala 735:91]
  wire  i0_rs2_depend_i0_x = _T_885 & _T_886; // @[dec_decode_ctl.scala 735:74]
  wire  _T_887 = io_decode_exu_dec_i0_rs2_en_d & r_d_bits_i0v; // @[dec_decode_ctl.scala 736:59]
  wire  _T_888 = r_d_bits_i0rd == i0r_rs2; // @[dec_decode_ctl.scala 736:91]
  wire  i0_rs2_depend_i0_r = _T_887 & _T_888; // @[dec_decode_ctl.scala 736:74]
  wire [1:0] _T_905 = i0_rs2_depend_i0_r ? 2'h2 : 2'h0; // @[dec_decode_ctl.scala 741:63]
  wire [1:0] i0_rs2_depth_d = i0_rs2_depend_i0_x ? 2'h1 : _T_905; // @[dec_decode_ctl.scala 741:24]
  wire  _T_912 = i0_dp_store & i0_rs2_depth_d[0]; // @[dec_decode_ctl.scala 753:43]
  wire  _T_901_load = i0_rs2_depend_i0_r & i0_r_c_load; // @[dec_decode_ctl.scala 740:61]
  wire  i0_rs2_class_d_load = i0_rs2_depend_i0_x ? i0_x_c_load : _T_901_load; // @[dec_decode_ctl.scala 740:24]
  wire  store_data_bypass_d = _T_912 & i0_rs2_class_d_load; // @[dec_decode_ctl.scala 753:63]
  wire  _T_349 = i0_dp_csr_clr | i0_dp_csr_set; // @[dec_decode_ctl.scala 427:42]
  reg  r_d_bits_csrwen; // @[lib.scala 384:16]
  reg  r_d_valid; // @[lib.scala 384:16]
  wire  _T_352 = r_d_bits_csrwen & r_d_valid; // @[dec_decode_ctl.scala 435:39]
  reg [11:0] r_d_bits_csrwaddr; // @[lib.scala 384:16]
  wire  _T_355 = r_d_bits_csrwaddr == 12'h300; // @[dec_decode_ctl.scala 438:50]
  wire  _T_356 = r_d_bits_csrwaddr == 12'h304; // @[dec_decode_ctl.scala 438:85]
  wire  _T_357 = _T_355 | _T_356; // @[dec_decode_ctl.scala 438:64]
  wire  _T_358 = _T_357 & r_d_bits_csrwen; // @[dec_decode_ctl.scala 438:100]
  wire  _T_359 = _T_358 & r_d_valid; // @[dec_decode_ctl.scala 438:118]
  wire  _T_360 = ~io_dec_tlu_i0_kill_writeb_wb; // @[dec_decode_ctl.scala 438:132]
  reg  csr_read_x; // @[dec_decode_ctl.scala 440:52]
  reg  csr_clr_x; // @[dec_decode_ctl.scala 441:51]
  reg  csr_set_x; // @[dec_decode_ctl.scala 442:51]
  reg  csr_write_x; // @[dec_decode_ctl.scala 443:53]
  reg  csr_imm_x; // @[dec_decode_ctl.scala 444:51]
  wire  i0_x_data_en = i0_pipe_en[3] | io_clk_override; // @[dec_decode_ctl.scala 621:50]
  reg [4:0] csrimm_x; // @[lib.scala 374:16]
  reg [31:0] csr_rddata_x; // @[lib.scala 374:16]
  wire [31:0] _T_394 = {27'h0,csrimm_x}; // @[Cat.scala 29:58]
  wire  _T_396 = ~csr_imm_x; // @[dec_decode_ctl.scala 452:5]
  wire [31:0] _T_397 = csr_imm_x ? _T_394 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_398 = _T_396 ? io_decode_exu_exu_csr_rs1_x : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] csr_mask_x = _T_397 | _T_398; // @[Mux.scala 27:72]
  wire [31:0] _T_400 = ~csr_mask_x; // @[dec_decode_ctl.scala 455:38]
  wire [31:0] _T_401 = csr_rddata_x & _T_400; // @[dec_decode_ctl.scala 455:35]
  wire [31:0] _T_402 = csr_rddata_x | csr_mask_x; // @[dec_decode_ctl.scala 456:35]
  wire [31:0] _T_403 = csr_clr_x ? _T_401 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_404 = csr_set_x ? _T_402 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_405 = csr_write_x ? csr_mask_x : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_406 = _T_403 | _T_404; // @[Mux.scala 27:72]
  wire [31:0] write_csr_data_x = _T_406 | _T_405; // @[Mux.scala 27:72]
  wire  _T_421 = ~tlu_wr_pause_r1; // @[dec_decode_ctl.scala 466:44]
  wire  _T_422 = ~tlu_wr_pause_r2; // @[dec_decode_ctl.scala 466:64]
  wire  _T_423 = _T_421 & _T_422; // @[dec_decode_ctl.scala 466:61]
  wire [31:0] _T_426 = write_csr_data - 32'h1; // @[dec_decode_ctl.scala 469:59]
  wire  _T_428 = csr_clr_x | csr_set_x; // @[dec_decode_ctl.scala 471:34]
  wire  _T_429 = _T_428 | csr_write_x; // @[dec_decode_ctl.scala 471:46]
  wire  _T_430 = _T_429 & csr_read_x; // @[dec_decode_ctl.scala 471:61]
  wire  _T_431 = _T_430 | io_dec_tlu_wr_pause_r; // @[dec_decode_ctl.scala 471:75]
  reg  r_d_bits_csrwonly; // @[lib.scala 384:16]
  wire  _T_769 = r_d_bits_i0v & r_d_bits_i0load; // @[dec_decode_ctl.scala 674:42]
  reg [31:0] i0_result_r_raw; // @[lib.scala 374:16]
  wire [31:0] i0_result_corr_r = _T_769 ? io_lsu_result_corr_r : i0_result_r_raw; // @[dec_decode_ctl.scala 674:27]
  reg  x_d_bits_csrwonly; // @[lib.scala 384:16]
  wire  _T_435 = x_d_bits_csrwonly | r_d_bits_csrwonly; // @[dec_decode_ctl.scala 480:43]
  reg  wbd_bits_csrwonly; // @[lib.scala 384:16]
  wire  prior_csr_write = _T_435 | wbd_bits_csrwonly; // @[dec_decode_ctl.scala 480:63]
  wire  debug_fence_raw = io_dec_debug_fence_d & io_dbg_dctl_dbg_cmd_wrdata[1]; // @[dec_decode_ctl.scala 483:48]
  wire  debug_fence = debug_fence_raw | debug_fence_i; // @[dec_decode_ctl.scala 484:40]
  wire  _T_439 = i0_dp_presync | io_dec_tlu_presync_d; // @[dec_decode_ctl.scala 487:34]
  wire  _T_440 = _T_439 | debug_fence_i; // @[dec_decode_ctl.scala 487:57]
  wire  _T_441 = _T_440 | debug_fence_raw; // @[dec_decode_ctl.scala 487:73]
  wire  i0_presync = _T_441 | io_dec_tlu_pipelining_disable; // @[dec_decode_ctl.scala 487:91]
  wire [31:0] _T_465 = {16'h0,io_dec_aln_ifu_i0_cinst}; // @[Cat.scala 29:58]
  wire  _T_467 = ~illegal_lockout; // @[dec_decode_ctl.scala 499:44]
  reg [31:0] _T_468; // @[lib.scala 374:16]
  wire  i0_div_prior_div_stall = i0_dp_div & io_dec_div_active; // @[dec_decode_ctl.scala 503:42]
  wire  _T_473 = i0_dp_csr_read & prior_csr_write; // @[dec_decode_ctl.scala 505:40]
  wire  _T_474 = _T_473 | io_decode_exu_dec_extint_stall; // @[dec_decode_ctl.scala 505:59]
  wire  _T_475 = _T_474 | pause_stall; // @[dec_decode_ctl.scala 505:92]
  wire  _T_476 = _T_475 | leak1_i0_stall; // @[dec_decode_ctl.scala 505:106]
  wire  _T_477 = _T_476 | io_dec_tlu_debug_stall; // @[dec_decode_ctl.scala 506:20]
  wire  _T_478 = _T_477 | postsync_stall; // @[dec_decode_ctl.scala 506:45]
  wire  prior_inflight = x_d_valid | r_d_valid; // @[dec_decode_ctl.scala 528:41]
  wire  prior_inflight_eff = i0_dp_div ? x_d_valid : prior_inflight; // @[dec_decode_ctl.scala 529:31]
  wire  presync_stall = i0_presync & prior_inflight_eff; // @[dec_decode_ctl.scala 531:37]
  wire  _T_479 = _T_478 | presync_stall; // @[dec_decode_ctl.scala 506:62]
  wire  _T_480 = i0_dp_fence | debug_fence; // @[dec_decode_ctl.scala 507:19]
  wire  _T_481 = ~lsu_idle; // @[dec_decode_ctl.scala 507:36]
  wire  _T_482 = _T_480 & _T_481; // @[dec_decode_ctl.scala 507:34]
  wire  _T_483 = _T_479 | _T_482; // @[dec_decode_ctl.scala 506:79]
  wire  _T_484 = _T_483 | i0_nonblock_load_stall; // @[dec_decode_ctl.scala 507:47]
  wire  _T_827 = io_decode_exu_dec_i0_rs1_en_d & io_dec_div_active; // @[dec_decode_ctl.scala 702:60]
  wire  _T_828 = io_div_waddr_wb == i0r_rs1; // @[dec_decode_ctl.scala 702:99]
  wire  _T_829 = _T_827 & _T_828; // @[dec_decode_ctl.scala 702:80]
  wire  _T_830 = io_decode_exu_dec_i0_rs2_en_d & io_dec_div_active; // @[dec_decode_ctl.scala 703:36]
  wire  _T_831 = io_div_waddr_wb == i0r_rs2; // @[dec_decode_ctl.scala 703:75]
  wire  _T_832 = _T_830 & _T_831; // @[dec_decode_ctl.scala 703:56]
  wire  i0_nonblock_div_stall = _T_829 | _T_832; // @[dec_decode_ctl.scala 702:113]
  wire  _T_486 = _T_484 | i0_nonblock_div_stall; // @[dec_decode_ctl.scala 508:21]
  wire  i0_block_raw_d = _T_486 | i0_div_prior_div_stall; // @[dec_decode_ctl.scala 508:45]
  wire  _T_487 = io_lsu_store_stall_any | io_dctl_dma_dma_dccm_stall_any; // @[dec_decode_ctl.scala 510:65]
  wire  i0_store_stall_d = i0_dp_store & _T_487; // @[dec_decode_ctl.scala 510:39]
  wire  _T_488 = io_lsu_load_stall_any | io_dctl_dma_dma_dccm_stall_any; // @[dec_decode_ctl.scala 511:63]
  wire  i0_load_stall_d = i0_dp_load & _T_488; // @[dec_decode_ctl.scala 511:38]
  wire  _T_489 = i0_block_raw_d | i0_store_stall_d; // @[dec_decode_ctl.scala 512:38]
  wire  i0_block_d = _T_489 | i0_load_stall_d; // @[dec_decode_ctl.scala 512:57]
  wire  _T_490 = ~i0_block_d; // @[dec_decode_ctl.scala 516:54]
  wire  _T_491 = io_dec_ib0_valid_d & _T_490; // @[dec_decode_ctl.scala 516:52]
  wire  _T_493 = _T_491 & _T_280; // @[dec_decode_ctl.scala 516:69]
  wire  _T_496 = ~i0_block_raw_d; // @[dec_decode_ctl.scala 517:46]
  wire  _T_497 = io_dec_ib0_valid_d & _T_496; // @[dec_decode_ctl.scala 517:44]
  wire  _T_499 = _T_497 & _T_280; // @[dec_decode_ctl.scala 517:61]
  wire  i0_exudecode_d = _T_499 & _T_470; // @[dec_decode_ctl.scala 517:89]
  wire  i0_exulegal_decode_d = i0_exudecode_d & i0_legal; // @[dec_decode_ctl.scala 518:46]
  wire  _T_501 = ~io_dec_aln_dec_i0_decode_d; // @[dec_decode_ctl.scala 522:51]
  wire  _T_520 = i0_dp_fence_i | debug_fence_i; // @[dec_decode_ctl.scala 550:44]
  wire [3:0] _T_525 = {io_dec_aln_dec_i0_decode_d,io_dec_aln_dec_i0_decode_d,io_dec_aln_dec_i0_decode_d,io_dec_aln_dec_i0_decode_d}; // @[Cat.scala 29:58]
  wire  _T_709 = |i0_pipe_en[3:2]; // @[dec_decode_ctl.scala 618:49]
  wire  i0_x_ctl_en = _T_709 | io_clk_override; // @[dec_decode_ctl.scala 618:53]
  reg  x_t_legal; // @[lib.scala 384:16]
  reg  x_t_icaf; // @[lib.scala 384:16]
  reg  x_t_icaf_f1; // @[lib.scala 384:16]
  reg [1:0] x_t_icaf_type; // @[lib.scala 384:16]
  reg  x_t_fence_i; // @[lib.scala 384:16]
  reg [3:0] x_t_i0trigger; // @[lib.scala 384:16]
  reg [3:0] x_t_pmu_i0_itype; // @[lib.scala 384:16]
  reg  x_t_pmu_i0_br_unpred; // @[lib.scala 384:16]
  wire [3:0] _T_533 = {io_dec_tlu_flush_lower_wb,io_dec_tlu_flush_lower_wb,io_dec_tlu_flush_lower_wb,io_dec_tlu_flush_lower_wb}; // @[Cat.scala 29:58]
  wire [3:0] _T_534 = ~_T_533; // @[dec_decode_ctl.scala 563:39]
  reg  r_t_legal; // @[lib.scala 384:16]
  reg  r_t_icaf; // @[lib.scala 384:16]
  reg  r_t_icaf_f1; // @[lib.scala 384:16]
  reg [1:0] r_t_icaf_type; // @[lib.scala 384:16]
  reg  r_t_fence_i; // @[lib.scala 384:16]
  reg [3:0] r_t_i0trigger; // @[lib.scala 384:16]
  reg [3:0] r_t_pmu_i0_itype; // @[lib.scala 384:16]
  reg  r_t_pmu_i0_br_unpred; // @[lib.scala 384:16]
  reg [3:0] lsu_trigger_match_r; // @[dec_decode_ctl.scala 566:36]
  reg  lsu_pmu_misaligned_r; // @[dec_decode_ctl.scala 567:37]
  reg  r_d_bits_i0store; // @[lib.scala 384:16]
  wire  _T_539 = r_d_bits_i0load | r_d_bits_i0store; // @[dec_decode_ctl.scala 571:61]
  wire [3:0] _T_543 = {_T_539,_T_539,_T_539,_T_539}; // @[Cat.scala 29:58]
  wire [3:0] _T_544 = _T_543 & lsu_trigger_match_r; // @[dec_decode_ctl.scala 571:82]
  wire [3:0] _T_545 = _T_544 | r_t_i0trigger; // @[dec_decode_ctl.scala 571:105]
  reg  r_d_bits_i0div; // @[lib.scala 384:16]
  wire  _T_548 = r_d_bits_i0div & r_d_valid; // @[dec_decode_ctl.scala 577:58]
  wire  _T_559 = i0r_rs1 != 5'h0; // @[dec_decode_ctl.scala 588:60]
  wire  _T_561 = i0r_rs2 != 5'h0; // @[dec_decode_ctl.scala 589:60]
  wire  _T_563 = i0r_rd != 5'h0; // @[dec_decode_ctl.scala 590:48]
  wire  i0_rd_en_d = i0_dp_rd & _T_563; // @[dec_decode_ctl.scala 590:37]
  wire  i0_jalimm20 = i0_dp_jal & i0_dp_imm20; // @[dec_decode_ctl.scala 594:38]
  wire  _T_564 = ~i0_dp_jal; // @[dec_decode_ctl.scala 595:27]
  wire  i0_uiimm20 = _T_564 & i0_dp_imm20; // @[dec_decode_ctl.scala 595:38]
  wire [31:0] _T_566 = i0_dp_csr_read ? io_dec_csr_rddata_d : 32'h0; // @[Mux.scala 27:72]
  wire [9:0] _T_580 = {io_dec_i0_instr_d[31],io_dec_i0_instr_d[31],io_dec_i0_instr_d[31],io_dec_i0_instr_d[31],io_dec_i0_instr_d[31],io_dec_i0_instr_d[31],io_dec_i0_instr_d[31],io_dec_i0_instr_d[31],io_dec_i0_instr_d[31],io_dec_i0_instr_d[31]}; // @[Cat.scala 29:58]
  wire [18:0] _T_589 = {_T_580,io_dec_i0_instr_d[31],io_dec_i0_instr_d[31],io_dec_i0_instr_d[31],io_dec_i0_instr_d[31],io_dec_i0_instr_d[31],io_dec_i0_instr_d[31],io_dec_i0_instr_d[31],io_dec_i0_instr_d[31],io_dec_i0_instr_d[31]}; // @[Cat.scala 29:58]
  wire [31:0] _T_592 = {_T_589,io_dec_i0_instr_d[31],io_dec_i0_instr_d[31:20]}; // @[Cat.scala 29:58]
  wire [31:0] _T_687 = i0_dp_imm12 ? _T_592 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_621 = {27'h0,i0r_rs2}; // @[Cat.scala 29:58]
  wire [31:0] _T_688 = i0_dp_shimm5 ? _T_621 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_692 = _T_687 | _T_688; // @[Mux.scala 27:72]
  wire [31:0] _T_641 = {_T_580,io_dec_i0_instr_d[31],io_dec_i0_instr_d[31],io_dec_i0_instr_d[19:12],io_dec_i0_instr_d[20],io_dec_i0_instr_d[30:21],1'h0}; // @[Cat.scala 29:58]
  wire [31:0] _T_689 = i0_jalimm20 ? _T_641 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_693 = _T_692 | _T_689; // @[Mux.scala 27:72]
  wire [31:0] _T_655 = {io_dec_i0_instr_d[31:12],12'h0}; // @[Cat.scala 29:58]
  wire [31:0] _T_690 = i0_uiimm20 ? _T_655 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_694 = _T_693 | _T_690; // @[Mux.scala 27:72]
  wire  _T_656 = i0_csr_write_only_d & i0_dp_csr_imm; // @[dec_decode_ctl.scala 606:26]
  wire [31:0] _T_686 = {27'h0,i0r_rs1}; // @[Cat.scala 29:58]
  wire [31:0] _T_691 = _T_656 ? _T_686 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] i0_immed_d = _T_694 | _T_691; // @[Mux.scala 27:72]
  wire [31:0] _T_567 = _T_347 ? i0_immed_d : 32'h0; // @[Mux.scala 27:72]
  wire  i0_d_c_mul = i0_dp_mul & i0_legal_decode_d; // @[dec_decode_ctl.scala 610:44]
  wire  i0_d_c_load = i0_dp_load & i0_legal_decode_d; // @[dec_decode_ctl.scala 611:44]
  wire  i0_d_c_alu = i0_dp_alu & i0_legal_decode_d; // @[dec_decode_ctl.scala 612:44]
  reg  i0_x_c_mul; // @[Reg.scala 27:20]
  reg  i0_x_c_alu; // @[Reg.scala 27:20]
  reg  i0_r_c_mul; // @[Reg.scala 27:20]
  reg  i0_r_c_alu; // @[Reg.scala 27:20]
  wire  _T_715 = |i0_pipe_en[1:0]; // @[dec_decode_ctl.scala 620:49]
  wire  i0_r_data_en = i0_pipe_en[2] | io_clk_override; // @[dec_decode_ctl.scala 622:50]
  reg  x_d_bits_i0store; // @[lib.scala 384:16]
  reg  x_d_bits_i0div; // @[lib.scala 384:16]
  reg  x_d_bits_csrwen; // @[lib.scala 384:16]
  reg [11:0] x_d_bits_csrwaddr; // @[lib.scala 384:16]
  wire  _T_738 = x_d_bits_i0v & _T_748; // @[dec_decode_ctl.scala 644:47]
  wire  _T_742 = x_d_valid & _T_748; // @[dec_decode_ctl.scala 645:33]
  wire  _T_761 = ~r_d_bits_i0div; // @[dec_decode_ctl.scala 660:49]
  wire  _T_762 = i0_wen_r & _T_761; // @[dec_decode_ctl.scala 660:47]
  wire  _T_763 = ~i0_load_kill_wen_r; // @[dec_decode_ctl.scala 660:70]
  wire  _T_766 = x_d_bits_i0v & x_d_bits_i0load; // @[dec_decode_ctl.scala 669:47]
  wire  _T_773 = io_decode_exu_i0_ap_predict_nt & _T_564; // @[dec_decode_ctl.scala 675:71]
  wire [11:0] _T_786 = {10'h0,io_dec_i0_pc4_d,i0_ap_pc2}; // @[Cat.scala 29:58]
  reg [11:0] last_br_immed_x; // @[lib.scala 374:16]
  wire  _T_804 = x_d_bits_i0div & x_d_valid; // @[dec_decode_ctl.scala 683:45]
  wire  div_e1_to_r = _T_804 | _T_548; // @[dec_decode_ctl.scala 683:58]
  wire  _T_807 = x_d_bits_i0rd == 5'h0; // @[dec_decode_ctl.scala 685:77]
  wire  _T_808 = _T_804 & _T_807; // @[dec_decode_ctl.scala 685:60]
  wire  _T_810 = _T_804 & io_dec_tlu_flush_lower_r; // @[dec_decode_ctl.scala 686:33]
  wire  _T_811 = _T_808 | _T_810; // @[dec_decode_ctl.scala 685:94]
  wire  _T_813 = _T_548 & io_dec_tlu_flush_lower_r; // @[dec_decode_ctl.scala 687:33]
  wire  _T_814 = _T_813 & io_dec_tlu_i0_kill_writeb_r; // @[dec_decode_ctl.scala 687:60]
  wire  div_flush = _T_811 | _T_814; // @[dec_decode_ctl.scala 686:62]
  wire  _T_815 = io_dec_div_active & div_flush; // @[dec_decode_ctl.scala 691:51]
  wire  _T_816 = ~div_e1_to_r; // @[dec_decode_ctl.scala 692:26]
  wire  _T_817 = io_dec_div_active & _T_816; // @[dec_decode_ctl.scala 692:24]
  wire  _T_818 = r_d_bits_i0rd == io_div_waddr_wb; // @[dec_decode_ctl.scala 692:56]
  wire  _T_819 = _T_817 & _T_818; // @[dec_decode_ctl.scala 692:39]
  wire  _T_820 = _T_819 & i0_wen_r; // @[dec_decode_ctl.scala 692:77]
  wire  nonblock_div_cancel = _T_815 | _T_820; // @[dec_decode_ctl.scala 691:65]
  wire  i0_div_decode_d = i0_legal_decode_d & i0_dp_div; // @[dec_decode_ctl.scala 695:55]
  wire  _T_822 = ~io_exu_div_wren; // @[dec_decode_ctl.scala 697:62]
  wire  _T_823 = io_dec_div_active & _T_822; // @[dec_decode_ctl.scala 697:60]
  wire  _T_824 = ~nonblock_div_cancel; // @[dec_decode_ctl.scala 697:81]
  wire  _T_825 = _T_823 & _T_824; // @[dec_decode_ctl.scala 697:79]
  reg  _T_826; // @[dec_decode_ctl.scala 699:54]
  reg [4:0] _T_835; // @[Reg.scala 27:20]
  reg [31:0] i0_inst_x; // @[lib.scala 374:16]
  reg [31:0] i0_inst_r; // @[lib.scala 374:16]
  reg [31:0] i0_inst_wb; // @[lib.scala 374:16]
  reg [31:0] _T_842; // @[lib.scala 374:16]
  reg [30:0] i0_pc_wb; // @[lib.scala 374:16]
  reg [30:0] _T_845; // @[lib.scala 374:16]
  reg [30:0] dec_i0_pc_r; // @[lib.scala 374:16]
  wire [31:0] _T_847 = {io_dec_alu_exu_i0_pc_x,1'h0}; // @[Cat.scala 29:58]
  wire [12:0] _T_848 = {last_br_immed_x,1'h0}; // @[Cat.scala 29:58]
  wire [12:0] _T_851 = _T_847[12:1] + _T_848[12:1]; // @[lib.scala 68:31]
  wire [18:0] _T_854 = _T_847[31:13] + 19'h1; // @[lib.scala 69:27]
  wire [18:0] _T_857 = _T_847[31:13] - 19'h1; // @[lib.scala 70:27]
  wire  _T_860 = ~_T_851[12]; // @[lib.scala 72:28]
  wire  _T_861 = _T_848[12] ^ _T_860; // @[lib.scala 72:26]
  wire  _T_864 = ~_T_848[12]; // @[lib.scala 73:20]
  wire  _T_866 = _T_864 & _T_851[12]; // @[lib.scala 73:26]
  wire  _T_870 = _T_848[12] & _T_860; // @[lib.scala 74:26]
  wire [18:0] _T_872 = _T_861 ? _T_847[31:13] : 19'h0; // @[Mux.scala 27:72]
  wire [18:0] _T_873 = _T_866 ? _T_854 : 19'h0; // @[Mux.scala 27:72]
  wire [18:0] _T_874 = _T_870 ? _T_857 : 19'h0; // @[Mux.scala 27:72]
  wire [18:0] _T_875 = _T_872 | _T_873; // @[Mux.scala 27:72]
  wire [18:0] _T_876 = _T_875 | _T_874; // @[Mux.scala 27:72]
  wire [31:0] temp_pred_correct_npc_x = {_T_876,_T_851[11:0],1'h0}; // @[Cat.scala 29:58]
  wire  _T_892_mul = i0_rs1_depend_i0_r & i0_r_c_mul; // @[dec_decode_ctl.scala 738:61]
  wire  _T_892_alu = i0_rs1_depend_i0_r & i0_r_c_alu; // @[dec_decode_ctl.scala 738:61]
  wire  i0_rs1_class_d_mul = i0_rs1_depend_i0_x ? i0_x_c_mul : _T_892_mul; // @[dec_decode_ctl.scala 738:24]
  wire  i0_rs1_class_d_alu = i0_rs1_depend_i0_x ? i0_x_c_alu : _T_892_alu; // @[dec_decode_ctl.scala 738:24]
  wire  _T_901_mul = i0_rs2_depend_i0_r & i0_r_c_mul; // @[dec_decode_ctl.scala 740:61]
  wire  _T_901_alu = i0_rs2_depend_i0_r & i0_r_c_alu; // @[dec_decode_ctl.scala 740:61]
  wire  i0_rs2_class_d_mul = i0_rs2_depend_i0_x ? i0_x_c_mul : _T_901_mul; // @[dec_decode_ctl.scala 740:24]
  wire  i0_rs2_class_d_alu = i0_rs2_depend_i0_x ? i0_x_c_alu : _T_901_alu; // @[dec_decode_ctl.scala 740:24]
  wire  _T_914 = io_decode_exu_dec_i0_rs1_en_d & io_dec_nonblock_load_wen; // @[dec_decode_ctl.scala 758:73]
  wire  _T_915 = io_dec_nonblock_load_waddr == i0r_rs1; // @[dec_decode_ctl.scala 758:130]
  wire  i0_rs1_nonblock_load_bypass_en_d = _T_914 & _T_915; // @[dec_decode_ctl.scala 758:100]
  wire  _T_916 = io_decode_exu_dec_i0_rs2_en_d & io_dec_nonblock_load_wen; // @[dec_decode_ctl.scala 760:73]
  wire  _T_917 = io_dec_nonblock_load_waddr == i0r_rs2; // @[dec_decode_ctl.scala 760:130]
  wire  i0_rs2_nonblock_load_bypass_en_d = _T_916 & _T_917; // @[dec_decode_ctl.scala 760:100]
  wire  _T_919 = i0_rs1_class_d_alu | i0_rs1_class_d_mul; // @[dec_decode_ctl.scala 763:66]
  wire  _T_920 = i0_rs1_depth_d[0] & _T_919; // @[dec_decode_ctl.scala 763:45]
  wire  _T_922 = i0_rs1_depth_d[0] & i0_rs1_class_d_load; // @[dec_decode_ctl.scala 763:108]
  wire  _T_925 = _T_919 | i0_rs1_class_d_load; // @[dec_decode_ctl.scala 763:196]
  wire  _T_926 = i0_rs1_depth_d[1] & _T_925; // @[dec_decode_ctl.scala 763:153]
  wire [2:0] i0_rs1bypass = {_T_920,_T_922,_T_926}; // @[Cat.scala 29:58]
  wire  _T_930 = i0_rs2_class_d_alu | i0_rs2_class_d_mul; // @[dec_decode_ctl.scala 765:67]
  wire  _T_931 = i0_rs2_depth_d[0] & _T_930; // @[dec_decode_ctl.scala 765:45]
  wire  _T_933 = i0_rs2_depth_d[0] & i0_rs2_class_d_load; // @[dec_decode_ctl.scala 765:109]
  wire  _T_936 = _T_930 | i0_rs2_class_d_load; // @[dec_decode_ctl.scala 765:196]
  wire  _T_937 = i0_rs2_depth_d[1] & _T_936; // @[dec_decode_ctl.scala 765:153]
  wire [2:0] i0_rs2bypass = {_T_931,_T_933,_T_937}; // @[Cat.scala 29:58]
  wire  _T_943 = i0_rs1bypass[1] | i0_rs1bypass[0]; // @[dec_decode_ctl.scala 767:86]
  wire  _T_945 = ~i0_rs1bypass[2]; // @[dec_decode_ctl.scala 767:107]
  wire  _T_946 = _T_945 & i0_rs1_nonblock_load_bypass_en_d; // @[dec_decode_ctl.scala 767:124]
  wire  _T_947 = _T_943 | _T_946; // @[dec_decode_ctl.scala 767:104]
  wire  _T_952 = i0_rs2bypass[1] | i0_rs2bypass[0]; // @[dec_decode_ctl.scala 768:86]
  wire  _T_954 = ~i0_rs2bypass[2]; // @[dec_decode_ctl.scala 768:107]
  wire  _T_955 = _T_954 & i0_rs2_nonblock_load_bypass_en_d; // @[dec_decode_ctl.scala 768:124]
  wire  _T_956 = _T_952 | _T_955; // @[dec_decode_ctl.scala 768:104]
  wire  _T_963 = ~i0_rs1bypass[1]; // @[dec_decode_ctl.scala 774:6]
  wire  _T_965 = ~i0_rs1bypass[0]; // @[dec_decode_ctl.scala 774:25]
  wire  _T_966 = _T_963 & _T_965; // @[dec_decode_ctl.scala 774:23]
  wire  _T_967 = _T_966 & i0_rs1_nonblock_load_bypass_en_d; // @[dec_decode_ctl.scala 774:42]
  wire [31:0] _T_969 = i0_rs1bypass[1] ? io_lsu_result_m : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_970 = i0_rs1bypass[0] ? i0_result_r_raw : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_971 = _T_967 ? io_dctl_busbuff_lsu_nonblock_load_data : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_972 = _T_969 | _T_970; // @[Mux.scala 27:72]
  wire  _T_980 = ~i0_rs2bypass[1]; // @[dec_decode_ctl.scala 779:6]
  wire  _T_982 = ~i0_rs2bypass[0]; // @[dec_decode_ctl.scala 779:25]
  wire  _T_983 = _T_980 & _T_982; // @[dec_decode_ctl.scala 779:23]
  wire  _T_984 = _T_983 & i0_rs2_nonblock_load_bypass_en_d; // @[dec_decode_ctl.scala 779:42]
  wire [31:0] _T_986 = i0_rs2bypass[1] ? io_lsu_result_m : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_987 = i0_rs2bypass[0] ? i0_result_r_raw : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_988 = _T_984 ? io_dctl_busbuff_lsu_nonblock_load_data : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_989 = _T_986 | _T_987; // @[Mux.scala 27:72]
  wire  _T_992 = i0_dp_raw_load | i0_dp_raw_store; // @[dec_decode_ctl.scala 781:68]
  wire  _T_993 = io_dec_ib0_valid_d & _T_992; // @[dec_decode_ctl.scala 781:50]
  wire  _T_994 = ~io_dctl_dma_dma_dccm_stall_any; // @[dec_decode_ctl.scala 781:89]
  wire  _T_995 = _T_993 & _T_994; // @[dec_decode_ctl.scala 781:87]
  wire  _T_997 = _T_995 & _T_496; // @[dec_decode_ctl.scala 781:121]
  wire  _T_999 = ~io_decode_exu_dec_extint_stall; // @[dec_decode_ctl.scala 783:6]
  wire  _T_1000 = _T_999 & i0_dp_lsu; // @[dec_decode_ctl.scala 783:38]
  wire  _T_1001 = _T_1000 & i0_dp_load; // @[dec_decode_ctl.scala 783:50]
  wire  _T_1006 = _T_1000 & i0_dp_store; // @[dec_decode_ctl.scala 784:50]
  wire [11:0] _T_1010 = {io_dec_i0_instr_d[31:25],i0r_rd}; // @[Cat.scala 29:58]
  wire [11:0] _T_1011 = _T_1001 ? io_dec_i0_instr_d[31:20] : 12'h0; // @[Mux.scala 27:72]
  wire [11:0] _T_1012 = _T_1006 ? _T_1010 : 12'h0; // @[Mux.scala 27:72]
  rvclkhdr rvclkhdr ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_io_l1clk),
    .io_clk(rvclkhdr_io_clk),
    .io_en(rvclkhdr_io_en),
    .io_scan_mode(rvclkhdr_io_scan_mode)
  );
  dec_dec_ctl i0_dec ( // @[dec_decode_ctl.scala 356:22]
    .io_ins(i0_dec_io_ins),
    .io_out_alu(i0_dec_io_out_alu),
    .io_out_rs1(i0_dec_io_out_rs1),
    .io_out_rs2(i0_dec_io_out_rs2),
    .io_out_imm12(i0_dec_io_out_imm12),
    .io_out_rd(i0_dec_io_out_rd),
    .io_out_shimm5(i0_dec_io_out_shimm5),
    .io_out_imm20(i0_dec_io_out_imm20),
    .io_out_pc(i0_dec_io_out_pc),
    .io_out_load(i0_dec_io_out_load),
    .io_out_store(i0_dec_io_out_store),
    .io_out_lsu(i0_dec_io_out_lsu),
    .io_out_add(i0_dec_io_out_add),
    .io_out_sub(i0_dec_io_out_sub),
    .io_out_land(i0_dec_io_out_land),
    .io_out_lor(i0_dec_io_out_lor),
    .io_out_lxor(i0_dec_io_out_lxor),
    .io_out_sll(i0_dec_io_out_sll),
    .io_out_sra(i0_dec_io_out_sra),
    .io_out_srl(i0_dec_io_out_srl),
    .io_out_slt(i0_dec_io_out_slt),
    .io_out_unsign(i0_dec_io_out_unsign),
    .io_out_condbr(i0_dec_io_out_condbr),
    .io_out_beq(i0_dec_io_out_beq),
    .io_out_bne(i0_dec_io_out_bne),
    .io_out_bge(i0_dec_io_out_bge),
    .io_out_blt(i0_dec_io_out_blt),
    .io_out_jal(i0_dec_io_out_jal),
    .io_out_by(i0_dec_io_out_by),
    .io_out_half(i0_dec_io_out_half),
    .io_out_word(i0_dec_io_out_word),
    .io_out_csr_read(i0_dec_io_out_csr_read),
    .io_out_csr_clr(i0_dec_io_out_csr_clr),
    .io_out_csr_set(i0_dec_io_out_csr_set),
    .io_out_csr_write(i0_dec_io_out_csr_write),
    .io_out_csr_imm(i0_dec_io_out_csr_imm),
    .io_out_presync(i0_dec_io_out_presync),
    .io_out_postsync(i0_dec_io_out_postsync),
    .io_out_ebreak(i0_dec_io_out_ebreak),
    .io_out_ecall(i0_dec_io_out_ecall),
    .io_out_mret(i0_dec_io_out_mret),
    .io_out_mul(i0_dec_io_out_mul),
    .io_out_rs1_sign(i0_dec_io_out_rs1_sign),
    .io_out_rs2_sign(i0_dec_io_out_rs2_sign),
    .io_out_low(i0_dec_io_out_low),
    .io_out_div(i0_dec_io_out_div),
    .io_out_rem(i0_dec_io_out_rem),
    .io_out_fence(i0_dec_io_out_fence),
    .io_out_fence_i(i0_dec_io_out_fence_i),
    .io_out_pm_alu(i0_dec_io_out_pm_alu),
    .io_out_legal(i0_dec_io_out_legal)
  );
  rvclkhdr rvclkhdr_1 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_1_io_l1clk),
    .io_clk(rvclkhdr_1_io_clk),
    .io_en(rvclkhdr_1_io_en),
    .io_scan_mode(rvclkhdr_1_io_scan_mode)
  );
  rvclkhdr rvclkhdr_2 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_2_io_l1clk),
    .io_clk(rvclkhdr_2_io_clk),
    .io_en(rvclkhdr_2_io_en),
    .io_scan_mode(rvclkhdr_2_io_scan_mode)
  );
  rvclkhdr rvclkhdr_3 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_3_io_l1clk),
    .io_clk(rvclkhdr_3_io_clk),
    .io_en(rvclkhdr_3_io_en),
    .io_scan_mode(rvclkhdr_3_io_scan_mode)
  );
  rvclkhdr rvclkhdr_4 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_4_io_l1clk),
    .io_clk(rvclkhdr_4_io_clk),
    .io_en(rvclkhdr_4_io_en),
    .io_scan_mode(rvclkhdr_4_io_scan_mode)
  );
  rvclkhdr rvclkhdr_5 ( // @[lib.scala 378:23]
    .io_l1clk(rvclkhdr_5_io_l1clk),
    .io_clk(rvclkhdr_5_io_clk),
    .io_en(rvclkhdr_5_io_en),
    .io_scan_mode(rvclkhdr_5_io_scan_mode)
  );
  rvclkhdr rvclkhdr_6 ( // @[lib.scala 378:23]
    .io_l1clk(rvclkhdr_6_io_l1clk),
    .io_clk(rvclkhdr_6_io_clk),
    .io_en(rvclkhdr_6_io_en),
    .io_scan_mode(rvclkhdr_6_io_scan_mode)
  );
  rvclkhdr rvclkhdr_7 ( // @[lib.scala 378:23]
    .io_l1clk(rvclkhdr_7_io_l1clk),
    .io_clk(rvclkhdr_7_io_clk),
    .io_en(rvclkhdr_7_io_en),
    .io_scan_mode(rvclkhdr_7_io_scan_mode)
  );
  rvclkhdr rvclkhdr_8 ( // @[lib.scala 378:23]
    .io_l1clk(rvclkhdr_8_io_l1clk),
    .io_clk(rvclkhdr_8_io_clk),
    .io_en(rvclkhdr_8_io_en),
    .io_scan_mode(rvclkhdr_8_io_scan_mode)
  );
  rvclkhdr rvclkhdr_9 ( // @[lib.scala 378:23]
    .io_l1clk(rvclkhdr_9_io_l1clk),
    .io_clk(rvclkhdr_9_io_clk),
    .io_en(rvclkhdr_9_io_en),
    .io_scan_mode(rvclkhdr_9_io_scan_mode)
  );
  rvclkhdr rvclkhdr_10 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_10_io_l1clk),
    .io_clk(rvclkhdr_10_io_clk),
    .io_en(rvclkhdr_10_io_en),
    .io_scan_mode(rvclkhdr_10_io_scan_mode)
  );
  rvclkhdr rvclkhdr_11 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_11_io_l1clk),
    .io_clk(rvclkhdr_11_io_clk),
    .io_en(rvclkhdr_11_io_en),
    .io_scan_mode(rvclkhdr_11_io_scan_mode)
  );
  rvclkhdr rvclkhdr_12 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_12_io_l1clk),
    .io_clk(rvclkhdr_12_io_clk),
    .io_en(rvclkhdr_12_io_en),
    .io_scan_mode(rvclkhdr_12_io_scan_mode)
  );
  rvclkhdr rvclkhdr_13 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_13_io_l1clk),
    .io_clk(rvclkhdr_13_io_clk),
    .io_en(rvclkhdr_13_io_en),
    .io_scan_mode(rvclkhdr_13_io_scan_mode)
  );
  rvclkhdr rvclkhdr_14 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_14_io_l1clk),
    .io_clk(rvclkhdr_14_io_clk),
    .io_en(rvclkhdr_14_io_en),
    .io_scan_mode(rvclkhdr_14_io_scan_mode)
  );
  rvclkhdr rvclkhdr_15 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_15_io_l1clk),
    .io_clk(rvclkhdr_15_io_clk),
    .io_en(rvclkhdr_15_io_en),
    .io_scan_mode(rvclkhdr_15_io_scan_mode)
  );
  rvclkhdr rvclkhdr_16 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_16_io_l1clk),
    .io_clk(rvclkhdr_16_io_clk),
    .io_en(rvclkhdr_16_io_en),
    .io_scan_mode(rvclkhdr_16_io_scan_mode)
  );
  rvclkhdr rvclkhdr_17 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_17_io_l1clk),
    .io_clk(rvclkhdr_17_io_clk),
    .io_en(rvclkhdr_17_io_en),
    .io_scan_mode(rvclkhdr_17_io_scan_mode)
  );
  rvclkhdr rvclkhdr_18 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_18_io_l1clk),
    .io_clk(rvclkhdr_18_io_clk),
    .io_en(rvclkhdr_18_io_en),
    .io_scan_mode(rvclkhdr_18_io_scan_mode)
  );
  rvclkhdr rvclkhdr_19 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_19_io_l1clk),
    .io_clk(rvclkhdr_19_io_clk),
    .io_en(rvclkhdr_19_io_en),
    .io_scan_mode(rvclkhdr_19_io_scan_mode)
  );
  assign io_decode_exu_dec_data_en = {i0_x_data_en,i0_r_data_en}; // @[dec_decode_ctl.scala 626:38]
  assign io_decode_exu_dec_ctl_en = {i0_x_ctl_en,i0_r_ctl_en}; // @[dec_decode_ctl.scala 627:38]
  assign io_decode_exu_i0_ap_land = _T_41 ? 1'h0 : i0_dp_raw_land; // @[dec_decode_ctl.scala 249:37]
  assign io_decode_exu_i0_ap_lor = _T_41 | i0_dp_raw_lor; // @[dec_decode_ctl.scala 250:37]
  assign io_decode_exu_i0_ap_lxor = _T_41 ? 1'h0 : i0_dp_raw_lxor; // @[dec_decode_ctl.scala 251:37]
  assign io_decode_exu_i0_ap_sll = _T_41 ? 1'h0 : i0_dp_raw_sll; // @[dec_decode_ctl.scala 252:37]
  assign io_decode_exu_i0_ap_srl = _T_41 ? 1'h0 : i0_dp_raw_srl; // @[dec_decode_ctl.scala 253:37]
  assign io_decode_exu_i0_ap_sra = _T_41 ? 1'h0 : i0_dp_raw_sra; // @[dec_decode_ctl.scala 254:37]
  assign io_decode_exu_i0_ap_beq = _T_41 ? 1'h0 : i0_dp_raw_beq; // @[dec_decode_ctl.scala 257:37]
  assign io_decode_exu_i0_ap_bne = _T_41 ? 1'h0 : i0_dp_raw_bne; // @[dec_decode_ctl.scala 258:37]
  assign io_decode_exu_i0_ap_blt = _T_41 ? 1'h0 : i0_dp_raw_blt; // @[dec_decode_ctl.scala 259:37]
  assign io_decode_exu_i0_ap_bge = _T_41 ? 1'h0 : i0_dp_raw_bge; // @[dec_decode_ctl.scala 260:37]
  assign io_decode_exu_i0_ap_add = _T_41 ? 1'h0 : i0_dp_raw_add; // @[dec_decode_ctl.scala 247:37]
  assign io_decode_exu_i0_ap_sub = _T_41 ? 1'h0 : i0_dp_raw_sub; // @[dec_decode_ctl.scala 248:37]
  assign io_decode_exu_i0_ap_slt = _T_41 ? 1'h0 : i0_dp_raw_slt; // @[dec_decode_ctl.scala 255:37]
  assign io_decode_exu_i0_ap_unsign = _T_41 ? 1'h0 : i0_dp_raw_unsign; // @[dec_decode_ctl.scala 256:37]
  assign io_decode_exu_i0_ap_jal = _T_336 & _T_337; // @[dec_decode_ctl.scala 263:37]
  assign io_decode_exu_i0_ap_predict_t = _T_47 & i0_predict_br; // @[dec_decode_ctl.scala 245:37]
  assign io_decode_exu_i0_ap_predict_nt = _T_48 & i0_predict_br; // @[dec_decode_ctl.scala 244:37]
  assign io_decode_exu_i0_ap_csr_write = i0_csr_write & _T_347; // @[dec_decode_ctl.scala 261:37]
  assign io_decode_exu_i0_ap_csr_imm = _T_41 ? 1'h0 : i0_dp_raw_csr_imm; // @[dec_decode_ctl.scala 262:37]
  assign io_decode_exu_dec_i0_predict_p_d_valid = i0_brp_valid & i0_legal_decode_d; // @[dec_decode_ctl.scala 202:55]
  assign io_decode_exu_dec_i0_predict_p_d_bits_pc4 = io_dec_i0_pc4_d; // @[dec_decode_ctl.scala 200:55]
  assign io_decode_exu_dec_i0_predict_p_d_bits_hist = io_dec_i0_brp_bits_hist; // @[dec_decode_ctl.scala 201:55]
  assign io_decode_exu_dec_i0_predict_p_d_bits_toffset = _T_314 ? i0_pcall_imm[11:0] : _T_323; // @[dec_decode_ctl.scala 214:56]
  assign io_decode_exu_dec_i0_predict_p_d_bits_br_error = _T_33 & _T_18; // @[dec_decode_ctl.scala 209:56]
  assign io_decode_exu_dec_i0_predict_p_d_bits_br_start_error = _T_36 & _T_18; // @[dec_decode_ctl.scala 210:56]
  assign io_decode_exu_dec_i0_predict_p_d_bits_prett = io_dec_i0_brp_bits_prett; // @[dec_decode_ctl.scala 199:55]
  assign io_decode_exu_dec_i0_predict_p_d_bits_pcall = i0_dp_jal & i0_pcall_case; // @[dec_decode_ctl.scala 196:55]
  assign io_decode_exu_dec_i0_predict_p_d_bits_pret = i0_dp_jal & i0_pret_case; // @[dec_decode_ctl.scala 198:55]
  assign io_decode_exu_dec_i0_predict_p_d_bits_pja = i0_dp_jal & i0_pja_case; // @[dec_decode_ctl.scala 197:55]
  assign io_decode_exu_dec_i0_predict_p_d_bits_way = io_dec_i0_brp_bits_way; // @[dec_decode_ctl.scala 216:56]
  assign io_decode_exu_i0_predict_fghr_d = io_dec_i0_bp_fghr; // @[dec_decode_ctl.scala 215:56]
  assign io_decode_exu_i0_predict_index_d = io_dec_i0_bp_index; // @[dec_decode_ctl.scala 211:56]
  assign io_decode_exu_i0_predict_btag_d = io_dec_i0_bp_btag; // @[dec_decode_ctl.scala 212:56]
  assign io_decode_exu_dec_i0_rs1_en_d = i0_dp_rs1 & _T_559; // @[dec_decode_ctl.scala 588:35]
  assign io_decode_exu_dec_i0_rs2_en_d = i0_dp_rs2 & _T_561; // @[dec_decode_ctl.scala 589:35]
  assign io_decode_exu_dec_i0_immed_d = _T_566 | _T_567; // @[dec_decode_ctl.scala 597:32]
  assign io_decode_exu_dec_i0_rs1_bypass_data_d = _T_972 | _T_971; // @[dec_decode_ctl.scala 771:42]
  assign io_decode_exu_dec_i0_rs2_bypass_data_d = _T_989 | _T_988; // @[dec_decode_ctl.scala 776:42]
  assign io_decode_exu_dec_i0_select_pc_d = _T_41 ? 1'h0 : i0_dp_raw_pc; // @[dec_decode_ctl.scala 236:36]
  assign io_decode_exu_dec_i0_rs1_bypass_en_d = {i0_rs1bypass[2],_T_947}; // @[dec_decode_ctl.scala 767:45]
  assign io_decode_exu_dec_i0_rs2_bypass_en_d = {i0_rs2bypass[2],_T_956}; // @[dec_decode_ctl.scala 768:45]
  assign io_decode_exu_mul_p_valid = i0_exulegal_decode_d & i0_dp_mul; // @[dec_decode_ctl.scala 95:25 dec_decode_ctl.scala 391:32]
  assign io_decode_exu_mul_p_bits_rs1_sign = _T_41 ? 1'h0 : i0_dp_raw_rs1_sign; // @[dec_decode_ctl.scala 95:25 dec_decode_ctl.scala 392:37]
  assign io_decode_exu_mul_p_bits_rs2_sign = _T_41 ? 1'h0 : i0_dp_raw_rs2_sign; // @[dec_decode_ctl.scala 95:25 dec_decode_ctl.scala 393:37]
  assign io_decode_exu_mul_p_bits_low = _T_41 ? 1'h0 : i0_dp_raw_low; // @[dec_decode_ctl.scala 95:25 dec_decode_ctl.scala 394:37]
  assign io_decode_exu_pred_correct_npc_x = temp_pred_correct_npc_x[31:1]; // @[dec_decode_ctl.scala 728:36]
  assign io_decode_exu_dec_extint_stall = _T_339; // @[dec_decode_ctl.scala 396:34]
  assign io_dec_alu_dec_i0_alu_decode_d = i0_exulegal_decode_d & i0_dp_alu; // @[dec_decode_ctl.scala 536:34]
  assign io_dec_alu_dec_csr_ren_d = _T_41 ? 1'h0 : i0_dp_raw_csr_read; // @[dec_decode_ctl.scala 418:29]
  assign io_dec_alu_dec_i0_br_immed_d = _T_773 ? i0_br_offset : _T_786; // @[dec_decode_ctl.scala 675:32]
  assign io_dec_div_div_p_valid = i0_exulegal_decode_d & i0_dp_div; // @[dec_decode_ctl.scala 387:29]
  assign io_dec_div_div_p_bits_unsign = _T_41 ? 1'h0 : i0_dp_raw_unsign; // @[dec_decode_ctl.scala 388:34]
  assign io_dec_div_div_p_bits_rem = _T_41 ? 1'h0 : i0_dp_raw_rem; // @[dec_decode_ctl.scala 389:34]
  assign io_dec_div_dec_div_cancel = _T_815 | _T_820; // @[dec_decode_ctl.scala 694:37]
  assign io_dec_aln_dec_i0_decode_d = _T_493 & _T_470; // @[dec_decode_ctl.scala 516:30 dec_decode_ctl.scala 582:30]
  assign io_dec_i0_inst_wb1 = _T_842; // @[dec_decode_ctl.scala 717:22]
  assign io_dec_i0_pc_wb1 = _T_845; // @[dec_decode_ctl.scala 720:20]
  assign io_dec_i0_rs1_d = io_dec_i0_instr_d[19:15]; // @[dec_decode_ctl.scala 591:19]
  assign io_dec_i0_rs2_d = io_dec_i0_instr_d[24:20]; // @[dec_decode_ctl.scala 592:19]
  assign io_dec_i0_waddr_r = r_d_bits_i0rd; // @[dec_decode_ctl.scala 658:27]
  assign io_dec_i0_wen_r = _T_762 & _T_763; // @[dec_decode_ctl.scala 660:32]
  assign io_dec_i0_wdata_r = _T_769 ? io_lsu_result_corr_r : i0_result_r_raw; // @[dec_decode_ctl.scala 661:26]
  assign io_lsu_p_valid = io_decode_exu_dec_extint_stall | lsu_decode_d; // @[dec_decode_ctl.scala 398:12 dec_decode_ctl.scala 403:24 dec_decode_ctl.scala 405:35]
  assign io_lsu_p_bits_fast_int = io_decode_exu_dec_extint_stall; // @[dec_decode_ctl.scala 398:12 dec_decode_ctl.scala 402:29]
  assign io_lsu_p_bits_by = io_decode_exu_dec_extint_stall ? 1'h0 : i0_dp_by; // @[dec_decode_ctl.scala 398:12 dec_decode_ctl.scala 408:40]
  assign io_lsu_p_bits_half = io_decode_exu_dec_extint_stall ? 1'h0 : i0_dp_half; // @[dec_decode_ctl.scala 398:12 dec_decode_ctl.scala 409:40]
  assign io_lsu_p_bits_word = io_decode_exu_dec_extint_stall | i0_dp_word; // @[dec_decode_ctl.scala 398:12 dec_decode_ctl.scala 401:29 dec_decode_ctl.scala 410:40]
  assign io_lsu_p_bits_load = io_decode_exu_dec_extint_stall | i0_dp_load; // @[dec_decode_ctl.scala 398:12 dec_decode_ctl.scala 400:29 dec_decode_ctl.scala 406:40]
  assign io_lsu_p_bits_store = io_decode_exu_dec_extint_stall ? 1'h0 : i0_dp_store; // @[dec_decode_ctl.scala 398:12 dec_decode_ctl.scala 407:40]
  assign io_lsu_p_bits_unsign = io_decode_exu_dec_extint_stall ? 1'h0 : i0_dp_unsign; // @[dec_decode_ctl.scala 398:12 dec_decode_ctl.scala 414:40]
  assign io_lsu_p_bits_store_data_bypass_d = io_decode_exu_dec_extint_stall ? 1'h0 : store_data_bypass_d; // @[dec_decode_ctl.scala 398:12 dec_decode_ctl.scala 412:40]
  assign io_lsu_p_bits_load_ldst_bypass_d = io_decode_exu_dec_extint_stall ? 1'h0 : load_ldst_bypass_d; // @[dec_decode_ctl.scala 398:12 dec_decode_ctl.scala 411:40]
  assign io_div_waddr_wb = _T_835; // @[dec_decode_ctl.scala 705:19]
  assign io_dec_lsu_valid_raw_d = _T_997 | io_decode_exu_dec_extint_stall; // @[dec_decode_ctl.scala 781:26]
  assign io_dec_lsu_offset_d = _T_1011 | _T_1012; // @[dec_decode_ctl.scala 782:23]
  assign io_dec_csr_wen_unq_d = _T_349 | i0_csr_write; // @[dec_decode_ctl.scala 427:24]
  assign io_dec_csr_any_unq_d = i0_dp_csr_read | i0_csr_write; // @[dec_decode_ctl.scala 493:24]
  assign io_dec_csr_rdaddr_d = io_dec_i0_instr_d[31:20]; // @[dec_decode_ctl.scala 430:24]
  assign io_dec_csr_wen_r = _T_352 & _T_759; // @[dec_decode_ctl.scala 435:20]
  assign io_dec_csr_wraddr_r = r_d_bits_csrwaddr; // @[dec_decode_ctl.scala 431:23]
  assign io_dec_csr_wrdata_r = r_d_bits_csrwonly ? i0_result_corr_r : write_csr_data; // @[dec_decode_ctl.scala 478:24]
  assign io_dec_csr_stall_int_ff = _T_359 & _T_360; // @[dec_decode_ctl.scala 438:27]
  assign io_dec_tlu_i0_valid_r = r_d_valid & _T_748; // @[dec_decode_ctl.scala 542:29]
  assign io_dec_tlu_packet_r_legal = io_dec_tlu_flush_lower_wb ? 1'h0 : r_t_legal; // @[dec_decode_ctl.scala 576:39]
  assign io_dec_tlu_packet_r_icaf = io_dec_tlu_flush_lower_wb ? 1'h0 : r_t_icaf; // @[dec_decode_ctl.scala 576:39]
  assign io_dec_tlu_packet_r_icaf_f1 = io_dec_tlu_flush_lower_wb ? 1'h0 : r_t_icaf_f1; // @[dec_decode_ctl.scala 576:39]
  assign io_dec_tlu_packet_r_icaf_type = io_dec_tlu_flush_lower_wb ? 2'h0 : r_t_icaf_type; // @[dec_decode_ctl.scala 576:39]
  assign io_dec_tlu_packet_r_fence_i = io_dec_tlu_flush_lower_wb ? 1'h0 : r_t_fence_i; // @[dec_decode_ctl.scala 576:39]
  assign io_dec_tlu_packet_r_i0trigger = io_dec_tlu_flush_lower_wb ? 4'h0 : _T_545; // @[dec_decode_ctl.scala 576:39]
  assign io_dec_tlu_packet_r_pmu_i0_itype = io_dec_tlu_flush_lower_wb ? 4'h0 : r_t_pmu_i0_itype; // @[dec_decode_ctl.scala 576:39]
  assign io_dec_tlu_packet_r_pmu_i0_br_unpred = io_dec_tlu_flush_lower_wb ? 1'h0 : r_t_pmu_i0_br_unpred; // @[dec_decode_ctl.scala 576:39]
  assign io_dec_tlu_packet_r_pmu_divide = r_d_bits_i0div & r_d_valid; // @[dec_decode_ctl.scala 576:39 dec_decode_ctl.scala 577:39]
  assign io_dec_tlu_packet_r_pmu_lsu_misaligned = io_dec_tlu_flush_lower_wb ? 1'h0 : lsu_pmu_misaligned_r; // @[dec_decode_ctl.scala 576:39]
  assign io_dec_tlu_i0_pc_r = dec_i0_pc_r; // @[dec_decode_ctl.scala 723:27]
  assign io_dec_illegal_inst = _T_468; // @[dec_decode_ctl.scala 500:23]
  assign io_dec_pmu_instr_decoded = io_dec_aln_dec_i0_decode_d; // @[dec_decode_ctl.scala 521:28]
  assign io_dec_pmu_decode_stall = io_dec_ib0_valid_d & _T_501; // @[dec_decode_ctl.scala 522:27]
  assign io_dec_pmu_presync_stall = i0_presync & prior_inflight_eff; // @[dec_decode_ctl.scala 524:29]
  assign io_dec_pmu_postsync_stall = postsync_stall; // @[dec_decode_ctl.scala 523:29]
  assign io_dec_nonblock_load_wen = _T_200 & _T_201; // @[dec_decode_ctl.scala 318:28]
  assign io_dec_nonblock_load_waddr = _T_246 | _T_238; // @[dec_decode_ctl.scala 315:29 dec_decode_ctl.scala 325:29]
  assign io_dec_pause_state = pause_stall; // @[dec_decode_ctl.scala 462:22]
  assign io_dec_pause_state_cg = pause_stall & _T_423; // @[dec_decode_ctl.scala 466:25]
  assign io_dec_div_active = _T_826; // @[dec_decode_ctl.scala 699:21]
  assign rvclkhdr_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_io_en = _T_15 | _T_16; // @[lib.scala 345:16]
  assign rvclkhdr_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign i0_dec_io_ins = io_dec_i0_instr_d; // @[dec_decode_ctl.scala 357:16]
  assign rvclkhdr_1_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_1_io_en = i0_pipe_en[3] | io_clk_override; // @[lib.scala 371:17]
  assign rvclkhdr_1_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_2_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_2_io_en = i0_pipe_en[3] | io_clk_override; // @[lib.scala 371:17]
  assign rvclkhdr_2_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_3_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_3_io_en = _T_431 | pause_stall; // @[lib.scala 371:17]
  assign rvclkhdr_3_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_4_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_4_io_en = shift_illegal & _T_467; // @[lib.scala 371:17]
  assign rvclkhdr_4_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_5_io_clk = clock; // @[lib.scala 380:18]
  assign rvclkhdr_5_io_en = _T_709 | io_clk_override; // @[lib.scala 381:17]
  assign rvclkhdr_5_io_scan_mode = io_scan_mode; // @[lib.scala 382:24]
  assign rvclkhdr_6_io_clk = clock; // @[lib.scala 380:18]
  assign rvclkhdr_6_io_en = _T_709 | io_clk_override; // @[lib.scala 381:17]
  assign rvclkhdr_6_io_scan_mode = io_scan_mode; // @[lib.scala 382:24]
  assign rvclkhdr_7_io_clk = clock; // @[lib.scala 380:18]
  assign rvclkhdr_7_io_en = _T_709 | io_clk_override; // @[lib.scala 381:17]
  assign rvclkhdr_7_io_scan_mode = io_scan_mode; // @[lib.scala 382:24]
  assign rvclkhdr_8_io_clk = clock; // @[lib.scala 380:18]
  assign rvclkhdr_8_io_en = _T_712 | io_clk_override; // @[lib.scala 381:17]
  assign rvclkhdr_8_io_scan_mode = io_scan_mode; // @[lib.scala 382:24]
  assign rvclkhdr_9_io_clk = clock; // @[lib.scala 380:18]
  assign rvclkhdr_9_io_en = _T_715 | io_clk_override; // @[lib.scala 381:17]
  assign rvclkhdr_9_io_scan_mode = io_scan_mode; // @[lib.scala 382:24]
  assign rvclkhdr_10_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_10_io_en = i0_pipe_en[2] | io_clk_override; // @[lib.scala 371:17]
  assign rvclkhdr_10_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_11_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_11_io_en = i0_pipe_en[3] | io_clk_override; // @[lib.scala 371:17]
  assign rvclkhdr_11_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_12_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_12_io_en = i0_legal_decode_d & i0_dp_div; // @[lib.scala 371:17]
  assign rvclkhdr_12_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_13_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_13_io_en = i0_pipe_en[3] | io_clk_override; // @[lib.scala 371:17]
  assign rvclkhdr_13_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_14_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_14_io_en = i0_pipe_en[2] | io_clk_override; // @[lib.scala 371:17]
  assign rvclkhdr_14_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_15_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_15_io_en = i0_pipe_en[1] | io_clk_override; // @[lib.scala 371:17]
  assign rvclkhdr_15_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_16_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_16_io_en = i0_pipe_en[0] | io_clk_override; // @[lib.scala 371:17]
  assign rvclkhdr_16_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_17_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_17_io_en = i0_pipe_en[1] | io_clk_override; // @[lib.scala 371:17]
  assign rvclkhdr_17_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_18_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_18_io_en = i0_pipe_en[0] | io_clk_override; // @[lib.scala 371:17]
  assign rvclkhdr_18_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_19_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_19_io_en = i0_pipe_en[2] | io_clk_override; // @[lib.scala 371:17]
  assign rvclkhdr_19_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  tlu_wr_pause_r1 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  tlu_wr_pause_r2 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  leak1_i1_stall = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  leak1_i0_stall = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  pause_stall = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  write_csr_data = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  postsync_stall = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  x_d_valid = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  flush_final_r = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  illegal_lockout = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  cam_raw_0_bits_tag = _RAND_10[2:0];
  _RAND_11 = {1{`RANDOM}};
  cam_raw_0_valid = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  cam_raw_1_bits_tag = _RAND_12[2:0];
  _RAND_13 = {1{`RANDOM}};
  cam_raw_1_valid = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  cam_raw_2_bits_tag = _RAND_14[2:0];
  _RAND_15 = {1{`RANDOM}};
  cam_raw_2_valid = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  cam_raw_3_bits_tag = _RAND_16[2:0];
  _RAND_17 = {1{`RANDOM}};
  cam_raw_3_valid = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  x_d_bits_i0load = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  x_d_bits_i0rd = _RAND_19[4:0];
  _RAND_20 = {1{`RANDOM}};
  _T_706 = _RAND_20[2:0];
  _RAND_21 = {1{`RANDOM}};
  nonblock_load_valid_m_delay = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  r_d_bits_i0load = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  r_d_bits_i0v = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  r_d_bits_i0rd = _RAND_24[4:0];
  _RAND_25 = {1{`RANDOM}};
  cam_raw_0_bits_rd = _RAND_25[4:0];
  _RAND_26 = {1{`RANDOM}};
  cam_raw_0_bits_wb = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  cam_raw_1_bits_rd = _RAND_27[4:0];
  _RAND_28 = {1{`RANDOM}};
  cam_raw_1_bits_wb = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  cam_raw_2_bits_rd = _RAND_29[4:0];
  _RAND_30 = {1{`RANDOM}};
  cam_raw_2_bits_wb = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  cam_raw_3_bits_rd = _RAND_31[4:0];
  _RAND_32 = {1{`RANDOM}};
  cam_raw_3_bits_wb = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  lsu_idle = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  _T_339 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  x_d_bits_i0v = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  i0_x_c_load = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  i0_r_c_load = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  r_d_bits_csrwen = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  r_d_valid = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  r_d_bits_csrwaddr = _RAND_40[11:0];
  _RAND_41 = {1{`RANDOM}};
  csr_read_x = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  csr_clr_x = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  csr_set_x = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  csr_write_x = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  csr_imm_x = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  csrimm_x = _RAND_46[4:0];
  _RAND_47 = {1{`RANDOM}};
  csr_rddata_x = _RAND_47[31:0];
  _RAND_48 = {1{`RANDOM}};
  r_d_bits_csrwonly = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  i0_result_r_raw = _RAND_49[31:0];
  _RAND_50 = {1{`RANDOM}};
  x_d_bits_csrwonly = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  wbd_bits_csrwonly = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  _T_468 = _RAND_52[31:0];
  _RAND_53 = {1{`RANDOM}};
  x_t_legal = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  x_t_icaf = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  x_t_icaf_f1 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  x_t_icaf_type = _RAND_56[1:0];
  _RAND_57 = {1{`RANDOM}};
  x_t_fence_i = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  x_t_i0trigger = _RAND_58[3:0];
  _RAND_59 = {1{`RANDOM}};
  x_t_pmu_i0_itype = _RAND_59[3:0];
  _RAND_60 = {1{`RANDOM}};
  x_t_pmu_i0_br_unpred = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  r_t_legal = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  r_t_icaf = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  r_t_icaf_f1 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  r_t_icaf_type = _RAND_64[1:0];
  _RAND_65 = {1{`RANDOM}};
  r_t_fence_i = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  r_t_i0trigger = _RAND_66[3:0];
  _RAND_67 = {1{`RANDOM}};
  r_t_pmu_i0_itype = _RAND_67[3:0];
  _RAND_68 = {1{`RANDOM}};
  r_t_pmu_i0_br_unpred = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  lsu_trigger_match_r = _RAND_69[3:0];
  _RAND_70 = {1{`RANDOM}};
  lsu_pmu_misaligned_r = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  r_d_bits_i0store = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  r_d_bits_i0div = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  i0_x_c_mul = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  i0_x_c_alu = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  i0_r_c_mul = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  i0_r_c_alu = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  x_d_bits_i0store = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  x_d_bits_i0div = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  x_d_bits_csrwen = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  x_d_bits_csrwaddr = _RAND_80[11:0];
  _RAND_81 = {1{`RANDOM}};
  last_br_immed_x = _RAND_81[11:0];
  _RAND_82 = {1{`RANDOM}};
  _T_826 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  _T_835 = _RAND_83[4:0];
  _RAND_84 = {1{`RANDOM}};
  i0_inst_x = _RAND_84[31:0];
  _RAND_85 = {1{`RANDOM}};
  i0_inst_r = _RAND_85[31:0];
  _RAND_86 = {1{`RANDOM}};
  i0_inst_wb = _RAND_86[31:0];
  _RAND_87 = {1{`RANDOM}};
  _T_842 = _RAND_87[31:0];
  _RAND_88 = {1{`RANDOM}};
  i0_pc_wb = _RAND_88[30:0];
  _RAND_89 = {1{`RANDOM}};
  _T_845 = _RAND_89[30:0];
  _RAND_90 = {1{`RANDOM}};
  dec_i0_pc_r = _RAND_90[30:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    tlu_wr_pause_r1 = 1'h0;
  end
  if (reset) begin
    tlu_wr_pause_r2 = 1'h0;
  end
  if (reset) begin
    leak1_i1_stall = 1'h0;
  end
  if (reset) begin
    leak1_i0_stall = 1'h0;
  end
  if (reset) begin
    pause_stall = 1'h0;
  end
  if (reset) begin
    write_csr_data = 32'h0;
  end
  if (reset) begin
    postsync_stall = 1'h0;
  end
  if (reset) begin
    x_d_valid = 1'h0;
  end
  if (reset) begin
    flush_final_r = 1'h0;
  end
  if (reset) begin
    illegal_lockout = 1'h0;
  end
  if (reset) begin
    cam_raw_0_bits_tag = 3'h0;
  end
  if (reset) begin
    cam_raw_0_valid = 1'h0;
  end
  if (reset) begin
    cam_raw_1_bits_tag = 3'h0;
  end
  if (reset) begin
    cam_raw_1_valid = 1'h0;
  end
  if (reset) begin
    cam_raw_2_bits_tag = 3'h0;
  end
  if (reset) begin
    cam_raw_2_valid = 1'h0;
  end
  if (reset) begin
    cam_raw_3_bits_tag = 3'h0;
  end
  if (reset) begin
    cam_raw_3_valid = 1'h0;
  end
  if (reset) begin
    x_d_bits_i0load = 1'h0;
  end
  if (reset) begin
    x_d_bits_i0rd = 5'h0;
  end
  if (reset) begin
    _T_706 = 3'h0;
  end
  if (reset) begin
    nonblock_load_valid_m_delay = 1'h0;
  end
  if (reset) begin
    r_d_bits_i0load = 1'h0;
  end
  if (reset) begin
    r_d_bits_i0v = 1'h0;
  end
  if (reset) begin
    r_d_bits_i0rd = 5'h0;
  end
  if (reset) begin
    cam_raw_0_bits_rd = 5'h0;
  end
  if (reset) begin
    cam_raw_0_bits_wb = 1'h0;
  end
  if (reset) begin
    cam_raw_1_bits_rd = 5'h0;
  end
  if (reset) begin
    cam_raw_1_bits_wb = 1'h0;
  end
  if (reset) begin
    cam_raw_2_bits_rd = 5'h0;
  end
  if (reset) begin
    cam_raw_2_bits_wb = 1'h0;
  end
  if (reset) begin
    cam_raw_3_bits_rd = 5'h0;
  end
  if (reset) begin
    cam_raw_3_bits_wb = 1'h0;
  end
  if (reset) begin
    lsu_idle = 1'h0;
  end
  if (reset) begin
    _T_339 = 1'h0;
  end
  if (reset) begin
    x_d_bits_i0v = 1'h0;
  end
  if (reset) begin
    i0_x_c_load = 1'h0;
  end
  if (reset) begin
    i0_r_c_load = 1'h0;
  end
  if (reset) begin
    r_d_bits_csrwen = 1'h0;
  end
  if (reset) begin
    r_d_valid = 1'h0;
  end
  if (reset) begin
    r_d_bits_csrwaddr = 12'h0;
  end
  if (reset) begin
    csr_read_x = 1'h0;
  end
  if (reset) begin
    csr_clr_x = 1'h0;
  end
  if (reset) begin
    csr_set_x = 1'h0;
  end
  if (reset) begin
    csr_write_x = 1'h0;
  end
  if (reset) begin
    csr_imm_x = 1'h0;
  end
  if (reset) begin
    csrimm_x = 5'h0;
  end
  if (reset) begin
    csr_rddata_x = 32'h0;
  end
  if (reset) begin
    r_d_bits_csrwonly = 1'h0;
  end
  if (reset) begin
    i0_result_r_raw = 32'h0;
  end
  if (reset) begin
    x_d_bits_csrwonly = 1'h0;
  end
  if (reset) begin
    wbd_bits_csrwonly = 1'h0;
  end
  if (reset) begin
    _T_468 = 32'h0;
  end
  if (reset) begin
    x_t_legal = 1'h0;
  end
  if (reset) begin
    x_t_icaf = 1'h0;
  end
  if (reset) begin
    x_t_icaf_f1 = 1'h0;
  end
  if (reset) begin
    x_t_icaf_type = 2'h0;
  end
  if (reset) begin
    x_t_fence_i = 1'h0;
  end
  if (reset) begin
    x_t_i0trigger = 4'h0;
  end
  if (reset) begin
    x_t_pmu_i0_itype = 4'h0;
  end
  if (reset) begin
    x_t_pmu_i0_br_unpred = 1'h0;
  end
  if (reset) begin
    r_t_legal = 1'h0;
  end
  if (reset) begin
    r_t_icaf = 1'h0;
  end
  if (reset) begin
    r_t_icaf_f1 = 1'h0;
  end
  if (reset) begin
    r_t_icaf_type = 2'h0;
  end
  if (reset) begin
    r_t_fence_i = 1'h0;
  end
  if (reset) begin
    r_t_i0trigger = 4'h0;
  end
  if (reset) begin
    r_t_pmu_i0_itype = 4'h0;
  end
  if (reset) begin
    r_t_pmu_i0_br_unpred = 1'h0;
  end
  if (reset) begin
    lsu_trigger_match_r = 4'h0;
  end
  if (reset) begin
    lsu_pmu_misaligned_r = 1'h0;
  end
  if (reset) begin
    r_d_bits_i0store = 1'h0;
  end
  if (reset) begin
    r_d_bits_i0div = 1'h0;
  end
  if (reset) begin
    i0_x_c_mul = 1'h0;
  end
  if (reset) begin
    i0_x_c_alu = 1'h0;
  end
  if (reset) begin
    i0_r_c_mul = 1'h0;
  end
  if (reset) begin
    i0_r_c_alu = 1'h0;
  end
  if (reset) begin
    x_d_bits_i0store = 1'h0;
  end
  if (reset) begin
    x_d_bits_i0div = 1'h0;
  end
  if (reset) begin
    x_d_bits_csrwen = 1'h0;
  end
  if (reset) begin
    x_d_bits_csrwaddr = 12'h0;
  end
  if (reset) begin
    last_br_immed_x = 12'h0;
  end
  if (reset) begin
    _T_826 = 1'h0;
  end
  if (reset) begin
    _T_835 = 5'h0;
  end
  if (reset) begin
    i0_inst_x = 32'h0;
  end
  if (reset) begin
    i0_inst_r = 32'h0;
  end
  if (reset) begin
    i0_inst_wb = 32'h0;
  end
  if (reset) begin
    _T_842 = 32'h0;
  end
  if (reset) begin
    i0_pc_wb = 31'h0;
  end
  if (reset) begin
    _T_845 = 31'h0;
  end
  if (reset) begin
    dec_i0_pc_r = 31'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge rvclkhdr_io_l1clk or posedge reset) begin
    if (reset) begin
      tlu_wr_pause_r1 <= 1'h0;
    end else begin
      tlu_wr_pause_r1 <= io_dec_tlu_wr_pause_r;
    end
  end
  always @(posedge rvclkhdr_io_l1clk or posedge reset) begin
    if (reset) begin
      tlu_wr_pause_r2 <= 1'h0;
    end else begin
      tlu_wr_pause_r2 <= tlu_wr_pause_r1;
    end
  end
  always @(posedge rvclkhdr_io_l1clk or posedge reset) begin
    if (reset) begin
      leak1_i1_stall <= 1'h0;
    end else begin
      leak1_i1_stall <= io_dec_tlu_flush_leak_one_r | _T_281;
    end
  end
  always @(posedge rvclkhdr_io_l1clk or posedge reset) begin
    if (reset) begin
      leak1_i0_stall <= 1'h0;
    end else begin
      leak1_i0_stall <= _T_284 | _T_286;
    end
  end
  always @(posedge rvclkhdr_io_l1clk or posedge reset) begin
    if (reset) begin
      pause_stall <= 1'h0;
    end else begin
      pause_stall <= _T_415 & _T_416;
    end
  end
  always @(posedge rvclkhdr_3_io_l1clk or posedge reset) begin
    if (reset) begin
      write_csr_data <= 32'h0;
    end else if (pause_stall) begin
      write_csr_data <= _T_426;
    end else if (io_dec_tlu_wr_pause_r) begin
      write_csr_data <= io_dec_csr_wrdata_r;
    end else begin
      write_csr_data <= write_csr_data_x;
    end
  end
  always @(posedge rvclkhdr_io_l1clk or posedge reset) begin
    if (reset) begin
      postsync_stall <= 1'h0;
    end else begin
      postsync_stall <= _T_509 | _T_510;
    end
  end
  always @(posedge rvclkhdr_7_io_l1clk or posedge reset) begin
    if (reset) begin
      x_d_valid <= 1'h0;
    end else begin
      x_d_valid <= io_dec_aln_dec_i0_decode_d;
    end
  end
  always @(posedge rvclkhdr_io_l1clk or posedge reset) begin
    if (reset) begin
      flush_final_r <= 1'h0;
    end else begin
      flush_final_r <= io_exu_flush_final;
    end
  end
  always @(posedge rvclkhdr_io_l1clk or posedge reset) begin
    if (reset) begin
      illegal_lockout <= 1'h0;
    end else begin
      illegal_lockout <= _T_469 & _T_470;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      cam_raw_0_bits_tag <= 3'h0;
    end else if (cam_wen[0]) begin
      cam_raw_0_bits_tag <= {{1'd0}, io_dctl_busbuff_lsu_nonblock_load_tag_m};
    end else if (_T_107) begin
      cam_raw_0_bits_tag <= 3'h0;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      cam_raw_0_valid <= 1'h0;
    end else if (io_dec_tlu_force_halt) begin
      cam_raw_0_valid <= 1'h0;
    end else begin
      cam_raw_0_valid <= _GEN_56;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      cam_raw_1_bits_tag <= 3'h0;
    end else if (cam_wen[1]) begin
      cam_raw_1_bits_tag <= {{1'd0}, io_dctl_busbuff_lsu_nonblock_load_tag_m};
    end else if (_T_133) begin
      cam_raw_1_bits_tag <= 3'h0;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      cam_raw_1_valid <= 1'h0;
    end else if (io_dec_tlu_force_halt) begin
      cam_raw_1_valid <= 1'h0;
    end else begin
      cam_raw_1_valid <= _GEN_67;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      cam_raw_2_bits_tag <= 3'h0;
    end else if (cam_wen[2]) begin
      cam_raw_2_bits_tag <= {{1'd0}, io_dctl_busbuff_lsu_nonblock_load_tag_m};
    end else if (_T_159) begin
      cam_raw_2_bits_tag <= 3'h0;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      cam_raw_2_valid <= 1'h0;
    end else if (io_dec_tlu_force_halt) begin
      cam_raw_2_valid <= 1'h0;
    end else begin
      cam_raw_2_valid <= _GEN_78;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      cam_raw_3_bits_tag <= 3'h0;
    end else if (cam_wen[3]) begin
      cam_raw_3_bits_tag <= {{1'd0}, io_dctl_busbuff_lsu_nonblock_load_tag_m};
    end else if (_T_185) begin
      cam_raw_3_bits_tag <= 3'h0;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      cam_raw_3_valid <= 1'h0;
    end else if (io_dec_tlu_force_halt) begin
      cam_raw_3_valid <= 1'h0;
    end else begin
      cam_raw_3_valid <= _GEN_89;
    end
  end
  always @(posedge rvclkhdr_7_io_l1clk or posedge reset) begin
    if (reset) begin
      x_d_bits_i0load <= 1'h0;
    end else begin
      x_d_bits_i0load <= i0_dp_load & i0_legal_decode_d;
    end
  end
  always @(posedge rvclkhdr_7_io_l1clk or posedge reset) begin
    if (reset) begin
      x_d_bits_i0rd <= 5'h0;
    end else begin
      x_d_bits_i0rd <= io_dec_i0_instr_d[11:7];
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      _T_706 <= 3'h0;
    end else begin
      _T_706 <= i0_pipe_en[3:1];
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      nonblock_load_valid_m_delay <= 1'h0;
    end else if (i0_r_ctl_en) begin
      nonblock_load_valid_m_delay <= io_dctl_busbuff_lsu_nonblock_load_valid_m;
    end
  end
  always @(posedge rvclkhdr_8_io_l1clk or posedge reset) begin
    if (reset) begin
      r_d_bits_i0load <= 1'h0;
    end else begin
      r_d_bits_i0load <= x_d_bits_i0load;
    end
  end
  always @(posedge rvclkhdr_8_io_l1clk or posedge reset) begin
    if (reset) begin
      r_d_bits_i0v <= 1'h0;
    end else begin
      r_d_bits_i0v <= _T_738 & _T_280;
    end
  end
  always @(posedge rvclkhdr_8_io_l1clk or posedge reset) begin
    if (reset) begin
      r_d_bits_i0rd <= 5'h0;
    end else begin
      r_d_bits_i0rd <= x_d_bits_i0rd;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      cam_raw_0_bits_rd <= 5'h0;
    end else if (cam_wen[0]) begin
      if (x_d_bits_i0load) begin
        cam_raw_0_bits_rd <= x_d_bits_i0rd;
      end else begin
        cam_raw_0_bits_rd <= 5'h0;
      end
    end else if (_T_107) begin
      cam_raw_0_bits_rd <= 5'h0;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      cam_raw_0_bits_wb <= 1'h0;
    end else begin
      cam_raw_0_bits_wb <= _T_112 | _GEN_57;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      cam_raw_1_bits_rd <= 5'h0;
    end else if (cam_wen[1]) begin
      if (x_d_bits_i0load) begin
        cam_raw_1_bits_rd <= x_d_bits_i0rd;
      end else begin
        cam_raw_1_bits_rd <= 5'h0;
      end
    end else if (_T_133) begin
      cam_raw_1_bits_rd <= 5'h0;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      cam_raw_1_bits_wb <= 1'h0;
    end else begin
      cam_raw_1_bits_wb <= _T_138 | _GEN_68;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      cam_raw_2_bits_rd <= 5'h0;
    end else if (cam_wen[2]) begin
      if (x_d_bits_i0load) begin
        cam_raw_2_bits_rd <= x_d_bits_i0rd;
      end else begin
        cam_raw_2_bits_rd <= 5'h0;
      end
    end else if (_T_159) begin
      cam_raw_2_bits_rd <= 5'h0;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      cam_raw_2_bits_wb <= 1'h0;
    end else begin
      cam_raw_2_bits_wb <= _T_164 | _GEN_79;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      cam_raw_3_bits_rd <= 5'h0;
    end else if (cam_wen[3]) begin
      if (x_d_bits_i0load) begin
        cam_raw_3_bits_rd <= x_d_bits_i0rd;
      end else begin
        cam_raw_3_bits_rd <= 5'h0;
      end
    end else if (_T_185) begin
      cam_raw_3_bits_rd <= 5'h0;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      cam_raw_3_bits_wb <= 1'h0;
    end else begin
      cam_raw_3_bits_wb <= _T_190 | _GEN_90;
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      lsu_idle <= 1'h0;
    end else begin
      lsu_idle <= io_lsu_idle_any;
    end
  end
  always @(posedge rvclkhdr_io_l1clk or posedge reset) begin
    if (reset) begin
      _T_339 <= 1'h0;
    end else begin
      _T_339 <= io_dec_tlu_flush_extint;
    end
  end
  always @(posedge rvclkhdr_7_io_l1clk or posedge reset) begin
    if (reset) begin
      x_d_bits_i0v <= 1'h0;
    end else begin
      x_d_bits_i0v <= i0_rd_en_d & i0_legal_decode_d;
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      i0_x_c_load <= 1'h0;
    end else if (i0_x_ctl_en) begin
      i0_x_c_load <= i0_d_c_load;
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      i0_r_c_load <= 1'h0;
    end else if (i0_r_ctl_en) begin
      i0_r_c_load <= i0_x_c_load;
    end
  end
  always @(posedge rvclkhdr_8_io_l1clk or posedge reset) begin
    if (reset) begin
      r_d_bits_csrwen <= 1'h0;
    end else begin
      r_d_bits_csrwen <= x_d_bits_csrwen;
    end
  end
  always @(posedge rvclkhdr_8_io_l1clk or posedge reset) begin
    if (reset) begin
      r_d_valid <= 1'h0;
    end else begin
      r_d_valid <= _T_742 & _T_280;
    end
  end
  always @(posedge rvclkhdr_8_io_l1clk or posedge reset) begin
    if (reset) begin
      r_d_bits_csrwaddr <= 12'h0;
    end else begin
      r_d_bits_csrwaddr <= x_d_bits_csrwaddr;
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      csr_read_x <= 1'h0;
    end else begin
      csr_read_x <= i0_dp_csr_read & i0_legal_decode_d;
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      csr_clr_x <= 1'h0;
    end else begin
      csr_clr_x <= i0_dp_csr_clr & i0_legal_decode_d;
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      csr_set_x <= 1'h0;
    end else begin
      csr_set_x <= i0_dp_csr_set & i0_legal_decode_d;
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      csr_write_x <= 1'h0;
    end else begin
      csr_write_x <= i0_csr_write & i0_legal_decode_d;
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      csr_imm_x <= 1'h0;
    end else if (_T_41) begin
      csr_imm_x <= 1'h0;
    end else begin
      csr_imm_x <= i0_dp_raw_csr_imm;
    end
  end
  always @(posedge rvclkhdr_1_io_l1clk or posedge reset) begin
    if (reset) begin
      csrimm_x <= 5'h0;
    end else begin
      csrimm_x <= io_dec_i0_instr_d[19:15];
    end
  end
  always @(posedge rvclkhdr_2_io_l1clk or posedge reset) begin
    if (reset) begin
      csr_rddata_x <= 32'h0;
    end else begin
      csr_rddata_x <= io_dec_csr_rddata_d;
    end
  end
  always @(posedge rvclkhdr_8_io_l1clk or posedge reset) begin
    if (reset) begin
      r_d_bits_csrwonly <= 1'h0;
    end else begin
      r_d_bits_csrwonly <= x_d_bits_csrwonly;
    end
  end
  always @(posedge rvclkhdr_10_io_l1clk or posedge reset) begin
    if (reset) begin
      i0_result_r_raw <= 32'h0;
    end else if (_T_766) begin
      i0_result_r_raw <= io_lsu_result_m;
    end else begin
      i0_result_r_raw <= io_decode_exu_exu_i0_result_x;
    end
  end
  always @(posedge rvclkhdr_7_io_l1clk or posedge reset) begin
    if (reset) begin
      x_d_bits_csrwonly <= 1'h0;
    end else begin
      x_d_bits_csrwonly <= i0_csr_write_only_d & io_dec_aln_dec_i0_decode_d;
    end
  end
  always @(posedge rvclkhdr_9_io_l1clk or posedge reset) begin
    if (reset) begin
      wbd_bits_csrwonly <= 1'h0;
    end else begin
      wbd_bits_csrwonly <= r_d_bits_csrwonly;
    end
  end
  always @(posedge rvclkhdr_4_io_l1clk or posedge reset) begin
    if (reset) begin
      _T_468 <= 32'h0;
    end else if (io_dec_i0_pc4_d) begin
      _T_468 <= io_dec_i0_instr_d;
    end else begin
      _T_468 <= _T_465;
    end
  end
  always @(posedge rvclkhdr_5_io_l1clk or posedge reset) begin
    if (reset) begin
      x_t_legal <= 1'h0;
    end else begin
      x_t_legal <= io_dec_aln_dec_i0_decode_d & i0_legal;
    end
  end
  always @(posedge rvclkhdr_5_io_l1clk or posedge reset) begin
    if (reset) begin
      x_t_icaf <= 1'h0;
    end else begin
      x_t_icaf <= i0_icaf_d & i0_legal_decode_d;
    end
  end
  always @(posedge rvclkhdr_5_io_l1clk or posedge reset) begin
    if (reset) begin
      x_t_icaf_f1 <= 1'h0;
    end else begin
      x_t_icaf_f1 <= io_dec_i0_icaf_f1_d & i0_legal_decode_d;
    end
  end
  always @(posedge rvclkhdr_5_io_l1clk or posedge reset) begin
    if (reset) begin
      x_t_icaf_type <= 2'h0;
    end else begin
      x_t_icaf_type <= io_dec_i0_icaf_type_d;
    end
  end
  always @(posedge rvclkhdr_5_io_l1clk or posedge reset) begin
    if (reset) begin
      x_t_fence_i <= 1'h0;
    end else begin
      x_t_fence_i <= _T_520 & i0_legal_decode_d;
    end
  end
  always @(posedge rvclkhdr_5_io_l1clk or posedge reset) begin
    if (reset) begin
      x_t_i0trigger <= 4'h0;
    end else begin
      x_t_i0trigger <= io_dec_i0_trigger_match_d & _T_525;
    end
  end
  always @(posedge rvclkhdr_5_io_l1clk or posedge reset) begin
    if (reset) begin
      x_t_pmu_i0_itype <= 4'h0;
    end else begin
      x_t_pmu_i0_itype <= _T_255 & _T_277;
    end
  end
  always @(posedge rvclkhdr_5_io_l1clk or posedge reset) begin
    if (reset) begin
      x_t_pmu_i0_br_unpred <= 1'h0;
    end else begin
      x_t_pmu_i0_br_unpred <= i0_dp_jal & _T_253;
    end
  end
  always @(posedge rvclkhdr_6_io_l1clk or posedge reset) begin
    if (reset) begin
      r_t_legal <= 1'h0;
    end else begin
      r_t_legal <= x_t_legal;
    end
  end
  always @(posedge rvclkhdr_6_io_l1clk or posedge reset) begin
    if (reset) begin
      r_t_icaf <= 1'h0;
    end else begin
      r_t_icaf <= x_t_icaf;
    end
  end
  always @(posedge rvclkhdr_6_io_l1clk or posedge reset) begin
    if (reset) begin
      r_t_icaf_f1 <= 1'h0;
    end else begin
      r_t_icaf_f1 <= x_t_icaf_f1;
    end
  end
  always @(posedge rvclkhdr_6_io_l1clk or posedge reset) begin
    if (reset) begin
      r_t_icaf_type <= 2'h0;
    end else begin
      r_t_icaf_type <= x_t_icaf_type;
    end
  end
  always @(posedge rvclkhdr_6_io_l1clk or posedge reset) begin
    if (reset) begin
      r_t_fence_i <= 1'h0;
    end else begin
      r_t_fence_i <= x_t_fence_i;
    end
  end
  always @(posedge rvclkhdr_6_io_l1clk or posedge reset) begin
    if (reset) begin
      r_t_i0trigger <= 4'h0;
    end else begin
      r_t_i0trigger <= x_t_i0trigger & _T_534;
    end
  end
  always @(posedge rvclkhdr_6_io_l1clk or posedge reset) begin
    if (reset) begin
      r_t_pmu_i0_itype <= 4'h0;
    end else begin
      r_t_pmu_i0_itype <= x_t_pmu_i0_itype;
    end
  end
  always @(posedge rvclkhdr_6_io_l1clk or posedge reset) begin
    if (reset) begin
      r_t_pmu_i0_br_unpred <= 1'h0;
    end else begin
      r_t_pmu_i0_br_unpred <= x_t_pmu_i0_br_unpred;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      lsu_trigger_match_r <= 4'h0;
    end else begin
      lsu_trigger_match_r <= io_lsu_trigger_match_m;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      lsu_pmu_misaligned_r <= 1'h0;
    end else begin
      lsu_pmu_misaligned_r <= io_lsu_pmu_misaligned_m;
    end
  end
  always @(posedge rvclkhdr_8_io_l1clk or posedge reset) begin
    if (reset) begin
      r_d_bits_i0store <= 1'h0;
    end else begin
      r_d_bits_i0store <= x_d_bits_i0store;
    end
  end
  always @(posedge rvclkhdr_8_io_l1clk or posedge reset) begin
    if (reset) begin
      r_d_bits_i0div <= 1'h0;
    end else begin
      r_d_bits_i0div <= x_d_bits_i0div;
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      i0_x_c_mul <= 1'h0;
    end else if (i0_x_ctl_en) begin
      i0_x_c_mul <= i0_d_c_mul;
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      i0_x_c_alu <= 1'h0;
    end else if (i0_x_ctl_en) begin
      i0_x_c_alu <= i0_d_c_alu;
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      i0_r_c_mul <= 1'h0;
    end else if (i0_r_ctl_en) begin
      i0_r_c_mul <= i0_x_c_mul;
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      i0_r_c_alu <= 1'h0;
    end else if (i0_r_ctl_en) begin
      i0_r_c_alu <= i0_x_c_alu;
    end
  end
  always @(posedge rvclkhdr_7_io_l1clk or posedge reset) begin
    if (reset) begin
      x_d_bits_i0store <= 1'h0;
    end else begin
      x_d_bits_i0store <= i0_dp_store & i0_legal_decode_d;
    end
  end
  always @(posedge rvclkhdr_7_io_l1clk or posedge reset) begin
    if (reset) begin
      x_d_bits_i0div <= 1'h0;
    end else begin
      x_d_bits_i0div <= i0_dp_div & i0_legal_decode_d;
    end
  end
  always @(posedge rvclkhdr_7_io_l1clk or posedge reset) begin
    if (reset) begin
      x_d_bits_csrwen <= 1'h0;
    end else begin
      x_d_bits_csrwen <= io_dec_csr_wen_unq_d & i0_legal_decode_d;
    end
  end
  always @(posedge rvclkhdr_7_io_l1clk or posedge reset) begin
    if (reset) begin
      x_d_bits_csrwaddr <= 12'h0;
    end else begin
      x_d_bits_csrwaddr <= io_dec_i0_instr_d[31:20];
    end
  end
  always @(posedge rvclkhdr_11_io_l1clk or posedge reset) begin
    if (reset) begin
      last_br_immed_x <= 12'h0;
    end else if (io_decode_exu_i0_ap_predict_nt) begin
      last_br_immed_x <= _T_786;
    end else if (_T_314) begin
      last_br_immed_x <= i0_pcall_imm[11:0];
    end else begin
      last_br_immed_x <= _T_323;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      _T_826 <= 1'h0;
    end else begin
      _T_826 <= i0_div_decode_d | _T_825;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_835 <= 5'h0;
    end else if (i0_div_decode_d) begin
      _T_835 <= i0r_rd;
    end
  end
  always @(posedge rvclkhdr_13_io_l1clk or posedge reset) begin
    if (reset) begin
      i0_inst_x <= 32'h0;
    end else if (io_dec_i0_pc4_d) begin
      i0_inst_x <= io_dec_i0_instr_d;
    end else begin
      i0_inst_x <= _T_465;
    end
  end
  always @(posedge rvclkhdr_14_io_l1clk or posedge reset) begin
    if (reset) begin
      i0_inst_r <= 32'h0;
    end else begin
      i0_inst_r <= i0_inst_x;
    end
  end
  always @(posedge rvclkhdr_15_io_l1clk or posedge reset) begin
    if (reset) begin
      i0_inst_wb <= 32'h0;
    end else begin
      i0_inst_wb <= i0_inst_r;
    end
  end
  always @(posedge rvclkhdr_16_io_l1clk or posedge reset) begin
    if (reset) begin
      _T_842 <= 32'h0;
    end else begin
      _T_842 <= i0_inst_wb;
    end
  end
  always @(posedge rvclkhdr_17_io_l1clk or posedge reset) begin
    if (reset) begin
      i0_pc_wb <= 31'h0;
    end else begin
      i0_pc_wb <= io_dec_tlu_i0_pc_r;
    end
  end
  always @(posedge rvclkhdr_18_io_l1clk or posedge reset) begin
    if (reset) begin
      _T_845 <= 31'h0;
    end else begin
      _T_845 <= i0_pc_wb;
    end
  end
  always @(posedge rvclkhdr_19_io_l1clk or posedge reset) begin
    if (reset) begin
      dec_i0_pc_r <= 31'h0;
    end else begin
      dec_i0_pc_r <= io_dec_alu_exu_i0_pc_x;
    end
  end
endmodule
module dec_gpr_ctl(
  input         clock,
  input         reset,
  input  [4:0]  io_raddr0,
  input  [4:0]  io_raddr1,
  input         io_wen0,
  input  [4:0]  io_waddr0,
  input  [31:0] io_wd0,
  input         io_wen1,
  input  [4:0]  io_waddr1,
  input  [31:0] io_wd1,
  input         io_wen2,
  input  [4:0]  io_waddr2,
  input  [31:0] io_wd2,
  input         io_scan_mode,
  output [31:0] io_gpr_exu_gpr_i0_rs1_d,
  output [31:0] io_gpr_exu_gpr_i0_rs2_d
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
`endif // RANDOMIZE_REG_INIT
  wire  rvclkhdr_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_1_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_1_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_1_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_1_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_2_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_2_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_2_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_2_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_3_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_3_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_3_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_3_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_4_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_4_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_4_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_4_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_5_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_5_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_5_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_5_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_6_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_6_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_6_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_6_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_7_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_7_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_7_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_7_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_8_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_8_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_8_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_8_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_9_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_9_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_9_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_9_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_10_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_10_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_10_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_10_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_11_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_11_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_11_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_11_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_12_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_12_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_12_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_12_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_13_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_13_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_13_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_13_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_14_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_14_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_14_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_14_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_15_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_15_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_15_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_15_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_16_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_16_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_16_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_16_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_17_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_17_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_17_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_17_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_18_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_18_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_18_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_18_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_19_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_19_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_19_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_19_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_20_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_20_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_20_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_20_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_21_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_21_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_21_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_21_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_22_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_22_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_22_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_22_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_23_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_23_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_23_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_23_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_24_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_24_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_24_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_24_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_25_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_25_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_25_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_25_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_26_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_26_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_26_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_26_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_27_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_27_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_27_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_27_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_28_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_28_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_28_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_28_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_29_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_29_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_29_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_29_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_30_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_30_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_30_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_30_io_scan_mode; // @[lib.scala 368:23]
  wire  _T = io_waddr0 == 5'h1; // @[dec_gpr_ctl.scala 52:45]
  wire  w0v_1 = io_wen0 & _T; // @[dec_gpr_ctl.scala 52:33]
  wire  _T_2 = io_waddr1 == 5'h1; // @[dec_gpr_ctl.scala 53:45]
  wire  w1v_1 = io_wen1 & _T_2; // @[dec_gpr_ctl.scala 53:33]
  wire  _T_4 = io_waddr2 == 5'h1; // @[dec_gpr_ctl.scala 54:45]
  wire  w2v_1 = io_wen2 & _T_4; // @[dec_gpr_ctl.scala 54:33]
  wire [31:0] _T_7 = w0v_1 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_8 = _T_7 & io_wd0; // @[dec_gpr_ctl.scala 55:42]
  wire [31:0] _T_10 = w1v_1 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_11 = _T_10 & io_wd1; // @[dec_gpr_ctl.scala 55:71]
  wire [31:0] _T_12 = _T_8 | _T_11; // @[dec_gpr_ctl.scala 55:52]
  wire [31:0] _T_14 = w2v_1 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_15 = _T_14 & io_wd2; // @[dec_gpr_ctl.scala 55:100]
  wire  _T_17 = io_waddr0 == 5'h2; // @[dec_gpr_ctl.scala 52:45]
  wire  w0v_2 = io_wen0 & _T_17; // @[dec_gpr_ctl.scala 52:33]
  wire  _T_19 = io_waddr1 == 5'h2; // @[dec_gpr_ctl.scala 53:45]
  wire  w1v_2 = io_wen1 & _T_19; // @[dec_gpr_ctl.scala 53:33]
  wire  _T_21 = io_waddr2 == 5'h2; // @[dec_gpr_ctl.scala 54:45]
  wire  w2v_2 = io_wen2 & _T_21; // @[dec_gpr_ctl.scala 54:33]
  wire [31:0] _T_24 = w0v_2 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_25 = _T_24 & io_wd0; // @[dec_gpr_ctl.scala 55:42]
  wire [31:0] _T_27 = w1v_2 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_28 = _T_27 & io_wd1; // @[dec_gpr_ctl.scala 55:71]
  wire [31:0] _T_29 = _T_25 | _T_28; // @[dec_gpr_ctl.scala 55:52]
  wire [31:0] _T_31 = w2v_2 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_32 = _T_31 & io_wd2; // @[dec_gpr_ctl.scala 55:100]
  wire  _T_34 = io_waddr0 == 5'h3; // @[dec_gpr_ctl.scala 52:45]
  wire  w0v_3 = io_wen0 & _T_34; // @[dec_gpr_ctl.scala 52:33]
  wire  _T_36 = io_waddr1 == 5'h3; // @[dec_gpr_ctl.scala 53:45]
  wire  w1v_3 = io_wen1 & _T_36; // @[dec_gpr_ctl.scala 53:33]
  wire  _T_38 = io_waddr2 == 5'h3; // @[dec_gpr_ctl.scala 54:45]
  wire  w2v_3 = io_wen2 & _T_38; // @[dec_gpr_ctl.scala 54:33]
  wire [31:0] _T_41 = w0v_3 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_42 = _T_41 & io_wd0; // @[dec_gpr_ctl.scala 55:42]
  wire [31:0] _T_44 = w1v_3 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_45 = _T_44 & io_wd1; // @[dec_gpr_ctl.scala 55:71]
  wire [31:0] _T_46 = _T_42 | _T_45; // @[dec_gpr_ctl.scala 55:52]
  wire [31:0] _T_48 = w2v_3 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_49 = _T_48 & io_wd2; // @[dec_gpr_ctl.scala 55:100]
  wire  _T_51 = io_waddr0 == 5'h4; // @[dec_gpr_ctl.scala 52:45]
  wire  w0v_4 = io_wen0 & _T_51; // @[dec_gpr_ctl.scala 52:33]
  wire  _T_53 = io_waddr1 == 5'h4; // @[dec_gpr_ctl.scala 53:45]
  wire  w1v_4 = io_wen1 & _T_53; // @[dec_gpr_ctl.scala 53:33]
  wire  _T_55 = io_waddr2 == 5'h4; // @[dec_gpr_ctl.scala 54:45]
  wire  w2v_4 = io_wen2 & _T_55; // @[dec_gpr_ctl.scala 54:33]
  wire [31:0] _T_58 = w0v_4 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_59 = _T_58 & io_wd0; // @[dec_gpr_ctl.scala 55:42]
  wire [31:0] _T_61 = w1v_4 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_62 = _T_61 & io_wd1; // @[dec_gpr_ctl.scala 55:71]
  wire [31:0] _T_63 = _T_59 | _T_62; // @[dec_gpr_ctl.scala 55:52]
  wire [31:0] _T_65 = w2v_4 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_66 = _T_65 & io_wd2; // @[dec_gpr_ctl.scala 55:100]
  wire  _T_68 = io_waddr0 == 5'h5; // @[dec_gpr_ctl.scala 52:45]
  wire  w0v_5 = io_wen0 & _T_68; // @[dec_gpr_ctl.scala 52:33]
  wire  _T_70 = io_waddr1 == 5'h5; // @[dec_gpr_ctl.scala 53:45]
  wire  w1v_5 = io_wen1 & _T_70; // @[dec_gpr_ctl.scala 53:33]
  wire  _T_72 = io_waddr2 == 5'h5; // @[dec_gpr_ctl.scala 54:45]
  wire  w2v_5 = io_wen2 & _T_72; // @[dec_gpr_ctl.scala 54:33]
  wire [31:0] _T_75 = w0v_5 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_76 = _T_75 & io_wd0; // @[dec_gpr_ctl.scala 55:42]
  wire [31:0] _T_78 = w1v_5 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_79 = _T_78 & io_wd1; // @[dec_gpr_ctl.scala 55:71]
  wire [31:0] _T_80 = _T_76 | _T_79; // @[dec_gpr_ctl.scala 55:52]
  wire [31:0] _T_82 = w2v_5 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_83 = _T_82 & io_wd2; // @[dec_gpr_ctl.scala 55:100]
  wire  _T_85 = io_waddr0 == 5'h6; // @[dec_gpr_ctl.scala 52:45]
  wire  w0v_6 = io_wen0 & _T_85; // @[dec_gpr_ctl.scala 52:33]
  wire  _T_87 = io_waddr1 == 5'h6; // @[dec_gpr_ctl.scala 53:45]
  wire  w1v_6 = io_wen1 & _T_87; // @[dec_gpr_ctl.scala 53:33]
  wire  _T_89 = io_waddr2 == 5'h6; // @[dec_gpr_ctl.scala 54:45]
  wire  w2v_6 = io_wen2 & _T_89; // @[dec_gpr_ctl.scala 54:33]
  wire [31:0] _T_92 = w0v_6 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_93 = _T_92 & io_wd0; // @[dec_gpr_ctl.scala 55:42]
  wire [31:0] _T_95 = w1v_6 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_96 = _T_95 & io_wd1; // @[dec_gpr_ctl.scala 55:71]
  wire [31:0] _T_97 = _T_93 | _T_96; // @[dec_gpr_ctl.scala 55:52]
  wire [31:0] _T_99 = w2v_6 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_100 = _T_99 & io_wd2; // @[dec_gpr_ctl.scala 55:100]
  wire  _T_102 = io_waddr0 == 5'h7; // @[dec_gpr_ctl.scala 52:45]
  wire  w0v_7 = io_wen0 & _T_102; // @[dec_gpr_ctl.scala 52:33]
  wire  _T_104 = io_waddr1 == 5'h7; // @[dec_gpr_ctl.scala 53:45]
  wire  w1v_7 = io_wen1 & _T_104; // @[dec_gpr_ctl.scala 53:33]
  wire  _T_106 = io_waddr2 == 5'h7; // @[dec_gpr_ctl.scala 54:45]
  wire  w2v_7 = io_wen2 & _T_106; // @[dec_gpr_ctl.scala 54:33]
  wire [31:0] _T_109 = w0v_7 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_110 = _T_109 & io_wd0; // @[dec_gpr_ctl.scala 55:42]
  wire [31:0] _T_112 = w1v_7 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_113 = _T_112 & io_wd1; // @[dec_gpr_ctl.scala 55:71]
  wire [31:0] _T_114 = _T_110 | _T_113; // @[dec_gpr_ctl.scala 55:52]
  wire [31:0] _T_116 = w2v_7 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_117 = _T_116 & io_wd2; // @[dec_gpr_ctl.scala 55:100]
  wire  _T_119 = io_waddr0 == 5'h8; // @[dec_gpr_ctl.scala 52:45]
  wire  w0v_8 = io_wen0 & _T_119; // @[dec_gpr_ctl.scala 52:33]
  wire  _T_121 = io_waddr1 == 5'h8; // @[dec_gpr_ctl.scala 53:45]
  wire  w1v_8 = io_wen1 & _T_121; // @[dec_gpr_ctl.scala 53:33]
  wire  _T_123 = io_waddr2 == 5'h8; // @[dec_gpr_ctl.scala 54:45]
  wire  w2v_8 = io_wen2 & _T_123; // @[dec_gpr_ctl.scala 54:33]
  wire [31:0] _T_126 = w0v_8 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_127 = _T_126 & io_wd0; // @[dec_gpr_ctl.scala 55:42]
  wire [31:0] _T_129 = w1v_8 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_130 = _T_129 & io_wd1; // @[dec_gpr_ctl.scala 55:71]
  wire [31:0] _T_131 = _T_127 | _T_130; // @[dec_gpr_ctl.scala 55:52]
  wire [31:0] _T_133 = w2v_8 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_134 = _T_133 & io_wd2; // @[dec_gpr_ctl.scala 55:100]
  wire  _T_136 = io_waddr0 == 5'h9; // @[dec_gpr_ctl.scala 52:45]
  wire  w0v_9 = io_wen0 & _T_136; // @[dec_gpr_ctl.scala 52:33]
  wire  _T_138 = io_waddr1 == 5'h9; // @[dec_gpr_ctl.scala 53:45]
  wire  w1v_9 = io_wen1 & _T_138; // @[dec_gpr_ctl.scala 53:33]
  wire  _T_140 = io_waddr2 == 5'h9; // @[dec_gpr_ctl.scala 54:45]
  wire  w2v_9 = io_wen2 & _T_140; // @[dec_gpr_ctl.scala 54:33]
  wire [31:0] _T_143 = w0v_9 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_144 = _T_143 & io_wd0; // @[dec_gpr_ctl.scala 55:42]
  wire [31:0] _T_146 = w1v_9 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_147 = _T_146 & io_wd1; // @[dec_gpr_ctl.scala 55:71]
  wire [31:0] _T_148 = _T_144 | _T_147; // @[dec_gpr_ctl.scala 55:52]
  wire [31:0] _T_150 = w2v_9 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_151 = _T_150 & io_wd2; // @[dec_gpr_ctl.scala 55:100]
  wire  _T_153 = io_waddr0 == 5'ha; // @[dec_gpr_ctl.scala 52:45]
  wire  w0v_10 = io_wen0 & _T_153; // @[dec_gpr_ctl.scala 52:33]
  wire  _T_155 = io_waddr1 == 5'ha; // @[dec_gpr_ctl.scala 53:45]
  wire  w1v_10 = io_wen1 & _T_155; // @[dec_gpr_ctl.scala 53:33]
  wire  _T_157 = io_waddr2 == 5'ha; // @[dec_gpr_ctl.scala 54:45]
  wire  w2v_10 = io_wen2 & _T_157; // @[dec_gpr_ctl.scala 54:33]
  wire [31:0] _T_160 = w0v_10 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_161 = _T_160 & io_wd0; // @[dec_gpr_ctl.scala 55:42]
  wire [31:0] _T_163 = w1v_10 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_164 = _T_163 & io_wd1; // @[dec_gpr_ctl.scala 55:71]
  wire [31:0] _T_165 = _T_161 | _T_164; // @[dec_gpr_ctl.scala 55:52]
  wire [31:0] _T_167 = w2v_10 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_168 = _T_167 & io_wd2; // @[dec_gpr_ctl.scala 55:100]
  wire  _T_170 = io_waddr0 == 5'hb; // @[dec_gpr_ctl.scala 52:45]
  wire  w0v_11 = io_wen0 & _T_170; // @[dec_gpr_ctl.scala 52:33]
  wire  _T_172 = io_waddr1 == 5'hb; // @[dec_gpr_ctl.scala 53:45]
  wire  w1v_11 = io_wen1 & _T_172; // @[dec_gpr_ctl.scala 53:33]
  wire  _T_174 = io_waddr2 == 5'hb; // @[dec_gpr_ctl.scala 54:45]
  wire  w2v_11 = io_wen2 & _T_174; // @[dec_gpr_ctl.scala 54:33]
  wire [31:0] _T_177 = w0v_11 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_178 = _T_177 & io_wd0; // @[dec_gpr_ctl.scala 55:42]
  wire [31:0] _T_180 = w1v_11 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_181 = _T_180 & io_wd1; // @[dec_gpr_ctl.scala 55:71]
  wire [31:0] _T_182 = _T_178 | _T_181; // @[dec_gpr_ctl.scala 55:52]
  wire [31:0] _T_184 = w2v_11 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_185 = _T_184 & io_wd2; // @[dec_gpr_ctl.scala 55:100]
  wire  _T_187 = io_waddr0 == 5'hc; // @[dec_gpr_ctl.scala 52:45]
  wire  w0v_12 = io_wen0 & _T_187; // @[dec_gpr_ctl.scala 52:33]
  wire  _T_189 = io_waddr1 == 5'hc; // @[dec_gpr_ctl.scala 53:45]
  wire  w1v_12 = io_wen1 & _T_189; // @[dec_gpr_ctl.scala 53:33]
  wire  _T_191 = io_waddr2 == 5'hc; // @[dec_gpr_ctl.scala 54:45]
  wire  w2v_12 = io_wen2 & _T_191; // @[dec_gpr_ctl.scala 54:33]
  wire [31:0] _T_194 = w0v_12 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_195 = _T_194 & io_wd0; // @[dec_gpr_ctl.scala 55:42]
  wire [31:0] _T_197 = w1v_12 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_198 = _T_197 & io_wd1; // @[dec_gpr_ctl.scala 55:71]
  wire [31:0] _T_199 = _T_195 | _T_198; // @[dec_gpr_ctl.scala 55:52]
  wire [31:0] _T_201 = w2v_12 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_202 = _T_201 & io_wd2; // @[dec_gpr_ctl.scala 55:100]
  wire  _T_204 = io_waddr0 == 5'hd; // @[dec_gpr_ctl.scala 52:45]
  wire  w0v_13 = io_wen0 & _T_204; // @[dec_gpr_ctl.scala 52:33]
  wire  _T_206 = io_waddr1 == 5'hd; // @[dec_gpr_ctl.scala 53:45]
  wire  w1v_13 = io_wen1 & _T_206; // @[dec_gpr_ctl.scala 53:33]
  wire  _T_208 = io_waddr2 == 5'hd; // @[dec_gpr_ctl.scala 54:45]
  wire  w2v_13 = io_wen2 & _T_208; // @[dec_gpr_ctl.scala 54:33]
  wire [31:0] _T_211 = w0v_13 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_212 = _T_211 & io_wd0; // @[dec_gpr_ctl.scala 55:42]
  wire [31:0] _T_214 = w1v_13 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_215 = _T_214 & io_wd1; // @[dec_gpr_ctl.scala 55:71]
  wire [31:0] _T_216 = _T_212 | _T_215; // @[dec_gpr_ctl.scala 55:52]
  wire [31:0] _T_218 = w2v_13 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_219 = _T_218 & io_wd2; // @[dec_gpr_ctl.scala 55:100]
  wire  _T_221 = io_waddr0 == 5'he; // @[dec_gpr_ctl.scala 52:45]
  wire  w0v_14 = io_wen0 & _T_221; // @[dec_gpr_ctl.scala 52:33]
  wire  _T_223 = io_waddr1 == 5'he; // @[dec_gpr_ctl.scala 53:45]
  wire  w1v_14 = io_wen1 & _T_223; // @[dec_gpr_ctl.scala 53:33]
  wire  _T_225 = io_waddr2 == 5'he; // @[dec_gpr_ctl.scala 54:45]
  wire  w2v_14 = io_wen2 & _T_225; // @[dec_gpr_ctl.scala 54:33]
  wire [31:0] _T_228 = w0v_14 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_229 = _T_228 & io_wd0; // @[dec_gpr_ctl.scala 55:42]
  wire [31:0] _T_231 = w1v_14 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_232 = _T_231 & io_wd1; // @[dec_gpr_ctl.scala 55:71]
  wire [31:0] _T_233 = _T_229 | _T_232; // @[dec_gpr_ctl.scala 55:52]
  wire [31:0] _T_235 = w2v_14 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_236 = _T_235 & io_wd2; // @[dec_gpr_ctl.scala 55:100]
  wire  _T_238 = io_waddr0 == 5'hf; // @[dec_gpr_ctl.scala 52:45]
  wire  w0v_15 = io_wen0 & _T_238; // @[dec_gpr_ctl.scala 52:33]
  wire  _T_240 = io_waddr1 == 5'hf; // @[dec_gpr_ctl.scala 53:45]
  wire  w1v_15 = io_wen1 & _T_240; // @[dec_gpr_ctl.scala 53:33]
  wire  _T_242 = io_waddr2 == 5'hf; // @[dec_gpr_ctl.scala 54:45]
  wire  w2v_15 = io_wen2 & _T_242; // @[dec_gpr_ctl.scala 54:33]
  wire [31:0] _T_245 = w0v_15 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_246 = _T_245 & io_wd0; // @[dec_gpr_ctl.scala 55:42]
  wire [31:0] _T_248 = w1v_15 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_249 = _T_248 & io_wd1; // @[dec_gpr_ctl.scala 55:71]
  wire [31:0] _T_250 = _T_246 | _T_249; // @[dec_gpr_ctl.scala 55:52]
  wire [31:0] _T_252 = w2v_15 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_253 = _T_252 & io_wd2; // @[dec_gpr_ctl.scala 55:100]
  wire  _T_255 = io_waddr0 == 5'h10; // @[dec_gpr_ctl.scala 52:45]
  wire  w0v_16 = io_wen0 & _T_255; // @[dec_gpr_ctl.scala 52:33]
  wire  _T_257 = io_waddr1 == 5'h10; // @[dec_gpr_ctl.scala 53:45]
  wire  w1v_16 = io_wen1 & _T_257; // @[dec_gpr_ctl.scala 53:33]
  wire  _T_259 = io_waddr2 == 5'h10; // @[dec_gpr_ctl.scala 54:45]
  wire  w2v_16 = io_wen2 & _T_259; // @[dec_gpr_ctl.scala 54:33]
  wire [31:0] _T_262 = w0v_16 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_263 = _T_262 & io_wd0; // @[dec_gpr_ctl.scala 55:42]
  wire [31:0] _T_265 = w1v_16 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_266 = _T_265 & io_wd1; // @[dec_gpr_ctl.scala 55:71]
  wire [31:0] _T_267 = _T_263 | _T_266; // @[dec_gpr_ctl.scala 55:52]
  wire [31:0] _T_269 = w2v_16 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_270 = _T_269 & io_wd2; // @[dec_gpr_ctl.scala 55:100]
  wire  _T_272 = io_waddr0 == 5'h11; // @[dec_gpr_ctl.scala 52:45]
  wire  w0v_17 = io_wen0 & _T_272; // @[dec_gpr_ctl.scala 52:33]
  wire  _T_274 = io_waddr1 == 5'h11; // @[dec_gpr_ctl.scala 53:45]
  wire  w1v_17 = io_wen1 & _T_274; // @[dec_gpr_ctl.scala 53:33]
  wire  _T_276 = io_waddr2 == 5'h11; // @[dec_gpr_ctl.scala 54:45]
  wire  w2v_17 = io_wen2 & _T_276; // @[dec_gpr_ctl.scala 54:33]
  wire [31:0] _T_279 = w0v_17 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_280 = _T_279 & io_wd0; // @[dec_gpr_ctl.scala 55:42]
  wire [31:0] _T_282 = w1v_17 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_283 = _T_282 & io_wd1; // @[dec_gpr_ctl.scala 55:71]
  wire [31:0] _T_284 = _T_280 | _T_283; // @[dec_gpr_ctl.scala 55:52]
  wire [31:0] _T_286 = w2v_17 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_287 = _T_286 & io_wd2; // @[dec_gpr_ctl.scala 55:100]
  wire  _T_289 = io_waddr0 == 5'h12; // @[dec_gpr_ctl.scala 52:45]
  wire  w0v_18 = io_wen0 & _T_289; // @[dec_gpr_ctl.scala 52:33]
  wire  _T_291 = io_waddr1 == 5'h12; // @[dec_gpr_ctl.scala 53:45]
  wire  w1v_18 = io_wen1 & _T_291; // @[dec_gpr_ctl.scala 53:33]
  wire  _T_293 = io_waddr2 == 5'h12; // @[dec_gpr_ctl.scala 54:45]
  wire  w2v_18 = io_wen2 & _T_293; // @[dec_gpr_ctl.scala 54:33]
  wire [31:0] _T_296 = w0v_18 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_297 = _T_296 & io_wd0; // @[dec_gpr_ctl.scala 55:42]
  wire [31:0] _T_299 = w1v_18 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_300 = _T_299 & io_wd1; // @[dec_gpr_ctl.scala 55:71]
  wire [31:0] _T_301 = _T_297 | _T_300; // @[dec_gpr_ctl.scala 55:52]
  wire [31:0] _T_303 = w2v_18 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_304 = _T_303 & io_wd2; // @[dec_gpr_ctl.scala 55:100]
  wire  _T_306 = io_waddr0 == 5'h13; // @[dec_gpr_ctl.scala 52:45]
  wire  w0v_19 = io_wen0 & _T_306; // @[dec_gpr_ctl.scala 52:33]
  wire  _T_308 = io_waddr1 == 5'h13; // @[dec_gpr_ctl.scala 53:45]
  wire  w1v_19 = io_wen1 & _T_308; // @[dec_gpr_ctl.scala 53:33]
  wire  _T_310 = io_waddr2 == 5'h13; // @[dec_gpr_ctl.scala 54:45]
  wire  w2v_19 = io_wen2 & _T_310; // @[dec_gpr_ctl.scala 54:33]
  wire [31:0] _T_313 = w0v_19 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_314 = _T_313 & io_wd0; // @[dec_gpr_ctl.scala 55:42]
  wire [31:0] _T_316 = w1v_19 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_317 = _T_316 & io_wd1; // @[dec_gpr_ctl.scala 55:71]
  wire [31:0] _T_318 = _T_314 | _T_317; // @[dec_gpr_ctl.scala 55:52]
  wire [31:0] _T_320 = w2v_19 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_321 = _T_320 & io_wd2; // @[dec_gpr_ctl.scala 55:100]
  wire  _T_323 = io_waddr0 == 5'h14; // @[dec_gpr_ctl.scala 52:45]
  wire  w0v_20 = io_wen0 & _T_323; // @[dec_gpr_ctl.scala 52:33]
  wire  _T_325 = io_waddr1 == 5'h14; // @[dec_gpr_ctl.scala 53:45]
  wire  w1v_20 = io_wen1 & _T_325; // @[dec_gpr_ctl.scala 53:33]
  wire  _T_327 = io_waddr2 == 5'h14; // @[dec_gpr_ctl.scala 54:45]
  wire  w2v_20 = io_wen2 & _T_327; // @[dec_gpr_ctl.scala 54:33]
  wire [31:0] _T_330 = w0v_20 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_331 = _T_330 & io_wd0; // @[dec_gpr_ctl.scala 55:42]
  wire [31:0] _T_333 = w1v_20 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_334 = _T_333 & io_wd1; // @[dec_gpr_ctl.scala 55:71]
  wire [31:0] _T_335 = _T_331 | _T_334; // @[dec_gpr_ctl.scala 55:52]
  wire [31:0] _T_337 = w2v_20 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_338 = _T_337 & io_wd2; // @[dec_gpr_ctl.scala 55:100]
  wire  _T_340 = io_waddr0 == 5'h15; // @[dec_gpr_ctl.scala 52:45]
  wire  w0v_21 = io_wen0 & _T_340; // @[dec_gpr_ctl.scala 52:33]
  wire  _T_342 = io_waddr1 == 5'h15; // @[dec_gpr_ctl.scala 53:45]
  wire  w1v_21 = io_wen1 & _T_342; // @[dec_gpr_ctl.scala 53:33]
  wire  _T_344 = io_waddr2 == 5'h15; // @[dec_gpr_ctl.scala 54:45]
  wire  w2v_21 = io_wen2 & _T_344; // @[dec_gpr_ctl.scala 54:33]
  wire [31:0] _T_347 = w0v_21 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_348 = _T_347 & io_wd0; // @[dec_gpr_ctl.scala 55:42]
  wire [31:0] _T_350 = w1v_21 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_351 = _T_350 & io_wd1; // @[dec_gpr_ctl.scala 55:71]
  wire [31:0] _T_352 = _T_348 | _T_351; // @[dec_gpr_ctl.scala 55:52]
  wire [31:0] _T_354 = w2v_21 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_355 = _T_354 & io_wd2; // @[dec_gpr_ctl.scala 55:100]
  wire  _T_357 = io_waddr0 == 5'h16; // @[dec_gpr_ctl.scala 52:45]
  wire  w0v_22 = io_wen0 & _T_357; // @[dec_gpr_ctl.scala 52:33]
  wire  _T_359 = io_waddr1 == 5'h16; // @[dec_gpr_ctl.scala 53:45]
  wire  w1v_22 = io_wen1 & _T_359; // @[dec_gpr_ctl.scala 53:33]
  wire  _T_361 = io_waddr2 == 5'h16; // @[dec_gpr_ctl.scala 54:45]
  wire  w2v_22 = io_wen2 & _T_361; // @[dec_gpr_ctl.scala 54:33]
  wire [31:0] _T_364 = w0v_22 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_365 = _T_364 & io_wd0; // @[dec_gpr_ctl.scala 55:42]
  wire [31:0] _T_367 = w1v_22 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_368 = _T_367 & io_wd1; // @[dec_gpr_ctl.scala 55:71]
  wire [31:0] _T_369 = _T_365 | _T_368; // @[dec_gpr_ctl.scala 55:52]
  wire [31:0] _T_371 = w2v_22 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_372 = _T_371 & io_wd2; // @[dec_gpr_ctl.scala 55:100]
  wire  _T_374 = io_waddr0 == 5'h17; // @[dec_gpr_ctl.scala 52:45]
  wire  w0v_23 = io_wen0 & _T_374; // @[dec_gpr_ctl.scala 52:33]
  wire  _T_376 = io_waddr1 == 5'h17; // @[dec_gpr_ctl.scala 53:45]
  wire  w1v_23 = io_wen1 & _T_376; // @[dec_gpr_ctl.scala 53:33]
  wire  _T_378 = io_waddr2 == 5'h17; // @[dec_gpr_ctl.scala 54:45]
  wire  w2v_23 = io_wen2 & _T_378; // @[dec_gpr_ctl.scala 54:33]
  wire [31:0] _T_381 = w0v_23 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_382 = _T_381 & io_wd0; // @[dec_gpr_ctl.scala 55:42]
  wire [31:0] _T_384 = w1v_23 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_385 = _T_384 & io_wd1; // @[dec_gpr_ctl.scala 55:71]
  wire [31:0] _T_386 = _T_382 | _T_385; // @[dec_gpr_ctl.scala 55:52]
  wire [31:0] _T_388 = w2v_23 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_389 = _T_388 & io_wd2; // @[dec_gpr_ctl.scala 55:100]
  wire  _T_391 = io_waddr0 == 5'h18; // @[dec_gpr_ctl.scala 52:45]
  wire  w0v_24 = io_wen0 & _T_391; // @[dec_gpr_ctl.scala 52:33]
  wire  _T_393 = io_waddr1 == 5'h18; // @[dec_gpr_ctl.scala 53:45]
  wire  w1v_24 = io_wen1 & _T_393; // @[dec_gpr_ctl.scala 53:33]
  wire  _T_395 = io_waddr2 == 5'h18; // @[dec_gpr_ctl.scala 54:45]
  wire  w2v_24 = io_wen2 & _T_395; // @[dec_gpr_ctl.scala 54:33]
  wire [31:0] _T_398 = w0v_24 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_399 = _T_398 & io_wd0; // @[dec_gpr_ctl.scala 55:42]
  wire [31:0] _T_401 = w1v_24 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_402 = _T_401 & io_wd1; // @[dec_gpr_ctl.scala 55:71]
  wire [31:0] _T_403 = _T_399 | _T_402; // @[dec_gpr_ctl.scala 55:52]
  wire [31:0] _T_405 = w2v_24 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_406 = _T_405 & io_wd2; // @[dec_gpr_ctl.scala 55:100]
  wire  _T_408 = io_waddr0 == 5'h19; // @[dec_gpr_ctl.scala 52:45]
  wire  w0v_25 = io_wen0 & _T_408; // @[dec_gpr_ctl.scala 52:33]
  wire  _T_410 = io_waddr1 == 5'h19; // @[dec_gpr_ctl.scala 53:45]
  wire  w1v_25 = io_wen1 & _T_410; // @[dec_gpr_ctl.scala 53:33]
  wire  _T_412 = io_waddr2 == 5'h19; // @[dec_gpr_ctl.scala 54:45]
  wire  w2v_25 = io_wen2 & _T_412; // @[dec_gpr_ctl.scala 54:33]
  wire [31:0] _T_415 = w0v_25 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_416 = _T_415 & io_wd0; // @[dec_gpr_ctl.scala 55:42]
  wire [31:0] _T_418 = w1v_25 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_419 = _T_418 & io_wd1; // @[dec_gpr_ctl.scala 55:71]
  wire [31:0] _T_420 = _T_416 | _T_419; // @[dec_gpr_ctl.scala 55:52]
  wire [31:0] _T_422 = w2v_25 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_423 = _T_422 & io_wd2; // @[dec_gpr_ctl.scala 55:100]
  wire  _T_425 = io_waddr0 == 5'h1a; // @[dec_gpr_ctl.scala 52:45]
  wire  w0v_26 = io_wen0 & _T_425; // @[dec_gpr_ctl.scala 52:33]
  wire  _T_427 = io_waddr1 == 5'h1a; // @[dec_gpr_ctl.scala 53:45]
  wire  w1v_26 = io_wen1 & _T_427; // @[dec_gpr_ctl.scala 53:33]
  wire  _T_429 = io_waddr2 == 5'h1a; // @[dec_gpr_ctl.scala 54:45]
  wire  w2v_26 = io_wen2 & _T_429; // @[dec_gpr_ctl.scala 54:33]
  wire [31:0] _T_432 = w0v_26 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_433 = _T_432 & io_wd0; // @[dec_gpr_ctl.scala 55:42]
  wire [31:0] _T_435 = w1v_26 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_436 = _T_435 & io_wd1; // @[dec_gpr_ctl.scala 55:71]
  wire [31:0] _T_437 = _T_433 | _T_436; // @[dec_gpr_ctl.scala 55:52]
  wire [31:0] _T_439 = w2v_26 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_440 = _T_439 & io_wd2; // @[dec_gpr_ctl.scala 55:100]
  wire  _T_442 = io_waddr0 == 5'h1b; // @[dec_gpr_ctl.scala 52:45]
  wire  w0v_27 = io_wen0 & _T_442; // @[dec_gpr_ctl.scala 52:33]
  wire  _T_444 = io_waddr1 == 5'h1b; // @[dec_gpr_ctl.scala 53:45]
  wire  w1v_27 = io_wen1 & _T_444; // @[dec_gpr_ctl.scala 53:33]
  wire  _T_446 = io_waddr2 == 5'h1b; // @[dec_gpr_ctl.scala 54:45]
  wire  w2v_27 = io_wen2 & _T_446; // @[dec_gpr_ctl.scala 54:33]
  wire [31:0] _T_449 = w0v_27 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_450 = _T_449 & io_wd0; // @[dec_gpr_ctl.scala 55:42]
  wire [31:0] _T_452 = w1v_27 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_453 = _T_452 & io_wd1; // @[dec_gpr_ctl.scala 55:71]
  wire [31:0] _T_454 = _T_450 | _T_453; // @[dec_gpr_ctl.scala 55:52]
  wire [31:0] _T_456 = w2v_27 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_457 = _T_456 & io_wd2; // @[dec_gpr_ctl.scala 55:100]
  wire  _T_459 = io_waddr0 == 5'h1c; // @[dec_gpr_ctl.scala 52:45]
  wire  w0v_28 = io_wen0 & _T_459; // @[dec_gpr_ctl.scala 52:33]
  wire  _T_461 = io_waddr1 == 5'h1c; // @[dec_gpr_ctl.scala 53:45]
  wire  w1v_28 = io_wen1 & _T_461; // @[dec_gpr_ctl.scala 53:33]
  wire  _T_463 = io_waddr2 == 5'h1c; // @[dec_gpr_ctl.scala 54:45]
  wire  w2v_28 = io_wen2 & _T_463; // @[dec_gpr_ctl.scala 54:33]
  wire [31:0] _T_466 = w0v_28 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_467 = _T_466 & io_wd0; // @[dec_gpr_ctl.scala 55:42]
  wire [31:0] _T_469 = w1v_28 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_470 = _T_469 & io_wd1; // @[dec_gpr_ctl.scala 55:71]
  wire [31:0] _T_471 = _T_467 | _T_470; // @[dec_gpr_ctl.scala 55:52]
  wire [31:0] _T_473 = w2v_28 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_474 = _T_473 & io_wd2; // @[dec_gpr_ctl.scala 55:100]
  wire  _T_476 = io_waddr0 == 5'h1d; // @[dec_gpr_ctl.scala 52:45]
  wire  w0v_29 = io_wen0 & _T_476; // @[dec_gpr_ctl.scala 52:33]
  wire  _T_478 = io_waddr1 == 5'h1d; // @[dec_gpr_ctl.scala 53:45]
  wire  w1v_29 = io_wen1 & _T_478; // @[dec_gpr_ctl.scala 53:33]
  wire  _T_480 = io_waddr2 == 5'h1d; // @[dec_gpr_ctl.scala 54:45]
  wire  w2v_29 = io_wen2 & _T_480; // @[dec_gpr_ctl.scala 54:33]
  wire [31:0] _T_483 = w0v_29 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_484 = _T_483 & io_wd0; // @[dec_gpr_ctl.scala 55:42]
  wire [31:0] _T_486 = w1v_29 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_487 = _T_486 & io_wd1; // @[dec_gpr_ctl.scala 55:71]
  wire [31:0] _T_488 = _T_484 | _T_487; // @[dec_gpr_ctl.scala 55:52]
  wire [31:0] _T_490 = w2v_29 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_491 = _T_490 & io_wd2; // @[dec_gpr_ctl.scala 55:100]
  wire  _T_493 = io_waddr0 == 5'h1e; // @[dec_gpr_ctl.scala 52:45]
  wire  w0v_30 = io_wen0 & _T_493; // @[dec_gpr_ctl.scala 52:33]
  wire  _T_495 = io_waddr1 == 5'h1e; // @[dec_gpr_ctl.scala 53:45]
  wire  w1v_30 = io_wen1 & _T_495; // @[dec_gpr_ctl.scala 53:33]
  wire  _T_497 = io_waddr2 == 5'h1e; // @[dec_gpr_ctl.scala 54:45]
  wire  w2v_30 = io_wen2 & _T_497; // @[dec_gpr_ctl.scala 54:33]
  wire [31:0] _T_500 = w0v_30 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_501 = _T_500 & io_wd0; // @[dec_gpr_ctl.scala 55:42]
  wire [31:0] _T_503 = w1v_30 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_504 = _T_503 & io_wd1; // @[dec_gpr_ctl.scala 55:71]
  wire [31:0] _T_505 = _T_501 | _T_504; // @[dec_gpr_ctl.scala 55:52]
  wire [31:0] _T_507 = w2v_30 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_508 = _T_507 & io_wd2; // @[dec_gpr_ctl.scala 55:100]
  wire  _T_510 = io_waddr0 == 5'h1f; // @[dec_gpr_ctl.scala 52:45]
  wire  w0v_31 = io_wen0 & _T_510; // @[dec_gpr_ctl.scala 52:33]
  wire  _T_512 = io_waddr1 == 5'h1f; // @[dec_gpr_ctl.scala 53:45]
  wire  w1v_31 = io_wen1 & _T_512; // @[dec_gpr_ctl.scala 53:33]
  wire  _T_514 = io_waddr2 == 5'h1f; // @[dec_gpr_ctl.scala 54:45]
  wire  w2v_31 = io_wen2 & _T_514; // @[dec_gpr_ctl.scala 54:33]
  wire [31:0] _T_517 = w0v_31 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_518 = _T_517 & io_wd0; // @[dec_gpr_ctl.scala 55:42]
  wire [31:0] _T_520 = w1v_31 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_521 = _T_520 & io_wd1; // @[dec_gpr_ctl.scala 55:71]
  wire [31:0] _T_522 = _T_518 | _T_521; // @[dec_gpr_ctl.scala 55:52]
  wire [31:0] _T_524 = w2v_31 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_525 = _T_524 & io_wd2; // @[dec_gpr_ctl.scala 55:100]
  wire [9:0] _T_535 = {w0v_9,w0v_8,w0v_7,w0v_6,w0v_5,w0v_4,w0v_3,w0v_2,w0v_1,1'h0}; // @[Cat.scala 29:58]
  wire [18:0] _T_544 = {w0v_18,w0v_17,w0v_16,w0v_15,w0v_14,w0v_13,w0v_12,w0v_11,w0v_10,_T_535}; // @[Cat.scala 29:58]
  wire [27:0] _T_553 = {w0v_27,w0v_26,w0v_25,w0v_24,w0v_23,w0v_22,w0v_21,w0v_20,w0v_19,_T_544}; // @[Cat.scala 29:58]
  wire [31:0] _T_557 = {w0v_31,w0v_30,w0v_29,w0v_28,_T_553}; // @[Cat.scala 29:58]
  wire [9:0] _T_566 = {w1v_9,w1v_8,w1v_7,w1v_6,w1v_5,w1v_4,w1v_3,w1v_2,w1v_1,1'h0}; // @[Cat.scala 29:58]
  wire [18:0] _T_575 = {w1v_18,w1v_17,w1v_16,w1v_15,w1v_14,w1v_13,w1v_12,w1v_11,w1v_10,_T_566}; // @[Cat.scala 29:58]
  wire [27:0] _T_584 = {w1v_27,w1v_26,w1v_25,w1v_24,w1v_23,w1v_22,w1v_21,w1v_20,w1v_19,_T_575}; // @[Cat.scala 29:58]
  wire [31:0] _T_588 = {w1v_31,w1v_30,w1v_29,w1v_28,_T_584}; // @[Cat.scala 29:58]
  wire [31:0] _T_589 = _T_557 | _T_588; // @[dec_gpr_ctl.scala 57:57]
  wire [9:0] _T_598 = {w2v_9,w2v_8,w2v_7,w2v_6,w2v_5,w2v_4,w2v_3,w2v_2,w2v_1,1'h0}; // @[Cat.scala 29:58]
  wire [18:0] _T_607 = {w2v_18,w2v_17,w2v_16,w2v_15,w2v_14,w2v_13,w2v_12,w2v_11,w2v_10,_T_598}; // @[Cat.scala 29:58]
  wire [27:0] _T_616 = {w2v_27,w2v_26,w2v_25,w2v_24,w2v_23,w2v_22,w2v_21,w2v_20,w2v_19,_T_607}; // @[Cat.scala 29:58]
  wire [31:0] _T_620 = {w2v_31,w2v_30,w2v_29,w2v_28,_T_616}; // @[Cat.scala 29:58]
  wire [31:0] gpr_wr_en = _T_589 | _T_620; // @[dec_gpr_ctl.scala 57:95]
  reg [31:0] gpr_out_1; // @[lib.scala 374:16]
  reg [31:0] gpr_out_2; // @[lib.scala 374:16]
  reg [31:0] gpr_out_3; // @[lib.scala 374:16]
  reg [31:0] gpr_out_4; // @[lib.scala 374:16]
  reg [31:0] gpr_out_5; // @[lib.scala 374:16]
  reg [31:0] gpr_out_6; // @[lib.scala 374:16]
  reg [31:0] gpr_out_7; // @[lib.scala 374:16]
  reg [31:0] gpr_out_8; // @[lib.scala 374:16]
  reg [31:0] gpr_out_9; // @[lib.scala 374:16]
  reg [31:0] gpr_out_10; // @[lib.scala 374:16]
  reg [31:0] gpr_out_11; // @[lib.scala 374:16]
  reg [31:0] gpr_out_12; // @[lib.scala 374:16]
  reg [31:0] gpr_out_13; // @[lib.scala 374:16]
  reg [31:0] gpr_out_14; // @[lib.scala 374:16]
  reg [31:0] gpr_out_15; // @[lib.scala 374:16]
  reg [31:0] gpr_out_16; // @[lib.scala 374:16]
  reg [31:0] gpr_out_17; // @[lib.scala 374:16]
  reg [31:0] gpr_out_18; // @[lib.scala 374:16]
  reg [31:0] gpr_out_19; // @[lib.scala 374:16]
  reg [31:0] gpr_out_20; // @[lib.scala 374:16]
  reg [31:0] gpr_out_21; // @[lib.scala 374:16]
  reg [31:0] gpr_out_22; // @[lib.scala 374:16]
  reg [31:0] gpr_out_23; // @[lib.scala 374:16]
  reg [31:0] gpr_out_24; // @[lib.scala 374:16]
  reg [31:0] gpr_out_25; // @[lib.scala 374:16]
  reg [31:0] gpr_out_26; // @[lib.scala 374:16]
  reg [31:0] gpr_out_27; // @[lib.scala 374:16]
  reg [31:0] gpr_out_28; // @[lib.scala 374:16]
  reg [31:0] gpr_out_29; // @[lib.scala 374:16]
  reg [31:0] gpr_out_30; // @[lib.scala 374:16]
  reg [31:0] gpr_out_31; // @[lib.scala 374:16]
  wire  _T_684 = io_raddr0 == 5'h1; // @[dec_gpr_ctl.scala 64:72]
  wire  _T_686 = io_raddr0 == 5'h2; // @[dec_gpr_ctl.scala 64:72]
  wire  _T_688 = io_raddr0 == 5'h3; // @[dec_gpr_ctl.scala 64:72]
  wire  _T_690 = io_raddr0 == 5'h4; // @[dec_gpr_ctl.scala 64:72]
  wire  _T_692 = io_raddr0 == 5'h5; // @[dec_gpr_ctl.scala 64:72]
  wire  _T_694 = io_raddr0 == 5'h6; // @[dec_gpr_ctl.scala 64:72]
  wire  _T_696 = io_raddr0 == 5'h7; // @[dec_gpr_ctl.scala 64:72]
  wire  _T_698 = io_raddr0 == 5'h8; // @[dec_gpr_ctl.scala 64:72]
  wire  _T_700 = io_raddr0 == 5'h9; // @[dec_gpr_ctl.scala 64:72]
  wire  _T_702 = io_raddr0 == 5'ha; // @[dec_gpr_ctl.scala 64:72]
  wire  _T_704 = io_raddr0 == 5'hb; // @[dec_gpr_ctl.scala 64:72]
  wire  _T_706 = io_raddr0 == 5'hc; // @[dec_gpr_ctl.scala 64:72]
  wire  _T_708 = io_raddr0 == 5'hd; // @[dec_gpr_ctl.scala 64:72]
  wire  _T_710 = io_raddr0 == 5'he; // @[dec_gpr_ctl.scala 64:72]
  wire  _T_712 = io_raddr0 == 5'hf; // @[dec_gpr_ctl.scala 64:72]
  wire  _T_714 = io_raddr0 == 5'h10; // @[dec_gpr_ctl.scala 64:72]
  wire  _T_716 = io_raddr0 == 5'h11; // @[dec_gpr_ctl.scala 64:72]
  wire  _T_718 = io_raddr0 == 5'h12; // @[dec_gpr_ctl.scala 64:72]
  wire  _T_720 = io_raddr0 == 5'h13; // @[dec_gpr_ctl.scala 64:72]
  wire  _T_722 = io_raddr0 == 5'h14; // @[dec_gpr_ctl.scala 64:72]
  wire  _T_724 = io_raddr0 == 5'h15; // @[dec_gpr_ctl.scala 64:72]
  wire  _T_726 = io_raddr0 == 5'h16; // @[dec_gpr_ctl.scala 64:72]
  wire  _T_728 = io_raddr0 == 5'h17; // @[dec_gpr_ctl.scala 64:72]
  wire  _T_730 = io_raddr0 == 5'h18; // @[dec_gpr_ctl.scala 64:72]
  wire  _T_732 = io_raddr0 == 5'h19; // @[dec_gpr_ctl.scala 64:72]
  wire  _T_734 = io_raddr0 == 5'h1a; // @[dec_gpr_ctl.scala 64:72]
  wire  _T_736 = io_raddr0 == 5'h1b; // @[dec_gpr_ctl.scala 64:72]
  wire  _T_738 = io_raddr0 == 5'h1c; // @[dec_gpr_ctl.scala 64:72]
  wire  _T_740 = io_raddr0 == 5'h1d; // @[dec_gpr_ctl.scala 64:72]
  wire  _T_742 = io_raddr0 == 5'h1e; // @[dec_gpr_ctl.scala 64:72]
  wire  _T_744 = io_raddr0 == 5'h1f; // @[dec_gpr_ctl.scala 64:72]
  wire [31:0] _T_746 = _T_684 ? gpr_out_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_747 = _T_686 ? gpr_out_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_748 = _T_688 ? gpr_out_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_749 = _T_690 ? gpr_out_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_750 = _T_692 ? gpr_out_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_751 = _T_694 ? gpr_out_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_752 = _T_696 ? gpr_out_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_753 = _T_698 ? gpr_out_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_754 = _T_700 ? gpr_out_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_755 = _T_702 ? gpr_out_10 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_756 = _T_704 ? gpr_out_11 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_757 = _T_706 ? gpr_out_12 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_758 = _T_708 ? gpr_out_13 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_759 = _T_710 ? gpr_out_14 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_760 = _T_712 ? gpr_out_15 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_761 = _T_714 ? gpr_out_16 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_762 = _T_716 ? gpr_out_17 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_763 = _T_718 ? gpr_out_18 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_764 = _T_720 ? gpr_out_19 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_765 = _T_722 ? gpr_out_20 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_766 = _T_724 ? gpr_out_21 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_767 = _T_726 ? gpr_out_22 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_768 = _T_728 ? gpr_out_23 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_769 = _T_730 ? gpr_out_24 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_770 = _T_732 ? gpr_out_25 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_771 = _T_734 ? gpr_out_26 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_772 = _T_736 ? gpr_out_27 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_773 = _T_738 ? gpr_out_28 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_774 = _T_740 ? gpr_out_29 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_775 = _T_742 ? gpr_out_30 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_776 = _T_744 ? gpr_out_31 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_777 = _T_746 | _T_747; // @[Mux.scala 27:72]
  wire [31:0] _T_778 = _T_777 | _T_748; // @[Mux.scala 27:72]
  wire [31:0] _T_779 = _T_778 | _T_749; // @[Mux.scala 27:72]
  wire [31:0] _T_780 = _T_779 | _T_750; // @[Mux.scala 27:72]
  wire [31:0] _T_781 = _T_780 | _T_751; // @[Mux.scala 27:72]
  wire [31:0] _T_782 = _T_781 | _T_752; // @[Mux.scala 27:72]
  wire [31:0] _T_783 = _T_782 | _T_753; // @[Mux.scala 27:72]
  wire [31:0] _T_784 = _T_783 | _T_754; // @[Mux.scala 27:72]
  wire [31:0] _T_785 = _T_784 | _T_755; // @[Mux.scala 27:72]
  wire [31:0] _T_786 = _T_785 | _T_756; // @[Mux.scala 27:72]
  wire [31:0] _T_787 = _T_786 | _T_757; // @[Mux.scala 27:72]
  wire [31:0] _T_788 = _T_787 | _T_758; // @[Mux.scala 27:72]
  wire [31:0] _T_789 = _T_788 | _T_759; // @[Mux.scala 27:72]
  wire [31:0] _T_790 = _T_789 | _T_760; // @[Mux.scala 27:72]
  wire [31:0] _T_791 = _T_790 | _T_761; // @[Mux.scala 27:72]
  wire [31:0] _T_792 = _T_791 | _T_762; // @[Mux.scala 27:72]
  wire [31:0] _T_793 = _T_792 | _T_763; // @[Mux.scala 27:72]
  wire [31:0] _T_794 = _T_793 | _T_764; // @[Mux.scala 27:72]
  wire [31:0] _T_795 = _T_794 | _T_765; // @[Mux.scala 27:72]
  wire [31:0] _T_796 = _T_795 | _T_766; // @[Mux.scala 27:72]
  wire [31:0] _T_797 = _T_796 | _T_767; // @[Mux.scala 27:72]
  wire [31:0] _T_798 = _T_797 | _T_768; // @[Mux.scala 27:72]
  wire [31:0] _T_799 = _T_798 | _T_769; // @[Mux.scala 27:72]
  wire [31:0] _T_800 = _T_799 | _T_770; // @[Mux.scala 27:72]
  wire [31:0] _T_801 = _T_800 | _T_771; // @[Mux.scala 27:72]
  wire [31:0] _T_802 = _T_801 | _T_772; // @[Mux.scala 27:72]
  wire [31:0] _T_803 = _T_802 | _T_773; // @[Mux.scala 27:72]
  wire [31:0] _T_804 = _T_803 | _T_774; // @[Mux.scala 27:72]
  wire [31:0] _T_805 = _T_804 | _T_775; // @[Mux.scala 27:72]
  wire  _T_808 = io_raddr1 == 5'h1; // @[dec_gpr_ctl.scala 65:72]
  wire  _T_810 = io_raddr1 == 5'h2; // @[dec_gpr_ctl.scala 65:72]
  wire  _T_812 = io_raddr1 == 5'h3; // @[dec_gpr_ctl.scala 65:72]
  wire  _T_814 = io_raddr1 == 5'h4; // @[dec_gpr_ctl.scala 65:72]
  wire  _T_816 = io_raddr1 == 5'h5; // @[dec_gpr_ctl.scala 65:72]
  wire  _T_818 = io_raddr1 == 5'h6; // @[dec_gpr_ctl.scala 65:72]
  wire  _T_820 = io_raddr1 == 5'h7; // @[dec_gpr_ctl.scala 65:72]
  wire  _T_822 = io_raddr1 == 5'h8; // @[dec_gpr_ctl.scala 65:72]
  wire  _T_824 = io_raddr1 == 5'h9; // @[dec_gpr_ctl.scala 65:72]
  wire  _T_826 = io_raddr1 == 5'ha; // @[dec_gpr_ctl.scala 65:72]
  wire  _T_828 = io_raddr1 == 5'hb; // @[dec_gpr_ctl.scala 65:72]
  wire  _T_830 = io_raddr1 == 5'hc; // @[dec_gpr_ctl.scala 65:72]
  wire  _T_832 = io_raddr1 == 5'hd; // @[dec_gpr_ctl.scala 65:72]
  wire  _T_834 = io_raddr1 == 5'he; // @[dec_gpr_ctl.scala 65:72]
  wire  _T_836 = io_raddr1 == 5'hf; // @[dec_gpr_ctl.scala 65:72]
  wire  _T_838 = io_raddr1 == 5'h10; // @[dec_gpr_ctl.scala 65:72]
  wire  _T_840 = io_raddr1 == 5'h11; // @[dec_gpr_ctl.scala 65:72]
  wire  _T_842 = io_raddr1 == 5'h12; // @[dec_gpr_ctl.scala 65:72]
  wire  _T_844 = io_raddr1 == 5'h13; // @[dec_gpr_ctl.scala 65:72]
  wire  _T_846 = io_raddr1 == 5'h14; // @[dec_gpr_ctl.scala 65:72]
  wire  _T_848 = io_raddr1 == 5'h15; // @[dec_gpr_ctl.scala 65:72]
  wire  _T_850 = io_raddr1 == 5'h16; // @[dec_gpr_ctl.scala 65:72]
  wire  _T_852 = io_raddr1 == 5'h17; // @[dec_gpr_ctl.scala 65:72]
  wire  _T_854 = io_raddr1 == 5'h18; // @[dec_gpr_ctl.scala 65:72]
  wire  _T_856 = io_raddr1 == 5'h19; // @[dec_gpr_ctl.scala 65:72]
  wire  _T_858 = io_raddr1 == 5'h1a; // @[dec_gpr_ctl.scala 65:72]
  wire  _T_860 = io_raddr1 == 5'h1b; // @[dec_gpr_ctl.scala 65:72]
  wire  _T_862 = io_raddr1 == 5'h1c; // @[dec_gpr_ctl.scala 65:72]
  wire  _T_864 = io_raddr1 == 5'h1d; // @[dec_gpr_ctl.scala 65:72]
  wire  _T_866 = io_raddr1 == 5'h1e; // @[dec_gpr_ctl.scala 65:72]
  wire  _T_868 = io_raddr1 == 5'h1f; // @[dec_gpr_ctl.scala 65:72]
  wire [31:0] _T_870 = _T_808 ? gpr_out_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_871 = _T_810 ? gpr_out_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_872 = _T_812 ? gpr_out_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_873 = _T_814 ? gpr_out_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_874 = _T_816 ? gpr_out_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_875 = _T_818 ? gpr_out_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_876 = _T_820 ? gpr_out_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_877 = _T_822 ? gpr_out_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_878 = _T_824 ? gpr_out_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_879 = _T_826 ? gpr_out_10 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_880 = _T_828 ? gpr_out_11 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_881 = _T_830 ? gpr_out_12 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_882 = _T_832 ? gpr_out_13 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_883 = _T_834 ? gpr_out_14 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_884 = _T_836 ? gpr_out_15 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_885 = _T_838 ? gpr_out_16 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_886 = _T_840 ? gpr_out_17 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_887 = _T_842 ? gpr_out_18 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_888 = _T_844 ? gpr_out_19 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_889 = _T_846 ? gpr_out_20 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_890 = _T_848 ? gpr_out_21 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_891 = _T_850 ? gpr_out_22 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_892 = _T_852 ? gpr_out_23 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_893 = _T_854 ? gpr_out_24 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_894 = _T_856 ? gpr_out_25 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_895 = _T_858 ? gpr_out_26 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_896 = _T_860 ? gpr_out_27 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_897 = _T_862 ? gpr_out_28 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_898 = _T_864 ? gpr_out_29 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_899 = _T_866 ? gpr_out_30 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_900 = _T_868 ? gpr_out_31 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_901 = _T_870 | _T_871; // @[Mux.scala 27:72]
  wire [31:0] _T_902 = _T_901 | _T_872; // @[Mux.scala 27:72]
  wire [31:0] _T_903 = _T_902 | _T_873; // @[Mux.scala 27:72]
  wire [31:0] _T_904 = _T_903 | _T_874; // @[Mux.scala 27:72]
  wire [31:0] _T_905 = _T_904 | _T_875; // @[Mux.scala 27:72]
  wire [31:0] _T_906 = _T_905 | _T_876; // @[Mux.scala 27:72]
  wire [31:0] _T_907 = _T_906 | _T_877; // @[Mux.scala 27:72]
  wire [31:0] _T_908 = _T_907 | _T_878; // @[Mux.scala 27:72]
  wire [31:0] _T_909 = _T_908 | _T_879; // @[Mux.scala 27:72]
  wire [31:0] _T_910 = _T_909 | _T_880; // @[Mux.scala 27:72]
  wire [31:0] _T_911 = _T_910 | _T_881; // @[Mux.scala 27:72]
  wire [31:0] _T_912 = _T_911 | _T_882; // @[Mux.scala 27:72]
  wire [31:0] _T_913 = _T_912 | _T_883; // @[Mux.scala 27:72]
  wire [31:0] _T_914 = _T_913 | _T_884; // @[Mux.scala 27:72]
  wire [31:0] _T_915 = _T_914 | _T_885; // @[Mux.scala 27:72]
  wire [31:0] _T_916 = _T_915 | _T_886; // @[Mux.scala 27:72]
  wire [31:0] _T_917 = _T_916 | _T_887; // @[Mux.scala 27:72]
  wire [31:0] _T_918 = _T_917 | _T_888; // @[Mux.scala 27:72]
  wire [31:0] _T_919 = _T_918 | _T_889; // @[Mux.scala 27:72]
  wire [31:0] _T_920 = _T_919 | _T_890; // @[Mux.scala 27:72]
  wire [31:0] _T_921 = _T_920 | _T_891; // @[Mux.scala 27:72]
  wire [31:0] _T_922 = _T_921 | _T_892; // @[Mux.scala 27:72]
  wire [31:0] _T_923 = _T_922 | _T_893; // @[Mux.scala 27:72]
  wire [31:0] _T_924 = _T_923 | _T_894; // @[Mux.scala 27:72]
  wire [31:0] _T_925 = _T_924 | _T_895; // @[Mux.scala 27:72]
  wire [31:0] _T_926 = _T_925 | _T_896; // @[Mux.scala 27:72]
  wire [31:0] _T_927 = _T_926 | _T_897; // @[Mux.scala 27:72]
  wire [31:0] _T_928 = _T_927 | _T_898; // @[Mux.scala 27:72]
  wire [31:0] _T_929 = _T_928 | _T_899; // @[Mux.scala 27:72]
  rvclkhdr rvclkhdr ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_io_l1clk),
    .io_clk(rvclkhdr_io_clk),
    .io_en(rvclkhdr_io_en),
    .io_scan_mode(rvclkhdr_io_scan_mode)
  );
  rvclkhdr rvclkhdr_1 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_1_io_l1clk),
    .io_clk(rvclkhdr_1_io_clk),
    .io_en(rvclkhdr_1_io_en),
    .io_scan_mode(rvclkhdr_1_io_scan_mode)
  );
  rvclkhdr rvclkhdr_2 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_2_io_l1clk),
    .io_clk(rvclkhdr_2_io_clk),
    .io_en(rvclkhdr_2_io_en),
    .io_scan_mode(rvclkhdr_2_io_scan_mode)
  );
  rvclkhdr rvclkhdr_3 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_3_io_l1clk),
    .io_clk(rvclkhdr_3_io_clk),
    .io_en(rvclkhdr_3_io_en),
    .io_scan_mode(rvclkhdr_3_io_scan_mode)
  );
  rvclkhdr rvclkhdr_4 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_4_io_l1clk),
    .io_clk(rvclkhdr_4_io_clk),
    .io_en(rvclkhdr_4_io_en),
    .io_scan_mode(rvclkhdr_4_io_scan_mode)
  );
  rvclkhdr rvclkhdr_5 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_5_io_l1clk),
    .io_clk(rvclkhdr_5_io_clk),
    .io_en(rvclkhdr_5_io_en),
    .io_scan_mode(rvclkhdr_5_io_scan_mode)
  );
  rvclkhdr rvclkhdr_6 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_6_io_l1clk),
    .io_clk(rvclkhdr_6_io_clk),
    .io_en(rvclkhdr_6_io_en),
    .io_scan_mode(rvclkhdr_6_io_scan_mode)
  );
  rvclkhdr rvclkhdr_7 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_7_io_l1clk),
    .io_clk(rvclkhdr_7_io_clk),
    .io_en(rvclkhdr_7_io_en),
    .io_scan_mode(rvclkhdr_7_io_scan_mode)
  );
  rvclkhdr rvclkhdr_8 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_8_io_l1clk),
    .io_clk(rvclkhdr_8_io_clk),
    .io_en(rvclkhdr_8_io_en),
    .io_scan_mode(rvclkhdr_8_io_scan_mode)
  );
  rvclkhdr rvclkhdr_9 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_9_io_l1clk),
    .io_clk(rvclkhdr_9_io_clk),
    .io_en(rvclkhdr_9_io_en),
    .io_scan_mode(rvclkhdr_9_io_scan_mode)
  );
  rvclkhdr rvclkhdr_10 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_10_io_l1clk),
    .io_clk(rvclkhdr_10_io_clk),
    .io_en(rvclkhdr_10_io_en),
    .io_scan_mode(rvclkhdr_10_io_scan_mode)
  );
  rvclkhdr rvclkhdr_11 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_11_io_l1clk),
    .io_clk(rvclkhdr_11_io_clk),
    .io_en(rvclkhdr_11_io_en),
    .io_scan_mode(rvclkhdr_11_io_scan_mode)
  );
  rvclkhdr rvclkhdr_12 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_12_io_l1clk),
    .io_clk(rvclkhdr_12_io_clk),
    .io_en(rvclkhdr_12_io_en),
    .io_scan_mode(rvclkhdr_12_io_scan_mode)
  );
  rvclkhdr rvclkhdr_13 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_13_io_l1clk),
    .io_clk(rvclkhdr_13_io_clk),
    .io_en(rvclkhdr_13_io_en),
    .io_scan_mode(rvclkhdr_13_io_scan_mode)
  );
  rvclkhdr rvclkhdr_14 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_14_io_l1clk),
    .io_clk(rvclkhdr_14_io_clk),
    .io_en(rvclkhdr_14_io_en),
    .io_scan_mode(rvclkhdr_14_io_scan_mode)
  );
  rvclkhdr rvclkhdr_15 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_15_io_l1clk),
    .io_clk(rvclkhdr_15_io_clk),
    .io_en(rvclkhdr_15_io_en),
    .io_scan_mode(rvclkhdr_15_io_scan_mode)
  );
  rvclkhdr rvclkhdr_16 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_16_io_l1clk),
    .io_clk(rvclkhdr_16_io_clk),
    .io_en(rvclkhdr_16_io_en),
    .io_scan_mode(rvclkhdr_16_io_scan_mode)
  );
  rvclkhdr rvclkhdr_17 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_17_io_l1clk),
    .io_clk(rvclkhdr_17_io_clk),
    .io_en(rvclkhdr_17_io_en),
    .io_scan_mode(rvclkhdr_17_io_scan_mode)
  );
  rvclkhdr rvclkhdr_18 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_18_io_l1clk),
    .io_clk(rvclkhdr_18_io_clk),
    .io_en(rvclkhdr_18_io_en),
    .io_scan_mode(rvclkhdr_18_io_scan_mode)
  );
  rvclkhdr rvclkhdr_19 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_19_io_l1clk),
    .io_clk(rvclkhdr_19_io_clk),
    .io_en(rvclkhdr_19_io_en),
    .io_scan_mode(rvclkhdr_19_io_scan_mode)
  );
  rvclkhdr rvclkhdr_20 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_20_io_l1clk),
    .io_clk(rvclkhdr_20_io_clk),
    .io_en(rvclkhdr_20_io_en),
    .io_scan_mode(rvclkhdr_20_io_scan_mode)
  );
  rvclkhdr rvclkhdr_21 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_21_io_l1clk),
    .io_clk(rvclkhdr_21_io_clk),
    .io_en(rvclkhdr_21_io_en),
    .io_scan_mode(rvclkhdr_21_io_scan_mode)
  );
  rvclkhdr rvclkhdr_22 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_22_io_l1clk),
    .io_clk(rvclkhdr_22_io_clk),
    .io_en(rvclkhdr_22_io_en),
    .io_scan_mode(rvclkhdr_22_io_scan_mode)
  );
  rvclkhdr rvclkhdr_23 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_23_io_l1clk),
    .io_clk(rvclkhdr_23_io_clk),
    .io_en(rvclkhdr_23_io_en),
    .io_scan_mode(rvclkhdr_23_io_scan_mode)
  );
  rvclkhdr rvclkhdr_24 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_24_io_l1clk),
    .io_clk(rvclkhdr_24_io_clk),
    .io_en(rvclkhdr_24_io_en),
    .io_scan_mode(rvclkhdr_24_io_scan_mode)
  );
  rvclkhdr rvclkhdr_25 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_25_io_l1clk),
    .io_clk(rvclkhdr_25_io_clk),
    .io_en(rvclkhdr_25_io_en),
    .io_scan_mode(rvclkhdr_25_io_scan_mode)
  );
  rvclkhdr rvclkhdr_26 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_26_io_l1clk),
    .io_clk(rvclkhdr_26_io_clk),
    .io_en(rvclkhdr_26_io_en),
    .io_scan_mode(rvclkhdr_26_io_scan_mode)
  );
  rvclkhdr rvclkhdr_27 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_27_io_l1clk),
    .io_clk(rvclkhdr_27_io_clk),
    .io_en(rvclkhdr_27_io_en),
    .io_scan_mode(rvclkhdr_27_io_scan_mode)
  );
  rvclkhdr rvclkhdr_28 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_28_io_l1clk),
    .io_clk(rvclkhdr_28_io_clk),
    .io_en(rvclkhdr_28_io_en),
    .io_scan_mode(rvclkhdr_28_io_scan_mode)
  );
  rvclkhdr rvclkhdr_29 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_29_io_l1clk),
    .io_clk(rvclkhdr_29_io_clk),
    .io_en(rvclkhdr_29_io_en),
    .io_scan_mode(rvclkhdr_29_io_scan_mode)
  );
  rvclkhdr rvclkhdr_30 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_30_io_l1clk),
    .io_clk(rvclkhdr_30_io_clk),
    .io_en(rvclkhdr_30_io_en),
    .io_scan_mode(rvclkhdr_30_io_scan_mode)
  );
  assign io_gpr_exu_gpr_i0_rs1_d = _T_805 | _T_776; // @[dec_gpr_ctl.scala 48:32 dec_gpr_ctl.scala 64:32]
  assign io_gpr_exu_gpr_i0_rs2_d = _T_929 | _T_900; // @[dec_gpr_ctl.scala 49:32 dec_gpr_ctl.scala 65:32]
  assign rvclkhdr_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_io_en = gpr_wr_en[1]; // @[lib.scala 371:17]
  assign rvclkhdr_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_1_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_1_io_en = gpr_wr_en[2]; // @[lib.scala 371:17]
  assign rvclkhdr_1_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_2_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_2_io_en = gpr_wr_en[3]; // @[lib.scala 371:17]
  assign rvclkhdr_2_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_3_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_3_io_en = gpr_wr_en[4]; // @[lib.scala 371:17]
  assign rvclkhdr_3_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_4_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_4_io_en = gpr_wr_en[5]; // @[lib.scala 371:17]
  assign rvclkhdr_4_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_5_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_5_io_en = gpr_wr_en[6]; // @[lib.scala 371:17]
  assign rvclkhdr_5_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_6_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_6_io_en = gpr_wr_en[7]; // @[lib.scala 371:17]
  assign rvclkhdr_6_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_7_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_7_io_en = gpr_wr_en[8]; // @[lib.scala 371:17]
  assign rvclkhdr_7_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_8_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_8_io_en = gpr_wr_en[9]; // @[lib.scala 371:17]
  assign rvclkhdr_8_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_9_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_9_io_en = gpr_wr_en[10]; // @[lib.scala 371:17]
  assign rvclkhdr_9_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_10_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_10_io_en = gpr_wr_en[11]; // @[lib.scala 371:17]
  assign rvclkhdr_10_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_11_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_11_io_en = gpr_wr_en[12]; // @[lib.scala 371:17]
  assign rvclkhdr_11_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_12_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_12_io_en = gpr_wr_en[13]; // @[lib.scala 371:17]
  assign rvclkhdr_12_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_13_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_13_io_en = gpr_wr_en[14]; // @[lib.scala 371:17]
  assign rvclkhdr_13_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_14_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_14_io_en = gpr_wr_en[15]; // @[lib.scala 371:17]
  assign rvclkhdr_14_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_15_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_15_io_en = gpr_wr_en[16]; // @[lib.scala 371:17]
  assign rvclkhdr_15_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_16_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_16_io_en = gpr_wr_en[17]; // @[lib.scala 371:17]
  assign rvclkhdr_16_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_17_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_17_io_en = gpr_wr_en[18]; // @[lib.scala 371:17]
  assign rvclkhdr_17_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_18_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_18_io_en = gpr_wr_en[19]; // @[lib.scala 371:17]
  assign rvclkhdr_18_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_19_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_19_io_en = gpr_wr_en[20]; // @[lib.scala 371:17]
  assign rvclkhdr_19_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_20_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_20_io_en = gpr_wr_en[21]; // @[lib.scala 371:17]
  assign rvclkhdr_20_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_21_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_21_io_en = gpr_wr_en[22]; // @[lib.scala 371:17]
  assign rvclkhdr_21_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_22_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_22_io_en = gpr_wr_en[23]; // @[lib.scala 371:17]
  assign rvclkhdr_22_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_23_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_23_io_en = gpr_wr_en[24]; // @[lib.scala 371:17]
  assign rvclkhdr_23_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_24_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_24_io_en = gpr_wr_en[25]; // @[lib.scala 371:17]
  assign rvclkhdr_24_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_25_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_25_io_en = gpr_wr_en[26]; // @[lib.scala 371:17]
  assign rvclkhdr_25_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_26_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_26_io_en = gpr_wr_en[27]; // @[lib.scala 371:17]
  assign rvclkhdr_26_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_27_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_27_io_en = gpr_wr_en[28]; // @[lib.scala 371:17]
  assign rvclkhdr_27_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_28_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_28_io_en = gpr_wr_en[29]; // @[lib.scala 371:17]
  assign rvclkhdr_28_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_29_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_29_io_en = gpr_wr_en[30]; // @[lib.scala 371:17]
  assign rvclkhdr_29_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_30_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_30_io_en = gpr_wr_en[31]; // @[lib.scala 371:17]
  assign rvclkhdr_30_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  gpr_out_1 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  gpr_out_2 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  gpr_out_3 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  gpr_out_4 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  gpr_out_5 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  gpr_out_6 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  gpr_out_7 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  gpr_out_8 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  gpr_out_9 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  gpr_out_10 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  gpr_out_11 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  gpr_out_12 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  gpr_out_13 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  gpr_out_14 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  gpr_out_15 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  gpr_out_16 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  gpr_out_17 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  gpr_out_18 = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  gpr_out_19 = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  gpr_out_20 = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  gpr_out_21 = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  gpr_out_22 = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  gpr_out_23 = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  gpr_out_24 = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  gpr_out_25 = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  gpr_out_26 = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  gpr_out_27 = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  gpr_out_28 = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  gpr_out_29 = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  gpr_out_30 = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  gpr_out_31 = _RAND_30[31:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    gpr_out_1 = 32'h0;
  end
  if (reset) begin
    gpr_out_2 = 32'h0;
  end
  if (reset) begin
    gpr_out_3 = 32'h0;
  end
  if (reset) begin
    gpr_out_4 = 32'h0;
  end
  if (reset) begin
    gpr_out_5 = 32'h0;
  end
  if (reset) begin
    gpr_out_6 = 32'h0;
  end
  if (reset) begin
    gpr_out_7 = 32'h0;
  end
  if (reset) begin
    gpr_out_8 = 32'h0;
  end
  if (reset) begin
    gpr_out_9 = 32'h0;
  end
  if (reset) begin
    gpr_out_10 = 32'h0;
  end
  if (reset) begin
    gpr_out_11 = 32'h0;
  end
  if (reset) begin
    gpr_out_12 = 32'h0;
  end
  if (reset) begin
    gpr_out_13 = 32'h0;
  end
  if (reset) begin
    gpr_out_14 = 32'h0;
  end
  if (reset) begin
    gpr_out_15 = 32'h0;
  end
  if (reset) begin
    gpr_out_16 = 32'h0;
  end
  if (reset) begin
    gpr_out_17 = 32'h0;
  end
  if (reset) begin
    gpr_out_18 = 32'h0;
  end
  if (reset) begin
    gpr_out_19 = 32'h0;
  end
  if (reset) begin
    gpr_out_20 = 32'h0;
  end
  if (reset) begin
    gpr_out_21 = 32'h0;
  end
  if (reset) begin
    gpr_out_22 = 32'h0;
  end
  if (reset) begin
    gpr_out_23 = 32'h0;
  end
  if (reset) begin
    gpr_out_24 = 32'h0;
  end
  if (reset) begin
    gpr_out_25 = 32'h0;
  end
  if (reset) begin
    gpr_out_26 = 32'h0;
  end
  if (reset) begin
    gpr_out_27 = 32'h0;
  end
  if (reset) begin
    gpr_out_28 = 32'h0;
  end
  if (reset) begin
    gpr_out_29 = 32'h0;
  end
  if (reset) begin
    gpr_out_30 = 32'h0;
  end
  if (reset) begin
    gpr_out_31 = 32'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge rvclkhdr_io_l1clk or posedge reset) begin
    if (reset) begin
      gpr_out_1 <= 32'h0;
    end else begin
      gpr_out_1 <= _T_12 | _T_15;
    end
  end
  always @(posedge rvclkhdr_1_io_l1clk or posedge reset) begin
    if (reset) begin
      gpr_out_2 <= 32'h0;
    end else begin
      gpr_out_2 <= _T_29 | _T_32;
    end
  end
  always @(posedge rvclkhdr_2_io_l1clk or posedge reset) begin
    if (reset) begin
      gpr_out_3 <= 32'h0;
    end else begin
      gpr_out_3 <= _T_46 | _T_49;
    end
  end
  always @(posedge rvclkhdr_3_io_l1clk or posedge reset) begin
    if (reset) begin
      gpr_out_4 <= 32'h0;
    end else begin
      gpr_out_4 <= _T_63 | _T_66;
    end
  end
  always @(posedge rvclkhdr_4_io_l1clk or posedge reset) begin
    if (reset) begin
      gpr_out_5 <= 32'h0;
    end else begin
      gpr_out_5 <= _T_80 | _T_83;
    end
  end
  always @(posedge rvclkhdr_5_io_l1clk or posedge reset) begin
    if (reset) begin
      gpr_out_6 <= 32'h0;
    end else begin
      gpr_out_6 <= _T_97 | _T_100;
    end
  end
  always @(posedge rvclkhdr_6_io_l1clk or posedge reset) begin
    if (reset) begin
      gpr_out_7 <= 32'h0;
    end else begin
      gpr_out_7 <= _T_114 | _T_117;
    end
  end
  always @(posedge rvclkhdr_7_io_l1clk or posedge reset) begin
    if (reset) begin
      gpr_out_8 <= 32'h0;
    end else begin
      gpr_out_8 <= _T_131 | _T_134;
    end
  end
  always @(posedge rvclkhdr_8_io_l1clk or posedge reset) begin
    if (reset) begin
      gpr_out_9 <= 32'h0;
    end else begin
      gpr_out_9 <= _T_148 | _T_151;
    end
  end
  always @(posedge rvclkhdr_9_io_l1clk or posedge reset) begin
    if (reset) begin
      gpr_out_10 <= 32'h0;
    end else begin
      gpr_out_10 <= _T_165 | _T_168;
    end
  end
  always @(posedge rvclkhdr_10_io_l1clk or posedge reset) begin
    if (reset) begin
      gpr_out_11 <= 32'h0;
    end else begin
      gpr_out_11 <= _T_182 | _T_185;
    end
  end
  always @(posedge rvclkhdr_11_io_l1clk or posedge reset) begin
    if (reset) begin
      gpr_out_12 <= 32'h0;
    end else begin
      gpr_out_12 <= _T_199 | _T_202;
    end
  end
  always @(posedge rvclkhdr_12_io_l1clk or posedge reset) begin
    if (reset) begin
      gpr_out_13 <= 32'h0;
    end else begin
      gpr_out_13 <= _T_216 | _T_219;
    end
  end
  always @(posedge rvclkhdr_13_io_l1clk or posedge reset) begin
    if (reset) begin
      gpr_out_14 <= 32'h0;
    end else begin
      gpr_out_14 <= _T_233 | _T_236;
    end
  end
  always @(posedge rvclkhdr_14_io_l1clk or posedge reset) begin
    if (reset) begin
      gpr_out_15 <= 32'h0;
    end else begin
      gpr_out_15 <= _T_250 | _T_253;
    end
  end
  always @(posedge rvclkhdr_15_io_l1clk or posedge reset) begin
    if (reset) begin
      gpr_out_16 <= 32'h0;
    end else begin
      gpr_out_16 <= _T_267 | _T_270;
    end
  end
  always @(posedge rvclkhdr_16_io_l1clk or posedge reset) begin
    if (reset) begin
      gpr_out_17 <= 32'h0;
    end else begin
      gpr_out_17 <= _T_284 | _T_287;
    end
  end
  always @(posedge rvclkhdr_17_io_l1clk or posedge reset) begin
    if (reset) begin
      gpr_out_18 <= 32'h0;
    end else begin
      gpr_out_18 <= _T_301 | _T_304;
    end
  end
  always @(posedge rvclkhdr_18_io_l1clk or posedge reset) begin
    if (reset) begin
      gpr_out_19 <= 32'h0;
    end else begin
      gpr_out_19 <= _T_318 | _T_321;
    end
  end
  always @(posedge rvclkhdr_19_io_l1clk or posedge reset) begin
    if (reset) begin
      gpr_out_20 <= 32'h0;
    end else begin
      gpr_out_20 <= _T_335 | _T_338;
    end
  end
  always @(posedge rvclkhdr_20_io_l1clk or posedge reset) begin
    if (reset) begin
      gpr_out_21 <= 32'h0;
    end else begin
      gpr_out_21 <= _T_352 | _T_355;
    end
  end
  always @(posedge rvclkhdr_21_io_l1clk or posedge reset) begin
    if (reset) begin
      gpr_out_22 <= 32'h0;
    end else begin
      gpr_out_22 <= _T_369 | _T_372;
    end
  end
  always @(posedge rvclkhdr_22_io_l1clk or posedge reset) begin
    if (reset) begin
      gpr_out_23 <= 32'h0;
    end else begin
      gpr_out_23 <= _T_386 | _T_389;
    end
  end
  always @(posedge rvclkhdr_23_io_l1clk or posedge reset) begin
    if (reset) begin
      gpr_out_24 <= 32'h0;
    end else begin
      gpr_out_24 <= _T_403 | _T_406;
    end
  end
  always @(posedge rvclkhdr_24_io_l1clk or posedge reset) begin
    if (reset) begin
      gpr_out_25 <= 32'h0;
    end else begin
      gpr_out_25 <= _T_420 | _T_423;
    end
  end
  always @(posedge rvclkhdr_25_io_l1clk or posedge reset) begin
    if (reset) begin
      gpr_out_26 <= 32'h0;
    end else begin
      gpr_out_26 <= _T_437 | _T_440;
    end
  end
  always @(posedge rvclkhdr_26_io_l1clk or posedge reset) begin
    if (reset) begin
      gpr_out_27 <= 32'h0;
    end else begin
      gpr_out_27 <= _T_454 | _T_457;
    end
  end
  always @(posedge rvclkhdr_27_io_l1clk or posedge reset) begin
    if (reset) begin
      gpr_out_28 <= 32'h0;
    end else begin
      gpr_out_28 <= _T_471 | _T_474;
    end
  end
  always @(posedge rvclkhdr_28_io_l1clk or posedge reset) begin
    if (reset) begin
      gpr_out_29 <= 32'h0;
    end else begin
      gpr_out_29 <= _T_488 | _T_491;
    end
  end
  always @(posedge rvclkhdr_29_io_l1clk or posedge reset) begin
    if (reset) begin
      gpr_out_30 <= 32'h0;
    end else begin
      gpr_out_30 <= _T_505 | _T_508;
    end
  end
  always @(posedge rvclkhdr_30_io_l1clk or posedge reset) begin
    if (reset) begin
      gpr_out_31 <= 32'h0;
    end else begin
      gpr_out_31 <= _T_522 | _T_525;
    end
  end
endmodule
module dec_timer_ctl(
  input         clock,
  input         reset,
  input         io_free_clk,
  input         io_scan_mode,
  input         io_dec_csr_wen_r_mod,
  input  [11:0] io_dec_csr_wraddr_r,
  input  [31:0] io_dec_csr_wrdata_r,
  input         io_csr_mitctl0,
  input         io_csr_mitctl1,
  input         io_csr_mitb0,
  input         io_csr_mitb1,
  input         io_csr_mitcnt0,
  input         io_csr_mitcnt1,
  input         io_dec_pause_state,
  input         io_dec_tlu_pmu_fw_halted,
  input         io_internal_dbg_halt_timers,
  output [31:0] io_dec_timer_rddata_d,
  output        io_dec_timer_read_d,
  output        io_dec_timer_t0_pulse,
  output        io_dec_timer_t1_pulse
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  wire  rvclkhdr_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_1_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_1_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_1_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_1_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_2_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_2_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_2_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_2_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_3_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_3_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_3_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_3_io_scan_mode; // @[lib.scala 368:23]
  reg [31:0] mitcnt0; // @[lib.scala 374:16]
  reg [31:0] mitb0_b; // @[lib.scala 374:16]
  wire [31:0] mitb0 = ~mitb0_b; // @[dec_tlu_ctl.scala 2713:22]
  wire  mit0_match_ns = mitcnt0 >= mitb0; // @[dec_tlu_ctl.scala 2674:36]
  reg [31:0] mitcnt1; // @[lib.scala 374:16]
  reg [31:0] mitb1_b; // @[lib.scala 374:16]
  wire [31:0] mitb1 = ~mitb1_b; // @[dec_tlu_ctl.scala 2722:18]
  wire  mit1_match_ns = mitcnt1 >= mitb1; // @[dec_tlu_ctl.scala 2675:36]
  wire  _T = io_dec_csr_wraddr_r == 12'h7d2; // @[dec_tlu_ctl.scala 2685:72]
  wire  wr_mitcnt0_r = io_dec_csr_wen_r_mod & _T; // @[dec_tlu_ctl.scala 2685:49]
  reg [1:0] _T_57; // @[dec_tlu_ctl.scala 2738:67]
  reg  mitctl0_0_b; // @[dec_tlu_ctl.scala 2737:60]
  wire  _T_58 = ~mitctl0_0_b; // @[dec_tlu_ctl.scala 2738:90]
  wire [2:0] mitctl0 = {_T_57,_T_58}; // @[Cat.scala 29:58]
  wire  _T_2 = ~io_dec_pause_state; // @[dec_tlu_ctl.scala 2687:56]
  wire  _T_4 = _T_2 | mitctl0[2]; // @[dec_tlu_ctl.scala 2687:76]
  wire  _T_5 = mitctl0[0] & _T_4; // @[dec_tlu_ctl.scala 2687:53]
  wire  _T_6 = ~io_dec_tlu_pmu_fw_halted; // @[dec_tlu_ctl.scala 2687:112]
  wire  _T_8 = _T_6 | mitctl0[1]; // @[dec_tlu_ctl.scala 2687:138]
  wire  _T_9 = _T_5 & _T_8; // @[dec_tlu_ctl.scala 2687:109]
  wire  _T_10 = ~io_internal_dbg_halt_timers; // @[dec_tlu_ctl.scala 2687:173]
  wire  mitcnt0_inc_ok = _T_9 & _T_10; // @[dec_tlu_ctl.scala 2687:171]
  wire [31:0] mitcnt0_inc = mitcnt0 + 32'h1; // @[dec_tlu_ctl.scala 2688:35]
  wire  _T_15 = wr_mitcnt0_r | mitcnt0_inc_ok; // @[dec_tlu_ctl.scala 2690:59]
  wire  _T_19 = io_dec_csr_wraddr_r == 12'h7d5; // @[dec_tlu_ctl.scala 2697:72]
  wire  wr_mitcnt1_r = io_dec_csr_wen_r_mod & _T_19; // @[dec_tlu_ctl.scala 2697:49]
  reg [2:0] _T_66; // @[dec_tlu_ctl.scala 2752:52]
  reg  mitctl1_0_b; // @[dec_tlu_ctl.scala 2751:55]
  wire  _T_67 = ~mitctl1_0_b; // @[dec_tlu_ctl.scala 2752:75]
  wire [3:0] mitctl1 = {_T_66,_T_67}; // @[Cat.scala 29:58]
  wire  _T_23 = _T_2 | mitctl1[2]; // @[dec_tlu_ctl.scala 2699:76]
  wire  _T_24 = mitctl1[0] & _T_23; // @[dec_tlu_ctl.scala 2699:53]
  wire  _T_27 = _T_6 | mitctl1[1]; // @[dec_tlu_ctl.scala 2699:138]
  wire  _T_28 = _T_24 & _T_27; // @[dec_tlu_ctl.scala 2699:109]
  wire  mitcnt1_inc_ok = _T_28 & _T_10; // @[dec_tlu_ctl.scala 2699:171]
  wire  _T_32 = ~mitctl1[3]; // @[dec_tlu_ctl.scala 2702:60]
  wire  _T_33 = _T_32 | mit0_match_ns; // @[dec_tlu_ctl.scala 2702:72]
  wire [31:0] _T_34 = {31'h0,_T_33}; // @[Cat.scala 29:58]
  wire [31:0] mitcnt1_inc = mitcnt1 + _T_34; // @[dec_tlu_ctl.scala 2702:35]
  wire  _T_39 = wr_mitcnt1_r | mitcnt1_inc_ok; // @[dec_tlu_ctl.scala 2704:60]
  wire  _T_43 = io_dec_csr_wraddr_r == 12'h7d3; // @[dec_tlu_ctl.scala 2711:70]
  wire  _T_47 = io_dec_csr_wraddr_r == 12'h7d6; // @[dec_tlu_ctl.scala 2720:69]
  wire  _T_51 = io_dec_csr_wraddr_r == 12'h7d4; // @[dec_tlu_ctl.scala 2733:72]
  wire  wr_mitctl0_r = io_dec_csr_wen_r_mod & _T_51; // @[dec_tlu_ctl.scala 2733:49]
  wire [2:0] mitctl0_ns = wr_mitctl0_r ? io_dec_csr_wrdata_r[2:0] : mitctl0; // @[dec_tlu_ctl.scala 2734:31]
  wire  _T_60 = io_dec_csr_wraddr_r == 12'h7d7; // @[dec_tlu_ctl.scala 2748:71]
  wire  wr_mitctl1_r = io_dec_csr_wen_r_mod & _T_60; // @[dec_tlu_ctl.scala 2748:49]
  wire [3:0] mitctl1_ns = wr_mitctl1_r ? io_dec_csr_wrdata_r[3:0] : mitctl1; // @[dec_tlu_ctl.scala 2749:31]
  wire  _T_69 = io_csr_mitcnt1 | io_csr_mitcnt0; // @[dec_tlu_ctl.scala 2754:51]
  wire  _T_70 = _T_69 | io_csr_mitb1; // @[dec_tlu_ctl.scala 2754:68]
  wire  _T_71 = _T_70 | io_csr_mitb0; // @[dec_tlu_ctl.scala 2754:83]
  wire  _T_72 = _T_71 | io_csr_mitctl0; // @[dec_tlu_ctl.scala 2754:98]
  wire [31:0] _T_81 = {29'h0,_T_57,_T_58}; // @[Cat.scala 29:58]
  wire [31:0] _T_84 = {28'h0,_T_66,_T_67}; // @[Cat.scala 29:58]
  wire [31:0] _T_85 = io_csr_mitcnt0 ? mitcnt0 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_86 = io_csr_mitcnt1 ? mitcnt1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_87 = io_csr_mitb0 ? mitb0 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_88 = io_csr_mitb1 ? mitb1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_89 = io_csr_mitctl0 ? _T_81 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_90 = io_csr_mitctl1 ? _T_84 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_91 = _T_85 | _T_86; // @[Mux.scala 27:72]
  wire [31:0] _T_92 = _T_91 | _T_87; // @[Mux.scala 27:72]
  wire [31:0] _T_93 = _T_92 | _T_88; // @[Mux.scala 27:72]
  wire [31:0] _T_94 = _T_93 | _T_89; // @[Mux.scala 27:72]
  rvclkhdr rvclkhdr ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_io_l1clk),
    .io_clk(rvclkhdr_io_clk),
    .io_en(rvclkhdr_io_en),
    .io_scan_mode(rvclkhdr_io_scan_mode)
  );
  rvclkhdr rvclkhdr_1 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_1_io_l1clk),
    .io_clk(rvclkhdr_1_io_clk),
    .io_en(rvclkhdr_1_io_en),
    .io_scan_mode(rvclkhdr_1_io_scan_mode)
  );
  rvclkhdr rvclkhdr_2 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_2_io_l1clk),
    .io_clk(rvclkhdr_2_io_clk),
    .io_en(rvclkhdr_2_io_en),
    .io_scan_mode(rvclkhdr_2_io_scan_mode)
  );
  rvclkhdr rvclkhdr_3 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_3_io_l1clk),
    .io_clk(rvclkhdr_3_io_clk),
    .io_en(rvclkhdr_3_io_en),
    .io_scan_mode(rvclkhdr_3_io_scan_mode)
  );
  assign io_dec_timer_rddata_d = _T_94 | _T_90; // @[dec_tlu_ctl.scala 2755:33]
  assign io_dec_timer_read_d = _T_72 | io_csr_mitctl1; // @[dec_tlu_ctl.scala 2754:33]
  assign io_dec_timer_t0_pulse = mitcnt0 >= mitb0; // @[dec_tlu_ctl.scala 2677:31]
  assign io_dec_timer_t1_pulse = mitcnt1 >= mitb1; // @[dec_tlu_ctl.scala 2678:31]
  assign rvclkhdr_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_io_en = _T_15 | mit0_match_ns; // @[lib.scala 371:17]
  assign rvclkhdr_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_1_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_1_io_en = _T_39 | mit1_match_ns; // @[lib.scala 371:17]
  assign rvclkhdr_1_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_2_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_2_io_en = io_dec_csr_wen_r_mod & _T_43; // @[lib.scala 371:17]
  assign rvclkhdr_2_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_3_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_3_io_en = io_dec_csr_wen_r_mod & _T_47; // @[lib.scala 371:17]
  assign rvclkhdr_3_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  mitcnt0 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  mitb0_b = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  mitcnt1 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  mitb1_b = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  _T_57 = _RAND_4[1:0];
  _RAND_5 = {1{`RANDOM}};
  mitctl0_0_b = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  _T_66 = _RAND_6[2:0];
  _RAND_7 = {1{`RANDOM}};
  mitctl1_0_b = _RAND_7[0:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    mitcnt0 = 32'h0;
  end
  if (reset) begin
    mitb0_b = 32'h0;
  end
  if (reset) begin
    mitcnt1 = 32'h0;
  end
  if (reset) begin
    mitb1_b = 32'h0;
  end
  if (reset) begin
    _T_57 = 2'h0;
  end
  if (reset) begin
    mitctl0_0_b = 1'h0;
  end
  if (reset) begin
    _T_66 = 3'h0;
  end
  if (reset) begin
    mitctl1_0_b = 1'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge rvclkhdr_io_l1clk or posedge reset) begin
    if (reset) begin
      mitcnt0 <= 32'h0;
    end else if (mit0_match_ns) begin
      mitcnt0 <= 32'h0;
    end else if (wr_mitcnt0_r) begin
      mitcnt0 <= io_dec_csr_wrdata_r;
    end else begin
      mitcnt0 <= mitcnt0_inc;
    end
  end
  always @(posedge rvclkhdr_2_io_l1clk or posedge reset) begin
    if (reset) begin
      mitb0_b <= 32'h0;
    end else begin
      mitb0_b <= ~io_dec_csr_wrdata_r;
    end
  end
  always @(posedge rvclkhdr_1_io_l1clk or posedge reset) begin
    if (reset) begin
      mitcnt1 <= 32'h0;
    end else if (mit1_match_ns) begin
      mitcnt1 <= 32'h0;
    end else if (wr_mitcnt1_r) begin
      mitcnt1 <= io_dec_csr_wrdata_r;
    end else begin
      mitcnt1 <= mitcnt1_inc;
    end
  end
  always @(posedge rvclkhdr_3_io_l1clk or posedge reset) begin
    if (reset) begin
      mitb1_b <= 32'h0;
    end else begin
      mitb1_b <= ~io_dec_csr_wrdata_r;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      _T_57 <= 2'h0;
    end else begin
      _T_57 <= mitctl0_ns[2:1];
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      mitctl0_0_b <= 1'h0;
    end else begin
      mitctl0_0_b <= ~mitctl0_ns[0];
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      _T_66 <= 3'h0;
    end else begin
      _T_66 <= mitctl1_ns[3:1];
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      mitctl1_0_b <= 1'h0;
    end else begin
      mitctl1_0_b <= ~mitctl1_ns[0];
    end
  end
endmodule
module csr_tlu(
  input         clock,
  input         reset,
  input         io_free_clk,
  input         io_active_clk,
  input         io_scan_mode,
  input  [31:0] io_dec_csr_wrdata_r,
  input  [11:0] io_dec_csr_wraddr_r,
  input  [11:0] io_dec_csr_rdaddr_d,
  input         io_dec_csr_wen_unq_d,
  input         io_dec_i0_decode_d,
  output [70:0] io_dec_tlu_ic_diag_pkt_icache_wrdata,
  output [16:0] io_dec_tlu_ic_diag_pkt_icache_dicawics,
  output        io_dec_tlu_ic_diag_pkt_icache_rd_valid,
  output        io_dec_tlu_ic_diag_pkt_icache_wr_valid,
  input         io_ifu_ic_debug_rd_data_valid,
  output        io_trigger_pkt_any_0_select,
  output        io_trigger_pkt_any_0_match_pkt,
  output        io_trigger_pkt_any_0_store,
  output        io_trigger_pkt_any_0_load,
  output        io_trigger_pkt_any_0_execute,
  output        io_trigger_pkt_any_0_m,
  output [31:0] io_trigger_pkt_any_0_tdata2,
  output        io_trigger_pkt_any_1_select,
  output        io_trigger_pkt_any_1_match_pkt,
  output        io_trigger_pkt_any_1_store,
  output        io_trigger_pkt_any_1_load,
  output        io_trigger_pkt_any_1_execute,
  output        io_trigger_pkt_any_1_m,
  output [31:0] io_trigger_pkt_any_1_tdata2,
  output        io_trigger_pkt_any_2_select,
  output        io_trigger_pkt_any_2_match_pkt,
  output        io_trigger_pkt_any_2_store,
  output        io_trigger_pkt_any_2_load,
  output        io_trigger_pkt_any_2_execute,
  output        io_trigger_pkt_any_2_m,
  output [31:0] io_trigger_pkt_any_2_tdata2,
  output        io_trigger_pkt_any_3_select,
  output        io_trigger_pkt_any_3_match_pkt,
  output        io_trigger_pkt_any_3_store,
  output        io_trigger_pkt_any_3_load,
  output        io_trigger_pkt_any_3_execute,
  output        io_trigger_pkt_any_3_m,
  output [31:0] io_trigger_pkt_any_3_tdata2,
  input         io_dma_iccm_stall_any,
  input         io_dma_dccm_stall_any,
  input         io_lsu_store_stall_any,
  input         io_dec_pmu_presync_stall,
  input         io_dec_pmu_postsync_stall,
  input         io_dec_pmu_decode_stall,
  input         io_ifu_pmu_fetch_stall,
  input  [1:0]  io_dec_tlu_packet_r_icaf_type,
  input  [3:0]  io_dec_tlu_packet_r_pmu_i0_itype,
  input         io_dec_tlu_packet_r_pmu_i0_br_unpred,
  input         io_dec_tlu_packet_r_pmu_divide,
  input         io_dec_tlu_packet_r_pmu_lsu_misaligned,
  input         io_exu_pmu_i0_br_ataken,
  input         io_exu_pmu_i0_br_misp,
  input         io_dec_pmu_instr_decoded,
  input         io_ifu_pmu_instr_aligned,
  input         io_exu_pmu_i0_pc4,
  input         io_ifu_pmu_ic_miss,
  input         io_ifu_pmu_ic_hit,
  output        io_dec_tlu_int_valid_wb1,
  output        io_dec_tlu_i0_exc_valid_wb1,
  output        io_dec_tlu_i0_valid_wb1,
  input         io_dec_csr_wen_r,
  output [31:0] io_dec_tlu_mtval_wb1,
  output [4:0]  io_dec_tlu_exc_cause_wb1,
  output        io_dec_tlu_perfcnt0,
  output        io_dec_tlu_perfcnt1,
  output        io_dec_tlu_perfcnt2,
  output        io_dec_tlu_perfcnt3,
  input         io_dec_tlu_dbg_halted,
  input         io_dma_pmu_dccm_write,
  input         io_dma_pmu_dccm_read,
  input         io_dma_pmu_any_write,
  input         io_dma_pmu_any_read,
  input         io_lsu_pmu_bus_busy,
  input  [30:0] io_dec_tlu_i0_pc_r,
  input         io_dec_tlu_i0_valid_r,
  input         io_dec_csr_any_unq_d,
  output        io_dec_tlu_misc_clk_override,
  output        io_dec_tlu_dec_clk_override,
  output        io_dec_tlu_lsu_clk_override,
  output        io_dec_tlu_bus_clk_override,
  output        io_dec_tlu_pic_clk_override,
  output        io_dec_tlu_dccm_clk_override,
  output        io_dec_tlu_icm_clk_override,
  output [31:0] io_dec_csr_rddata_d,
  output        io_dec_tlu_pipelining_disable,
  output        io_dec_tlu_wr_pause_r,
  input         io_ifu_pmu_bus_busy,
  input         io_lsu_pmu_bus_error,
  input         io_ifu_pmu_bus_error,
  input         io_lsu_pmu_bus_misaligned,
  input  [70:0] io_ifu_ic_debug_rd_data,
  output [3:0]  io_dec_tlu_meipt,
  input  [3:0]  io_pic_pl,
  output [3:0]  io_dec_tlu_meicurpl,
  output [29:0] io_dec_tlu_meihap,
  input  [7:0]  io_pic_claimid,
  input         io_iccm_dma_sb_error,
  input  [31:0] io_lsu_imprecise_error_addr_any,
  input         io_lsu_imprecise_error_load_any,
  input         io_lsu_imprecise_error_store_any,
  output [31:0] io_dec_tlu_mrac_ff,
  output        io_dec_tlu_wb_coalescing_disable,
  output        io_dec_tlu_bpred_disable,
  output        io_dec_tlu_sideeffect_posted_disable,
  output        io_dec_tlu_core_ecc_disable,
  output        io_dec_tlu_external_ldfwd_disable,
  output [2:0]  io_dec_tlu_dma_qos_prty,
  input  [31:0] io_dec_illegal_inst,
  input  [3:0]  io_lsu_error_pkt_r_bits_mscause,
  input         io_mexintpend,
  input  [30:0] io_exu_npc_r,
  input         io_mpc_reset_run_req,
  input  [30:0] io_rst_vec,
  input  [27:0] io_core_id,
  input  [31:0] io_dec_timer_rddata_d,
  input         io_dec_timer_read_d,
  output        io_dec_csr_wen_r_mod,
  input         io_rfpc_i0_r,
  input         io_i0_trigger_hit_r,
  output        io_fw_halt_req,
  output [1:0]  io_mstatus,
  input         io_exc_or_int_valid_r,
  input         io_mret_r,
  output        io_mstatus_mie_ns,
  input         io_dcsr_single_step_running_f,
  output [15:0] io_dcsr,
  output [30:0] io_mtvec,
  output [5:0]  io_mip,
  input         io_dec_timer_t0_pulse,
  input         io_dec_timer_t1_pulse,
  input         io_timer_int_sync,
  input         io_soft_int_sync,
  output [5:0]  io_mie_ns,
  input         io_csr_wr_clk,
  input         io_ebreak_to_debug_mode_r,
  input         io_dec_tlu_pmu_fw_halted,
  input  [1:0]  io_lsu_fir_error,
  output [30:0] io_npc_r,
  input         io_tlu_flush_lower_r_d1,
  input         io_dec_tlu_flush_noredir_r_d1,
  input  [30:0] io_tlu_flush_path_r_d1,
  output [30:0] io_npc_r_d1,
  input         io_reset_delayed,
  output [30:0] io_mepc,
  input         io_interrupt_valid_r,
  input         io_i0_exception_valid_r,
  input         io_lsu_exc_valid_r,
  input         io_mepc_trigger_hit_sel_pc_r,
  input         io_e4e5_int_clk,
  input         io_lsu_i0_exc_r,
  input         io_inst_acc_r,
  input         io_inst_acc_second_r,
  input         io_take_nmi,
  input  [31:0] io_lsu_error_pkt_addr_r,
  input  [4:0]  io_exc_cause_r,
  input         io_i0_valid_wb,
  input         io_exc_or_int_valid_r_d1,
  input         io_interrupt_valid_r_d1,
  input         io_clk_override,
  input         io_i0_exception_valid_r_d1,
  input         io_lsu_i0_exc_r_d1,
  input  [4:0]  io_exc_cause_wb,
  input         io_nmi_lsu_store_type,
  input         io_nmi_lsu_load_type,
  input         io_tlu_i0_commit_cmt,
  input         io_ebreak_r,
  input         io_ecall_r,
  input         io_illegal_r,
  output        io_mdseac_locked_ns,
  input         io_mdseac_locked_f,
  input         io_nmi_int_detected_f,
  input         io_internal_dbg_halt_mode_f2,
  input         io_ext_int_freeze_d1,
  input         io_ic_perr_r_d1,
  input         io_iccm_sbecc_r_d1,
  input         io_lsu_single_ecc_error_r_d1,
  input         io_ifu_miss_state_idle_f,
  input         io_lsu_idle_any_f,
  input         io_dbg_tlu_halted_f,
  input         io_dbg_tlu_halted,
  input         io_debug_halt_req_f,
  output        io_force_halt,
  input         io_take_ext_int_start,
  input         io_trigger_hit_dmode_r_d1,
  input         io_trigger_hit_r_d1,
  input         io_dcsr_single_step_done_f,
  input         io_ebreak_to_debug_mode_r_d1,
  input         io_debug_halt_req,
  input         io_allow_dbg_halt_csr_write,
  input         io_internal_dbg_halt_mode_f,
  input         io_enter_debug_halt_req,
  input         io_internal_dbg_halt_mode,
  input         io_request_debug_mode_done,
  input         io_request_debug_mode_r,
  output [30:0] io_dpc,
  input  [3:0]  io_update_hit_bit_r,
  input         io_take_timer_int,
  input         io_take_int_timer0_int,
  input         io_take_int_timer1_int,
  input         io_take_ext_int,
  input         io_tlu_flush_lower_r,
  input         io_dec_tlu_br0_error_r,
  input         io_dec_tlu_br0_start_error_r,
  input         io_lsu_pmu_load_external_r,
  input         io_lsu_pmu_store_external_r,
  input         io_csr_pkt_csr_misa,
  input         io_csr_pkt_csr_mvendorid,
  input         io_csr_pkt_csr_marchid,
  input         io_csr_pkt_csr_mimpid,
  input         io_csr_pkt_csr_mhartid,
  input         io_csr_pkt_csr_mstatus,
  input         io_csr_pkt_csr_mtvec,
  input         io_csr_pkt_csr_mip,
  input         io_csr_pkt_csr_mie,
  input         io_csr_pkt_csr_mcyclel,
  input         io_csr_pkt_csr_mcycleh,
  input         io_csr_pkt_csr_minstretl,
  input         io_csr_pkt_csr_minstreth,
  input         io_csr_pkt_csr_mscratch,
  input         io_csr_pkt_csr_mepc,
  input         io_csr_pkt_csr_mcause,
  input         io_csr_pkt_csr_mscause,
  input         io_csr_pkt_csr_mtval,
  input         io_csr_pkt_csr_mrac,
  input         io_csr_pkt_csr_mdseac,
  input         io_csr_pkt_csr_meihap,
  input         io_csr_pkt_csr_meivt,
  input         io_csr_pkt_csr_meipt,
  input         io_csr_pkt_csr_meicurpl,
  input         io_csr_pkt_csr_meicidpl,
  input         io_csr_pkt_csr_dcsr,
  input         io_csr_pkt_csr_mcgc,
  input         io_csr_pkt_csr_mfdc,
  input         io_csr_pkt_csr_dpc,
  input         io_csr_pkt_csr_mtsel,
  input         io_csr_pkt_csr_mtdata1,
  input         io_csr_pkt_csr_mtdata2,
  input         io_csr_pkt_csr_mhpmc3,
  input         io_csr_pkt_csr_mhpmc4,
  input         io_csr_pkt_csr_mhpmc5,
  input         io_csr_pkt_csr_mhpmc6,
  input         io_csr_pkt_csr_mhpmc3h,
  input         io_csr_pkt_csr_mhpmc4h,
  input         io_csr_pkt_csr_mhpmc5h,
  input         io_csr_pkt_csr_mhpmc6h,
  input         io_csr_pkt_csr_mhpme3,
  input         io_csr_pkt_csr_mhpme4,
  input         io_csr_pkt_csr_mhpme5,
  input         io_csr_pkt_csr_mhpme6,
  input         io_csr_pkt_csr_mcountinhibit,
  input         io_csr_pkt_csr_mpmc,
  input         io_csr_pkt_csr_micect,
  input         io_csr_pkt_csr_miccmect,
  input         io_csr_pkt_csr_mdccmect,
  input         io_csr_pkt_csr_mfdht,
  input         io_csr_pkt_csr_mfdhs,
  input         io_csr_pkt_csr_dicawics,
  input         io_csr_pkt_csr_dicad0h,
  input         io_csr_pkt_csr_dicad0,
  input         io_csr_pkt_csr_dicad1,
  output [9:0]  io_mtdata1_t_0,
  output [9:0]  io_mtdata1_t_1,
  output [9:0]  io_mtdata1_t_2,
  output [9:0]  io_mtdata1_t_3
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [95:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
`endif // RANDOMIZE_REG_INIT
  wire  rvclkhdr_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_1_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_1_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_1_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_1_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_2_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_2_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_2_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_2_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_3_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_3_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_3_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_3_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_4_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_4_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_4_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_4_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_5_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_5_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_5_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_5_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_6_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_6_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_6_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_6_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_7_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_7_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_7_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_7_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_8_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_8_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_8_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_8_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_9_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_9_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_9_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_9_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_10_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_10_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_10_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_10_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_11_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_11_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_11_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_11_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_12_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_12_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_12_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_12_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_13_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_13_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_13_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_13_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_14_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_14_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_14_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_14_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_15_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_15_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_15_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_15_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_16_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_16_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_16_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_16_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_17_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_17_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_17_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_17_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_18_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_18_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_18_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_18_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_19_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_19_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_19_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_19_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_20_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_20_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_20_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_20_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_21_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_21_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_21_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_21_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_22_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_22_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_22_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_22_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_23_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_23_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_23_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_23_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_24_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_24_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_24_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_24_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_25_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_25_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_25_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_25_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_26_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_26_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_26_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_26_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_27_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_27_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_27_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_27_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_28_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_28_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_28_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_28_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_29_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_29_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_29_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_29_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_30_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_30_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_30_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_30_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_31_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_31_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_31_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_31_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_32_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_32_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_32_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_32_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_33_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_33_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_33_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_33_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_34_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_34_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_34_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_34_io_scan_mode; // @[lib.scala 343:22]
  wire  _T = ~io_i0_trigger_hit_r; // @[dec_tlu_ctl.scala 1451:45]
  wire  _T_1 = io_dec_csr_wen_r & _T; // @[dec_tlu_ctl.scala 1451:43]
  wire  _T_2 = ~io_rfpc_i0_r; // @[dec_tlu_ctl.scala 1451:68]
  wire  _T_5 = io_dec_csr_wraddr_r == 12'h300; // @[dec_tlu_ctl.scala 1452:71]
  wire  wr_mstatus_r = io_dec_csr_wen_r_mod & _T_5; // @[dec_tlu_ctl.scala 1452:42]
  wire  _T_488 = io_dec_csr_wraddr_r == 12'h7c6; // @[dec_tlu_ctl.scala 1838:68]
  wire  wr_mpmc_r = io_dec_csr_wen_r_mod & _T_488; // @[dec_tlu_ctl.scala 1838:39]
  wire  _T_500 = ~io_dec_csr_wrdata_r[1]; // @[dec_tlu_ctl.scala 1846:37]
  reg  mpmc_b; // @[dec_tlu_ctl.scala 1848:44]
  wire  mpmc = ~mpmc_b; // @[dec_tlu_ctl.scala 1851:10]
  wire  _T_501 = ~mpmc; // @[dec_tlu_ctl.scala 1846:62]
  wire  mpmc_b_ns = wr_mpmc_r ? _T_500 : _T_501; // @[dec_tlu_ctl.scala 1846:18]
  wire  _T_6 = ~mpmc_b_ns; // @[dec_tlu_ctl.scala 1455:28]
  wire  set_mie_pmu_fw_halt = _T_6 & io_fw_halt_req; // @[dec_tlu_ctl.scala 1455:39]
  wire  _T_7 = ~wr_mstatus_r; // @[dec_tlu_ctl.scala 1458:5]
  wire  _T_8 = _T_7 & io_exc_or_int_valid_r; // @[dec_tlu_ctl.scala 1458:19]
  wire [1:0] _T_12 = {io_mstatus[0],1'h0}; // @[Cat.scala 29:58]
  wire  _T_13 = wr_mstatus_r & io_exc_or_int_valid_r; // @[dec_tlu_ctl.scala 1459:18]
  wire [1:0] _T_16 = {io_dec_csr_wrdata_r[3],1'h0}; // @[Cat.scala 29:58]
  wire  _T_17 = ~io_exc_or_int_valid_r; // @[dec_tlu_ctl.scala 1460:17]
  wire  _T_18 = io_mret_r & _T_17; // @[dec_tlu_ctl.scala 1460:15]
  wire [1:0] _T_21 = {1'h1,io_mstatus[1]}; // @[Cat.scala 29:58]
  wire [1:0] _T_24 = {io_mstatus[1],1'h1}; // @[Cat.scala 29:58]
  wire  _T_26 = wr_mstatus_r & _T_17; // @[dec_tlu_ctl.scala 1462:18]
  wire [1:0] _T_30 = {io_dec_csr_wrdata_r[7],io_dec_csr_wrdata_r[3]}; // @[Cat.scala 29:58]
  wire  _T_33 = _T_7 & _T_17; // @[dec_tlu_ctl.scala 1463:19]
  wire  _T_34 = ~io_mret_r; // @[dec_tlu_ctl.scala 1463:46]
  wire  _T_35 = _T_33 & _T_34; // @[dec_tlu_ctl.scala 1463:44]
  wire  _T_36 = ~set_mie_pmu_fw_halt; // @[dec_tlu_ctl.scala 1463:59]
  wire  _T_37 = _T_35 & _T_36; // @[dec_tlu_ctl.scala 1463:57]
  wire [1:0] _T_39 = _T_8 ? _T_12 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_40 = _T_13 ? _T_16 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_41 = _T_18 ? _T_21 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_42 = set_mie_pmu_fw_halt ? _T_24 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_43 = _T_26 ? _T_30 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_44 = _T_37 ? io_mstatus : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_45 = _T_39 | _T_40; // @[Mux.scala 27:72]
  wire [1:0] _T_46 = _T_45 | _T_41; // @[Mux.scala 27:72]
  wire [1:0] _T_47 = _T_46 | _T_42; // @[Mux.scala 27:72]
  wire [1:0] _T_48 = _T_47 | _T_43; // @[Mux.scala 27:72]
  wire  _T_52 = ~io_dcsr_single_step_running_f; // @[dec_tlu_ctl.scala 1466:50]
  wire  _T_54 = _T_52 | io_dcsr[11]; // @[dec_tlu_ctl.scala 1466:81]
  reg [1:0] _T_56; // @[dec_tlu_ctl.scala 1468:11]
  wire  _T_58 = io_dec_csr_wraddr_r == 12'h305; // @[dec_tlu_ctl.scala 1477:69]
  reg [30:0] _T_62; // @[lib.scala 374:16]
  reg [31:0] mdccmect; // @[lib.scala 374:16]
  wire [62:0] _T_564 = 63'hffffffff << mdccmect[31:27]; // @[dec_tlu_ctl.scala 1898:41]
  wire [31:0] _T_566 = {5'h0,mdccmect[26:0]}; // @[Cat.scala 29:58]
  wire [62:0] _GEN_9 = {{31'd0}, _T_566}; // @[dec_tlu_ctl.scala 1898:61]
  wire [62:0] _T_567 = _T_564 & _GEN_9; // @[dec_tlu_ctl.scala 1898:61]
  wire  mdccme_ce_req = |_T_567; // @[dec_tlu_ctl.scala 1898:94]
  reg [31:0] miccmect; // @[lib.scala 374:16]
  wire [62:0] _T_544 = 63'hffffffff << miccmect[31:27]; // @[dec_tlu_ctl.scala 1883:40]
  wire [31:0] _T_546 = {5'h0,miccmect[26:0]}; // @[Cat.scala 29:58]
  wire [62:0] _GEN_10 = {{31'd0}, _T_546}; // @[dec_tlu_ctl.scala 1883:60]
  wire [62:0] _T_547 = _T_544 & _GEN_10; // @[dec_tlu_ctl.scala 1883:60]
  wire  miccme_ce_req = |_T_547; // @[dec_tlu_ctl.scala 1883:93]
  wire  _T_63 = mdccme_ce_req | miccme_ce_req; // @[dec_tlu_ctl.scala 1491:30]
  reg [31:0] micect; // @[lib.scala 374:16]
  wire [62:0] _T_522 = 63'hffffffff << micect[31:27]; // @[dec_tlu_ctl.scala 1868:39]
  wire [31:0] _T_524 = {5'h0,micect[26:0]}; // @[Cat.scala 29:58]
  wire [62:0] _GEN_11 = {{31'd0}, _T_524}; // @[dec_tlu_ctl.scala 1868:57]
  wire [62:0] _T_525 = _T_522 & _GEN_11; // @[dec_tlu_ctl.scala 1868:57]
  wire  mice_ce_req = |_T_525; // @[dec_tlu_ctl.scala 1868:88]
  wire  ce_int = _T_63 | mice_ce_req; // @[dec_tlu_ctl.scala 1491:46]
  wire [2:0] _T_65 = {io_mexintpend,io_timer_int_sync,io_soft_int_sync}; // @[Cat.scala 29:58]
  wire [2:0] _T_67 = {ce_int,io_dec_timer_t0_pulse,io_dec_timer_t1_pulse}; // @[Cat.scala 29:58]
  reg [5:0] _T_68; // @[dec_tlu_ctl.scala 1495:11]
  wire  _T_70 = io_dec_csr_wraddr_r == 12'h304; // @[dec_tlu_ctl.scala 1507:67]
  wire  wr_mie_r = io_dec_csr_wen_r_mod & _T_70; // @[dec_tlu_ctl.scala 1507:38]
  wire [5:0] _T_78 = {io_dec_csr_wrdata_r[30:28],io_dec_csr_wrdata_r[11],io_dec_csr_wrdata_r[7],io_dec_csr_wrdata_r[3]}; // @[Cat.scala 29:58]
  reg [5:0] mie; // @[dec_tlu_ctl.scala 1510:11]
  wire  kill_ebreak_count_r = io_ebreak_to_debug_mode_r & io_dcsr[10]; // @[dec_tlu_ctl.scala 1517:54]
  wire  _T_83 = io_dec_csr_wraddr_r == 12'hb00; // @[dec_tlu_ctl.scala 1519:71]
  wire  wr_mcyclel_r = io_dec_csr_wen_r_mod & _T_83; // @[dec_tlu_ctl.scala 1519:42]
  wire  _T_85 = io_dec_tlu_dbg_halted & io_dcsr[10]; // @[dec_tlu_ctl.scala 1521:71]
  wire  _T_86 = kill_ebreak_count_r | _T_85; // @[dec_tlu_ctl.scala 1521:46]
  wire  _T_87 = _T_86 | io_dec_tlu_pmu_fw_halted; // @[dec_tlu_ctl.scala 1521:94]
  reg [4:0] temp_ncount6_2; // @[Reg.scala 27:20]
  reg  temp_ncount0; // @[Reg.scala 27:20]
  wire [6:0] mcountinhibit = {temp_ncount6_2,1'h0,temp_ncount0}; // @[Cat.scala 29:58]
  wire  _T_89 = _T_87 | mcountinhibit[0]; // @[dec_tlu_ctl.scala 1521:121]
  wire  mcyclel_cout_in = ~_T_89; // @[dec_tlu_ctl.scala 1521:24]
  wire [31:0] _T_90 = {31'h0,mcyclel_cout_in}; // @[Cat.scala 29:58]
  reg [31:0] mcyclel; // @[lib.scala 374:16]
  wire [32:0] mcyclel_inc = mcyclel + _T_90; // @[dec_tlu_ctl.scala 1525:25]
  wire  mcyclel_cout = mcyclel_inc[32]; // @[dec_tlu_ctl.scala 1527:32]
  wire  _T_101 = io_dec_csr_wraddr_r == 12'hb80; // @[dec_tlu_ctl.scala 1535:68]
  wire  wr_mcycleh_r = io_dec_csr_wen_r_mod & _T_101; // @[dec_tlu_ctl.scala 1535:39]
  wire  _T_98 = ~wr_mcycleh_r; // @[dec_tlu_ctl.scala 1529:71]
  reg  mcyclel_cout_f; // @[dec_tlu_ctl.scala 1529:54]
  wire [31:0] _T_103 = {31'h0,mcyclel_cout_f}; // @[Cat.scala 29:58]
  reg [31:0] mcycleh; // @[lib.scala 374:16]
  wire [31:0] mcycleh_inc = mcycleh + _T_103; // @[dec_tlu_ctl.scala 1537:28]
  wire  _T_109 = io_ebreak_r | io_ecall_r; // @[dec_tlu_ctl.scala 1554:72]
  wire  _T_110 = _T_109 | io_ebreak_to_debug_mode_r; // @[dec_tlu_ctl.scala 1554:85]
  wire  _T_111 = _T_110 | io_illegal_r; // @[dec_tlu_ctl.scala 1554:113]
  wire  _T_113 = _T_111 | mcountinhibit[2]; // @[dec_tlu_ctl.scala 1554:128]
  wire  _T_115 = ~_T_113; // @[dec_tlu_ctl.scala 1554:58]
  wire  i0_valid_no_ebreak_ecall_r = io_tlu_i0_commit_cmt & _T_115; // @[dec_tlu_ctl.scala 1554:56]
  wire  _T_117 = io_dec_csr_wraddr_r == 12'hb02; // @[dec_tlu_ctl.scala 1556:73]
  wire  wr_minstretl_r = io_dec_csr_wen_r_mod & _T_117; // @[dec_tlu_ctl.scala 1556:44]
  wire [31:0] _T_118 = {31'h0,i0_valid_no_ebreak_ecall_r}; // @[Cat.scala 29:58]
  reg [31:0] minstretl; // @[lib.scala 374:16]
  wire [32:0] minstretl_inc = minstretl + _T_118; // @[dec_tlu_ctl.scala 1558:29]
  wire  minstretl_cout = minstretl_inc[32]; // @[dec_tlu_ctl.scala 1559:36]
  reg  minstret_enable_f; // @[dec_tlu_ctl.scala 1564:56]
  wire  _T_128 = io_dec_csr_wraddr_r == 12'hb82; // @[dec_tlu_ctl.scala 1573:71]
  wire  wr_minstreth_r = io_dec_csr_wen_r_mod & _T_128; // @[dec_tlu_ctl.scala 1573:42]
  wire  _T_125 = ~wr_minstreth_r; // @[dec_tlu_ctl.scala 1565:75]
  reg  minstretl_cout_f; // @[dec_tlu_ctl.scala 1565:56]
  wire [31:0] _T_131 = {31'h0,minstretl_cout_f}; // @[Cat.scala 29:58]
  reg [31:0] minstreth; // @[lib.scala 374:16]
  wire [31:0] minstreth_inc = minstreth + _T_131; // @[dec_tlu_ctl.scala 1576:29]
  wire  _T_139 = io_dec_csr_wraddr_r == 12'h340; // @[dec_tlu_ctl.scala 1587:72]
  reg [31:0] mscratch; // @[lib.scala 374:16]
  wire  _T_142 = ~io_dec_tlu_dbg_halted; // @[dec_tlu_ctl.scala 1598:22]
  wire  _T_143 = ~io_tlu_flush_lower_r_d1; // @[dec_tlu_ctl.scala 1598:47]
  wire  _T_144 = _T_142 & _T_143; // @[dec_tlu_ctl.scala 1598:45]
  wire  sel_exu_npc_r = _T_144 & io_dec_tlu_i0_valid_r; // @[dec_tlu_ctl.scala 1598:72]
  wire  _T_146 = _T_142 & io_tlu_flush_lower_r_d1; // @[dec_tlu_ctl.scala 1599:47]
  wire  _T_147 = ~io_dec_tlu_flush_noredir_r_d1; // @[dec_tlu_ctl.scala 1599:75]
  wire  sel_flush_npc_r = _T_146 & _T_147; // @[dec_tlu_ctl.scala 1599:73]
  wire  _T_148 = ~sel_exu_npc_r; // @[dec_tlu_ctl.scala 1600:23]
  wire  _T_149 = ~sel_flush_npc_r; // @[dec_tlu_ctl.scala 1600:40]
  wire  sel_hold_npc_r = _T_148 & _T_149; // @[dec_tlu_ctl.scala 1600:38]
  wire  _T_151 = ~io_mpc_reset_run_req; // @[dec_tlu_ctl.scala 1604:13]
  wire  _T_152 = _T_151 & io_reset_delayed; // @[dec_tlu_ctl.scala 1604:35]
  wire [30:0] _T_156 = sel_exu_npc_r ? io_exu_npc_r : 31'h0; // @[Mux.scala 27:72]
  wire [30:0] _T_157 = _T_152 ? io_rst_vec : 31'h0; // @[Mux.scala 27:72]
  wire [30:0] _T_158 = sel_flush_npc_r ? io_tlu_flush_path_r_d1 : 31'h0; // @[Mux.scala 27:72]
  wire [30:0] _T_159 = sel_hold_npc_r ? io_npc_r_d1 : 31'h0; // @[Mux.scala 27:72]
  wire [30:0] _T_160 = _T_156 | _T_157; // @[Mux.scala 27:72]
  wire [30:0] _T_161 = _T_160 | _T_158; // @[Mux.scala 27:72]
  wire  _T_164 = sel_exu_npc_r | sel_flush_npc_r; // @[dec_tlu_ctl.scala 1608:48]
  reg [30:0] _T_167; // @[lib.scala 374:16]
  wire  pc0_valid_r = _T_142 & io_dec_tlu_i0_valid_r; // @[dec_tlu_ctl.scala 1611:44]
  wire  _T_170 = ~pc0_valid_r; // @[dec_tlu_ctl.scala 1615:22]
  wire [30:0] _T_171 = pc0_valid_r ? io_dec_tlu_i0_pc_r : 31'h0; // @[Mux.scala 27:72]
  reg [30:0] pc_r_d1; // @[lib.scala 374:16]
  wire [30:0] _T_172 = _T_170 ? pc_r_d1 : 31'h0; // @[Mux.scala 27:72]
  wire [30:0] pc_r = _T_171 | _T_172; // @[Mux.scala 27:72]
  wire  _T_176 = io_dec_csr_wraddr_r == 12'h341; // @[dec_tlu_ctl.scala 1619:68]
  wire  wr_mepc_r = io_dec_csr_wen_r_mod & _T_176; // @[dec_tlu_ctl.scala 1619:39]
  wire  _T_177 = io_i0_exception_valid_r | io_lsu_exc_valid_r; // @[dec_tlu_ctl.scala 1622:27]
  wire  _T_178 = _T_177 | io_mepc_trigger_hit_sel_pc_r; // @[dec_tlu_ctl.scala 1622:48]
  wire  _T_182 = wr_mepc_r & _T_17; // @[dec_tlu_ctl.scala 1624:13]
  wire  _T_185 = ~wr_mepc_r; // @[dec_tlu_ctl.scala 1625:3]
  wire  _T_187 = _T_185 & _T_17; // @[dec_tlu_ctl.scala 1625:14]
  wire [30:0] _T_189 = _T_178 ? pc_r : 31'h0; // @[Mux.scala 27:72]
  wire [30:0] _T_190 = io_interrupt_valid_r ? io_npc_r : 31'h0; // @[Mux.scala 27:72]
  wire [30:0] _T_191 = _T_182 ? io_dec_csr_wrdata_r[31:1] : 31'h0; // @[Mux.scala 27:72]
  wire [30:0] _T_192 = _T_187 ? io_mepc : 31'h0; // @[Mux.scala 27:72]
  wire [30:0] _T_193 = _T_189 | _T_190; // @[Mux.scala 27:72]
  wire [30:0] _T_194 = _T_193 | _T_191; // @[Mux.scala 27:72]
  reg [30:0] _T_196; // @[dec_tlu_ctl.scala 1627:47]
  wire  _T_198 = io_dec_csr_wraddr_r == 12'h342; // @[dec_tlu_ctl.scala 1634:72]
  wire  wr_mcause_r = io_dec_csr_wen_r_mod & _T_198; // @[dec_tlu_ctl.scala 1634:43]
  wire  _T_199 = io_exc_or_int_valid_r & io_take_nmi; // @[dec_tlu_ctl.scala 1635:53]
  wire  mcause_sel_nmi_store = _T_199 & io_nmi_lsu_store_type; // @[dec_tlu_ctl.scala 1635:67]
  wire  mcause_sel_nmi_load = _T_199 & io_nmi_lsu_load_type; // @[dec_tlu_ctl.scala 1636:66]
  wire  _T_202 = |io_lsu_fir_error; // @[dec_tlu_ctl.scala 1637:84]
  wire  mcause_sel_nmi_ext = _T_199 & _T_202; // @[dec_tlu_ctl.scala 1637:65]
  wire  _T_203 = &io_lsu_fir_error; // @[dec_tlu_ctl.scala 1643:53]
  wire  _T_206 = ~io_lsu_fir_error[0]; // @[dec_tlu_ctl.scala 1643:82]
  wire  _T_207 = io_lsu_fir_error[1] & _T_206; // @[dec_tlu_ctl.scala 1643:80]
  wire [31:0] _T_212 = {30'h3c000400,_T_203,_T_207}; // @[Cat.scala 29:58]
  wire  _T_213 = ~io_take_nmi; // @[dec_tlu_ctl.scala 1649:56]
  wire  _T_214 = io_exc_or_int_valid_r & _T_213; // @[dec_tlu_ctl.scala 1649:54]
  wire [31:0] _T_217 = {io_interrupt_valid_r,26'h0,io_exc_cause_r}; // @[Cat.scala 29:58]
  wire  _T_219 = wr_mcause_r & _T_17; // @[dec_tlu_ctl.scala 1650:44]
  wire  _T_221 = ~wr_mcause_r; // @[dec_tlu_ctl.scala 1651:32]
  wire  _T_223 = _T_221 & _T_17; // @[dec_tlu_ctl.scala 1651:45]
  wire [31:0] _T_225 = mcause_sel_nmi_store ? 32'hf0000000 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_226 = mcause_sel_nmi_load ? 32'hf0000001 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_227 = mcause_sel_nmi_ext ? _T_212 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_228 = _T_214 ? _T_217 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_229 = _T_219 ? io_dec_csr_wrdata_r : 32'h0; // @[Mux.scala 27:72]
  reg [31:0] mcause; // @[dec_tlu_ctl.scala 1653:49]
  wire [31:0] _T_230 = _T_223 ? mcause : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_231 = _T_225 | _T_226; // @[Mux.scala 27:72]
  wire [31:0] _T_232 = _T_231 | _T_227; // @[Mux.scala 27:72]
  wire [31:0] _T_233 = _T_232 | _T_228; // @[Mux.scala 27:72]
  wire [31:0] _T_234 = _T_233 | _T_229; // @[Mux.scala 27:72]
  wire  _T_238 = io_dec_csr_wraddr_r == 12'h7ff; // @[dec_tlu_ctl.scala 1660:71]
  wire  wr_mscause_r = io_dec_csr_wen_r_mod & _T_238; // @[dec_tlu_ctl.scala 1660:42]
  wire  _T_239 = io_dec_tlu_packet_r_icaf_type == 2'h0; // @[dec_tlu_ctl.scala 1662:56]
  wire [3:0] _T_240 = {2'h0,io_dec_tlu_packet_r_icaf_type}; // @[Cat.scala 29:58]
  wire [3:0] ifu_mscause = _T_239 ? 4'h9 : _T_240; // @[dec_tlu_ctl.scala 1662:24]
  wire [3:0] _T_245 = io_lsu_i0_exc_r ? io_lsu_error_pkt_r_bits_mscause : 4'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_247 = io_ebreak_r ? 2'h2 : 2'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_248 = io_inst_acc_r ? ifu_mscause : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _GEN_12 = {{3'd0}, io_i0_trigger_hit_r}; // @[Mux.scala 27:72]
  wire [3:0] _T_249 = _T_245 | _GEN_12; // @[Mux.scala 27:72]
  wire [3:0] _GEN_13 = {{2'd0}, _T_247}; // @[Mux.scala 27:72]
  wire [3:0] _T_250 = _T_249 | _GEN_13; // @[Mux.scala 27:72]
  wire [3:0] mscause_type = _T_250 | _T_248; // @[Mux.scala 27:72]
  wire  _T_254 = wr_mscause_r & _T_17; // @[dec_tlu_ctl.scala 1673:38]
  wire  _T_257 = ~wr_mscause_r; // @[dec_tlu_ctl.scala 1674:25]
  wire  _T_259 = _T_257 & _T_17; // @[dec_tlu_ctl.scala 1674:39]
  wire [3:0] _T_261 = io_exc_or_int_valid_r ? mscause_type : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_262 = _T_254 ? io_dec_csr_wrdata_r[3:0] : 4'h0; // @[Mux.scala 27:72]
  reg [3:0] mscause; // @[dec_tlu_ctl.scala 1676:47]
  wire [3:0] _T_263 = _T_259 ? mscause : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_264 = _T_261 | _T_262; // @[Mux.scala 27:72]
  wire  _T_268 = io_dec_csr_wraddr_r == 12'h343; // @[dec_tlu_ctl.scala 1683:69]
  wire  wr_mtval_r = io_dec_csr_wen_r_mod & _T_268; // @[dec_tlu_ctl.scala 1683:40]
  wire  _T_269 = ~io_inst_acc_second_r; // @[dec_tlu_ctl.scala 1684:83]
  wire  _T_270 = io_inst_acc_r & _T_269; // @[dec_tlu_ctl.scala 1684:81]
  wire  _T_271 = io_ebreak_r | _T_270; // @[dec_tlu_ctl.scala 1684:64]
  wire  _T_272 = _T_271 | io_mepc_trigger_hit_sel_pc_r; // @[dec_tlu_ctl.scala 1684:106]
  wire  _T_273 = io_exc_or_int_valid_r & _T_272; // @[dec_tlu_ctl.scala 1684:49]
  wire  mtval_capture_pc_r = _T_273 & _T_213; // @[dec_tlu_ctl.scala 1684:138]
  wire  _T_275 = io_inst_acc_r & io_inst_acc_second_r; // @[dec_tlu_ctl.scala 1685:72]
  wire  _T_276 = io_exc_or_int_valid_r & _T_275; // @[dec_tlu_ctl.scala 1685:55]
  wire  mtval_capture_pc_plus2_r = _T_276 & _T_213; // @[dec_tlu_ctl.scala 1685:96]
  wire  _T_278 = io_exc_or_int_valid_r & io_illegal_r; // @[dec_tlu_ctl.scala 1686:51]
  wire  mtval_capture_inst_r = _T_278 & _T_213; // @[dec_tlu_ctl.scala 1686:66]
  wire  _T_280 = io_exc_or_int_valid_r & io_lsu_exc_valid_r; // @[dec_tlu_ctl.scala 1687:50]
  wire  mtval_capture_lsu_r = _T_280 & _T_213; // @[dec_tlu_ctl.scala 1687:71]
  wire  _T_282 = ~mtval_capture_pc_r; // @[dec_tlu_ctl.scala 1688:46]
  wire  _T_283 = io_exc_or_int_valid_r & _T_282; // @[dec_tlu_ctl.scala 1688:44]
  wire  _T_284 = ~mtval_capture_inst_r; // @[dec_tlu_ctl.scala 1688:68]
  wire  _T_285 = _T_283 & _T_284; // @[dec_tlu_ctl.scala 1688:66]
  wire  _T_286 = ~mtval_capture_lsu_r; // @[dec_tlu_ctl.scala 1688:92]
  wire  _T_287 = _T_285 & _T_286; // @[dec_tlu_ctl.scala 1688:90]
  wire  _T_288 = ~io_mepc_trigger_hit_sel_pc_r; // @[dec_tlu_ctl.scala 1688:115]
  wire  mtval_clear_r = _T_287 & _T_288; // @[dec_tlu_ctl.scala 1688:113]
  wire [31:0] _T_290 = {pc_r,1'h0}; // @[Cat.scala 29:58]
  wire [30:0] _T_293 = pc_r + 31'h1; // @[dec_tlu_ctl.scala 1693:83]
  wire [31:0] _T_294 = {_T_293,1'h0}; // @[Cat.scala 29:58]
  wire  _T_297 = ~io_interrupt_valid_r; // @[dec_tlu_ctl.scala 1696:18]
  wire  _T_298 = wr_mtval_r & _T_297; // @[dec_tlu_ctl.scala 1696:16]
  wire  _T_301 = ~wr_mtval_r; // @[dec_tlu_ctl.scala 1697:20]
  wire  _T_302 = _T_213 & _T_301; // @[dec_tlu_ctl.scala 1697:18]
  wire  _T_304 = _T_302 & _T_282; // @[dec_tlu_ctl.scala 1697:32]
  wire  _T_306 = _T_304 & _T_284; // @[dec_tlu_ctl.scala 1697:54]
  wire  _T_307 = ~mtval_clear_r; // @[dec_tlu_ctl.scala 1697:80]
  wire  _T_308 = _T_306 & _T_307; // @[dec_tlu_ctl.scala 1697:78]
  wire  _T_310 = _T_308 & _T_286; // @[dec_tlu_ctl.scala 1697:95]
  wire [31:0] _T_312 = mtval_capture_pc_r ? _T_290 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_313 = mtval_capture_pc_plus2_r ? _T_294 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_314 = mtval_capture_inst_r ? io_dec_illegal_inst : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_315 = mtval_capture_lsu_r ? io_lsu_error_pkt_addr_r : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_316 = _T_298 ? io_dec_csr_wrdata_r : 32'h0; // @[Mux.scala 27:72]
  reg [31:0] mtval; // @[dec_tlu_ctl.scala 1699:46]
  wire [31:0] _T_317 = _T_310 ? mtval : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_318 = _T_312 | _T_313; // @[Mux.scala 27:72]
  wire [31:0] _T_319 = _T_318 | _T_314; // @[Mux.scala 27:72]
  wire [31:0] _T_320 = _T_319 | _T_315; // @[Mux.scala 27:72]
  wire [31:0] _T_321 = _T_320 | _T_316; // @[Mux.scala 27:72]
  wire  _T_325 = io_dec_csr_wraddr_r == 12'h7f8; // @[dec_tlu_ctl.scala 1714:68]
  reg [8:0] mcgc; // @[lib.scala 374:16]
  wire  _T_337 = io_dec_csr_wraddr_r == 12'h7f9; // @[dec_tlu_ctl.scala 1744:68]
  reg [14:0] mfdc_int; // @[lib.scala 374:16]
  wire [2:0] _T_341 = ~io_dec_csr_wrdata_r[18:16]; // @[dec_tlu_ctl.scala 1757:19]
  wire [2:0] _T_345 = ~mfdc_int[14:12]; // @[dec_tlu_ctl.scala 1758:19]
  wire [18:0] mfdc = {_T_345,4'h0,mfdc_int[11:0]}; // @[Cat.scala 29:58]
  wire  _T_357 = io_dec_csr_wraddr_r == 12'h7c2; // @[dec_tlu_ctl.scala 1777:77]
  wire  _T_358 = io_dec_csr_wen_r_mod & _T_357; // @[dec_tlu_ctl.scala 1777:48]
  wire  _T_360 = _T_358 & _T_297; // @[dec_tlu_ctl.scala 1777:87]
  wire  _T_361 = ~io_take_ext_int_start; // @[dec_tlu_ctl.scala 1777:113]
  wire  _T_364 = io_dec_csr_wraddr_r == 12'h7c0; // @[dec_tlu_ctl.scala 1784:68]
  wire  _T_368 = ~io_dec_csr_wrdata_r[31]; // @[dec_tlu_ctl.scala 1787:71]
  wire  _T_369 = io_dec_csr_wrdata_r[30] & _T_368; // @[dec_tlu_ctl.scala 1787:69]
  wire  _T_373 = ~io_dec_csr_wrdata_r[29]; // @[dec_tlu_ctl.scala 1788:73]
  wire  _T_374 = io_dec_csr_wrdata_r[28] & _T_373; // @[dec_tlu_ctl.scala 1788:71]
  wire  _T_378 = ~io_dec_csr_wrdata_r[27]; // @[dec_tlu_ctl.scala 1789:73]
  wire  _T_379 = io_dec_csr_wrdata_r[26] & _T_378; // @[dec_tlu_ctl.scala 1789:71]
  wire  _T_383 = ~io_dec_csr_wrdata_r[25]; // @[dec_tlu_ctl.scala 1790:73]
  wire  _T_384 = io_dec_csr_wrdata_r[24] & _T_383; // @[dec_tlu_ctl.scala 1790:71]
  wire  _T_388 = ~io_dec_csr_wrdata_r[23]; // @[dec_tlu_ctl.scala 1791:73]
  wire  _T_389 = io_dec_csr_wrdata_r[22] & _T_388; // @[dec_tlu_ctl.scala 1791:71]
  wire  _T_393 = ~io_dec_csr_wrdata_r[21]; // @[dec_tlu_ctl.scala 1792:73]
  wire  _T_394 = io_dec_csr_wrdata_r[20] & _T_393; // @[dec_tlu_ctl.scala 1792:71]
  wire  _T_398 = ~io_dec_csr_wrdata_r[19]; // @[dec_tlu_ctl.scala 1793:73]
  wire  _T_399 = io_dec_csr_wrdata_r[18] & _T_398; // @[dec_tlu_ctl.scala 1793:71]
  wire  _T_403 = ~io_dec_csr_wrdata_r[17]; // @[dec_tlu_ctl.scala 1794:73]
  wire  _T_404 = io_dec_csr_wrdata_r[16] & _T_403; // @[dec_tlu_ctl.scala 1794:71]
  wire  _T_408 = ~io_dec_csr_wrdata_r[15]; // @[dec_tlu_ctl.scala 1795:73]
  wire  _T_409 = io_dec_csr_wrdata_r[14] & _T_408; // @[dec_tlu_ctl.scala 1795:71]
  wire  _T_413 = ~io_dec_csr_wrdata_r[13]; // @[dec_tlu_ctl.scala 1796:73]
  wire  _T_414 = io_dec_csr_wrdata_r[12] & _T_413; // @[dec_tlu_ctl.scala 1796:71]
  wire  _T_418 = ~io_dec_csr_wrdata_r[11]; // @[dec_tlu_ctl.scala 1797:73]
  wire  _T_419 = io_dec_csr_wrdata_r[10] & _T_418; // @[dec_tlu_ctl.scala 1797:71]
  wire  _T_423 = ~io_dec_csr_wrdata_r[9]; // @[dec_tlu_ctl.scala 1798:73]
  wire  _T_424 = io_dec_csr_wrdata_r[8] & _T_423; // @[dec_tlu_ctl.scala 1798:70]
  wire  _T_428 = ~io_dec_csr_wrdata_r[7]; // @[dec_tlu_ctl.scala 1799:73]
  wire  _T_429 = io_dec_csr_wrdata_r[6] & _T_428; // @[dec_tlu_ctl.scala 1799:70]
  wire  _T_433 = ~io_dec_csr_wrdata_r[5]; // @[dec_tlu_ctl.scala 1800:73]
  wire  _T_434 = io_dec_csr_wrdata_r[4] & _T_433; // @[dec_tlu_ctl.scala 1800:70]
  wire  _T_438 = ~io_dec_csr_wrdata_r[3]; // @[dec_tlu_ctl.scala 1801:73]
  wire  _T_439 = io_dec_csr_wrdata_r[2] & _T_438; // @[dec_tlu_ctl.scala 1801:70]
  wire  _T_444 = io_dec_csr_wrdata_r[0] & _T_500; // @[dec_tlu_ctl.scala 1802:70]
  wire [7:0] _T_451 = {io_dec_csr_wrdata_r[7],_T_429,io_dec_csr_wrdata_r[5],_T_434,io_dec_csr_wrdata_r[3],_T_439,io_dec_csr_wrdata_r[1],_T_444}; // @[Cat.scala 29:58]
  wire [15:0] _T_459 = {io_dec_csr_wrdata_r[15],_T_409,io_dec_csr_wrdata_r[13],_T_414,io_dec_csr_wrdata_r[11],_T_419,io_dec_csr_wrdata_r[9],_T_424,_T_451}; // @[Cat.scala 29:58]
  wire [7:0] _T_466 = {io_dec_csr_wrdata_r[23],_T_389,io_dec_csr_wrdata_r[21],_T_394,io_dec_csr_wrdata_r[19],_T_399,io_dec_csr_wrdata_r[17],_T_404}; // @[Cat.scala 29:58]
  wire [15:0] _T_474 = {io_dec_csr_wrdata_r[31],_T_369,io_dec_csr_wrdata_r[29],_T_374,io_dec_csr_wrdata_r[27],_T_379,io_dec_csr_wrdata_r[25],_T_384,_T_466}; // @[Cat.scala 29:58]
  reg [31:0] mrac; // @[lib.scala 374:16]
  wire  _T_477 = io_dec_csr_wraddr_r == 12'hbc0; // @[dec_tlu_ctl.scala 1815:69]
  wire  wr_mdeau_r = io_dec_csr_wen_r_mod & _T_477; // @[dec_tlu_ctl.scala 1815:40]
  wire  _T_478 = ~wr_mdeau_r; // @[dec_tlu_ctl.scala 1825:59]
  wire  _T_479 = io_mdseac_locked_f & _T_478; // @[dec_tlu_ctl.scala 1825:57]
  wire  _T_481 = io_lsu_imprecise_error_store_any | io_lsu_imprecise_error_load_any; // @[dec_tlu_ctl.scala 1827:49]
  wire  _T_482 = ~io_nmi_int_detected_f; // @[dec_tlu_ctl.scala 1827:86]
  wire  _T_483 = _T_481 & _T_482; // @[dec_tlu_ctl.scala 1827:84]
  wire  _T_484 = ~io_mdseac_locked_f; // @[dec_tlu_ctl.scala 1827:111]
  wire  mdseac_en = _T_483 & _T_484; // @[dec_tlu_ctl.scala 1827:109]
  reg [31:0] mdseac; // @[lib.scala 374:16]
  wire  _T_490 = wr_mpmc_r & io_dec_csr_wrdata_r[0]; // @[dec_tlu_ctl.scala 1842:30]
  wire  _T_491 = ~io_internal_dbg_halt_mode_f2; // @[dec_tlu_ctl.scala 1842:57]
  wire  _T_492 = _T_490 & _T_491; // @[dec_tlu_ctl.scala 1842:55]
  wire  _T_493 = ~io_ext_int_freeze_d1; // @[dec_tlu_ctl.scala 1842:89]
  wire  _T_506 = io_dec_csr_wrdata_r[31:27] > 5'h1a; // @[dec_tlu_ctl.scala 1860:48]
  wire [4:0] csr_sat = _T_506 ? 5'h1a : io_dec_csr_wrdata_r[31:27]; // @[dec_tlu_ctl.scala 1860:19]
  wire  _T_509 = io_dec_csr_wraddr_r == 12'h7f0; // @[dec_tlu_ctl.scala 1862:70]
  wire  wr_micect_r = io_dec_csr_wen_r_mod & _T_509; // @[dec_tlu_ctl.scala 1862:41]
  wire [26:0] _T_510 = {26'h0,io_ic_perr_r_d1}; // @[Cat.scala 29:58]
  wire [31:0] _GEN_14 = {{5'd0}, _T_510}; // @[dec_tlu_ctl.scala 1863:23]
  wire [31:0] _T_512 = micect + _GEN_14; // @[dec_tlu_ctl.scala 1863:23]
  wire [31:0] _T_515 = {csr_sat,io_dec_csr_wrdata_r[26:0]}; // @[Cat.scala 29:58]
  wire [26:0] micect_inc = _T_512[26:0]; // @[dec_tlu_ctl.scala 1863:13]
  wire [31:0] _T_517 = {micect[31:27],micect_inc}; // @[Cat.scala 29:58]
  wire  _T_528 = io_dec_csr_wraddr_r == 12'h7f1; // @[dec_tlu_ctl.scala 1877:76]
  wire  wr_miccmect_r = io_dec_csr_wen_r_mod & _T_528; // @[dec_tlu_ctl.scala 1877:47]
  wire  _T_530 = io_iccm_sbecc_r_d1 | io_iccm_dma_sb_error; // @[dec_tlu_ctl.scala 1878:70]
  wire [26:0] _T_531 = {26'h0,_T_530}; // @[Cat.scala 29:58]
  wire [26:0] miccmect_inc = miccmect[26:0] + _T_531; // @[dec_tlu_ctl.scala 1878:33]
  wire [31:0] _T_538 = {miccmect[31:27],miccmect_inc}; // @[Cat.scala 29:58]
  wire  _T_539 = wr_miccmect_r | io_iccm_sbecc_r_d1; // @[dec_tlu_ctl.scala 1881:48]
  wire  _T_550 = io_dec_csr_wraddr_r == 12'h7f2; // @[dec_tlu_ctl.scala 1892:76]
  wire  wr_mdccmect_r = io_dec_csr_wen_r_mod & _T_550; // @[dec_tlu_ctl.scala 1892:47]
  wire [26:0] _T_552 = {26'h0,io_lsu_single_ecc_error_r_d1}; // @[Cat.scala 29:58]
  wire [26:0] mdccmect_inc = mdccmect[26:0] + _T_552; // @[dec_tlu_ctl.scala 1893:33]
  wire [31:0] _T_559 = {mdccmect[31:27],mdccmect_inc}; // @[Cat.scala 29:58]
  wire  _T_570 = io_dec_csr_wraddr_r == 12'h7ce; // @[dec_tlu_ctl.scala 1908:69]
  wire  wr_mfdht_r = io_dec_csr_wen_r_mod & _T_570; // @[dec_tlu_ctl.scala 1908:40]
  reg [5:0] mfdht; // @[dec_tlu_ctl.scala 1912:43]
  wire  _T_575 = io_dec_csr_wraddr_r == 12'h7cf; // @[dec_tlu_ctl.scala 1921:69]
  wire  wr_mfdhs_r = io_dec_csr_wen_r_mod & _T_575; // @[dec_tlu_ctl.scala 1921:40]
  wire  _T_578 = ~io_dbg_tlu_halted_f; // @[dec_tlu_ctl.scala 1924:43]
  wire  _T_579 = io_dbg_tlu_halted & _T_578; // @[dec_tlu_ctl.scala 1924:41]
  wire  _T_581 = ~io_lsu_idle_any_f; // @[dec_tlu_ctl.scala 1924:78]
  wire  _T_582 = ~io_ifu_miss_state_idle_f; // @[dec_tlu_ctl.scala 1924:98]
  wire [1:0] _T_583 = {_T_581,_T_582}; // @[Cat.scala 29:58]
  reg [1:0] mfdhs; // @[Reg.scala 27:20]
  wire  _T_585 = wr_mfdhs_r | io_dbg_tlu_halted; // @[dec_tlu_ctl.scala 1926:71]
  reg [31:0] force_halt_ctr_f; // @[Reg.scala 27:20]
  wire [31:0] _T_590 = force_halt_ctr_f + 32'h1; // @[dec_tlu_ctl.scala 1928:74]
  wire [62:0] _T_597 = 63'hffffffff << mfdht[5:1]; // @[dec_tlu_ctl.scala 1933:71]
  wire [62:0] _GEN_15 = {{31'd0}, force_halt_ctr_f}; // @[dec_tlu_ctl.scala 1933:48]
  wire [62:0] _T_598 = _GEN_15 & _T_597; // @[dec_tlu_ctl.scala 1933:48]
  wire  _T_599 = |_T_598; // @[dec_tlu_ctl.scala 1933:87]
  wire  _T_602 = io_dec_csr_wraddr_r == 12'hbc8; // @[dec_tlu_ctl.scala 1941:69]
  reg [21:0] meivt; // @[lib.scala 374:16]
  wire  _T_621 = io_dec_csr_wraddr_r == 12'hbca; // @[dec_tlu_ctl.scala 1992:69]
  wire  _T_622 = io_dec_csr_wen_r_mod & _T_621; // @[dec_tlu_ctl.scala 1992:40]
  wire  wr_meicpct_r = _T_622 | io_take_ext_int_start; // @[dec_tlu_ctl.scala 1992:83]
  reg [7:0] meihap; // @[lib.scala 374:16]
  wire  _T_608 = io_dec_csr_wraddr_r == 12'hbcc; // @[dec_tlu_ctl.scala 1965:72]
  wire  wr_meicurpl_r = io_dec_csr_wen_r_mod & _T_608; // @[dec_tlu_ctl.scala 1965:43]
  reg [3:0] meicurpl; // @[dec_tlu_ctl.scala 1968:46]
  wire  _T_613 = io_dec_csr_wraddr_r == 12'hbcb; // @[dec_tlu_ctl.scala 1980:73]
  wire  _T_614 = io_dec_csr_wen_r_mod & _T_613; // @[dec_tlu_ctl.scala 1980:44]
  wire  wr_meicidpl_r = _T_614 | io_take_ext_int_start; // @[dec_tlu_ctl.scala 1980:88]
  reg [3:0] meicidpl; // @[dec_tlu_ctl.scala 1985:44]
  wire  _T_625 = io_dec_csr_wraddr_r == 12'hbc9; // @[dec_tlu_ctl.scala 2001:69]
  wire  wr_meipt_r = io_dec_csr_wen_r_mod & _T_625; // @[dec_tlu_ctl.scala 2001:40]
  reg [3:0] meipt; // @[dec_tlu_ctl.scala 2004:43]
  wire  _T_629 = io_trigger_hit_r_d1 & io_dcsr_single_step_done_f; // @[dec_tlu_ctl.scala 2032:89]
  wire  trigger_hit_for_dscr_cause_r_d1 = io_trigger_hit_dmode_r_d1 | _T_629; // @[dec_tlu_ctl.scala 2032:66]
  wire  _T_630 = ~io_ebreak_to_debug_mode_r_d1; // @[dec_tlu_ctl.scala 2035:31]
  wire  _T_631 = io_dcsr_single_step_done_f & _T_630; // @[dec_tlu_ctl.scala 2035:29]
  wire  _T_632 = ~trigger_hit_for_dscr_cause_r_d1; // @[dec_tlu_ctl.scala 2035:63]
  wire  _T_633 = _T_631 & _T_632; // @[dec_tlu_ctl.scala 2035:61]
  wire  _T_634 = ~io_debug_halt_req; // @[dec_tlu_ctl.scala 2035:98]
  wire  _T_635 = _T_633 & _T_634; // @[dec_tlu_ctl.scala 2035:96]
  wire  _T_638 = io_debug_halt_req & _T_630; // @[dec_tlu_ctl.scala 2036:46]
  wire  _T_640 = _T_638 & _T_632; // @[dec_tlu_ctl.scala 2036:78]
  wire  _T_643 = io_ebreak_to_debug_mode_r_d1 & _T_632; // @[dec_tlu_ctl.scala 2037:75]
  wire [2:0] _T_646 = _T_635 ? 3'h4 : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_647 = _T_640 ? 3'h3 : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_648 = _T_643 ? 3'h1 : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_649 = trigger_hit_for_dscr_cause_r_d1 ? 3'h2 : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_650 = _T_646 | _T_647; // @[Mux.scala 27:72]
  wire [2:0] _T_651 = _T_650 | _T_648; // @[Mux.scala 27:72]
  wire [2:0] dcsr_cause = _T_651 | _T_649; // @[Mux.scala 27:72]
  wire  _T_653 = io_allow_dbg_halt_csr_write & io_dec_csr_wen_r_mod; // @[dec_tlu_ctl.scala 2040:46]
  wire  _T_655 = io_dec_csr_wraddr_r == 12'h7b0; // @[dec_tlu_ctl.scala 2040:98]
  wire  wr_dcsr_r = _T_653 & _T_655; // @[dec_tlu_ctl.scala 2040:69]
  wire  _T_657 = io_dcsr[8:6] == 3'h3; // @[dec_tlu_ctl.scala 2046:75]
  wire  dcsr_cause_upgradeable = io_internal_dbg_halt_mode_f & _T_657; // @[dec_tlu_ctl.scala 2046:59]
  wire  _T_658 = ~io_dbg_tlu_halted; // @[dec_tlu_ctl.scala 2047:59]
  wire  _T_659 = _T_658 | dcsr_cause_upgradeable; // @[dec_tlu_ctl.scala 2047:78]
  wire  enter_debug_halt_req_le = io_enter_debug_halt_req & _T_659; // @[dec_tlu_ctl.scala 2047:56]
  wire  nmi_in_debug_mode = io_nmi_int_detected_f & io_internal_dbg_halt_mode_f; // @[dec_tlu_ctl.scala 2049:48]
  wire [15:0] _T_665 = {io_dcsr[15:9],dcsr_cause,io_dcsr[5:2],2'h3}; // @[Cat.scala 29:58]
  wire  _T_671 = nmi_in_debug_mode | io_dcsr[3]; // @[dec_tlu_ctl.scala 2051:145]
  wire [15:0] _T_680 = {io_dec_csr_wrdata_r[15],3'h0,io_dec_csr_wrdata_r[11:10],1'h0,io_dcsr[8:6],2'h0,_T_671,io_dec_csr_wrdata_r[2],2'h3}; // @[Cat.scala 29:58]
  wire [15:0] _T_685 = {io_dcsr[15:4],nmi_in_debug_mode,io_dcsr[2],2'h3}; // @[Cat.scala 29:58]
  wire  _T_687 = enter_debug_halt_req_le | wr_dcsr_r; // @[dec_tlu_ctl.scala 2053:54]
  wire  _T_688 = _T_687 | io_internal_dbg_halt_mode; // @[dec_tlu_ctl.scala 2053:66]
  reg [15:0] _T_691; // @[lib.scala 374:16]
  wire  _T_694 = io_dec_csr_wraddr_r == 12'h7b1; // @[dec_tlu_ctl.scala 2061:97]
  wire  wr_dpc_r = _T_653 & _T_694; // @[dec_tlu_ctl.scala 2061:68]
  wire  _T_697 = ~io_request_debug_mode_done; // @[dec_tlu_ctl.scala 2062:67]
  wire  dpc_capture_npc = _T_579 & _T_697; // @[dec_tlu_ctl.scala 2062:65]
  wire  _T_698 = ~io_request_debug_mode_r; // @[dec_tlu_ctl.scala 2066:21]
  wire  _T_699 = ~dpc_capture_npc; // @[dec_tlu_ctl.scala 2066:39]
  wire  _T_700 = _T_698 & _T_699; // @[dec_tlu_ctl.scala 2066:37]
  wire  _T_701 = _T_700 & wr_dpc_r; // @[dec_tlu_ctl.scala 2066:56]
  wire  _T_706 = _T_698 & dpc_capture_npc; // @[dec_tlu_ctl.scala 2068:49]
  wire [30:0] _T_708 = _T_701 ? io_dec_csr_wrdata_r[31:1] : 31'h0; // @[Mux.scala 27:72]
  wire [30:0] _T_709 = io_request_debug_mode_r ? pc_r : 31'h0; // @[Mux.scala 27:72]
  wire [30:0] _T_710 = _T_706 ? io_npc_r : 31'h0; // @[Mux.scala 27:72]
  wire [30:0] _T_711 = _T_708 | _T_709; // @[Mux.scala 27:72]
  wire  _T_713 = wr_dpc_r | io_request_debug_mode_r; // @[dec_tlu_ctl.scala 2070:36]
  reg [30:0] _T_716; // @[lib.scala 374:16]
  wire [2:0] _T_720 = {io_dec_csr_wrdata_r[24],io_dec_csr_wrdata_r[21:20]}; // @[Cat.scala 29:58]
  wire  _T_723 = io_dec_csr_wraddr_r == 12'h7c8; // @[dec_tlu_ctl.scala 2085:102]
  reg [16:0] dicawics; // @[lib.scala 374:16]
  wire  _T_727 = io_dec_csr_wraddr_r == 12'h7c9; // @[dec_tlu_ctl.scala 2103:100]
  wire  wr_dicad0_r = _T_653 & _T_727; // @[dec_tlu_ctl.scala 2103:71]
  reg [70:0] dicad0; // @[lib.scala 374:16]
  wire  _T_733 = io_dec_csr_wraddr_r == 12'h7cc; // @[dec_tlu_ctl.scala 2116:101]
  wire  wr_dicad0h_r = _T_653 & _T_733; // @[dec_tlu_ctl.scala 2116:72]
  reg [31:0] dicad0h; // @[lib.scala 374:16]
  wire  _T_741 = io_dec_csr_wraddr_r == 12'h7ca; // @[dec_tlu_ctl.scala 2128:100]
  wire  _T_742 = _T_653 & _T_741; // @[dec_tlu_ctl.scala 2128:71]
  wire  _T_747 = _T_742 | io_ifu_ic_debug_rd_data_valid; // @[dec_tlu_ctl.scala 2132:78]
  reg [6:0] _T_749; // @[Reg.scala 27:20]
  wire [31:0] dicad1 = {25'h0,_T_749}; // @[Cat.scala 29:58]
  wire [38:0] _T_754 = {dicad1[6:0],dicad0h}; // @[Cat.scala 29:58]
  wire  _T_756 = io_allow_dbg_halt_csr_write & io_dec_csr_any_unq_d; // @[dec_tlu_ctl.scala 2160:52]
  wire  _T_757 = _T_756 & io_dec_i0_decode_d; // @[dec_tlu_ctl.scala 2160:75]
  wire  _T_758 = ~io_dec_csr_wen_unq_d; // @[dec_tlu_ctl.scala 2160:98]
  wire  _T_759 = _T_757 & _T_758; // @[dec_tlu_ctl.scala 2160:96]
  wire  _T_761 = io_dec_csr_rdaddr_d == 12'h7cb; // @[dec_tlu_ctl.scala 2160:149]
  wire  _T_764 = io_dec_csr_wraddr_r == 12'h7cb; // @[dec_tlu_ctl.scala 2161:104]
  reg  icache_rd_valid_f; // @[dec_tlu_ctl.scala 2163:58]
  reg  icache_wr_valid_f; // @[dec_tlu_ctl.scala 2164:58]
  wire  _T_766 = io_dec_csr_wraddr_r == 12'h7a0; // @[dec_tlu_ctl.scala 2175:69]
  wire  wr_mtsel_r = io_dec_csr_wen_r_mod & _T_766; // @[dec_tlu_ctl.scala 2175:40]
  reg [1:0] mtsel; // @[dec_tlu_ctl.scala 2178:43]
  wire  tdata_load = io_dec_csr_wrdata_r[0] & _T_398; // @[dec_tlu_ctl.scala 2213:42]
  wire  tdata_opcode = io_dec_csr_wrdata_r[2] & _T_398; // @[dec_tlu_ctl.scala 2215:44]
  wire  _T_777 = io_dec_csr_wrdata_r[27] & io_dbg_tlu_halted_f; // @[dec_tlu_ctl.scala 2217:46]
  wire  tdata_action = _T_777 & io_dec_csr_wrdata_r[12]; // @[dec_tlu_ctl.scala 2217:69]
  wire [9:0] tdata_wrdata_r = {_T_777,io_dec_csr_wrdata_r[20:19],tdata_action,io_dec_csr_wrdata_r[11],io_dec_csr_wrdata_r[7:6],tdata_opcode,io_dec_csr_wrdata_r[1],tdata_load}; // @[Cat.scala 29:58]
  wire  _T_792 = io_dec_csr_wraddr_r == 12'h7a1; // @[dec_tlu_ctl.scala 2223:99]
  wire  _T_793 = io_dec_csr_wen_r_mod & _T_792; // @[dec_tlu_ctl.scala 2223:70]
  wire  _T_794 = mtsel == 2'h0; // @[dec_tlu_ctl.scala 2223:121]
  wire  _T_795 = _T_793 & _T_794; // @[dec_tlu_ctl.scala 2223:112]
  wire  _T_797 = ~io_mtdata1_t_0[9]; // @[dec_tlu_ctl.scala 2223:138]
  wire  _T_798 = _T_797 | io_dbg_tlu_halted_f; // @[dec_tlu_ctl.scala 2223:170]
  wire  wr_mtdata1_t_r_0 = _T_795 & _T_798; // @[dec_tlu_ctl.scala 2223:135]
  wire  _T_803 = mtsel == 2'h1; // @[dec_tlu_ctl.scala 2223:121]
  wire  _T_804 = _T_793 & _T_803; // @[dec_tlu_ctl.scala 2223:112]
  wire  _T_806 = ~io_mtdata1_t_1[9]; // @[dec_tlu_ctl.scala 2223:138]
  wire  _T_807 = _T_806 | io_dbg_tlu_halted_f; // @[dec_tlu_ctl.scala 2223:170]
  wire  wr_mtdata1_t_r_1 = _T_804 & _T_807; // @[dec_tlu_ctl.scala 2223:135]
  wire  _T_812 = mtsel == 2'h2; // @[dec_tlu_ctl.scala 2223:121]
  wire  _T_813 = _T_793 & _T_812; // @[dec_tlu_ctl.scala 2223:112]
  wire  _T_815 = ~io_mtdata1_t_2[9]; // @[dec_tlu_ctl.scala 2223:138]
  wire  _T_816 = _T_815 | io_dbg_tlu_halted_f; // @[dec_tlu_ctl.scala 2223:170]
  wire  wr_mtdata1_t_r_2 = _T_813 & _T_816; // @[dec_tlu_ctl.scala 2223:135]
  wire  _T_821 = mtsel == 2'h3; // @[dec_tlu_ctl.scala 2223:121]
  wire  _T_822 = _T_793 & _T_821; // @[dec_tlu_ctl.scala 2223:112]
  wire  _T_824 = ~io_mtdata1_t_3[9]; // @[dec_tlu_ctl.scala 2223:138]
  wire  _T_825 = _T_824 | io_dbg_tlu_halted_f; // @[dec_tlu_ctl.scala 2223:170]
  wire  wr_mtdata1_t_r_3 = _T_822 & _T_825; // @[dec_tlu_ctl.scala 2223:135]
  wire  _T_831 = io_update_hit_bit_r[0] | io_mtdata1_t_0[8]; // @[dec_tlu_ctl.scala 2224:139]
  wire [9:0] _T_834 = {io_mtdata1_t_0[9],_T_831,io_mtdata1_t_0[7:0]}; // @[Cat.scala 29:58]
  wire  _T_840 = io_update_hit_bit_r[1] | io_mtdata1_t_1[8]; // @[dec_tlu_ctl.scala 2224:139]
  wire [9:0] _T_843 = {io_mtdata1_t_1[9],_T_840,io_mtdata1_t_1[7:0]}; // @[Cat.scala 29:58]
  wire  _T_849 = io_update_hit_bit_r[2] | io_mtdata1_t_2[8]; // @[dec_tlu_ctl.scala 2224:139]
  wire [9:0] _T_852 = {io_mtdata1_t_2[9],_T_849,io_mtdata1_t_2[7:0]}; // @[Cat.scala 29:58]
  wire  _T_858 = io_update_hit_bit_r[3] | io_mtdata1_t_3[8]; // @[dec_tlu_ctl.scala 2224:139]
  wire [9:0] _T_861 = {io_mtdata1_t_3[9],_T_858,io_mtdata1_t_3[7:0]}; // @[Cat.scala 29:58]
  reg [9:0] _T_863; // @[dec_tlu_ctl.scala 2226:74]
  reg [9:0] _T_864; // @[dec_tlu_ctl.scala 2226:74]
  reg [9:0] _T_865; // @[dec_tlu_ctl.scala 2226:74]
  reg [9:0] _T_866; // @[dec_tlu_ctl.scala 2226:74]
  wire [31:0] _T_881 = {4'h2,io_mtdata1_t_0[9],6'h1f,io_mtdata1_t_0[8:7],6'h0,io_mtdata1_t_0[6:5],3'h0,io_mtdata1_t_0[4:3],3'h0,io_mtdata1_t_0[2:0]}; // @[Cat.scala 29:58]
  wire [31:0] _T_896 = {4'h2,io_mtdata1_t_1[9],6'h1f,io_mtdata1_t_1[8:7],6'h0,io_mtdata1_t_1[6:5],3'h0,io_mtdata1_t_1[4:3],3'h0,io_mtdata1_t_1[2:0]}; // @[Cat.scala 29:58]
  wire [31:0] _T_911 = {4'h2,io_mtdata1_t_2[9],6'h1f,io_mtdata1_t_2[8:7],6'h0,io_mtdata1_t_2[6:5],3'h0,io_mtdata1_t_2[4:3],3'h0,io_mtdata1_t_2[2:0]}; // @[Cat.scala 29:58]
  wire [31:0] _T_926 = {4'h2,io_mtdata1_t_3[9],6'h1f,io_mtdata1_t_3[8:7],6'h0,io_mtdata1_t_3[6:5],3'h0,io_mtdata1_t_3[4:3],3'h0,io_mtdata1_t_3[2:0]}; // @[Cat.scala 29:58]
  wire [31:0] _T_927 = _T_794 ? _T_881 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_928 = _T_803 ? _T_896 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_929 = _T_812 ? _T_911 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_930 = _T_821 ? _T_926 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_931 = _T_927 | _T_928; // @[Mux.scala 27:72]
  wire [31:0] _T_932 = _T_931 | _T_929; // @[Mux.scala 27:72]
  wire [31:0] mtdata1_tsel_out = _T_932 | _T_930; // @[Mux.scala 27:72]
  wire  _T_959 = io_dec_csr_wraddr_r == 12'h7a2; // @[dec_tlu_ctl.scala 2243:98]
  wire  _T_960 = io_dec_csr_wen_r_mod & _T_959; // @[dec_tlu_ctl.scala 2243:69]
  wire  _T_962 = _T_960 & _T_794; // @[dec_tlu_ctl.scala 2243:111]
  wire  _T_971 = _T_960 & _T_803; // @[dec_tlu_ctl.scala 2243:111]
  wire  _T_980 = _T_960 & _T_812; // @[dec_tlu_ctl.scala 2243:111]
  wire  _T_989 = _T_960 & _T_821; // @[dec_tlu_ctl.scala 2243:111]
  reg [31:0] mtdata2_t_0; // @[lib.scala 374:16]
  reg [31:0] mtdata2_t_1; // @[lib.scala 374:16]
  reg [31:0] mtdata2_t_2; // @[lib.scala 374:16]
  reg [31:0] mtdata2_t_3; // @[lib.scala 374:16]
  wire [31:0] _T_1006 = _T_794 ? mtdata2_t_0 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1007 = _T_803 ? mtdata2_t_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1008 = _T_812 ? mtdata2_t_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1009 = _T_821 ? mtdata2_t_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1010 = _T_1006 | _T_1007; // @[Mux.scala 27:72]
  wire [31:0] _T_1011 = _T_1010 | _T_1008; // @[Mux.scala 27:72]
  wire [31:0] mtdata2_tsel_out = _T_1011 | _T_1009; // @[Mux.scala 27:72]
  wire [3:0] _T_1014 = io_tlu_i0_commit_cmt ? 4'hf : 4'h0; // @[Bitwise.scala 72:12]
  wire [3:0] pmu_i0_itype_qual = io_dec_tlu_packet_r_pmu_i0_itype & _T_1014; // @[dec_tlu_ctl.scala 2268:59]
  wire  _T_1016 = ~mcountinhibit[3]; // @[dec_tlu_ctl.scala 2274:24]
  reg [9:0] mhpme3; // @[Reg.scala 27:20]
  wire  _T_1017 = mhpme3 == 10'h1; // @[dec_tlu_ctl.scala 2275:34]
  wire  _T_1019 = mhpme3 == 10'h2; // @[dec_tlu_ctl.scala 2276:34]
  wire  _T_1021 = mhpme3 == 10'h3; // @[dec_tlu_ctl.scala 2277:34]
  wire  _T_1023 = mhpme3 == 10'h4; // @[dec_tlu_ctl.scala 2278:34]
  wire  _T_1025 = ~io_illegal_r; // @[dec_tlu_ctl.scala 2278:96]
  wire  _T_1026 = io_tlu_i0_commit_cmt & _T_1025; // @[dec_tlu_ctl.scala 2278:94]
  wire  _T_1027 = mhpme3 == 10'h5; // @[dec_tlu_ctl.scala 2279:34]
  wire  _T_1029 = ~io_exu_pmu_i0_pc4; // @[dec_tlu_ctl.scala 2279:96]
  wire  _T_1030 = io_tlu_i0_commit_cmt & _T_1029; // @[dec_tlu_ctl.scala 2279:94]
  wire  _T_1032 = _T_1030 & _T_1025; // @[dec_tlu_ctl.scala 2279:115]
  wire  _T_1033 = mhpme3 == 10'h6; // @[dec_tlu_ctl.scala 2280:34]
  wire  _T_1035 = io_tlu_i0_commit_cmt & io_exu_pmu_i0_pc4; // @[dec_tlu_ctl.scala 2280:94]
  wire  _T_1037 = _T_1035 & _T_1025; // @[dec_tlu_ctl.scala 2280:115]
  wire  _T_1038 = mhpme3 == 10'h7; // @[dec_tlu_ctl.scala 2281:34]
  wire  _T_1040 = mhpme3 == 10'h8; // @[dec_tlu_ctl.scala 2282:34]
  wire  _T_1042 = mhpme3 == 10'h1e; // @[dec_tlu_ctl.scala 2283:34]
  wire  _T_1044 = mhpme3 == 10'h9; // @[dec_tlu_ctl.scala 2284:34]
  wire  _T_1046 = pmu_i0_itype_qual == 4'h1; // @[dec_tlu_ctl.scala 2284:91]
  wire  _T_1047 = mhpme3 == 10'ha; // @[dec_tlu_ctl.scala 2285:34]
  wire  _T_1049 = io_dec_tlu_packet_r_pmu_divide & io_tlu_i0_commit_cmt; // @[dec_tlu_ctl.scala 2285:105]
  wire  _T_1050 = mhpme3 == 10'hb; // @[dec_tlu_ctl.scala 2286:34]
  wire  _T_1052 = pmu_i0_itype_qual == 4'h2; // @[dec_tlu_ctl.scala 2286:91]
  wire  _T_1053 = mhpme3 == 10'hc; // @[dec_tlu_ctl.scala 2287:34]
  wire  _T_1055 = pmu_i0_itype_qual == 4'h3; // @[dec_tlu_ctl.scala 2287:91]
  wire  _T_1056 = mhpme3 == 10'hd; // @[dec_tlu_ctl.scala 2288:34]
  wire  _T_1059 = _T_1052 & io_dec_tlu_packet_r_pmu_lsu_misaligned; // @[dec_tlu_ctl.scala 2288:100]
  wire  _T_1060 = mhpme3 == 10'he; // @[dec_tlu_ctl.scala 2289:34]
  wire  _T_1064 = _T_1055 & io_dec_tlu_packet_r_pmu_lsu_misaligned; // @[dec_tlu_ctl.scala 2289:101]
  wire  _T_1065 = mhpme3 == 10'hf; // @[dec_tlu_ctl.scala 2290:34]
  wire  _T_1067 = pmu_i0_itype_qual == 4'h4; // @[dec_tlu_ctl.scala 2290:89]
  wire  _T_1068 = mhpme3 == 10'h10; // @[dec_tlu_ctl.scala 2291:34]
  wire  _T_1070 = pmu_i0_itype_qual == 4'h5; // @[dec_tlu_ctl.scala 2291:89]
  wire  _T_1071 = mhpme3 == 10'h12; // @[dec_tlu_ctl.scala 2292:34]
  wire  _T_1073 = pmu_i0_itype_qual == 4'h6; // @[dec_tlu_ctl.scala 2292:89]
  wire  _T_1074 = mhpme3 == 10'h11; // @[dec_tlu_ctl.scala 2293:34]
  wire  _T_1076 = pmu_i0_itype_qual == 4'h7; // @[dec_tlu_ctl.scala 2293:89]
  wire  _T_1077 = mhpme3 == 10'h13; // @[dec_tlu_ctl.scala 2294:34]
  wire  _T_1079 = pmu_i0_itype_qual == 4'h8; // @[dec_tlu_ctl.scala 2294:89]
  wire  _T_1080 = mhpme3 == 10'h14; // @[dec_tlu_ctl.scala 2295:34]
  wire  _T_1082 = pmu_i0_itype_qual == 4'h9; // @[dec_tlu_ctl.scala 2295:89]
  wire  _T_1083 = mhpme3 == 10'h15; // @[dec_tlu_ctl.scala 2296:34]
  wire  _T_1085 = pmu_i0_itype_qual == 4'ha; // @[dec_tlu_ctl.scala 2296:89]
  wire  _T_1086 = mhpme3 == 10'h16; // @[dec_tlu_ctl.scala 2297:34]
  wire  _T_1088 = pmu_i0_itype_qual == 4'hb; // @[dec_tlu_ctl.scala 2297:89]
  wire  _T_1089 = mhpme3 == 10'h17; // @[dec_tlu_ctl.scala 2298:34]
  wire  _T_1091 = pmu_i0_itype_qual == 4'hc; // @[dec_tlu_ctl.scala 2298:89]
  wire  _T_1092 = mhpme3 == 10'h18; // @[dec_tlu_ctl.scala 2299:34]
  wire  _T_1094 = pmu_i0_itype_qual == 4'hd; // @[dec_tlu_ctl.scala 2299:89]
  wire  _T_1095 = pmu_i0_itype_qual == 4'he; // @[dec_tlu_ctl.scala 2299:122]
  wire  _T_1096 = _T_1094 | _T_1095; // @[dec_tlu_ctl.scala 2299:101]
  wire  _T_1097 = mhpme3 == 10'h19; // @[dec_tlu_ctl.scala 2300:34]
  wire  _T_1099 = io_exu_pmu_i0_br_misp & io_tlu_i0_commit_cmt; // @[dec_tlu_ctl.scala 2300:95]
  wire  _T_1100 = mhpme3 == 10'h1a; // @[dec_tlu_ctl.scala 2301:34]
  wire  _T_1102 = io_exu_pmu_i0_br_ataken & io_tlu_i0_commit_cmt; // @[dec_tlu_ctl.scala 2301:97]
  wire  _T_1103 = mhpme3 == 10'h1b; // @[dec_tlu_ctl.scala 2302:34]
  wire  _T_1105 = io_dec_tlu_packet_r_pmu_i0_br_unpred & io_tlu_i0_commit_cmt; // @[dec_tlu_ctl.scala 2302:110]
  wire  _T_1106 = mhpme3 == 10'h1c; // @[dec_tlu_ctl.scala 2303:34]
  wire  _T_1110 = mhpme3 == 10'h1f; // @[dec_tlu_ctl.scala 2305:34]
  wire  _T_1112 = mhpme3 == 10'h20; // @[dec_tlu_ctl.scala 2306:34]
  wire  _T_1114 = mhpme3 == 10'h22; // @[dec_tlu_ctl.scala 2307:34]
  wire  _T_1116 = mhpme3 == 10'h23; // @[dec_tlu_ctl.scala 2308:34]
  wire  _T_1118 = mhpme3 == 10'h24; // @[dec_tlu_ctl.scala 2309:34]
  wire  _T_1120 = mhpme3 == 10'h25; // @[dec_tlu_ctl.scala 2310:34]
  wire  _T_1122 = io_i0_exception_valid_r | io_i0_trigger_hit_r; // @[dec_tlu_ctl.scala 2310:98]
  wire  _T_1123 = _T_1122 | io_lsu_exc_valid_r; // @[dec_tlu_ctl.scala 2310:120]
  wire  _T_1124 = mhpme3 == 10'h26; // @[dec_tlu_ctl.scala 2311:34]
  wire  _T_1126 = io_take_timer_int | io_take_int_timer0_int; // @[dec_tlu_ctl.scala 2311:92]
  wire  _T_1127 = _T_1126 | io_take_int_timer1_int; // @[dec_tlu_ctl.scala 2311:117]
  wire  _T_1128 = mhpme3 == 10'h27; // @[dec_tlu_ctl.scala 2312:34]
  wire  _T_1130 = mhpme3 == 10'h28; // @[dec_tlu_ctl.scala 2313:34]
  wire  _T_1132 = mhpme3 == 10'h29; // @[dec_tlu_ctl.scala 2314:34]
  wire  _T_1134 = io_dec_tlu_br0_error_r | io_dec_tlu_br0_start_error_r; // @[dec_tlu_ctl.scala 2314:97]
  wire  _T_1135 = _T_1134 & io_rfpc_i0_r; // @[dec_tlu_ctl.scala 2314:129]
  wire  _T_1140 = mhpme3 == 10'h2c; // @[dec_tlu_ctl.scala 2317:34]
  wire  _T_1142 = mhpme3 == 10'h2d; // @[dec_tlu_ctl.scala 2318:34]
  wire  _T_1144 = mhpme3 == 10'h2e; // @[dec_tlu_ctl.scala 2319:34]
  wire  _T_1146 = mhpme3 == 10'h2f; // @[dec_tlu_ctl.scala 2320:34]
  wire  _T_1148 = mhpme3 == 10'h30; // @[dec_tlu_ctl.scala 2321:34]
  wire  _T_1150 = mhpme3 == 10'h31; // @[dec_tlu_ctl.scala 2322:34]
  wire  _T_1154 = ~io_mstatus[0]; // @[dec_tlu_ctl.scala 2322:73]
  wire  _T_1155 = mhpme3 == 10'h32; // @[dec_tlu_ctl.scala 2323:34]
  wire [5:0] _T_1162 = io_mip & mie; // @[dec_tlu_ctl.scala 2323:113]
  wire  _T_1163 = |_T_1162; // @[dec_tlu_ctl.scala 2323:125]
  wire  _T_1164 = _T_1154 & _T_1163; // @[dec_tlu_ctl.scala 2323:98]
  wire  _T_1165 = mhpme3 == 10'h36; // @[dec_tlu_ctl.scala 2324:34]
  wire  _T_1167 = pmu_i0_itype_qual == 4'hf; // @[dec_tlu_ctl.scala 2324:91]
  wire  _T_1168 = mhpme3 == 10'h37; // @[dec_tlu_ctl.scala 2325:34]
  wire  _T_1170 = io_tlu_i0_commit_cmt & io_lsu_pmu_load_external_r; // @[dec_tlu_ctl.scala 2325:94]
  wire  _T_1171 = mhpme3 == 10'h38; // @[dec_tlu_ctl.scala 2326:34]
  wire  _T_1173 = io_tlu_i0_commit_cmt & io_lsu_pmu_store_external_r; // @[dec_tlu_ctl.scala 2326:94]
  wire  _T_1174 = mhpme3 == 10'h200; // @[dec_tlu_ctl.scala 2328:34]
  wire  _T_1176 = mhpme3 == 10'h201; // @[dec_tlu_ctl.scala 2329:34]
  wire  _T_1178 = mhpme3 == 10'h202; // @[dec_tlu_ctl.scala 2330:34]
  wire  _T_1180 = mhpme3 == 10'h203; // @[dec_tlu_ctl.scala 2331:34]
  wire  _T_1182 = mhpme3 == 10'h204; // @[dec_tlu_ctl.scala 2332:34]
  wire  _T_1185 = _T_1019 & io_ifu_pmu_ic_hit; // @[Mux.scala 27:72]
  wire  _T_1186 = _T_1021 & io_ifu_pmu_ic_miss; // @[Mux.scala 27:72]
  wire  _T_1187 = _T_1023 & _T_1026; // @[Mux.scala 27:72]
  wire  _T_1188 = _T_1027 & _T_1032; // @[Mux.scala 27:72]
  wire  _T_1189 = _T_1033 & _T_1037; // @[Mux.scala 27:72]
  wire  _T_1190 = _T_1038 & io_ifu_pmu_instr_aligned; // @[Mux.scala 27:72]
  wire  _T_1191 = _T_1040 & io_dec_pmu_instr_decoded; // @[Mux.scala 27:72]
  wire  _T_1192 = _T_1042 & io_dec_pmu_decode_stall; // @[Mux.scala 27:72]
  wire  _T_1193 = _T_1044 & _T_1046; // @[Mux.scala 27:72]
  wire  _T_1194 = _T_1047 & _T_1049; // @[Mux.scala 27:72]
  wire  _T_1195 = _T_1050 & _T_1052; // @[Mux.scala 27:72]
  wire  _T_1196 = _T_1053 & _T_1055; // @[Mux.scala 27:72]
  wire  _T_1197 = _T_1056 & _T_1059; // @[Mux.scala 27:72]
  wire  _T_1198 = _T_1060 & _T_1064; // @[Mux.scala 27:72]
  wire  _T_1199 = _T_1065 & _T_1067; // @[Mux.scala 27:72]
  wire  _T_1200 = _T_1068 & _T_1070; // @[Mux.scala 27:72]
  wire  _T_1201 = _T_1071 & _T_1073; // @[Mux.scala 27:72]
  wire  _T_1202 = _T_1074 & _T_1076; // @[Mux.scala 27:72]
  wire  _T_1203 = _T_1077 & _T_1079; // @[Mux.scala 27:72]
  wire  _T_1204 = _T_1080 & _T_1082; // @[Mux.scala 27:72]
  wire  _T_1205 = _T_1083 & _T_1085; // @[Mux.scala 27:72]
  wire  _T_1206 = _T_1086 & _T_1088; // @[Mux.scala 27:72]
  wire  _T_1207 = _T_1089 & _T_1091; // @[Mux.scala 27:72]
  wire  _T_1208 = _T_1092 & _T_1096; // @[Mux.scala 27:72]
  wire  _T_1209 = _T_1097 & _T_1099; // @[Mux.scala 27:72]
  wire  _T_1210 = _T_1100 & _T_1102; // @[Mux.scala 27:72]
  wire  _T_1211 = _T_1103 & _T_1105; // @[Mux.scala 27:72]
  wire  _T_1212 = _T_1106 & io_ifu_pmu_fetch_stall; // @[Mux.scala 27:72]
  wire  _T_1214 = _T_1110 & io_dec_pmu_postsync_stall; // @[Mux.scala 27:72]
  wire  _T_1215 = _T_1112 & io_dec_pmu_presync_stall; // @[Mux.scala 27:72]
  wire  _T_1216 = _T_1114 & io_lsu_store_stall_any; // @[Mux.scala 27:72]
  wire  _T_1217 = _T_1116 & io_dma_dccm_stall_any; // @[Mux.scala 27:72]
  wire  _T_1218 = _T_1118 & io_dma_iccm_stall_any; // @[Mux.scala 27:72]
  wire  _T_1219 = _T_1120 & _T_1123; // @[Mux.scala 27:72]
  wire  _T_1220 = _T_1124 & _T_1127; // @[Mux.scala 27:72]
  wire  _T_1221 = _T_1128 & io_take_ext_int; // @[Mux.scala 27:72]
  wire  _T_1222 = _T_1130 & io_tlu_flush_lower_r; // @[Mux.scala 27:72]
  wire  _T_1223 = _T_1132 & _T_1135; // @[Mux.scala 27:72]
  wire  _T_1226 = _T_1140 & io_lsu_pmu_bus_misaligned; // @[Mux.scala 27:72]
  wire  _T_1227 = _T_1142 & io_ifu_pmu_bus_error; // @[Mux.scala 27:72]
  wire  _T_1228 = _T_1144 & io_lsu_pmu_bus_error; // @[Mux.scala 27:72]
  wire  _T_1229 = _T_1146 & io_ifu_pmu_bus_busy; // @[Mux.scala 27:72]
  wire  _T_1230 = _T_1148 & io_lsu_pmu_bus_busy; // @[Mux.scala 27:72]
  wire  _T_1231 = _T_1150 & _T_1154; // @[Mux.scala 27:72]
  wire  _T_1232 = _T_1155 & _T_1164; // @[Mux.scala 27:72]
  wire  _T_1233 = _T_1165 & _T_1167; // @[Mux.scala 27:72]
  wire  _T_1234 = _T_1168 & _T_1170; // @[Mux.scala 27:72]
  wire  _T_1235 = _T_1171 & _T_1173; // @[Mux.scala 27:72]
  wire  _T_1236 = _T_1174 & io_dec_tlu_pmu_fw_halted; // @[Mux.scala 27:72]
  wire  _T_1237 = _T_1176 & io_dma_pmu_any_read; // @[Mux.scala 27:72]
  wire  _T_1238 = _T_1178 & io_dma_pmu_any_write; // @[Mux.scala 27:72]
  wire  _T_1239 = _T_1180 & io_dma_pmu_dccm_read; // @[Mux.scala 27:72]
  wire  _T_1240 = _T_1182 & io_dma_pmu_dccm_write; // @[Mux.scala 27:72]
  wire  _T_1241 = _T_1017 | _T_1185; // @[Mux.scala 27:72]
  wire  _T_1242 = _T_1241 | _T_1186; // @[Mux.scala 27:72]
  wire  _T_1243 = _T_1242 | _T_1187; // @[Mux.scala 27:72]
  wire  _T_1244 = _T_1243 | _T_1188; // @[Mux.scala 27:72]
  wire  _T_1245 = _T_1244 | _T_1189; // @[Mux.scala 27:72]
  wire  _T_1246 = _T_1245 | _T_1190; // @[Mux.scala 27:72]
  wire  _T_1247 = _T_1246 | _T_1191; // @[Mux.scala 27:72]
  wire  _T_1248 = _T_1247 | _T_1192; // @[Mux.scala 27:72]
  wire  _T_1249 = _T_1248 | _T_1193; // @[Mux.scala 27:72]
  wire  _T_1250 = _T_1249 | _T_1194; // @[Mux.scala 27:72]
  wire  _T_1251 = _T_1250 | _T_1195; // @[Mux.scala 27:72]
  wire  _T_1252 = _T_1251 | _T_1196; // @[Mux.scala 27:72]
  wire  _T_1253 = _T_1252 | _T_1197; // @[Mux.scala 27:72]
  wire  _T_1254 = _T_1253 | _T_1198; // @[Mux.scala 27:72]
  wire  _T_1255 = _T_1254 | _T_1199; // @[Mux.scala 27:72]
  wire  _T_1256 = _T_1255 | _T_1200; // @[Mux.scala 27:72]
  wire  _T_1257 = _T_1256 | _T_1201; // @[Mux.scala 27:72]
  wire  _T_1258 = _T_1257 | _T_1202; // @[Mux.scala 27:72]
  wire  _T_1259 = _T_1258 | _T_1203; // @[Mux.scala 27:72]
  wire  _T_1260 = _T_1259 | _T_1204; // @[Mux.scala 27:72]
  wire  _T_1261 = _T_1260 | _T_1205; // @[Mux.scala 27:72]
  wire  _T_1262 = _T_1261 | _T_1206; // @[Mux.scala 27:72]
  wire  _T_1263 = _T_1262 | _T_1207; // @[Mux.scala 27:72]
  wire  _T_1264 = _T_1263 | _T_1208; // @[Mux.scala 27:72]
  wire  _T_1265 = _T_1264 | _T_1209; // @[Mux.scala 27:72]
  wire  _T_1266 = _T_1265 | _T_1210; // @[Mux.scala 27:72]
  wire  _T_1267 = _T_1266 | _T_1211; // @[Mux.scala 27:72]
  wire  _T_1268 = _T_1267 | _T_1212; // @[Mux.scala 27:72]
  wire  _T_1269 = _T_1268 | _T_1192; // @[Mux.scala 27:72]
  wire  _T_1270 = _T_1269 | _T_1214; // @[Mux.scala 27:72]
  wire  _T_1271 = _T_1270 | _T_1215; // @[Mux.scala 27:72]
  wire  _T_1272 = _T_1271 | _T_1216; // @[Mux.scala 27:72]
  wire  _T_1273 = _T_1272 | _T_1217; // @[Mux.scala 27:72]
  wire  _T_1274 = _T_1273 | _T_1218; // @[Mux.scala 27:72]
  wire  _T_1275 = _T_1274 | _T_1219; // @[Mux.scala 27:72]
  wire  _T_1276 = _T_1275 | _T_1220; // @[Mux.scala 27:72]
  wire  _T_1277 = _T_1276 | _T_1221; // @[Mux.scala 27:72]
  wire  _T_1278 = _T_1277 | _T_1222; // @[Mux.scala 27:72]
  wire  _T_1279 = _T_1278 | _T_1223; // @[Mux.scala 27:72]
  wire  _T_1282 = _T_1279 | _T_1226; // @[Mux.scala 27:72]
  wire  _T_1283 = _T_1282 | _T_1227; // @[Mux.scala 27:72]
  wire  _T_1284 = _T_1283 | _T_1228; // @[Mux.scala 27:72]
  wire  _T_1285 = _T_1284 | _T_1229; // @[Mux.scala 27:72]
  wire  _T_1286 = _T_1285 | _T_1230; // @[Mux.scala 27:72]
  wire  _T_1287 = _T_1286 | _T_1231; // @[Mux.scala 27:72]
  wire  _T_1288 = _T_1287 | _T_1232; // @[Mux.scala 27:72]
  wire  _T_1289 = _T_1288 | _T_1233; // @[Mux.scala 27:72]
  wire  _T_1290 = _T_1289 | _T_1234; // @[Mux.scala 27:72]
  wire  _T_1291 = _T_1290 | _T_1235; // @[Mux.scala 27:72]
  wire  _T_1292 = _T_1291 | _T_1236; // @[Mux.scala 27:72]
  wire  _T_1293 = _T_1292 | _T_1237; // @[Mux.scala 27:72]
  wire  _T_1294 = _T_1293 | _T_1238; // @[Mux.scala 27:72]
  wire  _T_1295 = _T_1294 | _T_1239; // @[Mux.scala 27:72]
  wire  _T_1296 = _T_1295 | _T_1240; // @[Mux.scala 27:72]
  wire  mhpmc_inc_r_0 = _T_1016 & _T_1296; // @[dec_tlu_ctl.scala 2274:44]
  wire  _T_1300 = ~mcountinhibit[4]; // @[dec_tlu_ctl.scala 2274:24]
  reg [9:0] mhpme4; // @[Reg.scala 27:20]
  wire  _T_1301 = mhpme4 == 10'h1; // @[dec_tlu_ctl.scala 2275:34]
  wire  _T_1303 = mhpme4 == 10'h2; // @[dec_tlu_ctl.scala 2276:34]
  wire  _T_1305 = mhpme4 == 10'h3; // @[dec_tlu_ctl.scala 2277:34]
  wire  _T_1307 = mhpme4 == 10'h4; // @[dec_tlu_ctl.scala 2278:34]
  wire  _T_1311 = mhpme4 == 10'h5; // @[dec_tlu_ctl.scala 2279:34]
  wire  _T_1317 = mhpme4 == 10'h6; // @[dec_tlu_ctl.scala 2280:34]
  wire  _T_1322 = mhpme4 == 10'h7; // @[dec_tlu_ctl.scala 2281:34]
  wire  _T_1324 = mhpme4 == 10'h8; // @[dec_tlu_ctl.scala 2282:34]
  wire  _T_1326 = mhpme4 == 10'h1e; // @[dec_tlu_ctl.scala 2283:34]
  wire  _T_1328 = mhpme4 == 10'h9; // @[dec_tlu_ctl.scala 2284:34]
  wire  _T_1331 = mhpme4 == 10'ha; // @[dec_tlu_ctl.scala 2285:34]
  wire  _T_1334 = mhpme4 == 10'hb; // @[dec_tlu_ctl.scala 2286:34]
  wire  _T_1337 = mhpme4 == 10'hc; // @[dec_tlu_ctl.scala 2287:34]
  wire  _T_1340 = mhpme4 == 10'hd; // @[dec_tlu_ctl.scala 2288:34]
  wire  _T_1344 = mhpme4 == 10'he; // @[dec_tlu_ctl.scala 2289:34]
  wire  _T_1349 = mhpme4 == 10'hf; // @[dec_tlu_ctl.scala 2290:34]
  wire  _T_1352 = mhpme4 == 10'h10; // @[dec_tlu_ctl.scala 2291:34]
  wire  _T_1355 = mhpme4 == 10'h12; // @[dec_tlu_ctl.scala 2292:34]
  wire  _T_1358 = mhpme4 == 10'h11; // @[dec_tlu_ctl.scala 2293:34]
  wire  _T_1361 = mhpme4 == 10'h13; // @[dec_tlu_ctl.scala 2294:34]
  wire  _T_1364 = mhpme4 == 10'h14; // @[dec_tlu_ctl.scala 2295:34]
  wire  _T_1367 = mhpme4 == 10'h15; // @[dec_tlu_ctl.scala 2296:34]
  wire  _T_1370 = mhpme4 == 10'h16; // @[dec_tlu_ctl.scala 2297:34]
  wire  _T_1373 = mhpme4 == 10'h17; // @[dec_tlu_ctl.scala 2298:34]
  wire  _T_1376 = mhpme4 == 10'h18; // @[dec_tlu_ctl.scala 2299:34]
  wire  _T_1381 = mhpme4 == 10'h19; // @[dec_tlu_ctl.scala 2300:34]
  wire  _T_1384 = mhpme4 == 10'h1a; // @[dec_tlu_ctl.scala 2301:34]
  wire  _T_1387 = mhpme4 == 10'h1b; // @[dec_tlu_ctl.scala 2302:34]
  wire  _T_1390 = mhpme4 == 10'h1c; // @[dec_tlu_ctl.scala 2303:34]
  wire  _T_1394 = mhpme4 == 10'h1f; // @[dec_tlu_ctl.scala 2305:34]
  wire  _T_1396 = mhpme4 == 10'h20; // @[dec_tlu_ctl.scala 2306:34]
  wire  _T_1398 = mhpme4 == 10'h22; // @[dec_tlu_ctl.scala 2307:34]
  wire  _T_1400 = mhpme4 == 10'h23; // @[dec_tlu_ctl.scala 2308:34]
  wire  _T_1402 = mhpme4 == 10'h24; // @[dec_tlu_ctl.scala 2309:34]
  wire  _T_1404 = mhpme4 == 10'h25; // @[dec_tlu_ctl.scala 2310:34]
  wire  _T_1408 = mhpme4 == 10'h26; // @[dec_tlu_ctl.scala 2311:34]
  wire  _T_1412 = mhpme4 == 10'h27; // @[dec_tlu_ctl.scala 2312:34]
  wire  _T_1414 = mhpme4 == 10'h28; // @[dec_tlu_ctl.scala 2313:34]
  wire  _T_1416 = mhpme4 == 10'h29; // @[dec_tlu_ctl.scala 2314:34]
  wire  _T_1424 = mhpme4 == 10'h2c; // @[dec_tlu_ctl.scala 2317:34]
  wire  _T_1426 = mhpme4 == 10'h2d; // @[dec_tlu_ctl.scala 2318:34]
  wire  _T_1428 = mhpme4 == 10'h2e; // @[dec_tlu_ctl.scala 2319:34]
  wire  _T_1430 = mhpme4 == 10'h2f; // @[dec_tlu_ctl.scala 2320:34]
  wire  _T_1432 = mhpme4 == 10'h30; // @[dec_tlu_ctl.scala 2321:34]
  wire  _T_1434 = mhpme4 == 10'h31; // @[dec_tlu_ctl.scala 2322:34]
  wire  _T_1439 = mhpme4 == 10'h32; // @[dec_tlu_ctl.scala 2323:34]
  wire  _T_1449 = mhpme4 == 10'h36; // @[dec_tlu_ctl.scala 2324:34]
  wire  _T_1452 = mhpme4 == 10'h37; // @[dec_tlu_ctl.scala 2325:34]
  wire  _T_1455 = mhpme4 == 10'h38; // @[dec_tlu_ctl.scala 2326:34]
  wire  _T_1458 = mhpme4 == 10'h200; // @[dec_tlu_ctl.scala 2328:34]
  wire  _T_1460 = mhpme4 == 10'h201; // @[dec_tlu_ctl.scala 2329:34]
  wire  _T_1462 = mhpme4 == 10'h202; // @[dec_tlu_ctl.scala 2330:34]
  wire  _T_1464 = mhpme4 == 10'h203; // @[dec_tlu_ctl.scala 2331:34]
  wire  _T_1466 = mhpme4 == 10'h204; // @[dec_tlu_ctl.scala 2332:34]
  wire  _T_1469 = _T_1303 & io_ifu_pmu_ic_hit; // @[Mux.scala 27:72]
  wire  _T_1470 = _T_1305 & io_ifu_pmu_ic_miss; // @[Mux.scala 27:72]
  wire  _T_1471 = _T_1307 & _T_1026; // @[Mux.scala 27:72]
  wire  _T_1472 = _T_1311 & _T_1032; // @[Mux.scala 27:72]
  wire  _T_1473 = _T_1317 & _T_1037; // @[Mux.scala 27:72]
  wire  _T_1474 = _T_1322 & io_ifu_pmu_instr_aligned; // @[Mux.scala 27:72]
  wire  _T_1475 = _T_1324 & io_dec_pmu_instr_decoded; // @[Mux.scala 27:72]
  wire  _T_1476 = _T_1326 & io_dec_pmu_decode_stall; // @[Mux.scala 27:72]
  wire  _T_1477 = _T_1328 & _T_1046; // @[Mux.scala 27:72]
  wire  _T_1478 = _T_1331 & _T_1049; // @[Mux.scala 27:72]
  wire  _T_1479 = _T_1334 & _T_1052; // @[Mux.scala 27:72]
  wire  _T_1480 = _T_1337 & _T_1055; // @[Mux.scala 27:72]
  wire  _T_1481 = _T_1340 & _T_1059; // @[Mux.scala 27:72]
  wire  _T_1482 = _T_1344 & _T_1064; // @[Mux.scala 27:72]
  wire  _T_1483 = _T_1349 & _T_1067; // @[Mux.scala 27:72]
  wire  _T_1484 = _T_1352 & _T_1070; // @[Mux.scala 27:72]
  wire  _T_1485 = _T_1355 & _T_1073; // @[Mux.scala 27:72]
  wire  _T_1486 = _T_1358 & _T_1076; // @[Mux.scala 27:72]
  wire  _T_1487 = _T_1361 & _T_1079; // @[Mux.scala 27:72]
  wire  _T_1488 = _T_1364 & _T_1082; // @[Mux.scala 27:72]
  wire  _T_1489 = _T_1367 & _T_1085; // @[Mux.scala 27:72]
  wire  _T_1490 = _T_1370 & _T_1088; // @[Mux.scala 27:72]
  wire  _T_1491 = _T_1373 & _T_1091; // @[Mux.scala 27:72]
  wire  _T_1492 = _T_1376 & _T_1096; // @[Mux.scala 27:72]
  wire  _T_1493 = _T_1381 & _T_1099; // @[Mux.scala 27:72]
  wire  _T_1494 = _T_1384 & _T_1102; // @[Mux.scala 27:72]
  wire  _T_1495 = _T_1387 & _T_1105; // @[Mux.scala 27:72]
  wire  _T_1496 = _T_1390 & io_ifu_pmu_fetch_stall; // @[Mux.scala 27:72]
  wire  _T_1498 = _T_1394 & io_dec_pmu_postsync_stall; // @[Mux.scala 27:72]
  wire  _T_1499 = _T_1396 & io_dec_pmu_presync_stall; // @[Mux.scala 27:72]
  wire  _T_1500 = _T_1398 & io_lsu_store_stall_any; // @[Mux.scala 27:72]
  wire  _T_1501 = _T_1400 & io_dma_dccm_stall_any; // @[Mux.scala 27:72]
  wire  _T_1502 = _T_1402 & io_dma_iccm_stall_any; // @[Mux.scala 27:72]
  wire  _T_1503 = _T_1404 & _T_1123; // @[Mux.scala 27:72]
  wire  _T_1504 = _T_1408 & _T_1127; // @[Mux.scala 27:72]
  wire  _T_1505 = _T_1412 & io_take_ext_int; // @[Mux.scala 27:72]
  wire  _T_1506 = _T_1414 & io_tlu_flush_lower_r; // @[Mux.scala 27:72]
  wire  _T_1507 = _T_1416 & _T_1135; // @[Mux.scala 27:72]
  wire  _T_1510 = _T_1424 & io_lsu_pmu_bus_misaligned; // @[Mux.scala 27:72]
  wire  _T_1511 = _T_1426 & io_ifu_pmu_bus_error; // @[Mux.scala 27:72]
  wire  _T_1512 = _T_1428 & io_lsu_pmu_bus_error; // @[Mux.scala 27:72]
  wire  _T_1513 = _T_1430 & io_ifu_pmu_bus_busy; // @[Mux.scala 27:72]
  wire  _T_1514 = _T_1432 & io_lsu_pmu_bus_busy; // @[Mux.scala 27:72]
  wire  _T_1515 = _T_1434 & _T_1154; // @[Mux.scala 27:72]
  wire  _T_1516 = _T_1439 & _T_1164; // @[Mux.scala 27:72]
  wire  _T_1517 = _T_1449 & _T_1167; // @[Mux.scala 27:72]
  wire  _T_1518 = _T_1452 & _T_1170; // @[Mux.scala 27:72]
  wire  _T_1519 = _T_1455 & _T_1173; // @[Mux.scala 27:72]
  wire  _T_1520 = _T_1458 & io_dec_tlu_pmu_fw_halted; // @[Mux.scala 27:72]
  wire  _T_1521 = _T_1460 & io_dma_pmu_any_read; // @[Mux.scala 27:72]
  wire  _T_1522 = _T_1462 & io_dma_pmu_any_write; // @[Mux.scala 27:72]
  wire  _T_1523 = _T_1464 & io_dma_pmu_dccm_read; // @[Mux.scala 27:72]
  wire  _T_1524 = _T_1466 & io_dma_pmu_dccm_write; // @[Mux.scala 27:72]
  wire  _T_1525 = _T_1301 | _T_1469; // @[Mux.scala 27:72]
  wire  _T_1526 = _T_1525 | _T_1470; // @[Mux.scala 27:72]
  wire  _T_1527 = _T_1526 | _T_1471; // @[Mux.scala 27:72]
  wire  _T_1528 = _T_1527 | _T_1472; // @[Mux.scala 27:72]
  wire  _T_1529 = _T_1528 | _T_1473; // @[Mux.scala 27:72]
  wire  _T_1530 = _T_1529 | _T_1474; // @[Mux.scala 27:72]
  wire  _T_1531 = _T_1530 | _T_1475; // @[Mux.scala 27:72]
  wire  _T_1532 = _T_1531 | _T_1476; // @[Mux.scala 27:72]
  wire  _T_1533 = _T_1532 | _T_1477; // @[Mux.scala 27:72]
  wire  _T_1534 = _T_1533 | _T_1478; // @[Mux.scala 27:72]
  wire  _T_1535 = _T_1534 | _T_1479; // @[Mux.scala 27:72]
  wire  _T_1536 = _T_1535 | _T_1480; // @[Mux.scala 27:72]
  wire  _T_1537 = _T_1536 | _T_1481; // @[Mux.scala 27:72]
  wire  _T_1538 = _T_1537 | _T_1482; // @[Mux.scala 27:72]
  wire  _T_1539 = _T_1538 | _T_1483; // @[Mux.scala 27:72]
  wire  _T_1540 = _T_1539 | _T_1484; // @[Mux.scala 27:72]
  wire  _T_1541 = _T_1540 | _T_1485; // @[Mux.scala 27:72]
  wire  _T_1542 = _T_1541 | _T_1486; // @[Mux.scala 27:72]
  wire  _T_1543 = _T_1542 | _T_1487; // @[Mux.scala 27:72]
  wire  _T_1544 = _T_1543 | _T_1488; // @[Mux.scala 27:72]
  wire  _T_1545 = _T_1544 | _T_1489; // @[Mux.scala 27:72]
  wire  _T_1546 = _T_1545 | _T_1490; // @[Mux.scala 27:72]
  wire  _T_1547 = _T_1546 | _T_1491; // @[Mux.scala 27:72]
  wire  _T_1548 = _T_1547 | _T_1492; // @[Mux.scala 27:72]
  wire  _T_1549 = _T_1548 | _T_1493; // @[Mux.scala 27:72]
  wire  _T_1550 = _T_1549 | _T_1494; // @[Mux.scala 27:72]
  wire  _T_1551 = _T_1550 | _T_1495; // @[Mux.scala 27:72]
  wire  _T_1552 = _T_1551 | _T_1496; // @[Mux.scala 27:72]
  wire  _T_1553 = _T_1552 | _T_1476; // @[Mux.scala 27:72]
  wire  _T_1554 = _T_1553 | _T_1498; // @[Mux.scala 27:72]
  wire  _T_1555 = _T_1554 | _T_1499; // @[Mux.scala 27:72]
  wire  _T_1556 = _T_1555 | _T_1500; // @[Mux.scala 27:72]
  wire  _T_1557 = _T_1556 | _T_1501; // @[Mux.scala 27:72]
  wire  _T_1558 = _T_1557 | _T_1502; // @[Mux.scala 27:72]
  wire  _T_1559 = _T_1558 | _T_1503; // @[Mux.scala 27:72]
  wire  _T_1560 = _T_1559 | _T_1504; // @[Mux.scala 27:72]
  wire  _T_1561 = _T_1560 | _T_1505; // @[Mux.scala 27:72]
  wire  _T_1562 = _T_1561 | _T_1506; // @[Mux.scala 27:72]
  wire  _T_1563 = _T_1562 | _T_1507; // @[Mux.scala 27:72]
  wire  _T_1566 = _T_1563 | _T_1510; // @[Mux.scala 27:72]
  wire  _T_1567 = _T_1566 | _T_1511; // @[Mux.scala 27:72]
  wire  _T_1568 = _T_1567 | _T_1512; // @[Mux.scala 27:72]
  wire  _T_1569 = _T_1568 | _T_1513; // @[Mux.scala 27:72]
  wire  _T_1570 = _T_1569 | _T_1514; // @[Mux.scala 27:72]
  wire  _T_1571 = _T_1570 | _T_1515; // @[Mux.scala 27:72]
  wire  _T_1572 = _T_1571 | _T_1516; // @[Mux.scala 27:72]
  wire  _T_1573 = _T_1572 | _T_1517; // @[Mux.scala 27:72]
  wire  _T_1574 = _T_1573 | _T_1518; // @[Mux.scala 27:72]
  wire  _T_1575 = _T_1574 | _T_1519; // @[Mux.scala 27:72]
  wire  _T_1576 = _T_1575 | _T_1520; // @[Mux.scala 27:72]
  wire  _T_1577 = _T_1576 | _T_1521; // @[Mux.scala 27:72]
  wire  _T_1578 = _T_1577 | _T_1522; // @[Mux.scala 27:72]
  wire  _T_1579 = _T_1578 | _T_1523; // @[Mux.scala 27:72]
  wire  _T_1580 = _T_1579 | _T_1524; // @[Mux.scala 27:72]
  wire  mhpmc_inc_r_1 = _T_1300 & _T_1580; // @[dec_tlu_ctl.scala 2274:44]
  wire  _T_1584 = ~mcountinhibit[5]; // @[dec_tlu_ctl.scala 2274:24]
  reg [9:0] mhpme5; // @[Reg.scala 27:20]
  wire  _T_1585 = mhpme5 == 10'h1; // @[dec_tlu_ctl.scala 2275:34]
  wire  _T_1587 = mhpme5 == 10'h2; // @[dec_tlu_ctl.scala 2276:34]
  wire  _T_1589 = mhpme5 == 10'h3; // @[dec_tlu_ctl.scala 2277:34]
  wire  _T_1591 = mhpme5 == 10'h4; // @[dec_tlu_ctl.scala 2278:34]
  wire  _T_1595 = mhpme5 == 10'h5; // @[dec_tlu_ctl.scala 2279:34]
  wire  _T_1601 = mhpme5 == 10'h6; // @[dec_tlu_ctl.scala 2280:34]
  wire  _T_1606 = mhpme5 == 10'h7; // @[dec_tlu_ctl.scala 2281:34]
  wire  _T_1608 = mhpme5 == 10'h8; // @[dec_tlu_ctl.scala 2282:34]
  wire  _T_1610 = mhpme5 == 10'h1e; // @[dec_tlu_ctl.scala 2283:34]
  wire  _T_1612 = mhpme5 == 10'h9; // @[dec_tlu_ctl.scala 2284:34]
  wire  _T_1615 = mhpme5 == 10'ha; // @[dec_tlu_ctl.scala 2285:34]
  wire  _T_1618 = mhpme5 == 10'hb; // @[dec_tlu_ctl.scala 2286:34]
  wire  _T_1621 = mhpme5 == 10'hc; // @[dec_tlu_ctl.scala 2287:34]
  wire  _T_1624 = mhpme5 == 10'hd; // @[dec_tlu_ctl.scala 2288:34]
  wire  _T_1628 = mhpme5 == 10'he; // @[dec_tlu_ctl.scala 2289:34]
  wire  _T_1633 = mhpme5 == 10'hf; // @[dec_tlu_ctl.scala 2290:34]
  wire  _T_1636 = mhpme5 == 10'h10; // @[dec_tlu_ctl.scala 2291:34]
  wire  _T_1639 = mhpme5 == 10'h12; // @[dec_tlu_ctl.scala 2292:34]
  wire  _T_1642 = mhpme5 == 10'h11; // @[dec_tlu_ctl.scala 2293:34]
  wire  _T_1645 = mhpme5 == 10'h13; // @[dec_tlu_ctl.scala 2294:34]
  wire  _T_1648 = mhpme5 == 10'h14; // @[dec_tlu_ctl.scala 2295:34]
  wire  _T_1651 = mhpme5 == 10'h15; // @[dec_tlu_ctl.scala 2296:34]
  wire  _T_1654 = mhpme5 == 10'h16; // @[dec_tlu_ctl.scala 2297:34]
  wire  _T_1657 = mhpme5 == 10'h17; // @[dec_tlu_ctl.scala 2298:34]
  wire  _T_1660 = mhpme5 == 10'h18; // @[dec_tlu_ctl.scala 2299:34]
  wire  _T_1665 = mhpme5 == 10'h19; // @[dec_tlu_ctl.scala 2300:34]
  wire  _T_1668 = mhpme5 == 10'h1a; // @[dec_tlu_ctl.scala 2301:34]
  wire  _T_1671 = mhpme5 == 10'h1b; // @[dec_tlu_ctl.scala 2302:34]
  wire  _T_1674 = mhpme5 == 10'h1c; // @[dec_tlu_ctl.scala 2303:34]
  wire  _T_1678 = mhpme5 == 10'h1f; // @[dec_tlu_ctl.scala 2305:34]
  wire  _T_1680 = mhpme5 == 10'h20; // @[dec_tlu_ctl.scala 2306:34]
  wire  _T_1682 = mhpme5 == 10'h22; // @[dec_tlu_ctl.scala 2307:34]
  wire  _T_1684 = mhpme5 == 10'h23; // @[dec_tlu_ctl.scala 2308:34]
  wire  _T_1686 = mhpme5 == 10'h24; // @[dec_tlu_ctl.scala 2309:34]
  wire  _T_1688 = mhpme5 == 10'h25; // @[dec_tlu_ctl.scala 2310:34]
  wire  _T_1692 = mhpme5 == 10'h26; // @[dec_tlu_ctl.scala 2311:34]
  wire  _T_1696 = mhpme5 == 10'h27; // @[dec_tlu_ctl.scala 2312:34]
  wire  _T_1698 = mhpme5 == 10'h28; // @[dec_tlu_ctl.scala 2313:34]
  wire  _T_1700 = mhpme5 == 10'h29; // @[dec_tlu_ctl.scala 2314:34]
  wire  _T_1708 = mhpme5 == 10'h2c; // @[dec_tlu_ctl.scala 2317:34]
  wire  _T_1710 = mhpme5 == 10'h2d; // @[dec_tlu_ctl.scala 2318:34]
  wire  _T_1712 = mhpme5 == 10'h2e; // @[dec_tlu_ctl.scala 2319:34]
  wire  _T_1714 = mhpme5 == 10'h2f; // @[dec_tlu_ctl.scala 2320:34]
  wire  _T_1716 = mhpme5 == 10'h30; // @[dec_tlu_ctl.scala 2321:34]
  wire  _T_1718 = mhpme5 == 10'h31; // @[dec_tlu_ctl.scala 2322:34]
  wire  _T_1723 = mhpme5 == 10'h32; // @[dec_tlu_ctl.scala 2323:34]
  wire  _T_1733 = mhpme5 == 10'h36; // @[dec_tlu_ctl.scala 2324:34]
  wire  _T_1736 = mhpme5 == 10'h37; // @[dec_tlu_ctl.scala 2325:34]
  wire  _T_1739 = mhpme5 == 10'h38; // @[dec_tlu_ctl.scala 2326:34]
  wire  _T_1742 = mhpme5 == 10'h200; // @[dec_tlu_ctl.scala 2328:34]
  wire  _T_1744 = mhpme5 == 10'h201; // @[dec_tlu_ctl.scala 2329:34]
  wire  _T_1746 = mhpme5 == 10'h202; // @[dec_tlu_ctl.scala 2330:34]
  wire  _T_1748 = mhpme5 == 10'h203; // @[dec_tlu_ctl.scala 2331:34]
  wire  _T_1750 = mhpme5 == 10'h204; // @[dec_tlu_ctl.scala 2332:34]
  wire  _T_1753 = _T_1587 & io_ifu_pmu_ic_hit; // @[Mux.scala 27:72]
  wire  _T_1754 = _T_1589 & io_ifu_pmu_ic_miss; // @[Mux.scala 27:72]
  wire  _T_1755 = _T_1591 & _T_1026; // @[Mux.scala 27:72]
  wire  _T_1756 = _T_1595 & _T_1032; // @[Mux.scala 27:72]
  wire  _T_1757 = _T_1601 & _T_1037; // @[Mux.scala 27:72]
  wire  _T_1758 = _T_1606 & io_ifu_pmu_instr_aligned; // @[Mux.scala 27:72]
  wire  _T_1759 = _T_1608 & io_dec_pmu_instr_decoded; // @[Mux.scala 27:72]
  wire  _T_1760 = _T_1610 & io_dec_pmu_decode_stall; // @[Mux.scala 27:72]
  wire  _T_1761 = _T_1612 & _T_1046; // @[Mux.scala 27:72]
  wire  _T_1762 = _T_1615 & _T_1049; // @[Mux.scala 27:72]
  wire  _T_1763 = _T_1618 & _T_1052; // @[Mux.scala 27:72]
  wire  _T_1764 = _T_1621 & _T_1055; // @[Mux.scala 27:72]
  wire  _T_1765 = _T_1624 & _T_1059; // @[Mux.scala 27:72]
  wire  _T_1766 = _T_1628 & _T_1064; // @[Mux.scala 27:72]
  wire  _T_1767 = _T_1633 & _T_1067; // @[Mux.scala 27:72]
  wire  _T_1768 = _T_1636 & _T_1070; // @[Mux.scala 27:72]
  wire  _T_1769 = _T_1639 & _T_1073; // @[Mux.scala 27:72]
  wire  _T_1770 = _T_1642 & _T_1076; // @[Mux.scala 27:72]
  wire  _T_1771 = _T_1645 & _T_1079; // @[Mux.scala 27:72]
  wire  _T_1772 = _T_1648 & _T_1082; // @[Mux.scala 27:72]
  wire  _T_1773 = _T_1651 & _T_1085; // @[Mux.scala 27:72]
  wire  _T_1774 = _T_1654 & _T_1088; // @[Mux.scala 27:72]
  wire  _T_1775 = _T_1657 & _T_1091; // @[Mux.scala 27:72]
  wire  _T_1776 = _T_1660 & _T_1096; // @[Mux.scala 27:72]
  wire  _T_1777 = _T_1665 & _T_1099; // @[Mux.scala 27:72]
  wire  _T_1778 = _T_1668 & _T_1102; // @[Mux.scala 27:72]
  wire  _T_1779 = _T_1671 & _T_1105; // @[Mux.scala 27:72]
  wire  _T_1780 = _T_1674 & io_ifu_pmu_fetch_stall; // @[Mux.scala 27:72]
  wire  _T_1782 = _T_1678 & io_dec_pmu_postsync_stall; // @[Mux.scala 27:72]
  wire  _T_1783 = _T_1680 & io_dec_pmu_presync_stall; // @[Mux.scala 27:72]
  wire  _T_1784 = _T_1682 & io_lsu_store_stall_any; // @[Mux.scala 27:72]
  wire  _T_1785 = _T_1684 & io_dma_dccm_stall_any; // @[Mux.scala 27:72]
  wire  _T_1786 = _T_1686 & io_dma_iccm_stall_any; // @[Mux.scala 27:72]
  wire  _T_1787 = _T_1688 & _T_1123; // @[Mux.scala 27:72]
  wire  _T_1788 = _T_1692 & _T_1127; // @[Mux.scala 27:72]
  wire  _T_1789 = _T_1696 & io_take_ext_int; // @[Mux.scala 27:72]
  wire  _T_1790 = _T_1698 & io_tlu_flush_lower_r; // @[Mux.scala 27:72]
  wire  _T_1791 = _T_1700 & _T_1135; // @[Mux.scala 27:72]
  wire  _T_1794 = _T_1708 & io_lsu_pmu_bus_misaligned; // @[Mux.scala 27:72]
  wire  _T_1795 = _T_1710 & io_ifu_pmu_bus_error; // @[Mux.scala 27:72]
  wire  _T_1796 = _T_1712 & io_lsu_pmu_bus_error; // @[Mux.scala 27:72]
  wire  _T_1797 = _T_1714 & io_ifu_pmu_bus_busy; // @[Mux.scala 27:72]
  wire  _T_1798 = _T_1716 & io_lsu_pmu_bus_busy; // @[Mux.scala 27:72]
  wire  _T_1799 = _T_1718 & _T_1154; // @[Mux.scala 27:72]
  wire  _T_1800 = _T_1723 & _T_1164; // @[Mux.scala 27:72]
  wire  _T_1801 = _T_1733 & _T_1167; // @[Mux.scala 27:72]
  wire  _T_1802 = _T_1736 & _T_1170; // @[Mux.scala 27:72]
  wire  _T_1803 = _T_1739 & _T_1173; // @[Mux.scala 27:72]
  wire  _T_1804 = _T_1742 & io_dec_tlu_pmu_fw_halted; // @[Mux.scala 27:72]
  wire  _T_1805 = _T_1744 & io_dma_pmu_any_read; // @[Mux.scala 27:72]
  wire  _T_1806 = _T_1746 & io_dma_pmu_any_write; // @[Mux.scala 27:72]
  wire  _T_1807 = _T_1748 & io_dma_pmu_dccm_read; // @[Mux.scala 27:72]
  wire  _T_1808 = _T_1750 & io_dma_pmu_dccm_write; // @[Mux.scala 27:72]
  wire  _T_1809 = _T_1585 | _T_1753; // @[Mux.scala 27:72]
  wire  _T_1810 = _T_1809 | _T_1754; // @[Mux.scala 27:72]
  wire  _T_1811 = _T_1810 | _T_1755; // @[Mux.scala 27:72]
  wire  _T_1812 = _T_1811 | _T_1756; // @[Mux.scala 27:72]
  wire  _T_1813 = _T_1812 | _T_1757; // @[Mux.scala 27:72]
  wire  _T_1814 = _T_1813 | _T_1758; // @[Mux.scala 27:72]
  wire  _T_1815 = _T_1814 | _T_1759; // @[Mux.scala 27:72]
  wire  _T_1816 = _T_1815 | _T_1760; // @[Mux.scala 27:72]
  wire  _T_1817 = _T_1816 | _T_1761; // @[Mux.scala 27:72]
  wire  _T_1818 = _T_1817 | _T_1762; // @[Mux.scala 27:72]
  wire  _T_1819 = _T_1818 | _T_1763; // @[Mux.scala 27:72]
  wire  _T_1820 = _T_1819 | _T_1764; // @[Mux.scala 27:72]
  wire  _T_1821 = _T_1820 | _T_1765; // @[Mux.scala 27:72]
  wire  _T_1822 = _T_1821 | _T_1766; // @[Mux.scala 27:72]
  wire  _T_1823 = _T_1822 | _T_1767; // @[Mux.scala 27:72]
  wire  _T_1824 = _T_1823 | _T_1768; // @[Mux.scala 27:72]
  wire  _T_1825 = _T_1824 | _T_1769; // @[Mux.scala 27:72]
  wire  _T_1826 = _T_1825 | _T_1770; // @[Mux.scala 27:72]
  wire  _T_1827 = _T_1826 | _T_1771; // @[Mux.scala 27:72]
  wire  _T_1828 = _T_1827 | _T_1772; // @[Mux.scala 27:72]
  wire  _T_1829 = _T_1828 | _T_1773; // @[Mux.scala 27:72]
  wire  _T_1830 = _T_1829 | _T_1774; // @[Mux.scala 27:72]
  wire  _T_1831 = _T_1830 | _T_1775; // @[Mux.scala 27:72]
  wire  _T_1832 = _T_1831 | _T_1776; // @[Mux.scala 27:72]
  wire  _T_1833 = _T_1832 | _T_1777; // @[Mux.scala 27:72]
  wire  _T_1834 = _T_1833 | _T_1778; // @[Mux.scala 27:72]
  wire  _T_1835 = _T_1834 | _T_1779; // @[Mux.scala 27:72]
  wire  _T_1836 = _T_1835 | _T_1780; // @[Mux.scala 27:72]
  wire  _T_1837 = _T_1836 | _T_1760; // @[Mux.scala 27:72]
  wire  _T_1838 = _T_1837 | _T_1782; // @[Mux.scala 27:72]
  wire  _T_1839 = _T_1838 | _T_1783; // @[Mux.scala 27:72]
  wire  _T_1840 = _T_1839 | _T_1784; // @[Mux.scala 27:72]
  wire  _T_1841 = _T_1840 | _T_1785; // @[Mux.scala 27:72]
  wire  _T_1842 = _T_1841 | _T_1786; // @[Mux.scala 27:72]
  wire  _T_1843 = _T_1842 | _T_1787; // @[Mux.scala 27:72]
  wire  _T_1844 = _T_1843 | _T_1788; // @[Mux.scala 27:72]
  wire  _T_1845 = _T_1844 | _T_1789; // @[Mux.scala 27:72]
  wire  _T_1846 = _T_1845 | _T_1790; // @[Mux.scala 27:72]
  wire  _T_1847 = _T_1846 | _T_1791; // @[Mux.scala 27:72]
  wire  _T_1850 = _T_1847 | _T_1794; // @[Mux.scala 27:72]
  wire  _T_1851 = _T_1850 | _T_1795; // @[Mux.scala 27:72]
  wire  _T_1852 = _T_1851 | _T_1796; // @[Mux.scala 27:72]
  wire  _T_1853 = _T_1852 | _T_1797; // @[Mux.scala 27:72]
  wire  _T_1854 = _T_1853 | _T_1798; // @[Mux.scala 27:72]
  wire  _T_1855 = _T_1854 | _T_1799; // @[Mux.scala 27:72]
  wire  _T_1856 = _T_1855 | _T_1800; // @[Mux.scala 27:72]
  wire  _T_1857 = _T_1856 | _T_1801; // @[Mux.scala 27:72]
  wire  _T_1858 = _T_1857 | _T_1802; // @[Mux.scala 27:72]
  wire  _T_1859 = _T_1858 | _T_1803; // @[Mux.scala 27:72]
  wire  _T_1860 = _T_1859 | _T_1804; // @[Mux.scala 27:72]
  wire  _T_1861 = _T_1860 | _T_1805; // @[Mux.scala 27:72]
  wire  _T_1862 = _T_1861 | _T_1806; // @[Mux.scala 27:72]
  wire  _T_1863 = _T_1862 | _T_1807; // @[Mux.scala 27:72]
  wire  _T_1864 = _T_1863 | _T_1808; // @[Mux.scala 27:72]
  wire  mhpmc_inc_r_2 = _T_1584 & _T_1864; // @[dec_tlu_ctl.scala 2274:44]
  wire  _T_1868 = ~mcountinhibit[6]; // @[dec_tlu_ctl.scala 2274:24]
  reg [9:0] mhpme6; // @[Reg.scala 27:20]
  wire  _T_1869 = mhpme6 == 10'h1; // @[dec_tlu_ctl.scala 2275:34]
  wire  _T_1871 = mhpme6 == 10'h2; // @[dec_tlu_ctl.scala 2276:34]
  wire  _T_1873 = mhpme6 == 10'h3; // @[dec_tlu_ctl.scala 2277:34]
  wire  _T_1875 = mhpme6 == 10'h4; // @[dec_tlu_ctl.scala 2278:34]
  wire  _T_1879 = mhpme6 == 10'h5; // @[dec_tlu_ctl.scala 2279:34]
  wire  _T_1885 = mhpme6 == 10'h6; // @[dec_tlu_ctl.scala 2280:34]
  wire  _T_1890 = mhpme6 == 10'h7; // @[dec_tlu_ctl.scala 2281:34]
  wire  _T_1892 = mhpme6 == 10'h8; // @[dec_tlu_ctl.scala 2282:34]
  wire  _T_1894 = mhpme6 == 10'h1e; // @[dec_tlu_ctl.scala 2283:34]
  wire  _T_1896 = mhpme6 == 10'h9; // @[dec_tlu_ctl.scala 2284:34]
  wire  _T_1899 = mhpme6 == 10'ha; // @[dec_tlu_ctl.scala 2285:34]
  wire  _T_1902 = mhpme6 == 10'hb; // @[dec_tlu_ctl.scala 2286:34]
  wire  _T_1905 = mhpme6 == 10'hc; // @[dec_tlu_ctl.scala 2287:34]
  wire  _T_1908 = mhpme6 == 10'hd; // @[dec_tlu_ctl.scala 2288:34]
  wire  _T_1912 = mhpme6 == 10'he; // @[dec_tlu_ctl.scala 2289:34]
  wire  _T_1917 = mhpme6 == 10'hf; // @[dec_tlu_ctl.scala 2290:34]
  wire  _T_1920 = mhpme6 == 10'h10; // @[dec_tlu_ctl.scala 2291:34]
  wire  _T_1923 = mhpme6 == 10'h12; // @[dec_tlu_ctl.scala 2292:34]
  wire  _T_1926 = mhpme6 == 10'h11; // @[dec_tlu_ctl.scala 2293:34]
  wire  _T_1929 = mhpme6 == 10'h13; // @[dec_tlu_ctl.scala 2294:34]
  wire  _T_1932 = mhpme6 == 10'h14; // @[dec_tlu_ctl.scala 2295:34]
  wire  _T_1935 = mhpme6 == 10'h15; // @[dec_tlu_ctl.scala 2296:34]
  wire  _T_1938 = mhpme6 == 10'h16; // @[dec_tlu_ctl.scala 2297:34]
  wire  _T_1941 = mhpme6 == 10'h17; // @[dec_tlu_ctl.scala 2298:34]
  wire  _T_1944 = mhpme6 == 10'h18; // @[dec_tlu_ctl.scala 2299:34]
  wire  _T_1949 = mhpme6 == 10'h19; // @[dec_tlu_ctl.scala 2300:34]
  wire  _T_1952 = mhpme6 == 10'h1a; // @[dec_tlu_ctl.scala 2301:34]
  wire  _T_1955 = mhpme6 == 10'h1b; // @[dec_tlu_ctl.scala 2302:34]
  wire  _T_1958 = mhpme6 == 10'h1c; // @[dec_tlu_ctl.scala 2303:34]
  wire  _T_1962 = mhpme6 == 10'h1f; // @[dec_tlu_ctl.scala 2305:34]
  wire  _T_1964 = mhpme6 == 10'h20; // @[dec_tlu_ctl.scala 2306:34]
  wire  _T_1966 = mhpme6 == 10'h22; // @[dec_tlu_ctl.scala 2307:34]
  wire  _T_1968 = mhpme6 == 10'h23; // @[dec_tlu_ctl.scala 2308:34]
  wire  _T_1970 = mhpme6 == 10'h24; // @[dec_tlu_ctl.scala 2309:34]
  wire  _T_1972 = mhpme6 == 10'h25; // @[dec_tlu_ctl.scala 2310:34]
  wire  _T_1976 = mhpme6 == 10'h26; // @[dec_tlu_ctl.scala 2311:34]
  wire  _T_1980 = mhpme6 == 10'h27; // @[dec_tlu_ctl.scala 2312:34]
  wire  _T_1982 = mhpme6 == 10'h28; // @[dec_tlu_ctl.scala 2313:34]
  wire  _T_1984 = mhpme6 == 10'h29; // @[dec_tlu_ctl.scala 2314:34]
  wire  _T_1992 = mhpme6 == 10'h2c; // @[dec_tlu_ctl.scala 2317:34]
  wire  _T_1994 = mhpme6 == 10'h2d; // @[dec_tlu_ctl.scala 2318:34]
  wire  _T_1996 = mhpme6 == 10'h2e; // @[dec_tlu_ctl.scala 2319:34]
  wire  _T_1998 = mhpme6 == 10'h2f; // @[dec_tlu_ctl.scala 2320:34]
  wire  _T_2000 = mhpme6 == 10'h30; // @[dec_tlu_ctl.scala 2321:34]
  wire  _T_2002 = mhpme6 == 10'h31; // @[dec_tlu_ctl.scala 2322:34]
  wire  _T_2007 = mhpme6 == 10'h32; // @[dec_tlu_ctl.scala 2323:34]
  wire  _T_2017 = mhpme6 == 10'h36; // @[dec_tlu_ctl.scala 2324:34]
  wire  _T_2020 = mhpme6 == 10'h37; // @[dec_tlu_ctl.scala 2325:34]
  wire  _T_2023 = mhpme6 == 10'h38; // @[dec_tlu_ctl.scala 2326:34]
  wire  _T_2026 = mhpme6 == 10'h200; // @[dec_tlu_ctl.scala 2328:34]
  wire  _T_2028 = mhpme6 == 10'h201; // @[dec_tlu_ctl.scala 2329:34]
  wire  _T_2030 = mhpme6 == 10'h202; // @[dec_tlu_ctl.scala 2330:34]
  wire  _T_2032 = mhpme6 == 10'h203; // @[dec_tlu_ctl.scala 2331:34]
  wire  _T_2034 = mhpme6 == 10'h204; // @[dec_tlu_ctl.scala 2332:34]
  wire  _T_2037 = _T_1871 & io_ifu_pmu_ic_hit; // @[Mux.scala 27:72]
  wire  _T_2038 = _T_1873 & io_ifu_pmu_ic_miss; // @[Mux.scala 27:72]
  wire  _T_2039 = _T_1875 & _T_1026; // @[Mux.scala 27:72]
  wire  _T_2040 = _T_1879 & _T_1032; // @[Mux.scala 27:72]
  wire  _T_2041 = _T_1885 & _T_1037; // @[Mux.scala 27:72]
  wire  _T_2042 = _T_1890 & io_ifu_pmu_instr_aligned; // @[Mux.scala 27:72]
  wire  _T_2043 = _T_1892 & io_dec_pmu_instr_decoded; // @[Mux.scala 27:72]
  wire  _T_2044 = _T_1894 & io_dec_pmu_decode_stall; // @[Mux.scala 27:72]
  wire  _T_2045 = _T_1896 & _T_1046; // @[Mux.scala 27:72]
  wire  _T_2046 = _T_1899 & _T_1049; // @[Mux.scala 27:72]
  wire  _T_2047 = _T_1902 & _T_1052; // @[Mux.scala 27:72]
  wire  _T_2048 = _T_1905 & _T_1055; // @[Mux.scala 27:72]
  wire  _T_2049 = _T_1908 & _T_1059; // @[Mux.scala 27:72]
  wire  _T_2050 = _T_1912 & _T_1064; // @[Mux.scala 27:72]
  wire  _T_2051 = _T_1917 & _T_1067; // @[Mux.scala 27:72]
  wire  _T_2052 = _T_1920 & _T_1070; // @[Mux.scala 27:72]
  wire  _T_2053 = _T_1923 & _T_1073; // @[Mux.scala 27:72]
  wire  _T_2054 = _T_1926 & _T_1076; // @[Mux.scala 27:72]
  wire  _T_2055 = _T_1929 & _T_1079; // @[Mux.scala 27:72]
  wire  _T_2056 = _T_1932 & _T_1082; // @[Mux.scala 27:72]
  wire  _T_2057 = _T_1935 & _T_1085; // @[Mux.scala 27:72]
  wire  _T_2058 = _T_1938 & _T_1088; // @[Mux.scala 27:72]
  wire  _T_2059 = _T_1941 & _T_1091; // @[Mux.scala 27:72]
  wire  _T_2060 = _T_1944 & _T_1096; // @[Mux.scala 27:72]
  wire  _T_2061 = _T_1949 & _T_1099; // @[Mux.scala 27:72]
  wire  _T_2062 = _T_1952 & _T_1102; // @[Mux.scala 27:72]
  wire  _T_2063 = _T_1955 & _T_1105; // @[Mux.scala 27:72]
  wire  _T_2064 = _T_1958 & io_ifu_pmu_fetch_stall; // @[Mux.scala 27:72]
  wire  _T_2066 = _T_1962 & io_dec_pmu_postsync_stall; // @[Mux.scala 27:72]
  wire  _T_2067 = _T_1964 & io_dec_pmu_presync_stall; // @[Mux.scala 27:72]
  wire  _T_2068 = _T_1966 & io_lsu_store_stall_any; // @[Mux.scala 27:72]
  wire  _T_2069 = _T_1968 & io_dma_dccm_stall_any; // @[Mux.scala 27:72]
  wire  _T_2070 = _T_1970 & io_dma_iccm_stall_any; // @[Mux.scala 27:72]
  wire  _T_2071 = _T_1972 & _T_1123; // @[Mux.scala 27:72]
  wire  _T_2072 = _T_1976 & _T_1127; // @[Mux.scala 27:72]
  wire  _T_2073 = _T_1980 & io_take_ext_int; // @[Mux.scala 27:72]
  wire  _T_2074 = _T_1982 & io_tlu_flush_lower_r; // @[Mux.scala 27:72]
  wire  _T_2075 = _T_1984 & _T_1135; // @[Mux.scala 27:72]
  wire  _T_2078 = _T_1992 & io_lsu_pmu_bus_misaligned; // @[Mux.scala 27:72]
  wire  _T_2079 = _T_1994 & io_ifu_pmu_bus_error; // @[Mux.scala 27:72]
  wire  _T_2080 = _T_1996 & io_lsu_pmu_bus_error; // @[Mux.scala 27:72]
  wire  _T_2081 = _T_1998 & io_ifu_pmu_bus_busy; // @[Mux.scala 27:72]
  wire  _T_2082 = _T_2000 & io_lsu_pmu_bus_busy; // @[Mux.scala 27:72]
  wire  _T_2083 = _T_2002 & _T_1154; // @[Mux.scala 27:72]
  wire  _T_2084 = _T_2007 & _T_1164; // @[Mux.scala 27:72]
  wire  _T_2085 = _T_2017 & _T_1167; // @[Mux.scala 27:72]
  wire  _T_2086 = _T_2020 & _T_1170; // @[Mux.scala 27:72]
  wire  _T_2087 = _T_2023 & _T_1173; // @[Mux.scala 27:72]
  wire  _T_2088 = _T_2026 & io_dec_tlu_pmu_fw_halted; // @[Mux.scala 27:72]
  wire  _T_2089 = _T_2028 & io_dma_pmu_any_read; // @[Mux.scala 27:72]
  wire  _T_2090 = _T_2030 & io_dma_pmu_any_write; // @[Mux.scala 27:72]
  wire  _T_2091 = _T_2032 & io_dma_pmu_dccm_read; // @[Mux.scala 27:72]
  wire  _T_2092 = _T_2034 & io_dma_pmu_dccm_write; // @[Mux.scala 27:72]
  wire  _T_2093 = _T_1869 | _T_2037; // @[Mux.scala 27:72]
  wire  _T_2094 = _T_2093 | _T_2038; // @[Mux.scala 27:72]
  wire  _T_2095 = _T_2094 | _T_2039; // @[Mux.scala 27:72]
  wire  _T_2096 = _T_2095 | _T_2040; // @[Mux.scala 27:72]
  wire  _T_2097 = _T_2096 | _T_2041; // @[Mux.scala 27:72]
  wire  _T_2098 = _T_2097 | _T_2042; // @[Mux.scala 27:72]
  wire  _T_2099 = _T_2098 | _T_2043; // @[Mux.scala 27:72]
  wire  _T_2100 = _T_2099 | _T_2044; // @[Mux.scala 27:72]
  wire  _T_2101 = _T_2100 | _T_2045; // @[Mux.scala 27:72]
  wire  _T_2102 = _T_2101 | _T_2046; // @[Mux.scala 27:72]
  wire  _T_2103 = _T_2102 | _T_2047; // @[Mux.scala 27:72]
  wire  _T_2104 = _T_2103 | _T_2048; // @[Mux.scala 27:72]
  wire  _T_2105 = _T_2104 | _T_2049; // @[Mux.scala 27:72]
  wire  _T_2106 = _T_2105 | _T_2050; // @[Mux.scala 27:72]
  wire  _T_2107 = _T_2106 | _T_2051; // @[Mux.scala 27:72]
  wire  _T_2108 = _T_2107 | _T_2052; // @[Mux.scala 27:72]
  wire  _T_2109 = _T_2108 | _T_2053; // @[Mux.scala 27:72]
  wire  _T_2110 = _T_2109 | _T_2054; // @[Mux.scala 27:72]
  wire  _T_2111 = _T_2110 | _T_2055; // @[Mux.scala 27:72]
  wire  _T_2112 = _T_2111 | _T_2056; // @[Mux.scala 27:72]
  wire  _T_2113 = _T_2112 | _T_2057; // @[Mux.scala 27:72]
  wire  _T_2114 = _T_2113 | _T_2058; // @[Mux.scala 27:72]
  wire  _T_2115 = _T_2114 | _T_2059; // @[Mux.scala 27:72]
  wire  _T_2116 = _T_2115 | _T_2060; // @[Mux.scala 27:72]
  wire  _T_2117 = _T_2116 | _T_2061; // @[Mux.scala 27:72]
  wire  _T_2118 = _T_2117 | _T_2062; // @[Mux.scala 27:72]
  wire  _T_2119 = _T_2118 | _T_2063; // @[Mux.scala 27:72]
  wire  _T_2120 = _T_2119 | _T_2064; // @[Mux.scala 27:72]
  wire  _T_2121 = _T_2120 | _T_2044; // @[Mux.scala 27:72]
  wire  _T_2122 = _T_2121 | _T_2066; // @[Mux.scala 27:72]
  wire  _T_2123 = _T_2122 | _T_2067; // @[Mux.scala 27:72]
  wire  _T_2124 = _T_2123 | _T_2068; // @[Mux.scala 27:72]
  wire  _T_2125 = _T_2124 | _T_2069; // @[Mux.scala 27:72]
  wire  _T_2126 = _T_2125 | _T_2070; // @[Mux.scala 27:72]
  wire  _T_2127 = _T_2126 | _T_2071; // @[Mux.scala 27:72]
  wire  _T_2128 = _T_2127 | _T_2072; // @[Mux.scala 27:72]
  wire  _T_2129 = _T_2128 | _T_2073; // @[Mux.scala 27:72]
  wire  _T_2130 = _T_2129 | _T_2074; // @[Mux.scala 27:72]
  wire  _T_2131 = _T_2130 | _T_2075; // @[Mux.scala 27:72]
  wire  _T_2134 = _T_2131 | _T_2078; // @[Mux.scala 27:72]
  wire  _T_2135 = _T_2134 | _T_2079; // @[Mux.scala 27:72]
  wire  _T_2136 = _T_2135 | _T_2080; // @[Mux.scala 27:72]
  wire  _T_2137 = _T_2136 | _T_2081; // @[Mux.scala 27:72]
  wire  _T_2138 = _T_2137 | _T_2082; // @[Mux.scala 27:72]
  wire  _T_2139 = _T_2138 | _T_2083; // @[Mux.scala 27:72]
  wire  _T_2140 = _T_2139 | _T_2084; // @[Mux.scala 27:72]
  wire  _T_2141 = _T_2140 | _T_2085; // @[Mux.scala 27:72]
  wire  _T_2142 = _T_2141 | _T_2086; // @[Mux.scala 27:72]
  wire  _T_2143 = _T_2142 | _T_2087; // @[Mux.scala 27:72]
  wire  _T_2144 = _T_2143 | _T_2088; // @[Mux.scala 27:72]
  wire  _T_2145 = _T_2144 | _T_2089; // @[Mux.scala 27:72]
  wire  _T_2146 = _T_2145 | _T_2090; // @[Mux.scala 27:72]
  wire  _T_2147 = _T_2146 | _T_2091; // @[Mux.scala 27:72]
  wire  _T_2148 = _T_2147 | _T_2092; // @[Mux.scala 27:72]
  wire  mhpmc_inc_r_3 = _T_1868 & _T_2148; // @[dec_tlu_ctl.scala 2274:44]
  reg  mhpmc_inc_r_d1_0; // @[dec_tlu_ctl.scala 2335:53]
  reg  mhpmc_inc_r_d1_1; // @[dec_tlu_ctl.scala 2336:53]
  reg  mhpmc_inc_r_d1_2; // @[dec_tlu_ctl.scala 2337:53]
  reg  mhpmc_inc_r_d1_3; // @[dec_tlu_ctl.scala 2338:53]
  reg  perfcnt_halted_d1; // @[dec_tlu_ctl.scala 2339:56]
  wire  perfcnt_halted = _T_85 | io_dec_tlu_pmu_fw_halted; // @[dec_tlu_ctl.scala 2342:67]
  wire  _T_2160 = ~_T_85; // @[dec_tlu_ctl.scala 2343:37]
  wire [3:0] _T_2162 = _T_2160 ? 4'hf : 4'h0; // @[Bitwise.scala 72:12]
  wire [3:0] _T_2169 = {mhpme6[9],mhpme5[9],mhpme4[9],mhpme3[9]}; // @[Cat.scala 29:58]
  wire [3:0] perfcnt_during_sleep = _T_2162 & _T_2169; // @[dec_tlu_ctl.scala 2343:86]
  wire  _T_2171 = ~perfcnt_during_sleep[0]; // @[dec_tlu_ctl.scala 2345:67]
  wire  _T_2172 = perfcnt_halted_d1 & _T_2171; // @[dec_tlu_ctl.scala 2345:65]
  wire  _T_2173 = ~_T_2172; // @[dec_tlu_ctl.scala 2345:45]
  wire  _T_2176 = ~perfcnt_during_sleep[1]; // @[dec_tlu_ctl.scala 2346:67]
  wire  _T_2177 = perfcnt_halted_d1 & _T_2176; // @[dec_tlu_ctl.scala 2346:65]
  wire  _T_2178 = ~_T_2177; // @[dec_tlu_ctl.scala 2346:45]
  wire  _T_2181 = ~perfcnt_during_sleep[2]; // @[dec_tlu_ctl.scala 2347:67]
  wire  _T_2182 = perfcnt_halted_d1 & _T_2181; // @[dec_tlu_ctl.scala 2347:65]
  wire  _T_2183 = ~_T_2182; // @[dec_tlu_ctl.scala 2347:45]
  wire  _T_2186 = ~perfcnt_during_sleep[3]; // @[dec_tlu_ctl.scala 2348:67]
  wire  _T_2187 = perfcnt_halted_d1 & _T_2186; // @[dec_tlu_ctl.scala 2348:65]
  wire  _T_2188 = ~_T_2187; // @[dec_tlu_ctl.scala 2348:45]
  wire  _T_2191 = io_dec_csr_wraddr_r == 12'hb03; // @[dec_tlu_ctl.scala 2354:72]
  wire  mhpmc3_wr_en0 = io_dec_csr_wen_r_mod & _T_2191; // @[dec_tlu_ctl.scala 2354:43]
  wire  _T_2192 = ~perfcnt_halted; // @[dec_tlu_ctl.scala 2355:23]
  wire  _T_2194 = _T_2192 | perfcnt_during_sleep[0]; // @[dec_tlu_ctl.scala 2355:39]
  wire  _T_2195 = |mhpmc_inc_r_0; // @[dec_tlu_ctl.scala 2355:86]
  wire  mhpmc3_wr_en1 = _T_2194 & _T_2195; // @[dec_tlu_ctl.scala 2355:66]
  reg [31:0] mhpmc3h; // @[lib.scala 374:16]
  reg [31:0] mhpmc3; // @[lib.scala 374:16]
  wire [63:0] _T_2198 = {mhpmc3h,mhpmc3}; // @[Cat.scala 29:58]
  wire [63:0] _T_2199 = {63'h0,mhpmc_inc_r_0}; // @[Cat.scala 29:58]
  wire [63:0] mhpmc3_incr = _T_2198 + _T_2199; // @[dec_tlu_ctl.scala 2359:49]
  wire  _T_2207 = io_dec_csr_wraddr_r == 12'hb83; // @[dec_tlu_ctl.scala 2364:73]
  wire  mhpmc3h_wr_en0 = io_dec_csr_wen_r_mod & _T_2207; // @[dec_tlu_ctl.scala 2364:44]
  wire  _T_2213 = io_dec_csr_wraddr_r == 12'hb04; // @[dec_tlu_ctl.scala 2373:72]
  wire  mhpmc4_wr_en0 = io_dec_csr_wen_r_mod & _T_2213; // @[dec_tlu_ctl.scala 2373:43]
  wire  _T_2216 = _T_2192 | perfcnt_during_sleep[1]; // @[dec_tlu_ctl.scala 2374:39]
  wire  _T_2217 = |mhpmc_inc_r_1; // @[dec_tlu_ctl.scala 2374:86]
  wire  mhpmc4_wr_en1 = _T_2216 & _T_2217; // @[dec_tlu_ctl.scala 2374:66]
  reg [31:0] mhpmc4h; // @[lib.scala 374:16]
  reg [31:0] mhpmc4; // @[lib.scala 374:16]
  wire [63:0] _T_2220 = {mhpmc4h,mhpmc4}; // @[Cat.scala 29:58]
  wire [63:0] _T_2221 = {63'h0,mhpmc_inc_r_1}; // @[Cat.scala 29:58]
  wire [63:0] mhpmc4_incr = _T_2220 + _T_2221; // @[dec_tlu_ctl.scala 2379:49]
  wire  _T_2230 = io_dec_csr_wraddr_r == 12'hb84; // @[dec_tlu_ctl.scala 2383:73]
  wire  mhpmc4h_wr_en0 = io_dec_csr_wen_r_mod & _T_2230; // @[dec_tlu_ctl.scala 2383:44]
  wire  _T_2236 = io_dec_csr_wraddr_r == 12'hb05; // @[dec_tlu_ctl.scala 2392:72]
  wire  mhpmc5_wr_en0 = io_dec_csr_wen_r_mod & _T_2236; // @[dec_tlu_ctl.scala 2392:43]
  wire  _T_2239 = _T_2192 | perfcnt_during_sleep[2]; // @[dec_tlu_ctl.scala 2393:39]
  wire  _T_2240 = |mhpmc_inc_r_2; // @[dec_tlu_ctl.scala 2393:86]
  wire  mhpmc5_wr_en1 = _T_2239 & _T_2240; // @[dec_tlu_ctl.scala 2393:66]
  reg [31:0] mhpmc5h; // @[lib.scala 374:16]
  reg [31:0] mhpmc5; // @[lib.scala 374:16]
  wire [63:0] _T_2243 = {mhpmc5h,mhpmc5}; // @[Cat.scala 29:58]
  wire [63:0] _T_2244 = {63'h0,mhpmc_inc_r_2}; // @[Cat.scala 29:58]
  wire [63:0] mhpmc5_incr = _T_2243 + _T_2244; // @[dec_tlu_ctl.scala 2396:49]
  wire  _T_2252 = io_dec_csr_wraddr_r == 12'hb85; // @[dec_tlu_ctl.scala 2401:73]
  wire  mhpmc5h_wr_en0 = io_dec_csr_wen_r_mod & _T_2252; // @[dec_tlu_ctl.scala 2401:44]
  wire  _T_2258 = io_dec_csr_wraddr_r == 12'hb06; // @[dec_tlu_ctl.scala 2410:72]
  wire  mhpmc6_wr_en0 = io_dec_csr_wen_r_mod & _T_2258; // @[dec_tlu_ctl.scala 2410:43]
  wire  _T_2261 = _T_2192 | perfcnt_during_sleep[3]; // @[dec_tlu_ctl.scala 2411:39]
  wire  _T_2262 = |mhpmc_inc_r_3; // @[dec_tlu_ctl.scala 2411:86]
  wire  mhpmc6_wr_en1 = _T_2261 & _T_2262; // @[dec_tlu_ctl.scala 2411:66]
  reg [31:0] mhpmc6h; // @[lib.scala 374:16]
  reg [31:0] mhpmc6; // @[lib.scala 374:16]
  wire [63:0] _T_2265 = {mhpmc6h,mhpmc6}; // @[Cat.scala 29:58]
  wire [63:0] _T_2266 = {63'h0,mhpmc_inc_r_3}; // @[Cat.scala 29:58]
  wire [63:0] mhpmc6_incr = _T_2265 + _T_2266; // @[dec_tlu_ctl.scala 2414:49]
  wire  _T_2274 = io_dec_csr_wraddr_r == 12'hb86; // @[dec_tlu_ctl.scala 2419:73]
  wire  mhpmc6h_wr_en0 = io_dec_csr_wen_r_mod & _T_2274; // @[dec_tlu_ctl.scala 2419:44]
  wire  _T_2280 = io_dec_csr_wrdata_r[9:0] > 10'h204; // @[dec_tlu_ctl.scala 2430:56]
  wire  _T_2282 = |io_dec_csr_wrdata_r[31:10]; // @[dec_tlu_ctl.scala 2430:102]
  wire  _T_2283 = _T_2280 | _T_2282; // @[dec_tlu_ctl.scala 2430:71]
  wire  _T_2286 = io_dec_csr_wraddr_r == 12'h323; // @[dec_tlu_ctl.scala 2432:70]
  wire  wr_mhpme3_r = io_dec_csr_wen_r_mod & _T_2286; // @[dec_tlu_ctl.scala 2432:41]
  wire  _T_2290 = io_dec_csr_wraddr_r == 12'h324; // @[dec_tlu_ctl.scala 2439:70]
  wire  wr_mhpme4_r = io_dec_csr_wen_r_mod & _T_2290; // @[dec_tlu_ctl.scala 2439:41]
  wire  _T_2294 = io_dec_csr_wraddr_r == 12'h325; // @[dec_tlu_ctl.scala 2446:70]
  wire  wr_mhpme5_r = io_dec_csr_wen_r_mod & _T_2294; // @[dec_tlu_ctl.scala 2446:41]
  wire  _T_2298 = io_dec_csr_wraddr_r == 12'h326; // @[dec_tlu_ctl.scala 2453:70]
  wire  wr_mhpme6_r = io_dec_csr_wen_r_mod & _T_2298; // @[dec_tlu_ctl.scala 2453:41]
  wire  _T_2302 = io_dec_csr_wraddr_r == 12'h320; // @[dec_tlu_ctl.scala 2470:77]
  wire  wr_mcountinhibit_r = io_dec_csr_wen_r_mod & _T_2302; // @[dec_tlu_ctl.scala 2470:48]
  wire  _T_2314 = io_i0_valid_wb | io_exc_or_int_valid_r_d1; // @[dec_tlu_ctl.scala 2485:51]
  wire  _T_2315 = _T_2314 | io_interrupt_valid_r_d1; // @[dec_tlu_ctl.scala 2485:78]
  wire  _T_2316 = _T_2315 | io_dec_tlu_i0_valid_wb1; // @[dec_tlu_ctl.scala 2485:104]
  wire  _T_2317 = _T_2316 | io_dec_tlu_i0_exc_valid_wb1; // @[dec_tlu_ctl.scala 2485:130]
  wire  _T_2318 = _T_2317 | io_dec_tlu_int_valid_wb1; // @[dec_tlu_ctl.scala 2486:32]
  reg  _T_2321; // @[dec_tlu_ctl.scala 2488:62]
  wire  _T_2322 = io_i0_exception_valid_r_d1 | io_lsu_i0_exc_r_d1; // @[dec_tlu_ctl.scala 2489:91]
  wire  _T_2323 = ~io_trigger_hit_dmode_r_d1; // @[dec_tlu_ctl.scala 2489:137]
  wire  _T_2324 = io_trigger_hit_r_d1 & _T_2323; // @[dec_tlu_ctl.scala 2489:135]
  reg  _T_2326; // @[dec_tlu_ctl.scala 2489:62]
  reg [4:0] _T_2327; // @[dec_tlu_ctl.scala 2490:62]
  reg  _T_2328; // @[dec_tlu_ctl.scala 2491:62]
  wire [31:0] _T_2334 = {io_core_id,4'h0}; // @[Cat.scala 29:58]
  wire [31:0] _T_2343 = {21'h3,3'h0,io_mstatus[1],3'h0,io_mstatus[0],3'h0}; // @[Cat.scala 29:58]
  wire [31:0] _T_2348 = {io_mtvec[30:1],1'h0,io_mtvec[0]}; // @[Cat.scala 29:58]
  wire [31:0] _T_2361 = {1'h0,io_mip[5:3],16'h0,io_mip[2],3'h0,io_mip[1],3'h0,io_mip[0],3'h0}; // @[Cat.scala 29:58]
  wire [31:0] _T_2374 = {1'h0,mie[5:3],16'h0,mie[2],3'h0,mie[1],3'h0,mie[0],3'h0}; // @[Cat.scala 29:58]
  wire [31:0] _T_2386 = {io_mepc,1'h0}; // @[Cat.scala 29:58]
  wire [31:0] _T_2391 = {28'h0,mscause}; // @[Cat.scala 29:58]
  wire [31:0] _T_2399 = {meivt,10'h0}; // @[Cat.scala 29:58]
  wire [31:0] _T_2402 = {meivt,meihap,2'h0}; // @[Cat.scala 29:58]
  wire [31:0] _T_2405 = {28'h0,meicurpl}; // @[Cat.scala 29:58]
  wire [31:0] _T_2408 = {28'h0,meicidpl}; // @[Cat.scala 29:58]
  wire [31:0] _T_2411 = {28'h0,meipt}; // @[Cat.scala 29:58]
  wire [31:0] _T_2414 = {23'h0,mcgc}; // @[Cat.scala 29:58]
  wire [31:0] _T_2417 = {13'h0,_T_345,4'h0,mfdc_int[11:0]}; // @[Cat.scala 29:58]
  wire [31:0] _T_2421 = {16'h4000,io_dcsr[15:2],2'h3}; // @[Cat.scala 29:58]
  wire [31:0] _T_2423 = {io_dpc,1'h0}; // @[Cat.scala 29:58]
  wire [31:0] _T_2439 = {7'h0,dicawics[16],2'h0,dicawics[15:14],3'h0,dicawics[13:0],3'h0}; // @[Cat.scala 29:58]
  wire [31:0] _T_2442 = {30'h0,mtsel}; // @[Cat.scala 29:58]
  wire [31:0] _T_2471 = {26'h0,mfdht}; // @[Cat.scala 29:58]
  wire [31:0] _T_2474 = {30'h0,mfdhs}; // @[Cat.scala 29:58]
  wire [31:0] _T_2477 = {22'h0,mhpme3}; // @[Cat.scala 29:58]
  wire [31:0] _T_2480 = {22'h0,mhpme4}; // @[Cat.scala 29:58]
  wire [31:0] _T_2483 = {22'h0,mhpme5}; // @[Cat.scala 29:58]
  wire [31:0] _T_2486 = {22'h0,mhpme6}; // @[Cat.scala 29:58]
  wire [31:0] _T_2489 = {25'h0,temp_ncount6_2,1'h0,temp_ncount0}; // @[Cat.scala 29:58]
  wire [31:0] _T_2492 = {30'h0,mpmc,1'h0}; // @[Cat.scala 29:58]
  wire [31:0] _T_2495 = io_csr_pkt_csr_misa ? 32'h40001104 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2496 = io_csr_pkt_csr_mvendorid ? 32'h45 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2497 = io_csr_pkt_csr_marchid ? 32'h10 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2498 = io_csr_pkt_csr_mimpid ? 32'h1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2499 = io_csr_pkt_csr_mhartid ? _T_2334 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2500 = io_csr_pkt_csr_mstatus ? _T_2343 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2501 = io_csr_pkt_csr_mtvec ? _T_2348 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2502 = io_csr_pkt_csr_mip ? _T_2361 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2503 = io_csr_pkt_csr_mie ? _T_2374 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2504 = io_csr_pkt_csr_mcyclel ? mcyclel : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2505 = io_csr_pkt_csr_mcycleh ? mcycleh_inc : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2506 = io_csr_pkt_csr_minstretl ? minstretl : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2507 = io_csr_pkt_csr_minstreth ? minstreth_inc : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2508 = io_csr_pkt_csr_mscratch ? mscratch : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2509 = io_csr_pkt_csr_mepc ? _T_2386 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2510 = io_csr_pkt_csr_mcause ? mcause : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2511 = io_csr_pkt_csr_mscause ? _T_2391 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2512 = io_csr_pkt_csr_mtval ? mtval : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2513 = io_csr_pkt_csr_mrac ? mrac : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2514 = io_csr_pkt_csr_mdseac ? mdseac : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2515 = io_csr_pkt_csr_meivt ? _T_2399 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2516 = io_csr_pkt_csr_meihap ? _T_2402 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2517 = io_csr_pkt_csr_meicurpl ? _T_2405 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2518 = io_csr_pkt_csr_meicidpl ? _T_2408 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2519 = io_csr_pkt_csr_meipt ? _T_2411 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2520 = io_csr_pkt_csr_mcgc ? _T_2414 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2521 = io_csr_pkt_csr_mfdc ? _T_2417 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2522 = io_csr_pkt_csr_dcsr ? _T_2421 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2523 = io_csr_pkt_csr_dpc ? _T_2423 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2524 = io_csr_pkt_csr_dicad0 ? dicad0[31:0] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2525 = io_csr_pkt_csr_dicad0h ? dicad0h : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2526 = io_csr_pkt_csr_dicad1 ? dicad1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2527 = io_csr_pkt_csr_dicawics ? _T_2439 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2528 = io_csr_pkt_csr_mtsel ? _T_2442 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2529 = io_csr_pkt_csr_mtdata1 ? mtdata1_tsel_out : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2530 = io_csr_pkt_csr_mtdata2 ? mtdata2_tsel_out : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2531 = io_csr_pkt_csr_micect ? micect : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2532 = io_csr_pkt_csr_miccmect ? miccmect : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2533 = io_csr_pkt_csr_mdccmect ? mdccmect : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2534 = io_csr_pkt_csr_mhpmc3 ? mhpmc3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2535 = io_csr_pkt_csr_mhpmc4 ? mhpmc4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2536 = io_csr_pkt_csr_mhpmc5 ? mhpmc5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2537 = io_csr_pkt_csr_mhpmc6 ? mhpmc6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2538 = io_csr_pkt_csr_mhpmc3h ? mhpmc3h : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2539 = io_csr_pkt_csr_mhpmc4h ? mhpmc4h : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2540 = io_csr_pkt_csr_mhpmc5h ? mhpmc5h : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2541 = io_csr_pkt_csr_mhpmc6h ? mhpmc6h : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2542 = io_csr_pkt_csr_mfdht ? _T_2471 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2543 = io_csr_pkt_csr_mfdhs ? _T_2474 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2544 = io_csr_pkt_csr_mhpme3 ? _T_2477 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2545 = io_csr_pkt_csr_mhpme4 ? _T_2480 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2546 = io_csr_pkt_csr_mhpme5 ? _T_2483 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2547 = io_csr_pkt_csr_mhpme6 ? _T_2486 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2548 = io_csr_pkt_csr_mcountinhibit ? _T_2489 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2549 = io_csr_pkt_csr_mpmc ? _T_2492 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2550 = io_dec_timer_read_d ? io_dec_timer_rddata_d : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2551 = _T_2495 | _T_2496; // @[Mux.scala 27:72]
  wire [31:0] _T_2552 = _T_2551 | _T_2497; // @[Mux.scala 27:72]
  wire [31:0] _T_2553 = _T_2552 | _T_2498; // @[Mux.scala 27:72]
  wire [31:0] _T_2554 = _T_2553 | _T_2499; // @[Mux.scala 27:72]
  wire [31:0] _T_2555 = _T_2554 | _T_2500; // @[Mux.scala 27:72]
  wire [31:0] _T_2556 = _T_2555 | _T_2501; // @[Mux.scala 27:72]
  wire [31:0] _T_2557 = _T_2556 | _T_2502; // @[Mux.scala 27:72]
  wire [31:0] _T_2558 = _T_2557 | _T_2503; // @[Mux.scala 27:72]
  wire [31:0] _T_2559 = _T_2558 | _T_2504; // @[Mux.scala 27:72]
  wire [31:0] _T_2560 = _T_2559 | _T_2505; // @[Mux.scala 27:72]
  wire [31:0] _T_2561 = _T_2560 | _T_2506; // @[Mux.scala 27:72]
  wire [31:0] _T_2562 = _T_2561 | _T_2507; // @[Mux.scala 27:72]
  wire [31:0] _T_2563 = _T_2562 | _T_2508; // @[Mux.scala 27:72]
  wire [31:0] _T_2564 = _T_2563 | _T_2509; // @[Mux.scala 27:72]
  wire [31:0] _T_2565 = _T_2564 | _T_2510; // @[Mux.scala 27:72]
  wire [31:0] _T_2566 = _T_2565 | _T_2511; // @[Mux.scala 27:72]
  wire [31:0] _T_2567 = _T_2566 | _T_2512; // @[Mux.scala 27:72]
  wire [31:0] _T_2568 = _T_2567 | _T_2513; // @[Mux.scala 27:72]
  wire [31:0] _T_2569 = _T_2568 | _T_2514; // @[Mux.scala 27:72]
  wire [31:0] _T_2570 = _T_2569 | _T_2515; // @[Mux.scala 27:72]
  wire [31:0] _T_2571 = _T_2570 | _T_2516; // @[Mux.scala 27:72]
  wire [31:0] _T_2572 = _T_2571 | _T_2517; // @[Mux.scala 27:72]
  wire [31:0] _T_2573 = _T_2572 | _T_2518; // @[Mux.scala 27:72]
  wire [31:0] _T_2574 = _T_2573 | _T_2519; // @[Mux.scala 27:72]
  wire [31:0] _T_2575 = _T_2574 | _T_2520; // @[Mux.scala 27:72]
  wire [31:0] _T_2576 = _T_2575 | _T_2521; // @[Mux.scala 27:72]
  wire [31:0] _T_2577 = _T_2576 | _T_2522; // @[Mux.scala 27:72]
  wire [31:0] _T_2578 = _T_2577 | _T_2523; // @[Mux.scala 27:72]
  wire [31:0] _T_2579 = _T_2578 | _T_2524; // @[Mux.scala 27:72]
  wire [31:0] _T_2580 = _T_2579 | _T_2525; // @[Mux.scala 27:72]
  wire [31:0] _T_2581 = _T_2580 | _T_2526; // @[Mux.scala 27:72]
  wire [31:0] _T_2582 = _T_2581 | _T_2527; // @[Mux.scala 27:72]
  wire [31:0] _T_2583 = _T_2582 | _T_2528; // @[Mux.scala 27:72]
  wire [31:0] _T_2584 = _T_2583 | _T_2529; // @[Mux.scala 27:72]
  wire [31:0] _T_2585 = _T_2584 | _T_2530; // @[Mux.scala 27:72]
  wire [31:0] _T_2586 = _T_2585 | _T_2531; // @[Mux.scala 27:72]
  wire [31:0] _T_2587 = _T_2586 | _T_2532; // @[Mux.scala 27:72]
  wire [31:0] _T_2588 = _T_2587 | _T_2533; // @[Mux.scala 27:72]
  wire [31:0] _T_2589 = _T_2588 | _T_2534; // @[Mux.scala 27:72]
  wire [31:0] _T_2590 = _T_2589 | _T_2535; // @[Mux.scala 27:72]
  wire [31:0] _T_2591 = _T_2590 | _T_2536; // @[Mux.scala 27:72]
  wire [31:0] _T_2592 = _T_2591 | _T_2537; // @[Mux.scala 27:72]
  wire [31:0] _T_2593 = _T_2592 | _T_2538; // @[Mux.scala 27:72]
  wire [31:0] _T_2594 = _T_2593 | _T_2539; // @[Mux.scala 27:72]
  wire [31:0] _T_2595 = _T_2594 | _T_2540; // @[Mux.scala 27:72]
  wire [31:0] _T_2596 = _T_2595 | _T_2541; // @[Mux.scala 27:72]
  wire [31:0] _T_2597 = _T_2596 | _T_2542; // @[Mux.scala 27:72]
  wire [31:0] _T_2598 = _T_2597 | _T_2543; // @[Mux.scala 27:72]
  wire [31:0] _T_2599 = _T_2598 | _T_2544; // @[Mux.scala 27:72]
  wire [31:0] _T_2600 = _T_2599 | _T_2545; // @[Mux.scala 27:72]
  wire [31:0] _T_2601 = _T_2600 | _T_2546; // @[Mux.scala 27:72]
  wire [31:0] _T_2602 = _T_2601 | _T_2547; // @[Mux.scala 27:72]
  wire [31:0] _T_2603 = _T_2602 | _T_2548; // @[Mux.scala 27:72]
  wire [31:0] _T_2604 = _T_2603 | _T_2549; // @[Mux.scala 27:72]
  rvclkhdr rvclkhdr ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_io_l1clk),
    .io_clk(rvclkhdr_io_clk),
    .io_en(rvclkhdr_io_en),
    .io_scan_mode(rvclkhdr_io_scan_mode)
  );
  rvclkhdr rvclkhdr_1 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_1_io_l1clk),
    .io_clk(rvclkhdr_1_io_clk),
    .io_en(rvclkhdr_1_io_en),
    .io_scan_mode(rvclkhdr_1_io_scan_mode)
  );
  rvclkhdr rvclkhdr_2 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_2_io_l1clk),
    .io_clk(rvclkhdr_2_io_clk),
    .io_en(rvclkhdr_2_io_en),
    .io_scan_mode(rvclkhdr_2_io_scan_mode)
  );
  rvclkhdr rvclkhdr_3 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_3_io_l1clk),
    .io_clk(rvclkhdr_3_io_clk),
    .io_en(rvclkhdr_3_io_en),
    .io_scan_mode(rvclkhdr_3_io_scan_mode)
  );
  rvclkhdr rvclkhdr_4 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_4_io_l1clk),
    .io_clk(rvclkhdr_4_io_clk),
    .io_en(rvclkhdr_4_io_en),
    .io_scan_mode(rvclkhdr_4_io_scan_mode)
  );
  rvclkhdr rvclkhdr_5 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_5_io_l1clk),
    .io_clk(rvclkhdr_5_io_clk),
    .io_en(rvclkhdr_5_io_en),
    .io_scan_mode(rvclkhdr_5_io_scan_mode)
  );
  rvclkhdr rvclkhdr_6 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_6_io_l1clk),
    .io_clk(rvclkhdr_6_io_clk),
    .io_en(rvclkhdr_6_io_en),
    .io_scan_mode(rvclkhdr_6_io_scan_mode)
  );
  rvclkhdr rvclkhdr_7 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_7_io_l1clk),
    .io_clk(rvclkhdr_7_io_clk),
    .io_en(rvclkhdr_7_io_en),
    .io_scan_mode(rvclkhdr_7_io_scan_mode)
  );
  rvclkhdr rvclkhdr_8 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_8_io_l1clk),
    .io_clk(rvclkhdr_8_io_clk),
    .io_en(rvclkhdr_8_io_en),
    .io_scan_mode(rvclkhdr_8_io_scan_mode)
  );
  rvclkhdr rvclkhdr_9 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_9_io_l1clk),
    .io_clk(rvclkhdr_9_io_clk),
    .io_en(rvclkhdr_9_io_en),
    .io_scan_mode(rvclkhdr_9_io_scan_mode)
  );
  rvclkhdr rvclkhdr_10 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_10_io_l1clk),
    .io_clk(rvclkhdr_10_io_clk),
    .io_en(rvclkhdr_10_io_en),
    .io_scan_mode(rvclkhdr_10_io_scan_mode)
  );
  rvclkhdr rvclkhdr_11 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_11_io_l1clk),
    .io_clk(rvclkhdr_11_io_clk),
    .io_en(rvclkhdr_11_io_en),
    .io_scan_mode(rvclkhdr_11_io_scan_mode)
  );
  rvclkhdr rvclkhdr_12 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_12_io_l1clk),
    .io_clk(rvclkhdr_12_io_clk),
    .io_en(rvclkhdr_12_io_en),
    .io_scan_mode(rvclkhdr_12_io_scan_mode)
  );
  rvclkhdr rvclkhdr_13 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_13_io_l1clk),
    .io_clk(rvclkhdr_13_io_clk),
    .io_en(rvclkhdr_13_io_en),
    .io_scan_mode(rvclkhdr_13_io_scan_mode)
  );
  rvclkhdr rvclkhdr_14 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_14_io_l1clk),
    .io_clk(rvclkhdr_14_io_clk),
    .io_en(rvclkhdr_14_io_en),
    .io_scan_mode(rvclkhdr_14_io_scan_mode)
  );
  rvclkhdr rvclkhdr_15 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_15_io_l1clk),
    .io_clk(rvclkhdr_15_io_clk),
    .io_en(rvclkhdr_15_io_en),
    .io_scan_mode(rvclkhdr_15_io_scan_mode)
  );
  rvclkhdr rvclkhdr_16 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_16_io_l1clk),
    .io_clk(rvclkhdr_16_io_clk),
    .io_en(rvclkhdr_16_io_en),
    .io_scan_mode(rvclkhdr_16_io_scan_mode)
  );
  rvclkhdr rvclkhdr_17 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_17_io_l1clk),
    .io_clk(rvclkhdr_17_io_clk),
    .io_en(rvclkhdr_17_io_en),
    .io_scan_mode(rvclkhdr_17_io_scan_mode)
  );
  rvclkhdr rvclkhdr_18 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_18_io_l1clk),
    .io_clk(rvclkhdr_18_io_clk),
    .io_en(rvclkhdr_18_io_en),
    .io_scan_mode(rvclkhdr_18_io_scan_mode)
  );
  rvclkhdr rvclkhdr_19 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_19_io_l1clk),
    .io_clk(rvclkhdr_19_io_clk),
    .io_en(rvclkhdr_19_io_en),
    .io_scan_mode(rvclkhdr_19_io_scan_mode)
  );
  rvclkhdr rvclkhdr_20 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_20_io_l1clk),
    .io_clk(rvclkhdr_20_io_clk),
    .io_en(rvclkhdr_20_io_en),
    .io_scan_mode(rvclkhdr_20_io_scan_mode)
  );
  rvclkhdr rvclkhdr_21 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_21_io_l1clk),
    .io_clk(rvclkhdr_21_io_clk),
    .io_en(rvclkhdr_21_io_en),
    .io_scan_mode(rvclkhdr_21_io_scan_mode)
  );
  rvclkhdr rvclkhdr_22 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_22_io_l1clk),
    .io_clk(rvclkhdr_22_io_clk),
    .io_en(rvclkhdr_22_io_en),
    .io_scan_mode(rvclkhdr_22_io_scan_mode)
  );
  rvclkhdr rvclkhdr_23 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_23_io_l1clk),
    .io_clk(rvclkhdr_23_io_clk),
    .io_en(rvclkhdr_23_io_en),
    .io_scan_mode(rvclkhdr_23_io_scan_mode)
  );
  rvclkhdr rvclkhdr_24 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_24_io_l1clk),
    .io_clk(rvclkhdr_24_io_clk),
    .io_en(rvclkhdr_24_io_en),
    .io_scan_mode(rvclkhdr_24_io_scan_mode)
  );
  rvclkhdr rvclkhdr_25 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_25_io_l1clk),
    .io_clk(rvclkhdr_25_io_clk),
    .io_en(rvclkhdr_25_io_en),
    .io_scan_mode(rvclkhdr_25_io_scan_mode)
  );
  rvclkhdr rvclkhdr_26 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_26_io_l1clk),
    .io_clk(rvclkhdr_26_io_clk),
    .io_en(rvclkhdr_26_io_en),
    .io_scan_mode(rvclkhdr_26_io_scan_mode)
  );
  rvclkhdr rvclkhdr_27 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_27_io_l1clk),
    .io_clk(rvclkhdr_27_io_clk),
    .io_en(rvclkhdr_27_io_en),
    .io_scan_mode(rvclkhdr_27_io_scan_mode)
  );
  rvclkhdr rvclkhdr_28 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_28_io_l1clk),
    .io_clk(rvclkhdr_28_io_clk),
    .io_en(rvclkhdr_28_io_en),
    .io_scan_mode(rvclkhdr_28_io_scan_mode)
  );
  rvclkhdr rvclkhdr_29 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_29_io_l1clk),
    .io_clk(rvclkhdr_29_io_clk),
    .io_en(rvclkhdr_29_io_en),
    .io_scan_mode(rvclkhdr_29_io_scan_mode)
  );
  rvclkhdr rvclkhdr_30 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_30_io_l1clk),
    .io_clk(rvclkhdr_30_io_clk),
    .io_en(rvclkhdr_30_io_en),
    .io_scan_mode(rvclkhdr_30_io_scan_mode)
  );
  rvclkhdr rvclkhdr_31 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_31_io_l1clk),
    .io_clk(rvclkhdr_31_io_clk),
    .io_en(rvclkhdr_31_io_en),
    .io_scan_mode(rvclkhdr_31_io_scan_mode)
  );
  rvclkhdr rvclkhdr_32 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_32_io_l1clk),
    .io_clk(rvclkhdr_32_io_clk),
    .io_en(rvclkhdr_32_io_en),
    .io_scan_mode(rvclkhdr_32_io_scan_mode)
  );
  rvclkhdr rvclkhdr_33 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_33_io_l1clk),
    .io_clk(rvclkhdr_33_io_clk),
    .io_en(rvclkhdr_33_io_en),
    .io_scan_mode(rvclkhdr_33_io_scan_mode)
  );
  rvclkhdr rvclkhdr_34 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_34_io_l1clk),
    .io_clk(rvclkhdr_34_io_clk),
    .io_en(rvclkhdr_34_io_en),
    .io_scan_mode(rvclkhdr_34_io_scan_mode)
  );
  assign io_dec_tlu_ic_diag_pkt_icache_wrdata = {_T_754,dicad0[31:0]}; // @[dec_tlu_ctl.scala 2155:56]
  assign io_dec_tlu_ic_diag_pkt_icache_dicawics = dicawics; // @[dec_tlu_ctl.scala 2158:41]
  assign io_dec_tlu_ic_diag_pkt_icache_rd_valid = icache_rd_valid_f; // @[dec_tlu_ctl.scala 2166:41]
  assign io_dec_tlu_ic_diag_pkt_icache_wr_valid = icache_wr_valid_f; // @[dec_tlu_ctl.scala 2167:41]
  assign io_trigger_pkt_any_0_select = io_mtdata1_t_0[7]; // @[dec_tlu_ctl.scala 2231:40]
  assign io_trigger_pkt_any_0_match_pkt = io_mtdata1_t_0[4]; // @[dec_tlu_ctl.scala 2232:43]
  assign io_trigger_pkt_any_0_store = io_mtdata1_t_0[1]; // @[dec_tlu_ctl.scala 2233:40]
  assign io_trigger_pkt_any_0_load = io_mtdata1_t_0[0]; // @[dec_tlu_ctl.scala 2234:40]
  assign io_trigger_pkt_any_0_execute = io_mtdata1_t_0[2]; // @[dec_tlu_ctl.scala 2235:40]
  assign io_trigger_pkt_any_0_m = io_mtdata1_t_0[3]; // @[dec_tlu_ctl.scala 2236:40]
  assign io_trigger_pkt_any_0_tdata2 = mtdata2_t_0; // @[dec_tlu_ctl.scala 2249:51]
  assign io_trigger_pkt_any_1_select = io_mtdata1_t_1[7]; // @[dec_tlu_ctl.scala 2231:40]
  assign io_trigger_pkt_any_1_match_pkt = io_mtdata1_t_1[4]; // @[dec_tlu_ctl.scala 2232:43]
  assign io_trigger_pkt_any_1_store = io_mtdata1_t_1[1]; // @[dec_tlu_ctl.scala 2233:40]
  assign io_trigger_pkt_any_1_load = io_mtdata1_t_1[0]; // @[dec_tlu_ctl.scala 2234:40]
  assign io_trigger_pkt_any_1_execute = io_mtdata1_t_1[2]; // @[dec_tlu_ctl.scala 2235:40]
  assign io_trigger_pkt_any_1_m = io_mtdata1_t_1[3]; // @[dec_tlu_ctl.scala 2236:40]
  assign io_trigger_pkt_any_1_tdata2 = mtdata2_t_1; // @[dec_tlu_ctl.scala 2249:51]
  assign io_trigger_pkt_any_2_select = io_mtdata1_t_2[7]; // @[dec_tlu_ctl.scala 2231:40]
  assign io_trigger_pkt_any_2_match_pkt = io_mtdata1_t_2[4]; // @[dec_tlu_ctl.scala 2232:43]
  assign io_trigger_pkt_any_2_store = io_mtdata1_t_2[1]; // @[dec_tlu_ctl.scala 2233:40]
  assign io_trigger_pkt_any_2_load = io_mtdata1_t_2[0]; // @[dec_tlu_ctl.scala 2234:40]
  assign io_trigger_pkt_any_2_execute = io_mtdata1_t_2[2]; // @[dec_tlu_ctl.scala 2235:40]
  assign io_trigger_pkt_any_2_m = io_mtdata1_t_2[3]; // @[dec_tlu_ctl.scala 2236:40]
  assign io_trigger_pkt_any_2_tdata2 = mtdata2_t_2; // @[dec_tlu_ctl.scala 2249:51]
  assign io_trigger_pkt_any_3_select = io_mtdata1_t_3[7]; // @[dec_tlu_ctl.scala 2231:40]
  assign io_trigger_pkt_any_3_match_pkt = io_mtdata1_t_3[4]; // @[dec_tlu_ctl.scala 2232:43]
  assign io_trigger_pkt_any_3_store = io_mtdata1_t_3[1]; // @[dec_tlu_ctl.scala 2233:40]
  assign io_trigger_pkt_any_3_load = io_mtdata1_t_3[0]; // @[dec_tlu_ctl.scala 2234:40]
  assign io_trigger_pkt_any_3_execute = io_mtdata1_t_3[2]; // @[dec_tlu_ctl.scala 2235:40]
  assign io_trigger_pkt_any_3_m = io_mtdata1_t_3[3]; // @[dec_tlu_ctl.scala 2236:40]
  assign io_trigger_pkt_any_3_tdata2 = mtdata2_t_3; // @[dec_tlu_ctl.scala 2249:51]
  assign io_dec_tlu_int_valid_wb1 = _T_2328; // @[dec_tlu_ctl.scala 2491:30]
  assign io_dec_tlu_i0_exc_valid_wb1 = _T_2326; // @[dec_tlu_ctl.scala 2489:30]
  assign io_dec_tlu_i0_valid_wb1 = _T_2321; // @[dec_tlu_ctl.scala 2488:30]
  assign io_dec_tlu_mtval_wb1 = mtval; // @[dec_tlu_ctl.scala 2493:24]
  assign io_dec_tlu_exc_cause_wb1 = _T_2327; // @[dec_tlu_ctl.scala 2490:30]
  assign io_dec_tlu_perfcnt0 = mhpmc_inc_r_d1_0 & _T_2173; // @[dec_tlu_ctl.scala 2345:22]
  assign io_dec_tlu_perfcnt1 = mhpmc_inc_r_d1_1 & _T_2178; // @[dec_tlu_ctl.scala 2346:22]
  assign io_dec_tlu_perfcnt2 = mhpmc_inc_r_d1_2 & _T_2183; // @[dec_tlu_ctl.scala 2347:22]
  assign io_dec_tlu_perfcnt3 = mhpmc_inc_r_d1_3 & _T_2188; // @[dec_tlu_ctl.scala 2348:22]
  assign io_dec_tlu_misc_clk_override = mcgc[8]; // @[dec_tlu_ctl.scala 1718:31]
  assign io_dec_tlu_dec_clk_override = mcgc[7]; // @[dec_tlu_ctl.scala 1719:31]
  assign io_dec_tlu_lsu_clk_override = mcgc[4]; // @[dec_tlu_ctl.scala 1721:31]
  assign io_dec_tlu_bus_clk_override = mcgc[3]; // @[dec_tlu_ctl.scala 1722:31]
  assign io_dec_tlu_pic_clk_override = mcgc[2]; // @[dec_tlu_ctl.scala 1723:31]
  assign io_dec_tlu_dccm_clk_override = mcgc[1]; // @[dec_tlu_ctl.scala 1724:31]
  assign io_dec_tlu_icm_clk_override = mcgc[0]; // @[dec_tlu_ctl.scala 1725:31]
  assign io_dec_csr_rddata_d = _T_2604 | _T_2550; // @[dec_tlu_ctl.scala 2498:21]
  assign io_dec_tlu_pipelining_disable = mfdc[0]; // @[dec_tlu_ctl.scala 1768:39]
  assign io_dec_tlu_wr_pause_r = _T_360 & _T_361; // @[dec_tlu_ctl.scala 1777:24]
  assign io_dec_tlu_meipt = meipt; // @[dec_tlu_ctl.scala 2006:19]
  assign io_dec_tlu_meicurpl = meicurpl; // @[dec_tlu_ctl.scala 1970:22]
  assign io_dec_tlu_meihap = {meivt,meihap}; // @[dec_tlu_ctl.scala 1956:20]
  assign io_dec_tlu_mrac_ff = mrac; // @[dec_tlu_ctl.scala 1807:21]
  assign io_dec_tlu_wb_coalescing_disable = mfdc[2]; // @[dec_tlu_ctl.scala 1767:39]
  assign io_dec_tlu_bpred_disable = mfdc[3]; // @[dec_tlu_ctl.scala 1766:39]
  assign io_dec_tlu_sideeffect_posted_disable = mfdc[6]; // @[dec_tlu_ctl.scala 1765:39]
  assign io_dec_tlu_core_ecc_disable = mfdc[8]; // @[dec_tlu_ctl.scala 1764:39]
  assign io_dec_tlu_external_ldfwd_disable = mfdc[11]; // @[dec_tlu_ctl.scala 1763:39]
  assign io_dec_tlu_dma_qos_prty = mfdc[18:16]; // @[dec_tlu_ctl.scala 1762:39]
  assign io_dec_csr_wen_r_mod = _T_1 & _T_2; // @[dec_tlu_ctl.scala 1451:23]
  assign io_fw_halt_req = _T_492 & _T_493; // @[dec_tlu_ctl.scala 1842:17]
  assign io_mstatus = _T_56; // @[dec_tlu_ctl.scala 1467:13]
  assign io_mstatus_mie_ns = io_mstatus[0] & _T_54; // @[dec_tlu_ctl.scala 1466:20]
  assign io_dcsr = _T_691; // @[dec_tlu_ctl.scala 2053:10]
  assign io_mtvec = _T_62; // @[dec_tlu_ctl.scala 1479:11]
  assign io_mip = _T_68; // @[dec_tlu_ctl.scala 1494:9]
  assign io_mie_ns = wr_mie_r ? _T_78 : mie; // @[dec_tlu_ctl.scala 1508:12]
  assign io_npc_r = _T_161 | _T_159; // @[dec_tlu_ctl.scala 1602:11]
  assign io_npc_r_d1 = _T_167; // @[dec_tlu_ctl.scala 1608:14]
  assign io_mepc = _T_196; // @[dec_tlu_ctl.scala 1627:10]
  assign io_mdseac_locked_ns = mdseac_en | _T_479; // @[dec_tlu_ctl.scala 1825:22]
  assign io_force_halt = mfdht[0] & _T_599; // @[dec_tlu_ctl.scala 1933:16]
  assign io_dpc = _T_716; // @[dec_tlu_ctl.scala 2070:9]
  assign io_mtdata1_t_0 = _T_863; // @[dec_tlu_ctl.scala 2226:39]
  assign io_mtdata1_t_1 = _T_864; // @[dec_tlu_ctl.scala 2226:39]
  assign io_mtdata1_t_2 = _T_865; // @[dec_tlu_ctl.scala 2226:39]
  assign io_mtdata1_t_3 = _T_866; // @[dec_tlu_ctl.scala 2226:39]
  assign rvclkhdr_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_io_en = io_dec_csr_wen_r_mod & _T_58; // @[lib.scala 371:17]
  assign rvclkhdr_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_1_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_1_io_en = wr_mcyclel_r | mcyclel_cout_in; // @[lib.scala 371:17]
  assign rvclkhdr_1_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_2_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_2_io_en = wr_mcycleh_r | mcyclel_cout_f; // @[lib.scala 371:17]
  assign rvclkhdr_2_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_3_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_3_io_en = i0_valid_no_ebreak_ecall_r | wr_minstretl_r; // @[lib.scala 371:17]
  assign rvclkhdr_3_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_4_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_4_io_en = minstret_enable_f | wr_minstreth_r; // @[lib.scala 371:17]
  assign rvclkhdr_4_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_5_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_5_io_en = io_dec_csr_wen_r_mod & _T_139; // @[lib.scala 371:17]
  assign rvclkhdr_5_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_6_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_6_io_en = _T_164 | io_reset_delayed; // @[lib.scala 371:17]
  assign rvclkhdr_6_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_7_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_7_io_en = _T_142 & io_dec_tlu_i0_valid_r; // @[lib.scala 371:17]
  assign rvclkhdr_7_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_8_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_8_io_en = io_dec_csr_wen_r_mod & _T_325; // @[lib.scala 371:17]
  assign rvclkhdr_8_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_9_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_9_io_en = io_dec_csr_wen_r_mod & _T_337; // @[lib.scala 371:17]
  assign rvclkhdr_9_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_10_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_10_io_en = io_dec_csr_wen_r_mod & _T_364; // @[lib.scala 371:17]
  assign rvclkhdr_10_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_11_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_11_io_en = _T_483 & _T_484; // @[lib.scala 371:17]
  assign rvclkhdr_11_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_12_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_12_io_en = wr_micect_r | io_ic_perr_r_d1; // @[lib.scala 371:17]
  assign rvclkhdr_12_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_13_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_13_io_en = _T_539 | io_iccm_dma_sb_error; // @[lib.scala 371:17]
  assign rvclkhdr_13_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_14_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_14_io_en = wr_mdccmect_r | io_lsu_single_ecc_error_r_d1; // @[lib.scala 371:17]
  assign rvclkhdr_14_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_15_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_15_io_en = io_dec_csr_wen_r_mod & _T_602; // @[lib.scala 371:17]
  assign rvclkhdr_15_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_16_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_16_io_en = _T_622 | io_take_ext_int_start; // @[lib.scala 371:17]
  assign rvclkhdr_16_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_17_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_17_io_en = _T_688 | io_take_nmi; // @[lib.scala 371:17]
  assign rvclkhdr_17_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_18_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_18_io_en = _T_713 | dpc_capture_npc; // @[lib.scala 371:17]
  assign rvclkhdr_18_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_19_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_19_io_en = _T_653 & _T_723; // @[lib.scala 371:17]
  assign rvclkhdr_19_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_20_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_20_io_en = wr_dicad0_r | io_ifu_ic_debug_rd_data_valid; // @[lib.scala 371:17]
  assign rvclkhdr_20_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_21_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_21_io_en = wr_dicad0h_r | io_ifu_ic_debug_rd_data_valid; // @[lib.scala 371:17]
  assign rvclkhdr_21_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_22_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_22_io_en = _T_962 & _T_798; // @[lib.scala 371:17]
  assign rvclkhdr_22_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_23_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_23_io_en = _T_971 & _T_807; // @[lib.scala 371:17]
  assign rvclkhdr_23_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_24_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_24_io_en = _T_980 & _T_816; // @[lib.scala 371:17]
  assign rvclkhdr_24_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_25_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_25_io_en = _T_989 & _T_825; // @[lib.scala 371:17]
  assign rvclkhdr_25_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_26_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_26_io_en = mhpmc3_wr_en0 | mhpmc3_wr_en1; // @[lib.scala 371:17]
  assign rvclkhdr_26_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_27_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_27_io_en = mhpmc3h_wr_en0 | mhpmc3_wr_en1; // @[lib.scala 371:17]
  assign rvclkhdr_27_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_28_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_28_io_en = mhpmc4_wr_en0 | mhpmc4_wr_en1; // @[lib.scala 371:17]
  assign rvclkhdr_28_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_29_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_29_io_en = mhpmc4h_wr_en0 | mhpmc4_wr_en1; // @[lib.scala 371:17]
  assign rvclkhdr_29_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_30_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_30_io_en = mhpmc5_wr_en0 | mhpmc5_wr_en1; // @[lib.scala 371:17]
  assign rvclkhdr_30_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_31_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_31_io_en = mhpmc5h_wr_en0 | mhpmc5_wr_en1; // @[lib.scala 371:17]
  assign rvclkhdr_31_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_32_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_32_io_en = mhpmc6_wr_en0 | mhpmc6_wr_en1; // @[lib.scala 371:17]
  assign rvclkhdr_32_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_33_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_33_io_en = mhpmc6h_wr_en0 | mhpmc6_wr_en1; // @[lib.scala 371:17]
  assign rvclkhdr_33_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_34_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_34_io_en = _T_2318 | io_clk_override; // @[lib.scala 345:16]
  assign rvclkhdr_34_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  mpmc_b = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  _T_56 = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  _T_62 = _RAND_2[30:0];
  _RAND_3 = {1{`RANDOM}};
  mdccmect = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  miccmect = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  micect = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  _T_68 = _RAND_6[5:0];
  _RAND_7 = {1{`RANDOM}};
  mie = _RAND_7[5:0];
  _RAND_8 = {1{`RANDOM}};
  temp_ncount6_2 = _RAND_8[4:0];
  _RAND_9 = {1{`RANDOM}};
  temp_ncount0 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  mcyclel = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  mcyclel_cout_f = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  mcycleh = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  minstretl = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  minstret_enable_f = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  minstretl_cout_f = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  minstreth = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  mscratch = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  _T_167 = _RAND_18[30:0];
  _RAND_19 = {1{`RANDOM}};
  pc_r_d1 = _RAND_19[30:0];
  _RAND_20 = {1{`RANDOM}};
  _T_196 = _RAND_20[30:0];
  _RAND_21 = {1{`RANDOM}};
  mcause = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  mscause = _RAND_22[3:0];
  _RAND_23 = {1{`RANDOM}};
  mtval = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  mcgc = _RAND_24[8:0];
  _RAND_25 = {1{`RANDOM}};
  mfdc_int = _RAND_25[14:0];
  _RAND_26 = {1{`RANDOM}};
  mrac = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  mdseac = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  mfdht = _RAND_28[5:0];
  _RAND_29 = {1{`RANDOM}};
  mfdhs = _RAND_29[1:0];
  _RAND_30 = {1{`RANDOM}};
  force_halt_ctr_f = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  meivt = _RAND_31[21:0];
  _RAND_32 = {1{`RANDOM}};
  meihap = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  meicurpl = _RAND_33[3:0];
  _RAND_34 = {1{`RANDOM}};
  meicidpl = _RAND_34[3:0];
  _RAND_35 = {1{`RANDOM}};
  meipt = _RAND_35[3:0];
  _RAND_36 = {1{`RANDOM}};
  _T_691 = _RAND_36[15:0];
  _RAND_37 = {1{`RANDOM}};
  _T_716 = _RAND_37[30:0];
  _RAND_38 = {1{`RANDOM}};
  dicawics = _RAND_38[16:0];
  _RAND_39 = {3{`RANDOM}};
  dicad0 = _RAND_39[70:0];
  _RAND_40 = {1{`RANDOM}};
  dicad0h = _RAND_40[31:0];
  _RAND_41 = {1{`RANDOM}};
  _T_749 = _RAND_41[6:0];
  _RAND_42 = {1{`RANDOM}};
  icache_rd_valid_f = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  icache_wr_valid_f = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  mtsel = _RAND_44[1:0];
  _RAND_45 = {1{`RANDOM}};
  _T_863 = _RAND_45[9:0];
  _RAND_46 = {1{`RANDOM}};
  _T_864 = _RAND_46[9:0];
  _RAND_47 = {1{`RANDOM}};
  _T_865 = _RAND_47[9:0];
  _RAND_48 = {1{`RANDOM}};
  _T_866 = _RAND_48[9:0];
  _RAND_49 = {1{`RANDOM}};
  mtdata2_t_0 = _RAND_49[31:0];
  _RAND_50 = {1{`RANDOM}};
  mtdata2_t_1 = _RAND_50[31:0];
  _RAND_51 = {1{`RANDOM}};
  mtdata2_t_2 = _RAND_51[31:0];
  _RAND_52 = {1{`RANDOM}};
  mtdata2_t_3 = _RAND_52[31:0];
  _RAND_53 = {1{`RANDOM}};
  mhpme3 = _RAND_53[9:0];
  _RAND_54 = {1{`RANDOM}};
  mhpme4 = _RAND_54[9:0];
  _RAND_55 = {1{`RANDOM}};
  mhpme5 = _RAND_55[9:0];
  _RAND_56 = {1{`RANDOM}};
  mhpme6 = _RAND_56[9:0];
  _RAND_57 = {1{`RANDOM}};
  mhpmc_inc_r_d1_0 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  mhpmc_inc_r_d1_1 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  mhpmc_inc_r_d1_2 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  mhpmc_inc_r_d1_3 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  perfcnt_halted_d1 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  mhpmc3h = _RAND_62[31:0];
  _RAND_63 = {1{`RANDOM}};
  mhpmc3 = _RAND_63[31:0];
  _RAND_64 = {1{`RANDOM}};
  mhpmc4h = _RAND_64[31:0];
  _RAND_65 = {1{`RANDOM}};
  mhpmc4 = _RAND_65[31:0];
  _RAND_66 = {1{`RANDOM}};
  mhpmc5h = _RAND_66[31:0];
  _RAND_67 = {1{`RANDOM}};
  mhpmc5 = _RAND_67[31:0];
  _RAND_68 = {1{`RANDOM}};
  mhpmc6h = _RAND_68[31:0];
  _RAND_69 = {1{`RANDOM}};
  mhpmc6 = _RAND_69[31:0];
  _RAND_70 = {1{`RANDOM}};
  _T_2321 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  _T_2326 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  _T_2327 = _RAND_72[4:0];
  _RAND_73 = {1{`RANDOM}};
  _T_2328 = _RAND_73[0:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    mpmc_b = 1'h0;
  end
  if (reset) begin
    _T_56 = 2'h0;
  end
  if (reset) begin
    _T_62 = 31'h0;
  end
  if (reset) begin
    mdccmect = 32'h0;
  end
  if (reset) begin
    miccmect = 32'h0;
  end
  if (reset) begin
    micect = 32'h0;
  end
  if (reset) begin
    _T_68 = 6'h0;
  end
  if (reset) begin
    mie = 6'h0;
  end
  if (reset) begin
    temp_ncount6_2 = 5'h0;
  end
  if (reset) begin
    temp_ncount0 = 1'h0;
  end
  if (reset) begin
    mcyclel = 32'h0;
  end
  if (reset) begin
    mcyclel_cout_f = 1'h0;
  end
  if (reset) begin
    mcycleh = 32'h0;
  end
  if (reset) begin
    minstretl = 32'h0;
  end
  if (reset) begin
    minstret_enable_f = 1'h0;
  end
  if (reset) begin
    minstretl_cout_f = 1'h0;
  end
  if (reset) begin
    minstreth = 32'h0;
  end
  if (reset) begin
    mscratch = 32'h0;
  end
  if (reset) begin
    _T_167 = 31'h0;
  end
  if (reset) begin
    pc_r_d1 = 31'h0;
  end
  if (reset) begin
    _T_196 = 31'h0;
  end
  if (reset) begin
    mcause = 32'h0;
  end
  if (reset) begin
    mscause = 4'h0;
  end
  if (reset) begin
    mtval = 32'h0;
  end
  if (reset) begin
    mcgc = 9'h0;
  end
  if (reset) begin
    mfdc_int = 15'h0;
  end
  if (reset) begin
    mrac = 32'h0;
  end
  if (reset) begin
    mdseac = 32'h0;
  end
  if (reset) begin
    mfdht = 6'h0;
  end
  if (reset) begin
    mfdhs = 2'h0;
  end
  if (reset) begin
    force_halt_ctr_f = 32'h0;
  end
  if (reset) begin
    meivt = 22'h0;
  end
  if (reset) begin
    meihap = 8'h0;
  end
  if (reset) begin
    meicurpl = 4'h0;
  end
  if (reset) begin
    meicidpl = 4'h0;
  end
  if (reset) begin
    meipt = 4'h0;
  end
  if (reset) begin
    _T_691 = 16'h0;
  end
  if (reset) begin
    _T_716 = 31'h0;
  end
  if (reset) begin
    dicawics = 17'h0;
  end
  if (reset) begin
    dicad0 = 71'h0;
  end
  if (reset) begin
    dicad0h = 32'h0;
  end
  if (reset) begin
    _T_749 = 7'h0;
  end
  if (reset) begin
    icache_rd_valid_f = 1'h0;
  end
  if (reset) begin
    icache_wr_valid_f = 1'h0;
  end
  if (reset) begin
    mtsel = 2'h0;
  end
  if (reset) begin
    _T_863 = 10'h0;
  end
  if (reset) begin
    _T_864 = 10'h0;
  end
  if (reset) begin
    _T_865 = 10'h0;
  end
  if (reset) begin
    _T_866 = 10'h0;
  end
  if (reset) begin
    mtdata2_t_0 = 32'h0;
  end
  if (reset) begin
    mtdata2_t_1 = 32'h0;
  end
  if (reset) begin
    mtdata2_t_2 = 32'h0;
  end
  if (reset) begin
    mtdata2_t_3 = 32'h0;
  end
  if (reset) begin
    mhpme3 = 10'h0;
  end
  if (reset) begin
    mhpme4 = 10'h0;
  end
  if (reset) begin
    mhpme5 = 10'h0;
  end
  if (reset) begin
    mhpme6 = 10'h0;
  end
  if (reset) begin
    mhpmc_inc_r_d1_0 = 1'h0;
  end
  if (reset) begin
    mhpmc_inc_r_d1_1 = 1'h0;
  end
  if (reset) begin
    mhpmc_inc_r_d1_2 = 1'h0;
  end
  if (reset) begin
    mhpmc_inc_r_d1_3 = 1'h0;
  end
  if (reset) begin
    perfcnt_halted_d1 = 1'h0;
  end
  if (reset) begin
    mhpmc3h = 32'h0;
  end
  if (reset) begin
    mhpmc3 = 32'h0;
  end
  if (reset) begin
    mhpmc4h = 32'h0;
  end
  if (reset) begin
    mhpmc4 = 32'h0;
  end
  if (reset) begin
    mhpmc5h = 32'h0;
  end
  if (reset) begin
    mhpmc5 = 32'h0;
  end
  if (reset) begin
    mhpmc6h = 32'h0;
  end
  if (reset) begin
    mhpmc6 = 32'h0;
  end
  if (reset) begin
    _T_2321 = 1'h0;
  end
  if (reset) begin
    _T_2326 = 1'h0;
  end
  if (reset) begin
    _T_2327 = 5'h0;
  end
  if (reset) begin
    _T_2328 = 1'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge io_csr_wr_clk or posedge reset) begin
    if (reset) begin
      mpmc_b <= 1'h0;
    end else if (wr_mpmc_r) begin
      mpmc_b <= _T_500;
    end else begin
      mpmc_b <= _T_501;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      _T_56 <= 2'h0;
    end else begin
      _T_56 <= _T_48 | _T_44;
    end
  end
  always @(posedge rvclkhdr_io_l1clk or posedge reset) begin
    if (reset) begin
      _T_62 <= 31'h0;
    end else begin
      _T_62 <= {io_dec_csr_wrdata_r[31:2],io_dec_csr_wrdata_r[0]};
    end
  end
  always @(posedge rvclkhdr_14_io_l1clk or posedge reset) begin
    if (reset) begin
      mdccmect <= 32'h0;
    end else if (wr_mdccmect_r) begin
      mdccmect <= _T_515;
    end else begin
      mdccmect <= _T_559;
    end
  end
  always @(posedge rvclkhdr_13_io_l1clk or posedge reset) begin
    if (reset) begin
      miccmect <= 32'h0;
    end else if (wr_miccmect_r) begin
      miccmect <= _T_515;
    end else begin
      miccmect <= _T_538;
    end
  end
  always @(posedge rvclkhdr_12_io_l1clk or posedge reset) begin
    if (reset) begin
      micect <= 32'h0;
    end else if (wr_micect_r) begin
      micect <= _T_515;
    end else begin
      micect <= _T_517;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      _T_68 <= 6'h0;
    end else begin
      _T_68 <= {_T_67,_T_65};
    end
  end
  always @(posedge io_csr_wr_clk or posedge reset) begin
    if (reset) begin
      mie <= 6'h0;
    end else begin
      mie <= io_mie_ns;
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      temp_ncount6_2 <= 5'h0;
    end else if (wr_mcountinhibit_r) begin
      temp_ncount6_2 <= io_dec_csr_wrdata_r[6:2];
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      temp_ncount0 <= 1'h0;
    end else if (wr_mcountinhibit_r) begin
      temp_ncount0 <= io_dec_csr_wrdata_r[0];
    end
  end
  always @(posedge rvclkhdr_1_io_l1clk or posedge reset) begin
    if (reset) begin
      mcyclel <= 32'h0;
    end else if (wr_mcyclel_r) begin
      mcyclel <= io_dec_csr_wrdata_r;
    end else begin
      mcyclel <= mcyclel_inc[31:0];
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      mcyclel_cout_f <= 1'h0;
    end else begin
      mcyclel_cout_f <= mcyclel_cout & _T_98;
    end
  end
  always @(posedge rvclkhdr_2_io_l1clk or posedge reset) begin
    if (reset) begin
      mcycleh <= 32'h0;
    end else if (wr_mcycleh_r) begin
      mcycleh <= io_dec_csr_wrdata_r;
    end else begin
      mcycleh <= mcycleh_inc;
    end
  end
  always @(posedge rvclkhdr_3_io_l1clk or posedge reset) begin
    if (reset) begin
      minstretl <= 32'h0;
    end else if (wr_minstretl_r) begin
      minstretl <= io_dec_csr_wrdata_r;
    end else begin
      minstretl <= minstretl_inc[31:0];
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      minstret_enable_f <= 1'h0;
    end else begin
      minstret_enable_f <= i0_valid_no_ebreak_ecall_r | wr_minstretl_r;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      minstretl_cout_f <= 1'h0;
    end else begin
      minstretl_cout_f <= minstretl_cout & _T_125;
    end
  end
  always @(posedge rvclkhdr_4_io_l1clk or posedge reset) begin
    if (reset) begin
      minstreth <= 32'h0;
    end else if (wr_minstreth_r) begin
      minstreth <= io_dec_csr_wrdata_r;
    end else begin
      minstreth <= minstreth_inc;
    end
  end
  always @(posedge rvclkhdr_5_io_l1clk or posedge reset) begin
    if (reset) begin
      mscratch <= 32'h0;
    end else begin
      mscratch <= io_dec_csr_wrdata_r;
    end
  end
  always @(posedge rvclkhdr_6_io_l1clk or posedge reset) begin
    if (reset) begin
      _T_167 <= 31'h0;
    end else begin
      _T_167 <= io_npc_r;
    end
  end
  always @(posedge rvclkhdr_7_io_l1clk or posedge reset) begin
    if (reset) begin
      pc_r_d1 <= 31'h0;
    end else begin
      pc_r_d1 <= _T_171 | _T_172;
    end
  end
  always @(posedge io_e4e5_int_clk or posedge reset) begin
    if (reset) begin
      _T_196 <= 31'h0;
    end else begin
      _T_196 <= _T_194 | _T_192;
    end
  end
  always @(posedge io_e4e5_int_clk or posedge reset) begin
    if (reset) begin
      mcause <= 32'h0;
    end else begin
      mcause <= _T_234 | _T_230;
    end
  end
  always @(posedge io_e4e5_int_clk or posedge reset) begin
    if (reset) begin
      mscause <= 4'h0;
    end else begin
      mscause <= _T_264 | _T_263;
    end
  end
  always @(posedge io_e4e5_int_clk or posedge reset) begin
    if (reset) begin
      mtval <= 32'h0;
    end else begin
      mtval <= _T_321 | _T_317;
    end
  end
  always @(posedge rvclkhdr_8_io_l1clk or posedge reset) begin
    if (reset) begin
      mcgc <= 9'h0;
    end else begin
      mcgc <= io_dec_csr_wrdata_r[8:0];
    end
  end
  always @(posedge rvclkhdr_9_io_l1clk or posedge reset) begin
    if (reset) begin
      mfdc_int <= 15'h0;
    end else begin
      mfdc_int <= {_T_341,io_dec_csr_wrdata_r[11:0]};
    end
  end
  always @(posedge rvclkhdr_10_io_l1clk or posedge reset) begin
    if (reset) begin
      mrac <= 32'h0;
    end else begin
      mrac <= {_T_474,_T_459};
    end
  end
  always @(posedge rvclkhdr_11_io_l1clk or posedge reset) begin
    if (reset) begin
      mdseac <= 32'h0;
    end else begin
      mdseac <= io_lsu_imprecise_error_addr_any;
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      mfdht <= 6'h0;
    end else if (wr_mfdht_r) begin
      mfdht <= io_dec_csr_wrdata_r[5:0];
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      mfdhs <= 2'h0;
    end else if (_T_585) begin
      if (wr_mfdhs_r) begin
        mfdhs <= io_dec_csr_wrdata_r[1:0];
      end else if (_T_579) begin
        mfdhs <= _T_583;
      end
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      force_halt_ctr_f <= 32'h0;
    end else if (mfdht[0]) begin
      if (io_debug_halt_req_f) begin
        force_halt_ctr_f <= _T_590;
      end else if (io_dbg_tlu_halted_f) begin
        force_halt_ctr_f <= 32'h0;
      end
    end
  end
  always @(posedge rvclkhdr_15_io_l1clk or posedge reset) begin
    if (reset) begin
      meivt <= 22'h0;
    end else begin
      meivt <= io_dec_csr_wrdata_r[31:10];
    end
  end
  always @(posedge rvclkhdr_16_io_l1clk or posedge reset) begin
    if (reset) begin
      meihap <= 8'h0;
    end else begin
      meihap <= io_pic_claimid;
    end
  end
  always @(posedge io_csr_wr_clk or posedge reset) begin
    if (reset) begin
      meicurpl <= 4'h0;
    end else if (wr_meicurpl_r) begin
      meicurpl <= io_dec_csr_wrdata_r[3:0];
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      meicidpl <= 4'h0;
    end else if (wr_meicpct_r) begin
      meicidpl <= io_pic_pl;
    end else if (wr_meicidpl_r) begin
      meicidpl <= io_dec_csr_wrdata_r[3:0];
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      meipt <= 4'h0;
    end else if (wr_meipt_r) begin
      meipt <= io_dec_csr_wrdata_r[3:0];
    end
  end
  always @(posedge rvclkhdr_17_io_l1clk or posedge reset) begin
    if (reset) begin
      _T_691 <= 16'h0;
    end else if (enter_debug_halt_req_le) begin
      _T_691 <= _T_665;
    end else if (wr_dcsr_r) begin
      _T_691 <= _T_680;
    end else begin
      _T_691 <= _T_685;
    end
  end
  always @(posedge rvclkhdr_18_io_l1clk or posedge reset) begin
    if (reset) begin
      _T_716 <= 31'h0;
    end else begin
      _T_716 <= _T_711 | _T_710;
    end
  end
  always @(posedge rvclkhdr_19_io_l1clk or posedge reset) begin
    if (reset) begin
      dicawics <= 17'h0;
    end else begin
      dicawics <= {_T_720,io_dec_csr_wrdata_r[16:3]};
    end
  end
  always @(posedge rvclkhdr_20_io_l1clk or posedge reset) begin
    if (reset) begin
      dicad0 <= 71'h0;
    end else if (wr_dicad0_r) begin
      dicad0 <= {{39'd0}, io_dec_csr_wrdata_r};
    end else begin
      dicad0 <= io_ifu_ic_debug_rd_data;
    end
  end
  always @(posedge rvclkhdr_21_io_l1clk or posedge reset) begin
    if (reset) begin
      dicad0h <= 32'h0;
    end else if (wr_dicad0h_r) begin
      dicad0h <= io_dec_csr_wrdata_r;
    end else begin
      dicad0h <= io_ifu_ic_debug_rd_data[63:32];
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      _T_749 <= 7'h0;
    end else if (_T_747) begin
      if (_T_742) begin
        _T_749 <= io_dec_csr_wrdata_r[6:0];
      end else begin
        _T_749 <= io_ifu_ic_debug_rd_data[70:64];
      end
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      icache_rd_valid_f <= 1'h0;
    end else begin
      icache_rd_valid_f <= _T_759 & _T_761;
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      icache_wr_valid_f <= 1'h0;
    end else begin
      icache_wr_valid_f <= _T_653 & _T_764;
    end
  end
  always @(posedge io_csr_wr_clk or posedge reset) begin
    if (reset) begin
      mtsel <= 2'h0;
    end else if (wr_mtsel_r) begin
      mtsel <= io_dec_csr_wrdata_r[1:0];
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      _T_863 <= 10'h0;
    end else if (wr_mtdata1_t_r_0) begin
      _T_863 <= tdata_wrdata_r;
    end else begin
      _T_863 <= _T_834;
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      _T_864 <= 10'h0;
    end else if (wr_mtdata1_t_r_1) begin
      _T_864 <= tdata_wrdata_r;
    end else begin
      _T_864 <= _T_843;
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      _T_865 <= 10'h0;
    end else if (wr_mtdata1_t_r_2) begin
      _T_865 <= tdata_wrdata_r;
    end else begin
      _T_865 <= _T_852;
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      _T_866 <= 10'h0;
    end else if (wr_mtdata1_t_r_3) begin
      _T_866 <= tdata_wrdata_r;
    end else begin
      _T_866 <= _T_861;
    end
  end
  always @(posedge rvclkhdr_22_io_l1clk or posedge reset) begin
    if (reset) begin
      mtdata2_t_0 <= 32'h0;
    end else begin
      mtdata2_t_0 <= io_dec_csr_wrdata_r;
    end
  end
  always @(posedge rvclkhdr_23_io_l1clk or posedge reset) begin
    if (reset) begin
      mtdata2_t_1 <= 32'h0;
    end else begin
      mtdata2_t_1 <= io_dec_csr_wrdata_r;
    end
  end
  always @(posedge rvclkhdr_24_io_l1clk or posedge reset) begin
    if (reset) begin
      mtdata2_t_2 <= 32'h0;
    end else begin
      mtdata2_t_2 <= io_dec_csr_wrdata_r;
    end
  end
  always @(posedge rvclkhdr_25_io_l1clk or posedge reset) begin
    if (reset) begin
      mtdata2_t_3 <= 32'h0;
    end else begin
      mtdata2_t_3 <= io_dec_csr_wrdata_r;
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      mhpme3 <= 10'h0;
    end else if (wr_mhpme3_r) begin
      if (_T_2283) begin
        mhpme3 <= 10'h204;
      end else begin
        mhpme3 <= io_dec_csr_wrdata_r[9:0];
      end
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      mhpme4 <= 10'h0;
    end else if (wr_mhpme4_r) begin
      if (_T_2283) begin
        mhpme4 <= 10'h204;
      end else begin
        mhpme4 <= io_dec_csr_wrdata_r[9:0];
      end
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      mhpme5 <= 10'h0;
    end else if (wr_mhpme5_r) begin
      if (_T_2283) begin
        mhpme5 <= 10'h204;
      end else begin
        mhpme5 <= io_dec_csr_wrdata_r[9:0];
      end
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      mhpme6 <= 10'h0;
    end else if (wr_mhpme6_r) begin
      if (_T_2283) begin
        mhpme6 <= 10'h204;
      end else begin
        mhpme6 <= io_dec_csr_wrdata_r[9:0];
      end
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      mhpmc_inc_r_d1_0 <= 1'h0;
    end else begin
      mhpmc_inc_r_d1_0 <= _T_1016 & _T_1296;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      mhpmc_inc_r_d1_1 <= 1'h0;
    end else begin
      mhpmc_inc_r_d1_1 <= _T_1300 & _T_1580;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      mhpmc_inc_r_d1_2 <= 1'h0;
    end else begin
      mhpmc_inc_r_d1_2 <= _T_1584 & _T_1864;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      mhpmc_inc_r_d1_3 <= 1'h0;
    end else begin
      mhpmc_inc_r_d1_3 <= _T_1868 & _T_2148;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      perfcnt_halted_d1 <= 1'h0;
    end else begin
      perfcnt_halted_d1 <= _T_85 | io_dec_tlu_pmu_fw_halted;
    end
  end
  always @(posedge rvclkhdr_27_io_l1clk or posedge reset) begin
    if (reset) begin
      mhpmc3h <= 32'h0;
    end else if (mhpmc3h_wr_en0) begin
      mhpmc3h <= io_dec_csr_wrdata_r;
    end else begin
      mhpmc3h <= mhpmc3_incr[63:32];
    end
  end
  always @(posedge rvclkhdr_26_io_l1clk or posedge reset) begin
    if (reset) begin
      mhpmc3 <= 32'h0;
    end else if (mhpmc3_wr_en0) begin
      mhpmc3 <= io_dec_csr_wrdata_r;
    end else begin
      mhpmc3 <= mhpmc3_incr[31:0];
    end
  end
  always @(posedge rvclkhdr_29_io_l1clk or posedge reset) begin
    if (reset) begin
      mhpmc4h <= 32'h0;
    end else if (mhpmc4h_wr_en0) begin
      mhpmc4h <= io_dec_csr_wrdata_r;
    end else begin
      mhpmc4h <= mhpmc4_incr[63:32];
    end
  end
  always @(posedge rvclkhdr_28_io_l1clk or posedge reset) begin
    if (reset) begin
      mhpmc4 <= 32'h0;
    end else if (mhpmc4_wr_en0) begin
      mhpmc4 <= io_dec_csr_wrdata_r;
    end else begin
      mhpmc4 <= mhpmc4_incr[31:0];
    end
  end
  always @(posedge rvclkhdr_31_io_l1clk or posedge reset) begin
    if (reset) begin
      mhpmc5h <= 32'h0;
    end else if (mhpmc5h_wr_en0) begin
      mhpmc5h <= io_dec_csr_wrdata_r;
    end else begin
      mhpmc5h <= mhpmc5_incr[63:32];
    end
  end
  always @(posedge rvclkhdr_30_io_l1clk or posedge reset) begin
    if (reset) begin
      mhpmc5 <= 32'h0;
    end else if (mhpmc5_wr_en0) begin
      mhpmc5 <= io_dec_csr_wrdata_r;
    end else begin
      mhpmc5 <= mhpmc5_incr[31:0];
    end
  end
  always @(posedge rvclkhdr_33_io_l1clk or posedge reset) begin
    if (reset) begin
      mhpmc6h <= 32'h0;
    end else if (mhpmc6h_wr_en0) begin
      mhpmc6h <= io_dec_csr_wrdata_r;
    end else begin
      mhpmc6h <= mhpmc6_incr[63:32];
    end
  end
  always @(posedge rvclkhdr_32_io_l1clk or posedge reset) begin
    if (reset) begin
      mhpmc6 <= 32'h0;
    end else if (mhpmc6_wr_en0) begin
      mhpmc6 <= io_dec_csr_wrdata_r;
    end else begin
      mhpmc6 <= mhpmc6_incr[31:0];
    end
  end
  always @(posedge rvclkhdr_34_io_l1clk or posedge reset) begin
    if (reset) begin
      _T_2321 <= 1'h0;
    end else begin
      _T_2321 <= io_i0_valid_wb;
    end
  end
  always @(posedge rvclkhdr_34_io_l1clk or posedge reset) begin
    if (reset) begin
      _T_2326 <= 1'h0;
    end else begin
      _T_2326 <= _T_2322 | _T_2324;
    end
  end
  always @(posedge rvclkhdr_34_io_l1clk or posedge reset) begin
    if (reset) begin
      _T_2327 <= 5'h0;
    end else begin
      _T_2327 <= io_exc_cause_wb;
    end
  end
  always @(posedge rvclkhdr_34_io_l1clk or posedge reset) begin
    if (reset) begin
      _T_2328 <= 1'h0;
    end else begin
      _T_2328 <= io_interrupt_valid_r_d1;
    end
  end
endmodule
module dec_decode_csr_read(
  input  [11:0] io_dec_csr_rdaddr_d,
  output        io_csr_pkt_csr_misa,
  output        io_csr_pkt_csr_mvendorid,
  output        io_csr_pkt_csr_marchid,
  output        io_csr_pkt_csr_mimpid,
  output        io_csr_pkt_csr_mhartid,
  output        io_csr_pkt_csr_mstatus,
  output        io_csr_pkt_csr_mtvec,
  output        io_csr_pkt_csr_mip,
  output        io_csr_pkt_csr_mie,
  output        io_csr_pkt_csr_mcyclel,
  output        io_csr_pkt_csr_mcycleh,
  output        io_csr_pkt_csr_minstretl,
  output        io_csr_pkt_csr_minstreth,
  output        io_csr_pkt_csr_mscratch,
  output        io_csr_pkt_csr_mepc,
  output        io_csr_pkt_csr_mcause,
  output        io_csr_pkt_csr_mscause,
  output        io_csr_pkt_csr_mtval,
  output        io_csr_pkt_csr_mrac,
  output        io_csr_pkt_csr_dmst,
  output        io_csr_pkt_csr_mdseac,
  output        io_csr_pkt_csr_meihap,
  output        io_csr_pkt_csr_meivt,
  output        io_csr_pkt_csr_meipt,
  output        io_csr_pkt_csr_meicurpl,
  output        io_csr_pkt_csr_meicidpl,
  output        io_csr_pkt_csr_dcsr,
  output        io_csr_pkt_csr_mcgc,
  output        io_csr_pkt_csr_mfdc,
  output        io_csr_pkt_csr_dpc,
  output        io_csr_pkt_csr_mtsel,
  output        io_csr_pkt_csr_mtdata1,
  output        io_csr_pkt_csr_mtdata2,
  output        io_csr_pkt_csr_mhpmc3,
  output        io_csr_pkt_csr_mhpmc4,
  output        io_csr_pkt_csr_mhpmc5,
  output        io_csr_pkt_csr_mhpmc6,
  output        io_csr_pkt_csr_mhpmc3h,
  output        io_csr_pkt_csr_mhpmc4h,
  output        io_csr_pkt_csr_mhpmc5h,
  output        io_csr_pkt_csr_mhpmc6h,
  output        io_csr_pkt_csr_mhpme3,
  output        io_csr_pkt_csr_mhpme4,
  output        io_csr_pkt_csr_mhpme5,
  output        io_csr_pkt_csr_mhpme6,
  output        io_csr_pkt_csr_mcountinhibit,
  output        io_csr_pkt_csr_mitctl0,
  output        io_csr_pkt_csr_mitctl1,
  output        io_csr_pkt_csr_mitb0,
  output        io_csr_pkt_csr_mitb1,
  output        io_csr_pkt_csr_mitcnt0,
  output        io_csr_pkt_csr_mitcnt1,
  output        io_csr_pkt_csr_mpmc,
  output        io_csr_pkt_csr_meicpct,
  output        io_csr_pkt_csr_micect,
  output        io_csr_pkt_csr_miccmect,
  output        io_csr_pkt_csr_mdccmect,
  output        io_csr_pkt_csr_mfdht,
  output        io_csr_pkt_csr_mfdhs,
  output        io_csr_pkt_csr_dicawics,
  output        io_csr_pkt_csr_dicad0h,
  output        io_csr_pkt_csr_dicad0,
  output        io_csr_pkt_csr_dicad1,
  output        io_csr_pkt_csr_dicago,
  output        io_csr_pkt_presync,
  output        io_csr_pkt_postsync,
  output        io_csr_pkt_legal
);
  wire  _T_1 = ~io_dec_csr_rdaddr_d[11]; // @[dec_tlu_ctl.scala 2570:129]
  wire  _T_3 = ~io_dec_csr_rdaddr_d[6]; // @[dec_tlu_ctl.scala 2570:129]
  wire  _T_5 = ~io_dec_csr_rdaddr_d[5]; // @[dec_tlu_ctl.scala 2570:129]
  wire  _T_7 = ~io_dec_csr_rdaddr_d[2]; // @[dec_tlu_ctl.scala 2570:129]
  wire  _T_9 = _T_1 & _T_3; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_10 = _T_9 & _T_5; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_11 = _T_10 & _T_7; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_15 = ~io_dec_csr_rdaddr_d[7]; // @[dec_tlu_ctl.scala 2570:129]
  wire  _T_17 = ~io_dec_csr_rdaddr_d[1]; // @[dec_tlu_ctl.scala 2570:129]
  wire  _T_19 = io_dec_csr_rdaddr_d[10] & _T_15; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_20 = _T_19 & _T_17; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_27 = ~io_dec_csr_rdaddr_d[0]; // @[dec_tlu_ctl.scala 2570:165]
  wire  _T_29 = _T_19 & io_dec_csr_rdaddr_d[1]; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_36 = io_dec_csr_rdaddr_d[10] & _T_3; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_37 = _T_36 & io_dec_csr_rdaddr_d[1]; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_69 = _T_10 & io_dec_csr_rdaddr_d[2]; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_70 = _T_69 & io_dec_csr_rdaddr_d[0]; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_75 = _T_15 & io_dec_csr_rdaddr_d[6]; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_94 = ~io_dec_csr_rdaddr_d[4]; // @[dec_tlu_ctl.scala 2570:129]
  wire  _T_96 = ~io_dec_csr_rdaddr_d[3]; // @[dec_tlu_ctl.scala 2570:129]
  wire  _T_101 = io_dec_csr_rdaddr_d[11] & _T_15; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_102 = _T_101 & _T_94; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_103 = _T_102 & _T_96; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_104 = _T_103 & _T_7; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_119 = io_dec_csr_rdaddr_d[7] & _T_3; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_120 = _T_119 & _T_5; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_121 = _T_120 & _T_94; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_122 = _T_121 & _T_96; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_123 = _T_122 & _T_7; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_138 = _T_15 & _T_3; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_139 = _T_138 & _T_94; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_140 = _T_139 & _T_96; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_141 = _T_140 & _T_7; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_142 = _T_141 & io_dec_csr_rdaddr_d[1]; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_145 = ~io_dec_csr_rdaddr_d[10]; // @[dec_tlu_ctl.scala 2570:129]
  wire  _T_156 = _T_145 & io_dec_csr_rdaddr_d[7]; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_157 = _T_156 & _T_94; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_158 = _T_157 & _T_96; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_159 = _T_158 & _T_7; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_160 = _T_159 & io_dec_csr_rdaddr_d[1]; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_172 = _T_75 & _T_7; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_173 = _T_172 & _T_17; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_182 = _T_75 & _T_17; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_183 = _T_182 & io_dec_csr_rdaddr_d[0]; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_191 = _T_75 & io_dec_csr_rdaddr_d[1]; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_196 = io_dec_csr_rdaddr_d[6] & io_dec_csr_rdaddr_d[5]; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_217 = _T_1 & io_dec_csr_rdaddr_d[7]; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_218 = _T_217 & _T_5; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_219 = _T_218 & _T_96; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_220 = _T_219 & _T_7; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_230 = io_dec_csr_rdaddr_d[10] & _T_94; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_231 = _T_230 & _T_96; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_232 = _T_231 & io_dec_csr_rdaddr_d[2]; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_240 = io_dec_csr_rdaddr_d[11] & io_dec_csr_rdaddr_d[10]; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_241 = _T_240 & _T_94; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_258 = _T_145 & io_dec_csr_rdaddr_d[6]; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_259 = _T_258 & io_dec_csr_rdaddr_d[3]; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_260 = _T_259 & _T_7; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_261 = _T_260 & _T_17; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_268 = io_dec_csr_rdaddr_d[11] & io_dec_csr_rdaddr_d[6]; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_269 = _T_268 & _T_17; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_281 = _T_268 & io_dec_csr_rdaddr_d[1]; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_291 = _T_36 & io_dec_csr_rdaddr_d[5]; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_292 = _T_291 & io_dec_csr_rdaddr_d[4]; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_299 = io_dec_csr_rdaddr_d[10] & io_dec_csr_rdaddr_d[4]; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_300 = _T_299 & io_dec_csr_rdaddr_d[3]; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_310 = _T_300 & _T_17; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_311 = _T_310 & io_dec_csr_rdaddr_d[0]; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_330 = io_dec_csr_rdaddr_d[10] & io_dec_csr_rdaddr_d[5]; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_331 = _T_330 & _T_94; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_332 = _T_331 & _T_17; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_342 = _T_231 & io_dec_csr_rdaddr_d[0]; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_381 = _T_103 & io_dec_csr_rdaddr_d[2]; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_382 = _T_381 & _T_17; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_397 = _T_103 & _T_17; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_411 = _T_15 & _T_5; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_412 = _T_411 & _T_94; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_413 = _T_412 & _T_96; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_414 = _T_413 & io_dec_csr_rdaddr_d[2]; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_415 = _T_414 & io_dec_csr_rdaddr_d[1]; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_426 = io_dec_csr_rdaddr_d[7] & _T_94; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_427 = _T_426 & _T_96; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_428 = _T_427 & _T_7; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_429 = _T_428 & io_dec_csr_rdaddr_d[1]; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_444 = _T_119 & _T_94; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_445 = _T_444 & _T_96; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_446 = _T_445 & io_dec_csr_rdaddr_d[2]; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_447 = _T_446 & _T_17; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_460 = _T_427 & io_dec_csr_rdaddr_d[2]; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_461 = _T_460 & _T_17; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_478 = _T_446 & io_dec_csr_rdaddr_d[1]; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_490 = _T_15 & io_dec_csr_rdaddr_d[5]; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_491 = _T_490 & _T_94; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_492 = _T_491 & _T_96; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_493 = _T_492 & _T_7; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_505 = io_dec_csr_rdaddr_d[5] & _T_94; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_506 = _T_505 & _T_96; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_507 = _T_506 & io_dec_csr_rdaddr_d[2]; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_508 = _T_507 & _T_17; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_536 = _T_507 & io_dec_csr_rdaddr_d[1]; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_553 = _T_493 & _T_27; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_562 = io_dec_csr_rdaddr_d[6] & _T_5; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_563 = _T_562 & io_dec_csr_rdaddr_d[4]; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_564 = _T_563 & _T_17; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_572 = io_dec_csr_rdaddr_d[6] & _T_96; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_573 = _T_572 & io_dec_csr_rdaddr_d[2]; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_574 = _T_573 & io_dec_csr_rdaddr_d[1]; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_585 = _T_563 & _T_7; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_593 = io_dec_csr_rdaddr_d[6] & io_dec_csr_rdaddr_d[4]; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_594 = _T_593 & io_dec_csr_rdaddr_d[2]; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_595 = _T_594 & io_dec_csr_rdaddr_d[1]; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_614 = io_dec_csr_rdaddr_d[6] & io_dec_csr_rdaddr_d[2]; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_615 = _T_614 & _T_17; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_624 = io_dec_csr_rdaddr_d[6] & _T_94; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_625 = _T_624 & _T_96; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_626 = _T_625 & io_dec_csr_rdaddr_d[2]; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_668 = _T_196 & _T_96; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_669 = _T_668 & _T_17; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_685 = _T_196 & io_dec_csr_rdaddr_d[1]; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_693 = io_dec_csr_rdaddr_d[6] & io_dec_csr_rdaddr_d[3]; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_694 = _T_693 & io_dec_csr_rdaddr_d[2]; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_695 = _T_694 & io_dec_csr_rdaddr_d[1]; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_703 = _T_624 & io_dec_csr_rdaddr_d[2]; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_716 = _T_1 & _T_5; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_717 = _T_716 & io_dec_csr_rdaddr_d[3]; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_718 = _T_717 & _T_7; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_719 = _T_718 & _T_17; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_726 = io_dec_csr_rdaddr_d[10] & io_dec_csr_rdaddr_d[3]; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_727 = _T_726 & io_dec_csr_rdaddr_d[2]; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_737 = _T_230 & io_dec_csr_rdaddr_d[3]; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_738 = _T_737 & _T_17; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_748 = _T_726 & _T_7; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_749 = _T_748 & io_dec_csr_rdaddr_d[1]; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_787 = _T_311 | _T_553; // @[dec_tlu_ctl.scala 2638:81]
  wire  _T_799 = _T_3 & _T_5; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_800 = _T_799 & _T_94; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_801 = _T_800 & _T_96; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_802 = _T_801 & _T_7; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_803 = _T_802 & io_dec_csr_rdaddr_d[1]; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_804 = _T_787 | _T_803; // @[dec_tlu_ctl.scala 2638:121]
  wire  _T_813 = io_dec_csr_rdaddr_d[11] & _T_94; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_814 = _T_813 & _T_96; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_815 = _T_814 & io_dec_csr_rdaddr_d[2]; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_816 = _T_815 & _T_17; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_817 = _T_804 | _T_816; // @[dec_tlu_ctl.scala 2638:155]
  wire  _T_828 = _T_814 & io_dec_csr_rdaddr_d[1]; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_829 = _T_828 & _T_27; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_830 = _T_817 | _T_829; // @[dec_tlu_ctl.scala 2639:97]
  wire  _T_841 = io_dec_csr_rdaddr_d[7] & _T_5; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_842 = _T_841 & _T_94; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_843 = _T_842 & _T_96; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_844 = _T_843 & _T_7; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_845 = _T_844 & io_dec_csr_rdaddr_d[1]; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_869 = _T_311 | _T_70; // @[dec_tlu_ctl.scala 2640:81]
  wire  _T_879 = _T_869 | _T_183; // @[dec_tlu_ctl.scala 2640:121]
  wire  _T_889 = _T_879 | _T_342; // @[dec_tlu_ctl.scala 2640:162]
  wire  _T_904 = _T_1 & _T_15; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_905 = _T_904 & _T_3; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_906 = _T_905 & _T_94; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_907 = _T_906 & _T_96; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_908 = _T_907 & _T_7; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_909 = _T_908 & _T_27; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_910 = _T_889 | _T_909; // @[dec_tlu_ctl.scala 2641:105]
  wire  _T_922 = _T_217 & io_dec_csr_rdaddr_d[6]; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_923 = _T_922 & _T_94; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_924 = _T_923 & _T_96; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_925 = _T_924 & _T_17; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_926 = _T_910 | _T_925; // @[dec_tlu_ctl.scala 2641:145]
  wire  _T_937 = _T_231 & _T_7; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_938 = _T_937 & io_dec_csr_rdaddr_d[1]; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_955 = _T_1 & io_dec_csr_rdaddr_d[10]; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_956 = _T_955 & io_dec_csr_rdaddr_d[9]; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_957 = _T_956 & io_dec_csr_rdaddr_d[8]; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_958 = _T_957 & io_dec_csr_rdaddr_d[7]; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_959 = _T_958 & io_dec_csr_rdaddr_d[6]; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_960 = _T_959 & io_dec_csr_rdaddr_d[4]; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_961 = _T_960 & _T_96; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_962 = _T_961 & _T_7; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_963 = _T_962 & io_dec_csr_rdaddr_d[1]; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_964 = _T_963 & _T_27; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_983 = _T_1 & _T_145; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_984 = _T_983 & io_dec_csr_rdaddr_d[9]; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_985 = _T_984 & io_dec_csr_rdaddr_d[8]; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_986 = _T_985 & _T_15; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_987 = _T_986 & _T_3; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_988 = _T_987 & _T_5; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_989 = _T_988 & _T_94; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_990 = _T_989 & _T_96; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_991 = _T_990 & _T_17; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_992 = _T_964 | _T_991; // @[dec_tlu_ctl.scala 2643:81]
  wire  _T_1013 = _T_987 & io_dec_csr_rdaddr_d[5]; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_1014 = _T_1013 & _T_17; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_1015 = _T_1014 & _T_27; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_1016 = _T_992 | _T_1015; // @[dec_tlu_ctl.scala 2643:129]
  wire  _T_1032 = io_dec_csr_rdaddr_d[11] & io_dec_csr_rdaddr_d[9]; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_1033 = _T_1032 & io_dec_csr_rdaddr_d[8]; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_1034 = _T_1033 & io_dec_csr_rdaddr_d[7]; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_1035 = _T_1034 & io_dec_csr_rdaddr_d[6]; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_1036 = _T_1035 & _T_5; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_1037 = _T_1036 & _T_94; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_1038 = _T_1037 & _T_7; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_1039 = _T_1038 & _T_17; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_1040 = _T_1039 & _T_27; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_1041 = _T_1016 | _T_1040; // @[dec_tlu_ctl.scala 2644:105]
  wire  _T_1053 = io_dec_csr_rdaddr_d[11] & _T_145; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_1054 = _T_1053 & io_dec_csr_rdaddr_d[9]; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_1055 = _T_1054 & io_dec_csr_rdaddr_d[8]; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_1056 = _T_1055 & _T_3; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_1057 = _T_1056 & _T_5; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_1058 = _T_1057 & _T_27; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_1059 = _T_1041 | _T_1058; // @[dec_tlu_ctl.scala 2644:153]
  wire  _T_1078 = _T_959 & io_dec_csr_rdaddr_d[5]; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_1079 = _T_1078 & io_dec_csr_rdaddr_d[4]; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_1080 = _T_1079 & io_dec_csr_rdaddr_d[3]; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_1081 = _T_1080 & io_dec_csr_rdaddr_d[2]; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_1082 = _T_1081 & io_dec_csr_rdaddr_d[1]; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_1083 = _T_1082 & io_dec_csr_rdaddr_d[0]; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_1084 = _T_1059 | _T_1083; // @[dec_tlu_ctl.scala 2645:105]
  wire  _T_1105 = _T_1079 & _T_7; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_1106 = _T_1105 & _T_17; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_1107 = _T_1084 | _T_1106; // @[dec_tlu_ctl.scala 2645:153]
  wire  _T_1125 = _T_1033 & _T_15; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_1126 = _T_1125 & _T_3; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_1127 = _T_1126 & _T_5; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_1128 = _T_1127 & io_dec_csr_rdaddr_d[4]; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_1129 = _T_1128 & _T_96; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_1130 = _T_1129 & _T_7; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_1131 = _T_1130 & io_dec_csr_rdaddr_d[0]; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_1132 = _T_1107 | _T_1131; // @[dec_tlu_ctl.scala 2646:105]
  wire  _T_1152 = _T_958 & _T_3; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_1153 = _T_1152 & io_dec_csr_rdaddr_d[5]; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_1154 = _T_1153 & _T_96; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_1155 = _T_1154 & _T_7; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_1156 = _T_1155 & _T_17; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_1157 = _T_1132 | _T_1156; // @[dec_tlu_ctl.scala 2646:161]
  wire  _T_1176 = _T_1013 & io_dec_csr_rdaddr_d[2]; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_1177 = _T_1157 | _T_1176; // @[dec_tlu_ctl.scala 2647:105]
  wire  _T_1202 = _T_1129 & io_dec_csr_rdaddr_d[2]; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_1203 = _T_1202 & _T_17; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_1204 = _T_1203 & _T_27; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_1205 = _T_1177 | _T_1204; // @[dec_tlu_ctl.scala 2647:161]
  wire  _T_1224 = _T_959 & _T_5; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_1225 = _T_1224 & _T_94; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_1226 = _T_1225 & io_dec_csr_rdaddr_d[3]; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_1227 = _T_1226 & io_dec_csr_rdaddr_d[1]; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_1228 = _T_1205 | _T_1227; // @[dec_tlu_ctl.scala 2648:97]
  wire  _T_1248 = _T_1224 & io_dec_csr_rdaddr_d[4]; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_1249 = _T_1248 & _T_96; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_1250 = _T_1249 & io_dec_csr_rdaddr_d[2]; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_1251 = _T_1228 | _T_1250; // @[dec_tlu_ctl.scala 2648:153]
  wire  _T_1275 = _T_1130 & io_dec_csr_rdaddr_d[1]; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_1276 = _T_1251 | _T_1275; // @[dec_tlu_ctl.scala 2649:105]
  wire  _T_1296 = _T_1013 & io_dec_csr_rdaddr_d[1]; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_1297 = _T_1296 & io_dec_csr_rdaddr_d[0]; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_1298 = _T_1276 | _T_1297; // @[dec_tlu_ctl.scala 2649:161]
  wire  _T_1315 = _T_1055 & io_dec_csr_rdaddr_d[7]; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_1316 = _T_1315 & _T_5; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_1317 = _T_1316 & _T_94; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_1318 = _T_1317 & io_dec_csr_rdaddr_d[3]; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_1319 = _T_1318 & _T_7; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_1320 = _T_1298 | _T_1319; // @[dec_tlu_ctl.scala 2650:105]
  wire  _T_1343 = _T_1318 & _T_17; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_1344 = _T_1343 & _T_27; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_1345 = _T_1320 | _T_1344; // @[dec_tlu_ctl.scala 2650:161]
  wire  _T_1361 = _T_1057 & io_dec_csr_rdaddr_d[2]; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_1362 = _T_1345 | _T_1361; // @[dec_tlu_ctl.scala 2651:105]
  wire  _T_1384 = _T_1249 & io_dec_csr_rdaddr_d[1]; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_1385 = _T_1362 | _T_1384; // @[dec_tlu_ctl.scala 2651:161]
  wire  _T_1406 = _T_1225 & _T_27; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_1407 = _T_1385 | _T_1406; // @[dec_tlu_ctl.scala 2652:105]
  wire  _T_1430 = _T_1226 & _T_7; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_1431 = _T_1407 | _T_1430; // @[dec_tlu_ctl.scala 2652:161]
  wire  _T_1455 = _T_1153 & _T_94; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_1456 = _T_1455 & _T_96; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_1457 = _T_1456 & _T_7; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_1458 = _T_1457 & _T_27; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_1459 = _T_1431 | _T_1458; // @[dec_tlu_ctl.scala 2653:105]
  wire  _T_1475 = _T_1057 & io_dec_csr_rdaddr_d[1]; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_1476 = _T_1459 | _T_1475; // @[dec_tlu_ctl.scala 2653:153]
  wire  _T_1498 = _T_986 & io_dec_csr_rdaddr_d[6]; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_1499 = _T_1498 & _T_5; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_1500 = _T_1499 & _T_94; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_1501 = _T_1500 & _T_96; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_1502 = _T_1501 & _T_7; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_1503 = _T_1476 | _T_1502; // @[dec_tlu_ctl.scala 2654:113]
  wire  _T_1526 = _T_986 & _T_5; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_1527 = _T_1526 & _T_94; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_1528 = _T_1527 & _T_96; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_1529 = _T_1528 & _T_17; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_1530 = _T_1529 & _T_27; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_1531 = _T_1503 | _T_1530; // @[dec_tlu_ctl.scala 2654:161]
  wire  _T_1550 = _T_1013 & io_dec_csr_rdaddr_d[3]; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_1551 = _T_1531 | _T_1550; // @[dec_tlu_ctl.scala 2655:97]
  wire  _T_1567 = _T_1057 & io_dec_csr_rdaddr_d[3]; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_1568 = _T_1551 | _T_1567; // @[dec_tlu_ctl.scala 2655:153]
  wire  _T_1587 = _T_1013 & io_dec_csr_rdaddr_d[4]; // @[dec_tlu_ctl.scala 2570:198]
  wire  _T_1588 = _T_1568 | _T_1587; // @[dec_tlu_ctl.scala 2656:113]
  wire  _T_1604 = _T_1057 & io_dec_csr_rdaddr_d[4]; // @[dec_tlu_ctl.scala 2570:198]
  assign io_csr_pkt_csr_misa = _T_11 & io_dec_csr_rdaddr_d[0]; // @[dec_tlu_ctl.scala 2572:57]
  assign io_csr_pkt_csr_mvendorid = _T_20 & io_dec_csr_rdaddr_d[0]; // @[dec_tlu_ctl.scala 2573:57]
  assign io_csr_pkt_csr_marchid = _T_29 & _T_27; // @[dec_tlu_ctl.scala 2574:57]
  assign io_csr_pkt_csr_mimpid = _T_37 & io_dec_csr_rdaddr_d[0]; // @[dec_tlu_ctl.scala 2575:57]
  assign io_csr_pkt_csr_mhartid = _T_19 & io_dec_csr_rdaddr_d[2]; // @[dec_tlu_ctl.scala 2576:57]
  assign io_csr_pkt_csr_mstatus = _T_11 & _T_27; // @[dec_tlu_ctl.scala 2577:57]
  assign io_csr_pkt_csr_mtvec = _T_69 & io_dec_csr_rdaddr_d[0]; // @[dec_tlu_ctl.scala 2578:57]
  assign io_csr_pkt_csr_mip = _T_75 & io_dec_csr_rdaddr_d[2]; // @[dec_tlu_ctl.scala 2579:65]
  assign io_csr_pkt_csr_mie = _T_69 & _T_27; // @[dec_tlu_ctl.scala 2580:65]
  assign io_csr_pkt_csr_mcyclel = _T_104 & _T_17; // @[dec_tlu_ctl.scala 2581:57]
  assign io_csr_pkt_csr_mcycleh = _T_123 & _T_17; // @[dec_tlu_ctl.scala 2582:57]
  assign io_csr_pkt_csr_minstretl = _T_142 & _T_27; // @[dec_tlu_ctl.scala 2583:57]
  assign io_csr_pkt_csr_minstreth = _T_160 & _T_27; // @[dec_tlu_ctl.scala 2584:57]
  assign io_csr_pkt_csr_mscratch = _T_173 & _T_27; // @[dec_tlu_ctl.scala 2585:57]
  assign io_csr_pkt_csr_mepc = _T_182 & io_dec_csr_rdaddr_d[0]; // @[dec_tlu_ctl.scala 2586:57]
  assign io_csr_pkt_csr_mcause = _T_191 & _T_27; // @[dec_tlu_ctl.scala 2587:57]
  assign io_csr_pkt_csr_mscause = _T_196 & io_dec_csr_rdaddr_d[2]; // @[dec_tlu_ctl.scala 2588:57]
  assign io_csr_pkt_csr_mtval = _T_191 & io_dec_csr_rdaddr_d[0]; // @[dec_tlu_ctl.scala 2589:57]
  assign io_csr_pkt_csr_mrac = _T_220 & _T_17; // @[dec_tlu_ctl.scala 2590:57]
  assign io_csr_pkt_csr_dmst = _T_232 & _T_17; // @[dec_tlu_ctl.scala 2591:57]
  assign io_csr_pkt_csr_mdseac = _T_241 & _T_96; // @[dec_tlu_ctl.scala 2592:57]
  assign io_csr_pkt_csr_meihap = _T_240 & io_dec_csr_rdaddr_d[3]; // @[dec_tlu_ctl.scala 2593:57]
  assign io_csr_pkt_csr_meivt = _T_261 & _T_27; // @[dec_tlu_ctl.scala 2594:57]
  assign io_csr_pkt_csr_meipt = _T_269 & io_dec_csr_rdaddr_d[0]; // @[dec_tlu_ctl.scala 2595:57]
  assign io_csr_pkt_csr_meicurpl = _T_268 & io_dec_csr_rdaddr_d[2]; // @[dec_tlu_ctl.scala 2596:57]
  assign io_csr_pkt_csr_meicidpl = _T_281 & io_dec_csr_rdaddr_d[0]; // @[dec_tlu_ctl.scala 2597:57]
  assign io_csr_pkt_csr_dcsr = _T_292 & _T_27; // @[dec_tlu_ctl.scala 2598:57]
  assign io_csr_pkt_csr_mcgc = _T_300 & _T_27; // @[dec_tlu_ctl.scala 2599:57]
  assign io_csr_pkt_csr_mfdc = _T_310 & io_dec_csr_rdaddr_d[0]; // @[dec_tlu_ctl.scala 2600:57]
  assign io_csr_pkt_csr_dpc = _T_292 & io_dec_csr_rdaddr_d[0]; // @[dec_tlu_ctl.scala 2601:65]
  assign io_csr_pkt_csr_mtsel = _T_332 & _T_27; // @[dec_tlu_ctl.scala 2602:57]
  assign io_csr_pkt_csr_mtdata1 = _T_231 & io_dec_csr_rdaddr_d[0]; // @[dec_tlu_ctl.scala 2603:57]
  assign io_csr_pkt_csr_mtdata2 = _T_331 & io_dec_csr_rdaddr_d[1]; // @[dec_tlu_ctl.scala 2604:57]
  assign io_csr_pkt_csr_mhpmc3 = _T_104 & io_dec_csr_rdaddr_d[0]; // @[dec_tlu_ctl.scala 2605:57]
  assign io_csr_pkt_csr_mhpmc4 = _T_382 & _T_27; // @[dec_tlu_ctl.scala 2606:57]
  assign io_csr_pkt_csr_mhpmc5 = _T_397 & io_dec_csr_rdaddr_d[0]; // @[dec_tlu_ctl.scala 2607:57]
  assign io_csr_pkt_csr_mhpmc6 = _T_415 & _T_27; // @[dec_tlu_ctl.scala 2608:57]
  assign io_csr_pkt_csr_mhpmc3h = _T_429 & io_dec_csr_rdaddr_d[0]; // @[dec_tlu_ctl.scala 2609:57]
  assign io_csr_pkt_csr_mhpmc4h = _T_447 & _T_27; // @[dec_tlu_ctl.scala 2610:57]
  assign io_csr_pkt_csr_mhpmc5h = _T_461 & io_dec_csr_rdaddr_d[0]; // @[dec_tlu_ctl.scala 2611:57]
  assign io_csr_pkt_csr_mhpmc6h = _T_478 & _T_27; // @[dec_tlu_ctl.scala 2612:57]
  assign io_csr_pkt_csr_mhpme3 = _T_493 & io_dec_csr_rdaddr_d[0]; // @[dec_tlu_ctl.scala 2613:57]
  assign io_csr_pkt_csr_mhpme4 = _T_508 & _T_27; // @[dec_tlu_ctl.scala 2614:57]
  assign io_csr_pkt_csr_mhpme5 = _T_508 & io_dec_csr_rdaddr_d[0]; // @[dec_tlu_ctl.scala 2615:57]
  assign io_csr_pkt_csr_mhpme6 = _T_536 & _T_27; // @[dec_tlu_ctl.scala 2616:57]
  assign io_csr_pkt_csr_mcountinhibit = _T_493 & _T_27; // @[dec_tlu_ctl.scala 2617:49]
  assign io_csr_pkt_csr_mitctl0 = _T_564 & _T_27; // @[dec_tlu_ctl.scala 2618:57]
  assign io_csr_pkt_csr_mitctl1 = _T_574 & io_dec_csr_rdaddr_d[0]; // @[dec_tlu_ctl.scala 2619:57]
  assign io_csr_pkt_csr_mitb0 = _T_585 & io_dec_csr_rdaddr_d[0]; // @[dec_tlu_ctl.scala 2620:57]
  assign io_csr_pkt_csr_mitb1 = _T_595 & _T_27; // @[dec_tlu_ctl.scala 2621:57]
  assign io_csr_pkt_csr_mitcnt0 = _T_585 & _T_27; // @[dec_tlu_ctl.scala 2622:57]
  assign io_csr_pkt_csr_mitcnt1 = _T_615 & io_dec_csr_rdaddr_d[0]; // @[dec_tlu_ctl.scala 2623:57]
  assign io_csr_pkt_csr_mpmc = _T_626 & io_dec_csr_rdaddr_d[1]; // @[dec_tlu_ctl.scala 2624:57]
  assign io_csr_pkt_csr_meicpct = _T_281 & _T_27; // @[dec_tlu_ctl.scala 2626:57]
  assign io_csr_pkt_csr_micect = _T_669 & _T_27; // @[dec_tlu_ctl.scala 2628:57]
  assign io_csr_pkt_csr_miccmect = _T_668 & io_dec_csr_rdaddr_d[0]; // @[dec_tlu_ctl.scala 2629:57]
  assign io_csr_pkt_csr_mdccmect = _T_685 & _T_27; // @[dec_tlu_ctl.scala 2630:57]
  assign io_csr_pkt_csr_mfdht = _T_695 & _T_27; // @[dec_tlu_ctl.scala 2631:57]
  assign io_csr_pkt_csr_mfdhs = _T_703 & io_dec_csr_rdaddr_d[0]; // @[dec_tlu_ctl.scala 2632:57]
  assign io_csr_pkt_csr_dicawics = _T_719 & _T_27; // @[dec_tlu_ctl.scala 2633:57]
  assign io_csr_pkt_csr_dicad0h = _T_727 & _T_17; // @[dec_tlu_ctl.scala 2634:57]
  assign io_csr_pkt_csr_dicad0 = _T_738 & io_dec_csr_rdaddr_d[0]; // @[dec_tlu_ctl.scala 2635:57]
  assign io_csr_pkt_csr_dicad1 = _T_749 & _T_27; // @[dec_tlu_ctl.scala 2636:57]
  assign io_csr_pkt_csr_dicago = _T_749 & io_dec_csr_rdaddr_d[0]; // @[dec_tlu_ctl.scala 2637:57]
  assign io_csr_pkt_presync = _T_830 | _T_845; // @[dec_tlu_ctl.scala 2638:34]
  assign io_csr_pkt_postsync = _T_926 | _T_938; // @[dec_tlu_ctl.scala 2640:30]
  assign io_csr_pkt_legal = _T_1588 | _T_1604; // @[dec_tlu_ctl.scala 2643:26]
endmodule
module dec_tlu_ctl(
  input         clock,
  input         reset,
  output [29:0] io_tlu_exu_dec_tlu_meihap,
  output        io_tlu_exu_dec_tlu_flush_lower_r,
  output [30:0] io_tlu_exu_dec_tlu_flush_path_r,
  input  [1:0]  io_tlu_exu_exu_i0_br_hist_r,
  input         io_tlu_exu_exu_i0_br_error_r,
  input         io_tlu_exu_exu_i0_br_start_error_r,
  input         io_tlu_exu_exu_i0_br_valid_r,
  input         io_tlu_exu_exu_i0_br_mp_r,
  input         io_tlu_exu_exu_i0_br_middle_r,
  input         io_tlu_exu_exu_pmu_i0_br_misp,
  input         io_tlu_exu_exu_pmu_i0_br_ataken,
  input         io_tlu_exu_exu_pmu_i0_pc4,
  input  [30:0] io_tlu_exu_exu_npc_r,
  input         io_tlu_dma_dma_pmu_dccm_read,
  input         io_tlu_dma_dma_pmu_dccm_write,
  input         io_tlu_dma_dma_pmu_any_read,
  input         io_tlu_dma_dma_pmu_any_write,
  output [2:0]  io_tlu_dma_dec_tlu_dma_qos_prty,
  input         io_tlu_dma_dma_dccm_stall_any,
  input         io_tlu_dma_dma_iccm_stall_any,
  input         io_active_clk,
  input         io_free_clk,
  input         io_scan_mode,
  input  [30:0] io_rst_vec,
  input         io_nmi_int,
  input  [30:0] io_nmi_vec,
  input         io_i_cpu_halt_req,
  input         io_i_cpu_run_req,
  input         io_lsu_fastint_stall_any,
  input         io_lsu_idle_any,
  input         io_dec_pmu_instr_decoded,
  input         io_dec_pmu_decode_stall,
  input         io_dec_pmu_presync_stall,
  input         io_dec_pmu_postsync_stall,
  input         io_lsu_store_stall_any,
  input  [30:0] io_lsu_fir_addr,
  input  [1:0]  io_lsu_fir_error,
  input         io_iccm_dma_sb_error,
  input         io_lsu_error_pkt_r_valid,
  input         io_lsu_error_pkt_r_bits_single_ecc_error,
  input         io_lsu_error_pkt_r_bits_inst_type,
  input         io_lsu_error_pkt_r_bits_exc_type,
  input  [3:0]  io_lsu_error_pkt_r_bits_mscause,
  input  [31:0] io_lsu_error_pkt_r_bits_addr,
  input         io_lsu_single_ecc_error_incr,
  input         io_dec_pause_state,
  input         io_dec_csr_wen_unq_d,
  input         io_dec_csr_any_unq_d,
  input  [11:0] io_dec_csr_rdaddr_d,
  input         io_dec_csr_wen_r,
  input  [11:0] io_dec_csr_wraddr_r,
  input  [31:0] io_dec_csr_wrdata_r,
  input         io_dec_csr_stall_int_ff,
  input         io_dec_tlu_i0_valid_r,
  input  [30:0] io_dec_tlu_i0_pc_r,
  input         io_dec_tlu_packet_r_legal,
  input         io_dec_tlu_packet_r_icaf,
  input         io_dec_tlu_packet_r_icaf_f1,
  input  [1:0]  io_dec_tlu_packet_r_icaf_type,
  input         io_dec_tlu_packet_r_fence_i,
  input  [3:0]  io_dec_tlu_packet_r_i0trigger,
  input  [3:0]  io_dec_tlu_packet_r_pmu_i0_itype,
  input         io_dec_tlu_packet_r_pmu_i0_br_unpred,
  input         io_dec_tlu_packet_r_pmu_divide,
  input         io_dec_tlu_packet_r_pmu_lsu_misaligned,
  input  [31:0] io_dec_illegal_inst,
  input         io_dec_i0_decode_d,
  input         io_exu_i0_br_way_r,
  output        io_dec_dbg_cmd_done,
  output        io_dec_dbg_cmd_fail,
  output        io_dec_tlu_dbg_halted,
  output        io_dec_tlu_debug_mode,
  output        io_dec_tlu_resume_ack,
  output        io_dec_tlu_debug_stall,
  output        io_dec_tlu_mpc_halted_only,
  output        io_dec_tlu_flush_extint,
  input         io_dbg_halt_req,
  input         io_dbg_resume_req,
  input         io_dec_div_active,
  output        io_trigger_pkt_any_0_select,
  output        io_trigger_pkt_any_0_match_pkt,
  output        io_trigger_pkt_any_0_store,
  output        io_trigger_pkt_any_0_load,
  output        io_trigger_pkt_any_0_execute,
  output        io_trigger_pkt_any_0_m,
  output [31:0] io_trigger_pkt_any_0_tdata2,
  output        io_trigger_pkt_any_1_select,
  output        io_trigger_pkt_any_1_match_pkt,
  output        io_trigger_pkt_any_1_store,
  output        io_trigger_pkt_any_1_load,
  output        io_trigger_pkt_any_1_execute,
  output        io_trigger_pkt_any_1_m,
  output [31:0] io_trigger_pkt_any_1_tdata2,
  output        io_trigger_pkt_any_2_select,
  output        io_trigger_pkt_any_2_match_pkt,
  output        io_trigger_pkt_any_2_store,
  output        io_trigger_pkt_any_2_load,
  output        io_trigger_pkt_any_2_execute,
  output        io_trigger_pkt_any_2_m,
  output [31:0] io_trigger_pkt_any_2_tdata2,
  output        io_trigger_pkt_any_3_select,
  output        io_trigger_pkt_any_3_match_pkt,
  output        io_trigger_pkt_any_3_store,
  output        io_trigger_pkt_any_3_load,
  output        io_trigger_pkt_any_3_execute,
  output        io_trigger_pkt_any_3_m,
  output [31:0] io_trigger_pkt_any_3_tdata2,
  input         io_timer_int,
  input         io_soft_int,
  output        io_o_cpu_halt_status,
  output        io_o_cpu_halt_ack,
  output        io_o_cpu_run_ack,
  output        io_o_debug_mode_status,
  input  [27:0] io_core_id,
  input         io_mpc_debug_halt_req,
  input         io_mpc_debug_run_req,
  input         io_mpc_reset_run_req,
  output        io_mpc_debug_halt_ack,
  output        io_mpc_debug_run_ack,
  output        io_debug_brkpt_status,
  output [31:0] io_dec_csr_rddata_d,
  output        io_dec_csr_legal_d,
  output        io_dec_tlu_i0_kill_writeb_wb,
  output        io_dec_tlu_i0_kill_writeb_r,
  output        io_dec_tlu_wr_pause_r,
  output        io_dec_tlu_flush_pause_r,
  output        io_dec_tlu_presync_d,
  output        io_dec_tlu_postsync_d,
  output        io_dec_tlu_perfcnt0,
  output        io_dec_tlu_perfcnt1,
  output        io_dec_tlu_perfcnt2,
  output        io_dec_tlu_perfcnt3,
  output        io_dec_tlu_i0_exc_valid_wb1,
  output        io_dec_tlu_i0_valid_wb1,
  output        io_dec_tlu_int_valid_wb1,
  output [4:0]  io_dec_tlu_exc_cause_wb1,
  output [31:0] io_dec_tlu_mtval_wb1,
  output        io_dec_tlu_pipelining_disable,
  output        io_dec_tlu_misc_clk_override,
  output        io_dec_tlu_dec_clk_override,
  output        io_dec_tlu_lsu_clk_override,
  output        io_dec_tlu_bus_clk_override,
  output        io_dec_tlu_pic_clk_override,
  output        io_dec_tlu_dccm_clk_override,
  output        io_dec_tlu_icm_clk_override,
  output        io_dec_tlu_flush_lower_wb,
  input         io_ifu_pmu_instr_aligned,
  output        io_tlu_bp_dec_tlu_br0_r_pkt_valid,
  output [1:0]  io_tlu_bp_dec_tlu_br0_r_pkt_bits_hist,
  output        io_tlu_bp_dec_tlu_br0_r_pkt_bits_br_error,
  output        io_tlu_bp_dec_tlu_br0_r_pkt_bits_br_start_error,
  output        io_tlu_bp_dec_tlu_br0_r_pkt_bits_way,
  output        io_tlu_bp_dec_tlu_br0_r_pkt_bits_middle,
  output        io_tlu_bp_dec_tlu_flush_leak_one_wb,
  output        io_tlu_bp_dec_tlu_bpred_disable,
  output        io_tlu_ifc_dec_tlu_flush_noredir_wb,
  output [31:0] io_tlu_ifc_dec_tlu_mrac_ff,
  input         io_tlu_ifc_ifu_pmu_fetch_stall,
  output        io_tlu_mem_dec_tlu_flush_err_wb,
  output        io_tlu_mem_dec_tlu_i0_commit_cmt,
  output        io_tlu_mem_dec_tlu_force_halt,
  output        io_tlu_mem_dec_tlu_fence_i_wb,
  output [70:0] io_tlu_mem_dec_tlu_ic_diag_pkt_icache_wrdata,
  output [16:0] io_tlu_mem_dec_tlu_ic_diag_pkt_icache_dicawics,
  output        io_tlu_mem_dec_tlu_ic_diag_pkt_icache_rd_valid,
  output        io_tlu_mem_dec_tlu_ic_diag_pkt_icache_wr_valid,
  output        io_tlu_mem_dec_tlu_core_ecc_disable,
  input         io_tlu_mem_ifu_pmu_ic_miss,
  input         io_tlu_mem_ifu_pmu_ic_hit,
  input         io_tlu_mem_ifu_pmu_bus_error,
  input         io_tlu_mem_ifu_pmu_bus_busy,
  input         io_tlu_mem_ifu_ic_error_start,
  input         io_tlu_mem_ifu_iccm_rd_ecc_single_err,
  input  [70:0] io_tlu_mem_ifu_ic_debug_rd_data,
  input         io_tlu_mem_ifu_ic_debug_rd_data_valid,
  input         io_tlu_mem_ifu_miss_state_idle,
  input         io_tlu_busbuff_lsu_pmu_bus_misaligned,
  input         io_tlu_busbuff_lsu_pmu_bus_error,
  input         io_tlu_busbuff_lsu_pmu_bus_busy,
  output        io_tlu_busbuff_dec_tlu_external_ldfwd_disable,
  output        io_tlu_busbuff_dec_tlu_wb_coalescing_disable,
  output        io_tlu_busbuff_dec_tlu_sideeffect_posted_disable,
  input         io_tlu_busbuff_lsu_imprecise_error_load_any,
  input         io_tlu_busbuff_lsu_imprecise_error_store_any,
  input  [31:0] io_tlu_busbuff_lsu_imprecise_error_addr_any,
  input         io_lsu_tlu_lsu_pmu_load_external_m,
  input         io_lsu_tlu_lsu_pmu_store_external_m,
  input  [7:0]  io_dec_pic_pic_claimid,
  input  [3:0]  io_dec_pic_pic_pl,
  input         io_dec_pic_mhwakeup,
  output [3:0]  io_dec_pic_dec_tlu_meicurpl,
  output [3:0]  io_dec_pic_dec_tlu_meipt,
  input         io_dec_pic_mexintpend
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
`endif // RANDOMIZE_REG_INIT
  wire  int_timers_clock; // @[dec_tlu_ctl.scala 275:30]
  wire  int_timers_reset; // @[dec_tlu_ctl.scala 275:30]
  wire  int_timers_io_free_clk; // @[dec_tlu_ctl.scala 275:30]
  wire  int_timers_io_scan_mode; // @[dec_tlu_ctl.scala 275:30]
  wire  int_timers_io_dec_csr_wen_r_mod; // @[dec_tlu_ctl.scala 275:30]
  wire [11:0] int_timers_io_dec_csr_wraddr_r; // @[dec_tlu_ctl.scala 275:30]
  wire [31:0] int_timers_io_dec_csr_wrdata_r; // @[dec_tlu_ctl.scala 275:30]
  wire  int_timers_io_csr_mitctl0; // @[dec_tlu_ctl.scala 275:30]
  wire  int_timers_io_csr_mitctl1; // @[dec_tlu_ctl.scala 275:30]
  wire  int_timers_io_csr_mitb0; // @[dec_tlu_ctl.scala 275:30]
  wire  int_timers_io_csr_mitb1; // @[dec_tlu_ctl.scala 275:30]
  wire  int_timers_io_csr_mitcnt0; // @[dec_tlu_ctl.scala 275:30]
  wire  int_timers_io_csr_mitcnt1; // @[dec_tlu_ctl.scala 275:30]
  wire  int_timers_io_dec_pause_state; // @[dec_tlu_ctl.scala 275:30]
  wire  int_timers_io_dec_tlu_pmu_fw_halted; // @[dec_tlu_ctl.scala 275:30]
  wire  int_timers_io_internal_dbg_halt_timers; // @[dec_tlu_ctl.scala 275:30]
  wire [31:0] int_timers_io_dec_timer_rddata_d; // @[dec_tlu_ctl.scala 275:30]
  wire  int_timers_io_dec_timer_read_d; // @[dec_tlu_ctl.scala 275:30]
  wire  int_timers_io_dec_timer_t0_pulse; // @[dec_tlu_ctl.scala 275:30]
  wire  int_timers_io_dec_timer_t1_pulse; // @[dec_tlu_ctl.scala 275:30]
  wire  rvclkhdr_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_1_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_1_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_1_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_1_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_2_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_2_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_2_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_2_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_3_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_3_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_3_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_3_io_scan_mode; // @[lib.scala 343:22]
  wire  csr_clock; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_reset; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_free_clk; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_active_clk; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_scan_mode; // @[dec_tlu_ctl.scala 818:15]
  wire [31:0] csr_io_dec_csr_wrdata_r; // @[dec_tlu_ctl.scala 818:15]
  wire [11:0] csr_io_dec_csr_wraddr_r; // @[dec_tlu_ctl.scala 818:15]
  wire [11:0] csr_io_dec_csr_rdaddr_d; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_dec_csr_wen_unq_d; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_dec_i0_decode_d; // @[dec_tlu_ctl.scala 818:15]
  wire [70:0] csr_io_dec_tlu_ic_diag_pkt_icache_wrdata; // @[dec_tlu_ctl.scala 818:15]
  wire [16:0] csr_io_dec_tlu_ic_diag_pkt_icache_dicawics; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_dec_tlu_ic_diag_pkt_icache_rd_valid; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_dec_tlu_ic_diag_pkt_icache_wr_valid; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_ifu_ic_debug_rd_data_valid; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_trigger_pkt_any_0_select; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_trigger_pkt_any_0_match_pkt; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_trigger_pkt_any_0_store; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_trigger_pkt_any_0_load; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_trigger_pkt_any_0_execute; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_trigger_pkt_any_0_m; // @[dec_tlu_ctl.scala 818:15]
  wire [31:0] csr_io_trigger_pkt_any_0_tdata2; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_trigger_pkt_any_1_select; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_trigger_pkt_any_1_match_pkt; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_trigger_pkt_any_1_store; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_trigger_pkt_any_1_load; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_trigger_pkt_any_1_execute; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_trigger_pkt_any_1_m; // @[dec_tlu_ctl.scala 818:15]
  wire [31:0] csr_io_trigger_pkt_any_1_tdata2; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_trigger_pkt_any_2_select; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_trigger_pkt_any_2_match_pkt; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_trigger_pkt_any_2_store; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_trigger_pkt_any_2_load; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_trigger_pkt_any_2_execute; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_trigger_pkt_any_2_m; // @[dec_tlu_ctl.scala 818:15]
  wire [31:0] csr_io_trigger_pkt_any_2_tdata2; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_trigger_pkt_any_3_select; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_trigger_pkt_any_3_match_pkt; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_trigger_pkt_any_3_store; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_trigger_pkt_any_3_load; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_trigger_pkt_any_3_execute; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_trigger_pkt_any_3_m; // @[dec_tlu_ctl.scala 818:15]
  wire [31:0] csr_io_trigger_pkt_any_3_tdata2; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_dma_iccm_stall_any; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_dma_dccm_stall_any; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_lsu_store_stall_any; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_dec_pmu_presync_stall; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_dec_pmu_postsync_stall; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_dec_pmu_decode_stall; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_ifu_pmu_fetch_stall; // @[dec_tlu_ctl.scala 818:15]
  wire [1:0] csr_io_dec_tlu_packet_r_icaf_type; // @[dec_tlu_ctl.scala 818:15]
  wire [3:0] csr_io_dec_tlu_packet_r_pmu_i0_itype; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_dec_tlu_packet_r_pmu_i0_br_unpred; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_dec_tlu_packet_r_pmu_divide; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_dec_tlu_packet_r_pmu_lsu_misaligned; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_exu_pmu_i0_br_ataken; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_exu_pmu_i0_br_misp; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_dec_pmu_instr_decoded; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_ifu_pmu_instr_aligned; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_exu_pmu_i0_pc4; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_ifu_pmu_ic_miss; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_ifu_pmu_ic_hit; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_dec_tlu_int_valid_wb1; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_dec_tlu_i0_exc_valid_wb1; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_dec_tlu_i0_valid_wb1; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_dec_csr_wen_r; // @[dec_tlu_ctl.scala 818:15]
  wire [31:0] csr_io_dec_tlu_mtval_wb1; // @[dec_tlu_ctl.scala 818:15]
  wire [4:0] csr_io_dec_tlu_exc_cause_wb1; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_dec_tlu_perfcnt0; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_dec_tlu_perfcnt1; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_dec_tlu_perfcnt2; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_dec_tlu_perfcnt3; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_dec_tlu_dbg_halted; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_dma_pmu_dccm_write; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_dma_pmu_dccm_read; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_dma_pmu_any_write; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_dma_pmu_any_read; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_lsu_pmu_bus_busy; // @[dec_tlu_ctl.scala 818:15]
  wire [30:0] csr_io_dec_tlu_i0_pc_r; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_dec_tlu_i0_valid_r; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_dec_csr_any_unq_d; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_dec_tlu_misc_clk_override; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_dec_tlu_dec_clk_override; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_dec_tlu_lsu_clk_override; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_dec_tlu_bus_clk_override; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_dec_tlu_pic_clk_override; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_dec_tlu_dccm_clk_override; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_dec_tlu_icm_clk_override; // @[dec_tlu_ctl.scala 818:15]
  wire [31:0] csr_io_dec_csr_rddata_d; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_dec_tlu_pipelining_disable; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_dec_tlu_wr_pause_r; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_ifu_pmu_bus_busy; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_lsu_pmu_bus_error; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_ifu_pmu_bus_error; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_lsu_pmu_bus_misaligned; // @[dec_tlu_ctl.scala 818:15]
  wire [70:0] csr_io_ifu_ic_debug_rd_data; // @[dec_tlu_ctl.scala 818:15]
  wire [3:0] csr_io_dec_tlu_meipt; // @[dec_tlu_ctl.scala 818:15]
  wire [3:0] csr_io_pic_pl; // @[dec_tlu_ctl.scala 818:15]
  wire [3:0] csr_io_dec_tlu_meicurpl; // @[dec_tlu_ctl.scala 818:15]
  wire [29:0] csr_io_dec_tlu_meihap; // @[dec_tlu_ctl.scala 818:15]
  wire [7:0] csr_io_pic_claimid; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_iccm_dma_sb_error; // @[dec_tlu_ctl.scala 818:15]
  wire [31:0] csr_io_lsu_imprecise_error_addr_any; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_lsu_imprecise_error_load_any; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_lsu_imprecise_error_store_any; // @[dec_tlu_ctl.scala 818:15]
  wire [31:0] csr_io_dec_tlu_mrac_ff; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_dec_tlu_wb_coalescing_disable; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_dec_tlu_bpred_disable; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_dec_tlu_sideeffect_posted_disable; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_dec_tlu_core_ecc_disable; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_dec_tlu_external_ldfwd_disable; // @[dec_tlu_ctl.scala 818:15]
  wire [2:0] csr_io_dec_tlu_dma_qos_prty; // @[dec_tlu_ctl.scala 818:15]
  wire [31:0] csr_io_dec_illegal_inst; // @[dec_tlu_ctl.scala 818:15]
  wire [3:0] csr_io_lsu_error_pkt_r_bits_mscause; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_mexintpend; // @[dec_tlu_ctl.scala 818:15]
  wire [30:0] csr_io_exu_npc_r; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_mpc_reset_run_req; // @[dec_tlu_ctl.scala 818:15]
  wire [30:0] csr_io_rst_vec; // @[dec_tlu_ctl.scala 818:15]
  wire [27:0] csr_io_core_id; // @[dec_tlu_ctl.scala 818:15]
  wire [31:0] csr_io_dec_timer_rddata_d; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_dec_timer_read_d; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_dec_csr_wen_r_mod; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_rfpc_i0_r; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_i0_trigger_hit_r; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_fw_halt_req; // @[dec_tlu_ctl.scala 818:15]
  wire [1:0] csr_io_mstatus; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_exc_or_int_valid_r; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_mret_r; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_mstatus_mie_ns; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_dcsr_single_step_running_f; // @[dec_tlu_ctl.scala 818:15]
  wire [15:0] csr_io_dcsr; // @[dec_tlu_ctl.scala 818:15]
  wire [30:0] csr_io_mtvec; // @[dec_tlu_ctl.scala 818:15]
  wire [5:0] csr_io_mip; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_dec_timer_t0_pulse; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_dec_timer_t1_pulse; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_timer_int_sync; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_soft_int_sync; // @[dec_tlu_ctl.scala 818:15]
  wire [5:0] csr_io_mie_ns; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_csr_wr_clk; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_ebreak_to_debug_mode_r; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_dec_tlu_pmu_fw_halted; // @[dec_tlu_ctl.scala 818:15]
  wire [1:0] csr_io_lsu_fir_error; // @[dec_tlu_ctl.scala 818:15]
  wire [30:0] csr_io_npc_r; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_tlu_flush_lower_r_d1; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_dec_tlu_flush_noredir_r_d1; // @[dec_tlu_ctl.scala 818:15]
  wire [30:0] csr_io_tlu_flush_path_r_d1; // @[dec_tlu_ctl.scala 818:15]
  wire [30:0] csr_io_npc_r_d1; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_reset_delayed; // @[dec_tlu_ctl.scala 818:15]
  wire [30:0] csr_io_mepc; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_interrupt_valid_r; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_i0_exception_valid_r; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_lsu_exc_valid_r; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_mepc_trigger_hit_sel_pc_r; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_e4e5_int_clk; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_lsu_i0_exc_r; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_inst_acc_r; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_inst_acc_second_r; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_take_nmi; // @[dec_tlu_ctl.scala 818:15]
  wire [31:0] csr_io_lsu_error_pkt_addr_r; // @[dec_tlu_ctl.scala 818:15]
  wire [4:0] csr_io_exc_cause_r; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_i0_valid_wb; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_exc_or_int_valid_r_d1; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_interrupt_valid_r_d1; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_clk_override; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_i0_exception_valid_r_d1; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_lsu_i0_exc_r_d1; // @[dec_tlu_ctl.scala 818:15]
  wire [4:0] csr_io_exc_cause_wb; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_nmi_lsu_store_type; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_nmi_lsu_load_type; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_tlu_i0_commit_cmt; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_ebreak_r; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_ecall_r; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_illegal_r; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_mdseac_locked_ns; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_mdseac_locked_f; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_nmi_int_detected_f; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_internal_dbg_halt_mode_f2; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_ext_int_freeze_d1; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_ic_perr_r_d1; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_iccm_sbecc_r_d1; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_lsu_single_ecc_error_r_d1; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_ifu_miss_state_idle_f; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_lsu_idle_any_f; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_dbg_tlu_halted_f; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_dbg_tlu_halted; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_debug_halt_req_f; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_force_halt; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_take_ext_int_start; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_trigger_hit_dmode_r_d1; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_trigger_hit_r_d1; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_dcsr_single_step_done_f; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_ebreak_to_debug_mode_r_d1; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_debug_halt_req; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_allow_dbg_halt_csr_write; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_internal_dbg_halt_mode_f; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_enter_debug_halt_req; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_internal_dbg_halt_mode; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_request_debug_mode_done; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_request_debug_mode_r; // @[dec_tlu_ctl.scala 818:15]
  wire [30:0] csr_io_dpc; // @[dec_tlu_ctl.scala 818:15]
  wire [3:0] csr_io_update_hit_bit_r; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_take_timer_int; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_take_int_timer0_int; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_take_int_timer1_int; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_take_ext_int; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_tlu_flush_lower_r; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_dec_tlu_br0_error_r; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_dec_tlu_br0_start_error_r; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_lsu_pmu_load_external_r; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_lsu_pmu_store_external_r; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_csr_pkt_csr_misa; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_csr_pkt_csr_mvendorid; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_csr_pkt_csr_marchid; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_csr_pkt_csr_mimpid; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_csr_pkt_csr_mhartid; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_csr_pkt_csr_mstatus; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_csr_pkt_csr_mtvec; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_csr_pkt_csr_mip; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_csr_pkt_csr_mie; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_csr_pkt_csr_mcyclel; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_csr_pkt_csr_mcycleh; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_csr_pkt_csr_minstretl; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_csr_pkt_csr_minstreth; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_csr_pkt_csr_mscratch; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_csr_pkt_csr_mepc; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_csr_pkt_csr_mcause; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_csr_pkt_csr_mscause; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_csr_pkt_csr_mtval; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_csr_pkt_csr_mrac; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_csr_pkt_csr_mdseac; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_csr_pkt_csr_meihap; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_csr_pkt_csr_meivt; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_csr_pkt_csr_meipt; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_csr_pkt_csr_meicurpl; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_csr_pkt_csr_meicidpl; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_csr_pkt_csr_dcsr; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_csr_pkt_csr_mcgc; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_csr_pkt_csr_mfdc; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_csr_pkt_csr_dpc; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_csr_pkt_csr_mtsel; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_csr_pkt_csr_mtdata1; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_csr_pkt_csr_mtdata2; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_csr_pkt_csr_mhpmc3; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_csr_pkt_csr_mhpmc4; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_csr_pkt_csr_mhpmc5; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_csr_pkt_csr_mhpmc6; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_csr_pkt_csr_mhpmc3h; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_csr_pkt_csr_mhpmc4h; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_csr_pkt_csr_mhpmc5h; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_csr_pkt_csr_mhpmc6h; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_csr_pkt_csr_mhpme3; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_csr_pkt_csr_mhpme4; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_csr_pkt_csr_mhpme5; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_csr_pkt_csr_mhpme6; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_csr_pkt_csr_mcountinhibit; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_csr_pkt_csr_mpmc; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_csr_pkt_csr_micect; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_csr_pkt_csr_miccmect; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_csr_pkt_csr_mdccmect; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_csr_pkt_csr_mfdht; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_csr_pkt_csr_mfdhs; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_csr_pkt_csr_dicawics; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_csr_pkt_csr_dicad0h; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_csr_pkt_csr_dicad0; // @[dec_tlu_ctl.scala 818:15]
  wire  csr_io_csr_pkt_csr_dicad1; // @[dec_tlu_ctl.scala 818:15]
  wire [9:0] csr_io_mtdata1_t_0; // @[dec_tlu_ctl.scala 818:15]
  wire [9:0] csr_io_mtdata1_t_1; // @[dec_tlu_ctl.scala 818:15]
  wire [9:0] csr_io_mtdata1_t_2; // @[dec_tlu_ctl.scala 818:15]
  wire [9:0] csr_io_mtdata1_t_3; // @[dec_tlu_ctl.scala 818:15]
  wire [11:0] csr_read_io_dec_csr_rdaddr_d; // @[dec_tlu_ctl.scala 1011:22]
  wire  csr_read_io_csr_pkt_csr_misa; // @[dec_tlu_ctl.scala 1011:22]
  wire  csr_read_io_csr_pkt_csr_mvendorid; // @[dec_tlu_ctl.scala 1011:22]
  wire  csr_read_io_csr_pkt_csr_marchid; // @[dec_tlu_ctl.scala 1011:22]
  wire  csr_read_io_csr_pkt_csr_mimpid; // @[dec_tlu_ctl.scala 1011:22]
  wire  csr_read_io_csr_pkt_csr_mhartid; // @[dec_tlu_ctl.scala 1011:22]
  wire  csr_read_io_csr_pkt_csr_mstatus; // @[dec_tlu_ctl.scala 1011:22]
  wire  csr_read_io_csr_pkt_csr_mtvec; // @[dec_tlu_ctl.scala 1011:22]
  wire  csr_read_io_csr_pkt_csr_mip; // @[dec_tlu_ctl.scala 1011:22]
  wire  csr_read_io_csr_pkt_csr_mie; // @[dec_tlu_ctl.scala 1011:22]
  wire  csr_read_io_csr_pkt_csr_mcyclel; // @[dec_tlu_ctl.scala 1011:22]
  wire  csr_read_io_csr_pkt_csr_mcycleh; // @[dec_tlu_ctl.scala 1011:22]
  wire  csr_read_io_csr_pkt_csr_minstretl; // @[dec_tlu_ctl.scala 1011:22]
  wire  csr_read_io_csr_pkt_csr_minstreth; // @[dec_tlu_ctl.scala 1011:22]
  wire  csr_read_io_csr_pkt_csr_mscratch; // @[dec_tlu_ctl.scala 1011:22]
  wire  csr_read_io_csr_pkt_csr_mepc; // @[dec_tlu_ctl.scala 1011:22]
  wire  csr_read_io_csr_pkt_csr_mcause; // @[dec_tlu_ctl.scala 1011:22]
  wire  csr_read_io_csr_pkt_csr_mscause; // @[dec_tlu_ctl.scala 1011:22]
  wire  csr_read_io_csr_pkt_csr_mtval; // @[dec_tlu_ctl.scala 1011:22]
  wire  csr_read_io_csr_pkt_csr_mrac; // @[dec_tlu_ctl.scala 1011:22]
  wire  csr_read_io_csr_pkt_csr_dmst; // @[dec_tlu_ctl.scala 1011:22]
  wire  csr_read_io_csr_pkt_csr_mdseac; // @[dec_tlu_ctl.scala 1011:22]
  wire  csr_read_io_csr_pkt_csr_meihap; // @[dec_tlu_ctl.scala 1011:22]
  wire  csr_read_io_csr_pkt_csr_meivt; // @[dec_tlu_ctl.scala 1011:22]
  wire  csr_read_io_csr_pkt_csr_meipt; // @[dec_tlu_ctl.scala 1011:22]
  wire  csr_read_io_csr_pkt_csr_meicurpl; // @[dec_tlu_ctl.scala 1011:22]
  wire  csr_read_io_csr_pkt_csr_meicidpl; // @[dec_tlu_ctl.scala 1011:22]
  wire  csr_read_io_csr_pkt_csr_dcsr; // @[dec_tlu_ctl.scala 1011:22]
  wire  csr_read_io_csr_pkt_csr_mcgc; // @[dec_tlu_ctl.scala 1011:22]
  wire  csr_read_io_csr_pkt_csr_mfdc; // @[dec_tlu_ctl.scala 1011:22]
  wire  csr_read_io_csr_pkt_csr_dpc; // @[dec_tlu_ctl.scala 1011:22]
  wire  csr_read_io_csr_pkt_csr_mtsel; // @[dec_tlu_ctl.scala 1011:22]
  wire  csr_read_io_csr_pkt_csr_mtdata1; // @[dec_tlu_ctl.scala 1011:22]
  wire  csr_read_io_csr_pkt_csr_mtdata2; // @[dec_tlu_ctl.scala 1011:22]
  wire  csr_read_io_csr_pkt_csr_mhpmc3; // @[dec_tlu_ctl.scala 1011:22]
  wire  csr_read_io_csr_pkt_csr_mhpmc4; // @[dec_tlu_ctl.scala 1011:22]
  wire  csr_read_io_csr_pkt_csr_mhpmc5; // @[dec_tlu_ctl.scala 1011:22]
  wire  csr_read_io_csr_pkt_csr_mhpmc6; // @[dec_tlu_ctl.scala 1011:22]
  wire  csr_read_io_csr_pkt_csr_mhpmc3h; // @[dec_tlu_ctl.scala 1011:22]
  wire  csr_read_io_csr_pkt_csr_mhpmc4h; // @[dec_tlu_ctl.scala 1011:22]
  wire  csr_read_io_csr_pkt_csr_mhpmc5h; // @[dec_tlu_ctl.scala 1011:22]
  wire  csr_read_io_csr_pkt_csr_mhpmc6h; // @[dec_tlu_ctl.scala 1011:22]
  wire  csr_read_io_csr_pkt_csr_mhpme3; // @[dec_tlu_ctl.scala 1011:22]
  wire  csr_read_io_csr_pkt_csr_mhpme4; // @[dec_tlu_ctl.scala 1011:22]
  wire  csr_read_io_csr_pkt_csr_mhpme5; // @[dec_tlu_ctl.scala 1011:22]
  wire  csr_read_io_csr_pkt_csr_mhpme6; // @[dec_tlu_ctl.scala 1011:22]
  wire  csr_read_io_csr_pkt_csr_mcountinhibit; // @[dec_tlu_ctl.scala 1011:22]
  wire  csr_read_io_csr_pkt_csr_mitctl0; // @[dec_tlu_ctl.scala 1011:22]
  wire  csr_read_io_csr_pkt_csr_mitctl1; // @[dec_tlu_ctl.scala 1011:22]
  wire  csr_read_io_csr_pkt_csr_mitb0; // @[dec_tlu_ctl.scala 1011:22]
  wire  csr_read_io_csr_pkt_csr_mitb1; // @[dec_tlu_ctl.scala 1011:22]
  wire  csr_read_io_csr_pkt_csr_mitcnt0; // @[dec_tlu_ctl.scala 1011:22]
  wire  csr_read_io_csr_pkt_csr_mitcnt1; // @[dec_tlu_ctl.scala 1011:22]
  wire  csr_read_io_csr_pkt_csr_mpmc; // @[dec_tlu_ctl.scala 1011:22]
  wire  csr_read_io_csr_pkt_csr_meicpct; // @[dec_tlu_ctl.scala 1011:22]
  wire  csr_read_io_csr_pkt_csr_micect; // @[dec_tlu_ctl.scala 1011:22]
  wire  csr_read_io_csr_pkt_csr_miccmect; // @[dec_tlu_ctl.scala 1011:22]
  wire  csr_read_io_csr_pkt_csr_mdccmect; // @[dec_tlu_ctl.scala 1011:22]
  wire  csr_read_io_csr_pkt_csr_mfdht; // @[dec_tlu_ctl.scala 1011:22]
  wire  csr_read_io_csr_pkt_csr_mfdhs; // @[dec_tlu_ctl.scala 1011:22]
  wire  csr_read_io_csr_pkt_csr_dicawics; // @[dec_tlu_ctl.scala 1011:22]
  wire  csr_read_io_csr_pkt_csr_dicad0h; // @[dec_tlu_ctl.scala 1011:22]
  wire  csr_read_io_csr_pkt_csr_dicad0; // @[dec_tlu_ctl.scala 1011:22]
  wire  csr_read_io_csr_pkt_csr_dicad1; // @[dec_tlu_ctl.scala 1011:22]
  wire  csr_read_io_csr_pkt_csr_dicago; // @[dec_tlu_ctl.scala 1011:22]
  wire  csr_read_io_csr_pkt_presync; // @[dec_tlu_ctl.scala 1011:22]
  wire  csr_read_io_csr_pkt_postsync; // @[dec_tlu_ctl.scala 1011:22]
  wire  csr_read_io_csr_pkt_legal; // @[dec_tlu_ctl.scala 1011:22]
  reg  dbg_halt_state_f; // @[dec_tlu_ctl.scala 367:89]
  wire  _T = ~dbg_halt_state_f; // @[dec_tlu_ctl.scala 274:39]
  reg  mpc_halt_state_f; // @[dec_tlu_ctl.scala 362:89]
  wire [2:0] _T_3 = {io_i_cpu_run_req,io_mpc_debug_halt_req,io_mpc_debug_run_req}; // @[Cat.scala 29:58]
  wire [3:0] _T_6 = {io_nmi_int,io_timer_int,io_soft_int,io_i_cpu_halt_req}; // @[Cat.scala 29:58]
  reg [6:0] _T_8; // @[lib.scala 37:81]
  reg [6:0] syncro_ff; // @[lib.scala 37:58]
  wire  nmi_int_sync = syncro_ff[6]; // @[dec_tlu_ctl.scala 302:67]
  wire  i_cpu_halt_req_sync = syncro_ff[3]; // @[dec_tlu_ctl.scala 305:59]
  wire  i_cpu_run_req_sync = syncro_ff[2]; // @[dec_tlu_ctl.scala 306:59]
  wire  mpc_debug_halt_req_sync_raw = syncro_ff[1]; // @[dec_tlu_ctl.scala 307:51]
  wire  mpc_debug_run_req_sync = syncro_ff[0]; // @[dec_tlu_ctl.scala 308:51]
  wire  dec_csr_wen_r_mod = csr_io_dec_csr_wen_r_mod; // @[dec_tlu_ctl.scala 1004:31]
  reg  lsu_exc_valid_r_d1; // @[dec_tlu_ctl.scala 613:74]
  wire  _T_11 = io_lsu_error_pkt_r_valid | lsu_exc_valid_r_d1; // @[dec_tlu_ctl.scala 312:67]
  reg  e5_valid; // @[dec_tlu_ctl.scala 324:97]
  wire  e4e5_valid = io_dec_tlu_i0_valid_r | e5_valid; // @[dec_tlu_ctl.scala 315:30]
  reg  debug_mode_status; // @[dec_tlu_ctl.scala 325:81]
  reg  i_cpu_run_req_d1_raw; // @[dec_tlu_ctl.scala 573:80]
  reg  nmi_int_delayed; // @[dec_tlu_ctl.scala 340:72]
  wire  _T_37 = ~nmi_int_delayed; // @[dec_tlu_ctl.scala 349:45]
  wire  _T_38 = nmi_int_sync & _T_37; // @[dec_tlu_ctl.scala 349:43]
  reg  mdseac_locked_f; // @[dec_tlu_ctl.scala 606:89]
  wire  _T_35 = ~mdseac_locked_f; // @[dec_tlu_ctl.scala 347:32]
  wire  _T_36 = io_tlu_busbuff_lsu_imprecise_error_load_any | io_tlu_busbuff_lsu_imprecise_error_store_any; // @[dec_tlu_ctl.scala 347:96]
  wire  nmi_lsu_detected = _T_35 & _T_36; // @[dec_tlu_ctl.scala 347:49]
  wire  _T_39 = _T_38 | nmi_lsu_detected; // @[dec_tlu_ctl.scala 349:63]
  reg  nmi_int_detected_f; // @[dec_tlu_ctl.scala 341:72]
  reg  take_nmi_r_d1; // @[dec_tlu_ctl.scala 815:98]
  wire  _T_40 = ~take_nmi_r_d1; // @[dec_tlu_ctl.scala 349:106]
  wire  _T_41 = nmi_int_detected_f & _T_40; // @[dec_tlu_ctl.scala 349:104]
  wire  _T_42 = _T_39 | _T_41; // @[dec_tlu_ctl.scala 349:82]
  reg  take_ext_int_start_d3; // @[dec_tlu_ctl.scala 746:62]
  wire  _T_43 = |io_lsu_fir_error; // @[dec_tlu_ctl.scala 349:165]
  wire  _T_44 = take_ext_int_start_d3 & _T_43; // @[dec_tlu_ctl.scala 349:146]
  wire  nmi_int_detected = _T_42 | _T_44; // @[dec_tlu_ctl.scala 349:122]
  wire  _T_631 = ~io_dec_csr_stall_int_ff; // @[dec_tlu_ctl.scala 723:23]
  wire  mstatus_mie_ns = csr_io_mstatus_mie_ns; // @[dec_tlu_ctl.scala 1003:31]
  wire  _T_632 = _T_631 & mstatus_mie_ns; // @[dec_tlu_ctl.scala 723:48]
  wire [5:0] mip = csr_io_mip; // @[dec_tlu_ctl.scala 1009:31]
  wire  _T_634 = _T_632 & mip[1]; // @[dec_tlu_ctl.scala 723:65]
  wire [5:0] mie_ns = csr_io_mie_ns; // @[dec_tlu_ctl.scala 998:31]
  wire  timer_int_ready = _T_634 & mie_ns[1]; // @[dec_tlu_ctl.scala 723:83]
  wire  _T_391 = nmi_int_detected | timer_int_ready; // @[dec_tlu_ctl.scala 600:66]
  wire  _T_628 = _T_632 & mip[0]; // @[dec_tlu_ctl.scala 722:65]
  wire  soft_int_ready = _T_628 & mie_ns[0]; // @[dec_tlu_ctl.scala 722:83]
  wire  _T_392 = _T_391 | soft_int_ready; // @[dec_tlu_ctl.scala 600:84]
  reg  int_timer0_int_hold_f; // @[dec_tlu_ctl.scala 580:73]
  wire  _T_393 = _T_392 | int_timer0_int_hold_f; // @[dec_tlu_ctl.scala 600:101]
  reg  int_timer1_int_hold_f; // @[dec_tlu_ctl.scala 581:73]
  wire  _T_394 = _T_393 | int_timer1_int_hold_f; // @[dec_tlu_ctl.scala 600:125]
  wire  _T_608 = _T_632 & mip[2]; // @[dec_tlu_ctl.scala 719:66]
  wire  mhwakeup_ready = _T_608 & mie_ns[2]; // @[dec_tlu_ctl.scala 719:84]
  wire  _T_395 = io_dec_pic_mhwakeup & mhwakeup_ready; // @[dec_tlu_ctl.scala 600:172]
  wire  _T_396 = _T_394 | _T_395; // @[dec_tlu_ctl.scala 600:149]
  wire  _T_397 = _T_396 & io_o_cpu_halt_status; // @[dec_tlu_ctl.scala 600:191]
  reg  i_cpu_halt_req_d1; // @[dec_tlu_ctl.scala 572:80]
  wire  _T_398 = ~i_cpu_halt_req_d1; // @[dec_tlu_ctl.scala 600:216]
  wire  _T_399 = _T_397 & _T_398; // @[dec_tlu_ctl.scala 600:214]
  wire  i_cpu_run_req_d1 = i_cpu_run_req_d1_raw | _T_399; // @[dec_tlu_ctl.scala 600:45]
  wire  _T_14 = debug_mode_status | i_cpu_run_req_d1; // @[dec_tlu_ctl.scala 316:50]
  wire  _T_685 = ~_T_43; // @[dec_tlu_ctl.scala 751:49]
  wire  take_ext_int = take_ext_int_start_d3 & _T_685; // @[dec_tlu_ctl.scala 751:47]
  wire  _T_698 = ~soft_int_ready; // @[dec_tlu_ctl.scala 768:40]
  wire  _T_699 = timer_int_ready & _T_698; // @[dec_tlu_ctl.scala 768:38]
  wire  _T_617 = ~io_lsu_fastint_stall_any; // @[dec_tlu_ctl.scala 720:104]
  wire  ext_int_ready = mhwakeup_ready & _T_617; // @[dec_tlu_ctl.scala 720:102]
  wire  _T_700 = ~ext_int_ready; // @[dec_tlu_ctl.scala 768:58]
  wire  _T_701 = _T_699 & _T_700; // @[dec_tlu_ctl.scala 768:56]
  wire  _T_622 = _T_632 & mip[5]; // @[dec_tlu_ctl.scala 721:65]
  wire  ce_int_ready = _T_622 & mie_ns[5]; // @[dec_tlu_ctl.scala 721:83]
  wire  _T_702 = ~ce_int_ready; // @[dec_tlu_ctl.scala 768:75]
  wire  _T_703 = _T_701 & _T_702; // @[dec_tlu_ctl.scala 768:73]
  wire  _T_152 = ~debug_mode_status; // @[dec_tlu_ctl.scala 423:37]
  reg  dbg_halt_req_held; // @[dec_tlu_ctl.scala 466:81]
  wire  _T_106 = io_dbg_halt_req | dbg_halt_req_held; // @[dec_tlu_ctl.scala 400:48]
  reg  ext_int_freeze_d1; // @[dec_tlu_ctl.scala 747:66]
  wire  _T_107 = ~ext_int_freeze_d1; // @[dec_tlu_ctl.scala 400:71]
  wire  dbg_halt_req_final = _T_106 & _T_107; // @[dec_tlu_ctl.scala 400:69]
  wire  mpc_debug_halt_req_sync = mpc_debug_halt_req_sync_raw & _T_107; // @[dec_tlu_ctl.scala 359:67]
  wire  _T_109 = dbg_halt_req_final | mpc_debug_halt_req_sync; // @[dec_tlu_ctl.scala 403:50]
  reg  reset_detect; // @[dec_tlu_ctl.scala 336:88]
  reg  reset_detected; // @[dec_tlu_ctl.scala 337:88]
  wire  reset_delayed = reset_detect ^ reset_detected; // @[dec_tlu_ctl.scala 338:64]
  wire  _T_110 = ~io_mpc_reset_run_req; // @[dec_tlu_ctl.scala 403:95]
  wire  _T_111 = reset_delayed & _T_110; // @[dec_tlu_ctl.scala 403:93]
  wire  _T_112 = _T_109 | _T_111; // @[dec_tlu_ctl.scala 403:76]
  wire  _T_114 = _T_112 & _T_152; // @[dec_tlu_ctl.scala 403:119]
  wire  debug_halt_req = _T_114 & _T_107; // @[dec_tlu_ctl.scala 403:147]
  wire  _T_153 = _T_152 & debug_halt_req; // @[dec_tlu_ctl.scala 423:63]
  reg  dcsr_single_step_done_f; // @[dec_tlu_ctl.scala 458:81]
  wire  _T_154 = _T_153 | dcsr_single_step_done_f; // @[dec_tlu_ctl.scala 423:81]
  reg  trigger_hit_dmode_r_d1; // @[dec_tlu_ctl.scala 457:81]
  wire  _T_155 = _T_154 | trigger_hit_dmode_r_d1; // @[dec_tlu_ctl.scala 423:107]
  reg  ebreak_to_debug_mode_r_d1; // @[dec_tlu_ctl.scala 672:64]
  wire  enter_debug_halt_req = _T_155 | ebreak_to_debug_mode_r_d1; // @[dec_tlu_ctl.scala 423:132]
  reg  debug_halt_req_f; // @[dec_tlu_ctl.scala 455:89]
  wire  force_halt = csr_io_force_halt; // @[dec_tlu_ctl.scala 1001:31]
  reg  lsu_idle_any_f; // @[dec_tlu_ctl.scala 451:89]
  wire  _T_142 = io_lsu_idle_any & lsu_idle_any_f; // @[dec_tlu_ctl.scala 417:53]
  wire  _T_143 = _T_142 & io_tlu_mem_ifu_miss_state_idle; // @[dec_tlu_ctl.scala 417:70]
  reg  ifu_miss_state_idle_f; // @[dec_tlu_ctl.scala 452:81]
  wire  _T_144 = _T_143 & ifu_miss_state_idle_f; // @[dec_tlu_ctl.scala 417:103]
  wire  _T_145 = ~debug_halt_req; // @[dec_tlu_ctl.scala 417:129]
  wire  _T_146 = _T_144 & _T_145; // @[dec_tlu_ctl.scala 417:127]
  reg  debug_halt_req_d1; // @[dec_tlu_ctl.scala 459:89]
  wire  _T_147 = ~debug_halt_req_d1; // @[dec_tlu_ctl.scala 417:147]
  wire  _T_148 = _T_146 & _T_147; // @[dec_tlu_ctl.scala 417:145]
  wire  _T_149 = ~io_dec_div_active; // @[dec_tlu_ctl.scala 417:168]
  wire  _T_150 = _T_148 & _T_149; // @[dec_tlu_ctl.scala 417:166]
  wire  core_empty = force_halt | _T_150; // @[dec_tlu_ctl.scala 417:34]
  wire  _T_163 = debug_halt_req_f & core_empty; // @[dec_tlu_ctl.scala 433:48]
  reg  dec_tlu_flush_noredir_r_d1; // @[dec_tlu_ctl.scala 449:81]
  reg  dec_tlu_flush_pause_r_d1; // @[dec_tlu_ctl.scala 465:73]
  wire  _T_132 = ~dec_tlu_flush_pause_r_d1; // @[dec_tlu_ctl.scala 413:56]
  wire  _T_133 = dec_tlu_flush_noredir_r_d1 & _T_132; // @[dec_tlu_ctl.scala 413:54]
  reg  take_ext_int_start_d1; // @[dec_tlu_ctl.scala 744:62]
  wire  _T_134 = ~take_ext_int_start_d1; // @[dec_tlu_ctl.scala 413:84]
  wire  _T_135 = _T_133 & _T_134; // @[dec_tlu_ctl.scala 413:82]
  reg  halt_taken_f; // @[dec_tlu_ctl.scala 450:89]
  reg  dbg_tlu_halted_f; // @[dec_tlu_ctl.scala 453:89]
  wire  _T_136 = ~dbg_tlu_halted_f; // @[dec_tlu_ctl.scala 413:126]
  wire  _T_137 = halt_taken_f & _T_136; // @[dec_tlu_ctl.scala 413:124]
  reg  pmu_fw_tlu_halted_f; // @[dec_tlu_ctl.scala 579:73]
  wire  _T_138 = ~pmu_fw_tlu_halted_f; // @[dec_tlu_ctl.scala 413:146]
  wire  _T_139 = _T_137 & _T_138; // @[dec_tlu_ctl.scala 413:144]
  reg  interrupt_valid_r_d1; // @[dec_tlu_ctl.scala 809:90]
  wire  _T_140 = ~interrupt_valid_r_d1; // @[dec_tlu_ctl.scala 413:169]
  wire  _T_141 = _T_139 & _T_140; // @[dec_tlu_ctl.scala 413:167]
  wire  halt_taken = _T_135 | _T_141; // @[dec_tlu_ctl.scala 413:108]
  wire  _T_164 = _T_163 & halt_taken; // @[dec_tlu_ctl.scala 433:61]
  reg  debug_resume_req_f; // @[dec_tlu_ctl.scala 456:89]
  wire  _T_165 = ~debug_resume_req_f; // @[dec_tlu_ctl.scala 433:97]
  wire  _T_166 = dbg_tlu_halted_f & _T_165; // @[dec_tlu_ctl.scala 433:95]
  wire  dbg_tlu_halted = _T_164 | _T_166; // @[dec_tlu_ctl.scala 433:75]
  wire  _T_167 = ~dbg_tlu_halted; // @[dec_tlu_ctl.scala 434:73]
  wire  _T_168 = debug_halt_req_f & _T_167; // @[dec_tlu_ctl.scala 434:71]
  wire  debug_halt_req_ns = enter_debug_halt_req | _T_168; // @[dec_tlu_ctl.scala 434:51]
  wire [15:0] dcsr = csr_io_dcsr; // @[dec_tlu_ctl.scala 1007:31]
  wire  _T_157 = ~dcsr[2]; // @[dec_tlu_ctl.scala 426:106]
  wire  _T_158 = debug_resume_req_f & _T_157; // @[dec_tlu_ctl.scala 426:104]
  wire  _T_159 = ~_T_158; // @[dec_tlu_ctl.scala 426:83]
  wire  _T_160 = debug_mode_status & _T_159; // @[dec_tlu_ctl.scala 426:81]
  wire  internal_dbg_halt_mode = debug_halt_req_ns | _T_160; // @[dec_tlu_ctl.scala 426:53]
  wire  _T_177 = debug_resume_req_f & dcsr[2]; // @[dec_tlu_ctl.scala 439:60]
  reg  dcsr_single_step_running_f; // @[dec_tlu_ctl.scala 464:73]
  wire  _T_178 = ~dcsr_single_step_done_f; // @[dec_tlu_ctl.scala 439:111]
  wire  _T_179 = dcsr_single_step_running_f & _T_178; // @[dec_tlu_ctl.scala 439:109]
  wire  dcsr_single_step_running = _T_177 | _T_179; // @[dec_tlu_ctl.scala 439:79]
  wire  _T_665 = ~dcsr_single_step_running; // @[dec_tlu_ctl.scala 740:55]
  wire  _T_666 = _T_665 | io_dec_tlu_i0_valid_r; // @[dec_tlu_ctl.scala 740:81]
  wire  _T_667 = internal_dbg_halt_mode & _T_666; // @[dec_tlu_ctl.scala 740:52]
  wire  _T_346 = ~io_dec_tlu_debug_mode; // @[dec_tlu_ctl.scala 569:62]
  wire  _T_347 = i_cpu_halt_req_sync & _T_346; // @[dec_tlu_ctl.scala 569:60]
  wire  i_cpu_halt_req_sync_qual = _T_347 & _T_107; // @[dec_tlu_ctl.scala 569:85]
  wire  ext_halt_pulse = i_cpu_halt_req_sync_qual & _T_398; // @[dec_tlu_ctl.scala 585:50]
  wire  fw_halt_req = csr_io_fw_halt_req; // @[dec_tlu_ctl.scala 1005:31]
  wire  enter_pmu_fw_halt_req = ext_halt_pulse | fw_halt_req; // @[dec_tlu_ctl.scala 586:48]
  reg  pmu_fw_halt_req_f; // @[dec_tlu_ctl.scala 578:73]
  wire  _T_371 = pmu_fw_halt_req_f & core_empty; // @[dec_tlu_ctl.scala 591:45]
  wire  _T_372 = _T_371 & halt_taken; // @[dec_tlu_ctl.scala 591:58]
  wire  _T_373 = ~enter_debug_halt_req; // @[dec_tlu_ctl.scala 591:73]
  wire  _T_374 = _T_372 & _T_373; // @[dec_tlu_ctl.scala 591:71]
  wire  _T_375 = ~i_cpu_run_req_d1; // @[dec_tlu_ctl.scala 591:121]
  wire  _T_376 = pmu_fw_tlu_halted_f & _T_375; // @[dec_tlu_ctl.scala 591:119]
  wire  _T_377 = _T_374 | _T_376; // @[dec_tlu_ctl.scala 591:96]
  wire  _T_378 = ~debug_halt_req_f; // @[dec_tlu_ctl.scala 591:143]
  wire  pmu_fw_tlu_halted = _T_377 & _T_378; // @[dec_tlu_ctl.scala 591:141]
  wire  _T_361 = ~pmu_fw_tlu_halted; // @[dec_tlu_ctl.scala 587:72]
  wire  _T_362 = pmu_fw_halt_req_f & _T_361; // @[dec_tlu_ctl.scala 587:70]
  wire  _T_363 = enter_pmu_fw_halt_req | _T_362; // @[dec_tlu_ctl.scala 587:49]
  wire  pmu_fw_halt_req_ns = _T_363 & _T_378; // @[dec_tlu_ctl.scala 587:93]
  reg  internal_pmu_fw_halt_mode_f; // @[dec_tlu_ctl.scala 577:68]
  wire  _T_367 = internal_pmu_fw_halt_mode_f & _T_375; // @[dec_tlu_ctl.scala 588:83]
  wire  _T_369 = _T_367 & _T_378; // @[dec_tlu_ctl.scala 588:103]
  wire  internal_pmu_fw_halt_mode = pmu_fw_halt_req_ns | _T_369; // @[dec_tlu_ctl.scala 588:52]
  wire  _T_668 = _T_667 | internal_pmu_fw_halt_mode; // @[dec_tlu_ctl.scala 740:107]
  wire  _T_669 = _T_668 | i_cpu_halt_req_d1; // @[dec_tlu_ctl.scala 740:135]
  wire  _T_738 = ~internal_pmu_fw_halt_mode; // @[dec_tlu_ctl.scala 772:35]
  wire  _T_739 = nmi_int_detected & _T_738; // @[dec_tlu_ctl.scala 772:33]
  wire  _T_740 = ~internal_dbg_halt_mode; // @[dec_tlu_ctl.scala 772:65]
  wire  _T_742 = dcsr_single_step_running_f & dcsr[11]; // @[dec_tlu_ctl.scala 772:119]
  wire  _T_743 = ~io_dec_tlu_i0_valid_r; // @[dec_tlu_ctl.scala 772:141]
  wire  _T_744 = _T_742 & _T_743; // @[dec_tlu_ctl.scala 772:139]
  wire  _T_746 = _T_744 & _T_178; // @[dec_tlu_ctl.scala 772:164]
  wire  _T_747 = _T_740 | _T_746; // @[dec_tlu_ctl.scala 772:89]
  wire  _T_748 = _T_739 & _T_747; // @[dec_tlu_ctl.scala 772:62]
  wire  _T_463 = io_dec_tlu_packet_r_pmu_i0_itype == 4'h8; // @[dec_tlu_ctl.scala 658:51]
  wire  _T_464 = _T_463 & io_dec_tlu_i0_valid_r; // @[dec_tlu_ctl.scala 658:64]
  wire  _T_297 = io_dec_tlu_flush_lower_wb | io_dec_tlu_dbg_halted; // @[dec_tlu_ctl.scala 520:58]
  wire [3:0] _T_299 = _T_297 ? 4'hf : 4'h0; // @[Bitwise.scala 72:12]
  wire [3:0] _T_300 = ~_T_299; // @[dec_tlu_ctl.scala 520:23]
  wire [3:0] _T_292 = io_dec_tlu_i0_valid_r ? 4'hf : 4'h0; // @[Bitwise.scala 72:12]
  wire [3:0] _T_294 = _T_292 & io_dec_tlu_packet_r_i0trigger; // @[dec_tlu_ctl.scala 518:53]
  wire [9:0] mtdata1_t_3 = csr_io_mtdata1_t_3; // @[dec_tlu_ctl.scala 156:67 dec_tlu_ctl.scala 1010:33]
  wire [9:0] mtdata1_t_2 = csr_io_mtdata1_t_2; // @[dec_tlu_ctl.scala 156:67 dec_tlu_ctl.scala 1010:33]
  wire [9:0] mtdata1_t_1 = csr_io_mtdata1_t_1; // @[dec_tlu_ctl.scala 156:67 dec_tlu_ctl.scala 1010:33]
  wire [9:0] mtdata1_t_0 = csr_io_mtdata1_t_0; // @[dec_tlu_ctl.scala 156:67 dec_tlu_ctl.scala 1010:33]
  wire [3:0] trigger_execute = {mtdata1_t_3[2],mtdata1_t_2[2],mtdata1_t_1[2],mtdata1_t_0[2]}; // @[Cat.scala 29:58]
  wire [3:0] trigger_data = {mtdata1_t_3[7],mtdata1_t_2[7],mtdata1_t_1[7],mtdata1_t_0[7]}; // @[Cat.scala 29:58]
  wire [3:0] _T_279 = trigger_execute & trigger_data; // @[dec_tlu_ctl.scala 510:57]
  wire  inst_acc_r_raw = io_dec_tlu_packet_r_icaf & io_dec_tlu_i0_valid_r; // @[dec_tlu_ctl.scala 666:49]
  wire [3:0] _T_281 = inst_acc_r_raw ? 4'hf : 4'h0; // @[Bitwise.scala 72:12]
  wire [3:0] _T_282 = _T_279 & _T_281; // @[dec_tlu_ctl.scala 510:72]
  wire  _T_283 = io_tlu_exu_exu_i0_br_error_r | io_tlu_exu_exu_i0_br_start_error_r; // @[dec_tlu_ctl.scala 510:137]
  wire [3:0] _T_285 = _T_283 ? 4'hf : 4'h0; // @[Bitwise.scala 72:12]
  wire [3:0] _T_286 = _T_282 | _T_285; // @[dec_tlu_ctl.scala 510:98]
  wire [3:0] i0_iside_trigger_has_pri_r = ~_T_286; // @[dec_tlu_ctl.scala 510:38]
  wire [3:0] _T_295 = _T_294 & i0_iside_trigger_has_pri_r; // @[dec_tlu_ctl.scala 518:90]
  wire [3:0] trigger_store = {mtdata1_t_3[1],mtdata1_t_2[1],mtdata1_t_1[1],mtdata1_t_0[1]}; // @[Cat.scala 29:58]
  wire [3:0] _T_287 = trigger_store & trigger_data; // @[dec_tlu_ctl.scala 513:51]
  wire [3:0] _T_289 = io_lsu_error_pkt_r_valid ? 4'hf : 4'h0; // @[Bitwise.scala 72:12]
  wire [3:0] _T_290 = _T_287 & _T_289; // @[dec_tlu_ctl.scala 513:66]
  wire [3:0] i0_lsu_trigger_has_pri_r = ~_T_290; // @[dec_tlu_ctl.scala 513:35]
  wire [3:0] _T_296 = _T_295 & i0_lsu_trigger_has_pri_r; // @[dec_tlu_ctl.scala 518:119]
  wire [1:0] mstatus = csr_io_mstatus; // @[dec_tlu_ctl.scala 1006:31]
  wire  _T_259 = mtdata1_t_3[6] | mstatus[0]; // @[dec_tlu_ctl.scala 507:62]
  wire  _T_261 = _T_259 & mtdata1_t_3[3]; // @[dec_tlu_ctl.scala 507:86]
  wire  _T_264 = mtdata1_t_2[6] | mstatus[0]; // @[dec_tlu_ctl.scala 507:150]
  wire  _T_266 = _T_264 & mtdata1_t_2[3]; // @[dec_tlu_ctl.scala 507:174]
  wire  _T_269 = mtdata1_t_1[6] | mstatus[0]; // @[dec_tlu_ctl.scala 507:239]
  wire  _T_271 = _T_269 & mtdata1_t_1[3]; // @[dec_tlu_ctl.scala 507:263]
  wire  _T_274 = mtdata1_t_0[6] | mstatus[0]; // @[dec_tlu_ctl.scala 507:328]
  wire  _T_276 = _T_274 & mtdata1_t_0[3]; // @[dec_tlu_ctl.scala 507:352]
  wire [3:0] trigger_enabled = {_T_261,_T_266,_T_271,_T_276}; // @[Cat.scala 29:58]
  wire [3:0] i0trigger_qual_r = _T_296 & trigger_enabled; // @[dec_tlu_ctl.scala 518:146]
  wire [3:0] i0_trigger_r = _T_300 & i0trigger_qual_r; // @[dec_tlu_ctl.scala 520:84]
  wire  _T_303 = ~mtdata1_t_2[5]; // @[dec_tlu_ctl.scala 523:60]
  wire  _T_305 = _T_303 | i0_trigger_r[2]; // @[dec_tlu_ctl.scala 523:89]
  wire  _T_306 = i0_trigger_r[3] & _T_305; // @[dec_tlu_ctl.scala 523:57]
  wire  _T_311 = _T_303 | i0_trigger_r[3]; // @[dec_tlu_ctl.scala 523:157]
  wire  _T_312 = i0_trigger_r[2] & _T_311; // @[dec_tlu_ctl.scala 523:125]
  wire  _T_315 = ~mtdata1_t_0[5]; // @[dec_tlu_ctl.scala 523:196]
  wire  _T_317 = _T_315 | i0_trigger_r[0]; // @[dec_tlu_ctl.scala 523:225]
  wire  _T_318 = i0_trigger_r[1] & _T_317; // @[dec_tlu_ctl.scala 523:193]
  wire  _T_323 = _T_315 | i0_trigger_r[1]; // @[dec_tlu_ctl.scala 523:293]
  wire  _T_324 = i0_trigger_r[0] & _T_323; // @[dec_tlu_ctl.scala 523:261]
  wire [3:0] i0_trigger_chain_masked_r = {_T_306,_T_312,_T_318,_T_324}; // @[Cat.scala 29:58]
  wire  i0_trigger_hit_raw_r = |i0_trigger_chain_masked_r; // @[dec_tlu_ctl.scala 526:57]
  wire  _T_465 = ~i0_trigger_hit_raw_r; // @[dec_tlu_ctl.scala 658:90]
  wire  _T_466 = _T_464 & _T_465; // @[dec_tlu_ctl.scala 658:88]
  wire  _T_468 = ~dcsr[15]; // @[dec_tlu_ctl.scala 658:110]
  wire  _T_469 = _T_466 & _T_468; // @[dec_tlu_ctl.scala 658:108]
  reg  tlu_flush_lower_r_d1; // @[dec_tlu_ctl.scala 328:80]
  wire  _T_429 = ~tlu_flush_lower_r_d1; // @[dec_tlu_ctl.scala 633:44]
  wire  _T_430 = io_dec_tlu_i0_valid_r & _T_429; // @[dec_tlu_ctl.scala 633:42]
  wire  _T_432 = _T_430 & _T_283; // @[dec_tlu_ctl.scala 633:66]
  reg  ic_perr_r_d1; // @[dec_tlu_ctl.scala 322:89]
  reg  iccm_sbecc_r_d1; // @[dec_tlu_ctl.scala 323:89]
  wire  _T_433 = ic_perr_r_d1 | iccm_sbecc_r_d1; // @[dec_tlu_ctl.scala 633:154]
  wire  _T_435 = _T_433 & _T_107; // @[dec_tlu_ctl.scala 633:173]
  wire  _T_436 = _T_432 | _T_435; // @[dec_tlu_ctl.scala 633:137]
  wire  _T_438 = _T_436 & _T_465; // @[dec_tlu_ctl.scala 633:196]
  wire  _T_410 = io_dec_tlu_i0_valid_r & _T_465; // @[dec_tlu_ctl.scala 621:47]
  wire  _T_411 = ~io_lsu_error_pkt_r_bits_inst_type; // @[dec_tlu_ctl.scala 621:70]
  wire  _T_412 = _T_411 & io_lsu_error_pkt_r_bits_single_ecc_error; // @[dec_tlu_ctl.scala 621:105]
  wire  lsu_i0_rfnpc_r = _T_410 & _T_412; // @[dec_tlu_ctl.scala 621:67]
  wire  _T_439 = ~lsu_i0_rfnpc_r; // @[dec_tlu_ctl.scala 633:220]
  wire  rfpc_i0_r = _T_438 & _T_439; // @[dec_tlu_ctl.scala 633:217]
  wire  _T_470 = ~rfpc_i0_r; // @[dec_tlu_ctl.scala 658:132]
  wire  ebreak_r = _T_469 & _T_470; // @[dec_tlu_ctl.scala 658:130]
  wire  _T_472 = io_dec_tlu_packet_r_pmu_i0_itype == 4'h9; // @[dec_tlu_ctl.scala 659:51]
  wire  _T_473 = _T_472 & io_dec_tlu_i0_valid_r; // @[dec_tlu_ctl.scala 659:64]
  wire  _T_475 = _T_473 & _T_465; // @[dec_tlu_ctl.scala 659:88]
  wire  ecall_r = _T_475 & _T_470; // @[dec_tlu_ctl.scala 659:108]
  wire  _T_523 = ebreak_r | ecall_r; // @[dec_tlu_ctl.scala 686:41]
  wire  _T_478 = ~io_dec_tlu_packet_r_legal; // @[dec_tlu_ctl.scala 660:17]
  wire  _T_479 = _T_478 & io_dec_tlu_i0_valid_r; // @[dec_tlu_ctl.scala 660:46]
  wire  _T_481 = _T_479 & _T_465; // @[dec_tlu_ctl.scala 660:70]
  wire  illegal_r = _T_481 & _T_470; // @[dec_tlu_ctl.scala 660:90]
  wire  _T_524 = _T_523 | illegal_r; // @[dec_tlu_ctl.scala 686:51]
  wire  _T_511 = inst_acc_r_raw & _T_470; // @[dec_tlu_ctl.scala 667:33]
  wire  inst_acc_r = _T_511 & _T_465; // @[dec_tlu_ctl.scala 667:46]
  wire  _T_525 = _T_524 | inst_acc_r; // @[dec_tlu_ctl.scala 686:63]
  wire  _T_527 = _T_525 & _T_470; // @[dec_tlu_ctl.scala 686:77]
  wire  _T_528 = ~io_dec_tlu_dbg_halted; // @[dec_tlu_ctl.scala 686:92]
  wire  i0_exception_valid_r = _T_527 & _T_528; // @[dec_tlu_ctl.scala 686:90]
  wire  _T_789 = i0_exception_valid_r | rfpc_i0_r; // @[dec_tlu_ctl.scala 785:49]
  wire  _T_402 = ~io_dec_tlu_flush_lower_wb; // @[dec_tlu_ctl.scala 609:57]
  wire  lsu_exc_valid_r_raw = io_lsu_error_pkt_r_valid & _T_402; // @[dec_tlu_ctl.scala 609:55]
  wire  _T_403 = io_lsu_error_pkt_r_valid & lsu_exc_valid_r_raw; // @[dec_tlu_ctl.scala 611:40]
  wire  _T_405 = _T_403 & _T_465; // @[dec_tlu_ctl.scala 611:62]
  wire  lsu_exc_valid_r = _T_405 & _T_470; // @[dec_tlu_ctl.scala 611:82]
  wire  _T_790 = _T_789 | lsu_exc_valid_r; // @[dec_tlu_ctl.scala 785:61]
  wire  _T_490 = io_dec_tlu_packet_r_fence_i & io_dec_tlu_i0_valid_r; // @[dec_tlu_ctl.scala 663:50]
  wire  _T_492 = _T_490 & _T_465; // @[dec_tlu_ctl.scala 663:74]
  wire  fence_i_r = _T_492 & _T_470; // @[dec_tlu_ctl.scala 663:95]
  wire  _T_791 = _T_790 | fence_i_r; // @[dec_tlu_ctl.scala 785:79]
  wire  _T_792 = _T_791 | lsu_i0_rfnpc_r; // @[dec_tlu_ctl.scala 785:91]
  wire  _T_414 = io_dec_tlu_i0_valid_r & _T_470; // @[dec_tlu_ctl.scala 624:50]
  wire  _T_415 = ~lsu_exc_valid_r; // @[dec_tlu_ctl.scala 624:65]
  wire  _T_416 = _T_414 & _T_415; // @[dec_tlu_ctl.scala 624:63]
  wire  _T_417 = ~inst_acc_r; // @[dec_tlu_ctl.scala 624:82]
  wire  _T_418 = _T_416 & _T_417; // @[dec_tlu_ctl.scala 624:79]
  wire  _T_420 = _T_418 & _T_528; // @[dec_tlu_ctl.scala 624:94]
  reg  request_debug_mode_r_d1; // @[dec_tlu_ctl.scala 462:81]
  wire  _T_421 = ~request_debug_mode_r_d1; // @[dec_tlu_ctl.scala 624:121]
  wire  _T_422 = _T_420 & _T_421; // @[dec_tlu_ctl.scala 624:119]
  wire  tlu_i0_commit_cmt = _T_422 & _T_465; // @[dec_tlu_ctl.scala 624:146]
  reg  iccm_repair_state_d1; // @[dec_tlu_ctl.scala 321:80]
  wire  _T_444 = tlu_i0_commit_cmt & iccm_repair_state_d1; // @[dec_tlu_ctl.scala 642:52]
  wire  _T_484 = io_dec_tlu_packet_r_pmu_i0_itype == 4'hc; // @[dec_tlu_ctl.scala 661:51]
  wire  _T_485 = _T_484 & io_dec_tlu_i0_valid_r; // @[dec_tlu_ctl.scala 661:64]
  wire  _T_487 = _T_485 & _T_465; // @[dec_tlu_ctl.scala 661:88]
  wire  mret_r = _T_487 & _T_470; // @[dec_tlu_ctl.scala 661:108]
  wire  _T_446 = _T_523 | mret_r; // @[dec_tlu_ctl.scala 642:98]
  wire  take_reset = reset_delayed & io_mpc_reset_run_req; // @[dec_tlu_ctl.scala 771:32]
  wire  _T_447 = _T_446 | take_reset; // @[dec_tlu_ctl.scala 642:107]
  wire  _T_448 = _T_447 | illegal_r; // @[dec_tlu_ctl.scala 642:120]
  wire  _T_449 = io_dec_csr_wraddr_r == 12'h7c2; // @[dec_tlu_ctl.scala 642:176]
  wire  _T_450 = dec_csr_wen_r_mod & _T_449; // @[dec_tlu_ctl.scala 642:153]
  wire  _T_451 = _T_448 | _T_450; // @[dec_tlu_ctl.scala 642:132]
  wire  _T_452 = ~_T_451; // @[dec_tlu_ctl.scala 642:77]
  wire  iccm_repair_state_rfnpc = _T_444 & _T_452; // @[dec_tlu_ctl.scala 642:75]
  wire  _T_793 = _T_792 | iccm_repair_state_rfnpc; // @[dec_tlu_ctl.scala 785:108]
  wire  _T_794 = _T_793 | debug_resume_req_f; // @[dec_tlu_ctl.scala 785:135]
  wire  _T_786 = i_cpu_run_req_d1 & pmu_fw_tlu_halted_f; // @[dec_tlu_ctl.scala 783:43]
  wire  _T_211 = ~io_dec_pause_state; // @[dec_tlu_ctl.scala 482:28]
  reg  dec_pause_state_f; // @[dec_tlu_ctl.scala 461:81]
  wire  _T_212 = _T_211 & dec_pause_state_f; // @[dec_tlu_ctl.scala 482:48]
  wire  _T_213 = ext_int_ready | ce_int_ready; // @[dec_tlu_ctl.scala 482:86]
  wire  _T_214 = _T_213 | timer_int_ready; // @[dec_tlu_ctl.scala 482:101]
  wire  _T_215 = _T_214 | soft_int_ready; // @[dec_tlu_ctl.scala 482:119]
  wire  _T_216 = _T_215 | int_timer0_int_hold_f; // @[dec_tlu_ctl.scala 482:136]
  wire  _T_217 = _T_216 | int_timer1_int_hold_f; // @[dec_tlu_ctl.scala 482:160]
  wire  _T_218 = _T_217 | nmi_int_detected; // @[dec_tlu_ctl.scala 482:184]
  wire  _T_219 = _T_218 | ext_int_freeze_d1; // @[dec_tlu_ctl.scala 482:203]
  wire  _T_220 = ~_T_219; // @[dec_tlu_ctl.scala 482:70]
  wire  _T_221 = _T_212 & _T_220; // @[dec_tlu_ctl.scala 482:68]
  wire  _T_223 = _T_221 & _T_140; // @[dec_tlu_ctl.scala 482:224]
  wire  _T_225 = _T_223 & _T_378; // @[dec_tlu_ctl.scala 482:248]
  wire  _T_226 = ~pmu_fw_halt_req_f; // @[dec_tlu_ctl.scala 482:270]
  wire  _T_227 = _T_225 & _T_226; // @[dec_tlu_ctl.scala 482:268]
  wire  _T_228 = ~halt_taken_f; // @[dec_tlu_ctl.scala 482:291]
  wire  pause_expired_r = _T_227 & _T_228; // @[dec_tlu_ctl.scala 482:289]
  wire  sel_npc_resume = _T_786 | pause_expired_r; // @[dec_tlu_ctl.scala 783:66]
  wire  _T_795 = _T_794 | sel_npc_resume; // @[dec_tlu_ctl.scala 785:157]
  reg  dec_tlu_wr_pause_r_d1; // @[dec_tlu_ctl.scala 460:81]
  wire  _T_796 = _T_795 | dec_tlu_wr_pause_r_d1; // @[dec_tlu_ctl.scala 785:175]
  wire  synchronous_flush_r = _T_796 | i0_trigger_hit_raw_r; // @[dec_tlu_ctl.scala 785:201]
  wire  _T_749 = ~synchronous_flush_r; // @[dec_tlu_ctl.scala 772:195]
  wire  _T_750 = _T_748 & _T_749; // @[dec_tlu_ctl.scala 772:193]
  wire  _T_751 = ~mret_r; // @[dec_tlu_ctl.scala 772:218]
  wire  _T_752 = _T_750 & _T_751; // @[dec_tlu_ctl.scala 772:216]
  wire  _T_753 = ~take_reset; // @[dec_tlu_ctl.scala 772:228]
  wire  _T_754 = _T_752 & _T_753; // @[dec_tlu_ctl.scala 772:226]
  wire  _T_519 = _T_466 & dcsr[15]; // @[dec_tlu_ctl.scala 670:121]
  wire  ebreak_to_debug_mode_r = _T_519 & _T_470; // @[dec_tlu_ctl.scala 670:142]
  wire  _T_755 = ~ebreak_to_debug_mode_r; // @[dec_tlu_ctl.scala 772:242]
  wire  _T_756 = _T_754 & _T_755; // @[dec_tlu_ctl.scala 772:240]
  wire  _T_760 = _T_107 | _T_44; // @[dec_tlu_ctl.scala 772:288]
  wire  take_nmi = _T_756 & _T_760; // @[dec_tlu_ctl.scala 772:266]
  wire  _T_670 = _T_669 | take_nmi; // @[dec_tlu_ctl.scala 740:155]
  wire  _T_671 = _T_670 | ebreak_to_debug_mode_r; // @[dec_tlu_ctl.scala 740:166]
  wire  _T_672 = _T_671 | synchronous_flush_r; // @[dec_tlu_ctl.scala 740:191]
  reg  exc_or_int_valid_r_d1; // @[dec_tlu_ctl.scala 811:90]
  wire  _T_673 = _T_672 | exc_or_int_valid_r_d1; // @[dec_tlu_ctl.scala 740:214]
  wire  _T_674 = _T_673 | mret_r; // @[dec_tlu_ctl.scala 740:238]
  wire  block_interrupts = _T_674 | ext_int_freeze_d1; // @[dec_tlu_ctl.scala 740:247]
  wire  _T_704 = ~block_interrupts; // @[dec_tlu_ctl.scala 768:91]
  wire  take_timer_int = _T_703 & _T_704; // @[dec_tlu_ctl.scala 768:89]
  wire  _T_762 = take_ext_int | take_timer_int; // @[dec_tlu_ctl.scala 775:38]
  wire  _T_693 = soft_int_ready & _T_700; // @[dec_tlu_ctl.scala 767:36]
  wire  _T_695 = _T_693 & _T_702; // @[dec_tlu_ctl.scala 767:53]
  wire  take_soft_int = _T_695 & _T_704; // @[dec_tlu_ctl.scala 767:69]
  wire  _T_763 = _T_762 | take_soft_int; // @[dec_tlu_ctl.scala 775:55]
  wire  _T_764 = _T_763 | take_nmi; // @[dec_tlu_ctl.scala 775:71]
  wire  _T_689 = ce_int_ready & _T_700; // @[dec_tlu_ctl.scala 766:33]
  wire  take_ce_int = _T_689 & _T_704; // @[dec_tlu_ctl.scala 766:50]
  wire  _T_765 = _T_764 | take_ce_int; // @[dec_tlu_ctl.scala 775:82]
  wire  int_timer0_int_possible = mstatus_mie_ns & mie_ns[4]; // @[dec_tlu_ctl.scala 726:49]
  wire  int_timer0_int_ready = mip[4] & int_timer0_int_possible; // @[dec_tlu_ctl.scala 727:47]
  wire  _T_706 = int_timer0_int_ready | int_timer0_int_hold_f; // @[dec_tlu_ctl.scala 769:49]
  wire  _T_707 = _T_706 & int_timer0_int_possible; // @[dec_tlu_ctl.scala 769:74]
  wire  _T_709 = _T_707 & _T_631; // @[dec_tlu_ctl.scala 769:100]
  wire  _T_710 = ~timer_int_ready; // @[dec_tlu_ctl.scala 769:129]
  wire  _T_711 = _T_709 & _T_710; // @[dec_tlu_ctl.scala 769:127]
  wire  _T_713 = _T_711 & _T_698; // @[dec_tlu_ctl.scala 769:146]
  wire  _T_715 = _T_713 & _T_700; // @[dec_tlu_ctl.scala 769:164]
  wire  _T_717 = _T_715 & _T_702; // @[dec_tlu_ctl.scala 769:181]
  wire  take_int_timer0_int = _T_717 & _T_704; // @[dec_tlu_ctl.scala 769:197]
  wire  _T_766 = _T_765 | take_int_timer0_int; // @[dec_tlu_ctl.scala 775:96]
  wire  int_timer1_int_possible = mstatus_mie_ns & mie_ns[3]; // @[dec_tlu_ctl.scala 728:49]
  wire  int_timer1_int_ready = mip[3] & int_timer1_int_possible; // @[dec_tlu_ctl.scala 729:47]
  wire  _T_720 = int_timer1_int_ready | int_timer1_int_hold_f; // @[dec_tlu_ctl.scala 770:49]
  wire  _T_721 = _T_720 & int_timer1_int_possible; // @[dec_tlu_ctl.scala 770:74]
  wire  _T_723 = _T_721 & _T_631; // @[dec_tlu_ctl.scala 770:100]
  wire  _T_725 = ~_T_706; // @[dec_tlu_ctl.scala 770:129]
  wire  _T_726 = _T_723 & _T_725; // @[dec_tlu_ctl.scala 770:127]
  wire  _T_728 = _T_726 & _T_710; // @[dec_tlu_ctl.scala 770:177]
  wire  _T_730 = _T_728 & _T_698; // @[dec_tlu_ctl.scala 770:196]
  wire  _T_732 = _T_730 & _T_700; // @[dec_tlu_ctl.scala 770:214]
  wire  _T_734 = _T_732 & _T_702; // @[dec_tlu_ctl.scala 770:231]
  wire  take_int_timer1_int = _T_734 & _T_704; // @[dec_tlu_ctl.scala 770:247]
  wire  interrupt_valid_r = _T_766 | take_int_timer1_int; // @[dec_tlu_ctl.scala 775:118]
  wire  _T_15 = _T_14 | interrupt_valid_r; // @[dec_tlu_ctl.scala 316:69]
  wire  _T_16 = _T_15 | interrupt_valid_r_d1; // @[dec_tlu_ctl.scala 316:89]
  wire  _T_17 = _T_16 | reset_delayed; // @[dec_tlu_ctl.scala 316:112]
  wire  _T_18 = _T_17 | pause_expired_r; // @[dec_tlu_ctl.scala 316:128]
  reg  pause_expired_wb; // @[dec_tlu_ctl.scala 816:90]
  wire  _T_19 = _T_18 | pause_expired_wb; // @[dec_tlu_ctl.scala 316:146]
  wire  _T_496 = io_tlu_mem_ifu_ic_error_start & _T_107; // @[dec_tlu_ctl.scala 664:51]
  wire  _T_498 = _T_152 | dcsr_single_step_running; // @[dec_tlu_ctl.scala 664:101]
  wire  _T_499 = _T_496 & _T_498; // @[dec_tlu_ctl.scala 664:72]
  wire  _T_500 = ~internal_pmu_fw_halt_mode_f; // @[dec_tlu_ctl.scala 664:131]
  wire  ic_perr_r = _T_499 & _T_500; // @[dec_tlu_ctl.scala 664:129]
  wire  _T_20 = _T_19 | ic_perr_r; // @[dec_tlu_ctl.scala 316:165]
  wire  _T_21 = _T_20 | ic_perr_r_d1; // @[dec_tlu_ctl.scala 316:177]
  wire  _T_503 = io_tlu_mem_ifu_iccm_rd_ecc_single_err & _T_107; // @[dec_tlu_ctl.scala 665:59]
  wire  _T_506 = _T_503 & _T_498; // @[dec_tlu_ctl.scala 665:80]
  wire  iccm_sbecc_r = _T_506 & _T_500; // @[dec_tlu_ctl.scala 665:137]
  wire  _T_22 = _T_21 | iccm_sbecc_r; // @[dec_tlu_ctl.scala 316:192]
  wire  _T_23 = _T_22 | iccm_sbecc_r_d1; // @[dec_tlu_ctl.scala 316:207]
  wire  flush_clkvalid = _T_23 | io_dec_tlu_dec_clk_override; // @[dec_tlu_ctl.scala 316:225]
  reg  lsu_pmu_load_external_r; // @[dec_tlu_ctl.scala 326:80]
  reg  lsu_pmu_store_external_r; // @[dec_tlu_ctl.scala 327:72]
  reg  _T_32; // @[dec_tlu_ctl.scala 329:73]
  reg  internal_dbg_halt_mode_f2; // @[dec_tlu_ctl.scala 330:72]
  reg  _T_33; // @[dec_tlu_ctl.scala 331:89]
  reg  nmi_lsu_load_type_f; // @[dec_tlu_ctl.scala 342:72]
  reg  nmi_lsu_store_type_f; // @[dec_tlu_ctl.scala 343:72]
  wire  _T_46 = nmi_lsu_detected & io_tlu_busbuff_lsu_imprecise_error_load_any; // @[dec_tlu_ctl.scala 351:48]
  wire  _T_49 = ~_T_41; // @[dec_tlu_ctl.scala 351:96]
  wire  _T_50 = _T_46 & _T_49; // @[dec_tlu_ctl.scala 351:94]
  wire  _T_52 = nmi_lsu_load_type_f & _T_40; // @[dec_tlu_ctl.scala 351:159]
  wire  _T_54 = nmi_lsu_detected & io_tlu_busbuff_lsu_imprecise_error_store_any; // @[dec_tlu_ctl.scala 352:49]
  wire  _T_58 = _T_54 & _T_49; // @[dec_tlu_ctl.scala 352:96]
  wire  _T_60 = nmi_lsu_store_type_f & _T_40; // @[dec_tlu_ctl.scala 352:162]
  reg  mpc_debug_halt_req_sync_f; // @[dec_tlu_ctl.scala 360:72]
  reg  mpc_debug_run_req_sync_f; // @[dec_tlu_ctl.scala 361:72]
  reg  mpc_run_state_f; // @[dec_tlu_ctl.scala 363:88]
  reg  debug_brkpt_status_f; // @[dec_tlu_ctl.scala 364:80]
  reg  mpc_debug_halt_ack_f; // @[dec_tlu_ctl.scala 365:80]
  reg  mpc_debug_run_ack_f; // @[dec_tlu_ctl.scala 366:80]
  reg  dbg_run_state_f; // @[dec_tlu_ctl.scala 368:88]
  reg  _T_65; // @[dec_tlu_ctl.scala 369:81]
  wire  _T_66 = ~mpc_debug_halt_req_sync_f; // @[dec_tlu_ctl.scala 373:71]
  wire  mpc_debug_halt_req_sync_pulse = mpc_debug_halt_req_sync & _T_66; // @[dec_tlu_ctl.scala 373:69]
  wire  _T_67 = ~mpc_debug_run_req_sync_f; // @[dec_tlu_ctl.scala 374:70]
  wire  mpc_debug_run_req_sync_pulse = mpc_debug_run_req_sync & _T_67; // @[dec_tlu_ctl.scala 374:68]
  wire  _T_68 = mpc_halt_state_f | mpc_debug_halt_req_sync_pulse; // @[dec_tlu_ctl.scala 376:48]
  wire  _T_71 = _T_68 | _T_111; // @[dec_tlu_ctl.scala 376:80]
  wire  _T_72 = ~mpc_debug_run_req_sync; // @[dec_tlu_ctl.scala 376:125]
  wire  mpc_halt_state_ns = _T_71 & _T_72; // @[dec_tlu_ctl.scala 376:123]
  wire  _T_74 = ~mpc_debug_run_ack_f; // @[dec_tlu_ctl.scala 377:80]
  wire  _T_75 = mpc_debug_run_req_sync_pulse & _T_74; // @[dec_tlu_ctl.scala 377:78]
  wire  _T_76 = mpc_run_state_f | _T_75; // @[dec_tlu_ctl.scala 377:46]
  wire  _T_77 = ~dcsr_single_step_running_f; // @[dec_tlu_ctl.scala 377:133]
  wire  _T_78 = debug_mode_status & _T_77; // @[dec_tlu_ctl.scala 377:131]
  wire  mpc_run_state_ns = _T_76 & _T_78; // @[dec_tlu_ctl.scala 377:103]
  wire  _T_80 = dbg_halt_req_final | dcsr_single_step_done_f; // @[dec_tlu_ctl.scala 379:70]
  wire  _T_81 = _T_80 | trigger_hit_dmode_r_d1; // @[dec_tlu_ctl.scala 379:96]
  wire  _T_82 = _T_81 | ebreak_to_debug_mode_r_d1; // @[dec_tlu_ctl.scala 379:121]
  wire  _T_83 = dbg_halt_state_f | _T_82; // @[dec_tlu_ctl.scala 379:48]
  wire  _T_84 = ~io_dbg_resume_req; // @[dec_tlu_ctl.scala 379:153]
  wire  dbg_halt_state_ns = _T_83 & _T_84; // @[dec_tlu_ctl.scala 379:151]
  wire  _T_86 = dbg_run_state_f | io_dbg_resume_req; // @[dec_tlu_ctl.scala 380:46]
  wire  dbg_run_state_ns = _T_86 & _T_78; // @[dec_tlu_ctl.scala 380:67]
  wire  debug_brkpt_valid = ebreak_to_debug_mode_r_d1 | trigger_hit_dmode_r_d1; // @[dec_tlu_ctl.scala 386:59]
  wire  _T_92 = debug_brkpt_valid | debug_brkpt_status_f; // @[dec_tlu_ctl.scala 387:53]
  wire  _T_94 = internal_dbg_halt_mode & _T_77; // @[dec_tlu_ctl.scala 387:103]
  wire  _T_96 = mpc_halt_state_f & debug_mode_status; // @[dec_tlu_ctl.scala 390:51]
  wire  _T_97 = _T_96 & mpc_debug_halt_req_sync; // @[dec_tlu_ctl.scala 390:78]
  wire  _T_99 = ~dbg_halt_state_ns; // @[dec_tlu_ctl.scala 391:59]
  wire  _T_100 = mpc_debug_run_req_sync & _T_99; // @[dec_tlu_ctl.scala 391:57]
  wire  _T_101 = ~mpc_debug_halt_req_sync; // @[dec_tlu_ctl.scala 391:80]
  wire  _T_102 = _T_100 & _T_101; // @[dec_tlu_ctl.scala 391:78]
  wire  _T_103 = mpc_debug_run_ack_f & mpc_debug_run_req_sync; // @[dec_tlu_ctl.scala 391:129]
  wire  _T_118 = mpc_run_state_ns & _T_99; // @[dec_tlu_ctl.scala 405:73]
  wire  _T_119 = ~mpc_halt_state_ns; // @[dec_tlu_ctl.scala 405:117]
  wire  _T_120 = dbg_run_state_ns & _T_119; // @[dec_tlu_ctl.scala 405:115]
  wire  _T_121 = _T_118 | _T_120; // @[dec_tlu_ctl.scala 405:95]
  wire  _T_122 = debug_halt_req_f | pmu_fw_halt_req_f; // @[dec_tlu_ctl.scala 410:43]
  wire  _T_124 = _T_122 & _T_749; // @[dec_tlu_ctl.scala 410:64]
  wire  _T_126 = _T_124 & _T_751; // @[dec_tlu_ctl.scala 410:87]
  wire  _T_128 = _T_126 & _T_228; // @[dec_tlu_ctl.scala 410:97]
  wire  _T_129 = ~dec_tlu_flush_noredir_r_d1; // @[dec_tlu_ctl.scala 410:115]
  wire  _T_130 = _T_128 & _T_129; // @[dec_tlu_ctl.scala 410:113]
  wire  take_halt = _T_130 & _T_753; // @[dec_tlu_ctl.scala 410:143]
  wire  _T_170 = debug_resume_req_f & dbg_tlu_halted_f; // @[dec_tlu_ctl.scala 435:49]
  wire  _T_172 = io_dec_tlu_i0_valid_r & _T_528; // @[dec_tlu_ctl.scala 437:59]
  wire  _T_174 = _T_172 & dcsr[2]; // @[dec_tlu_ctl.scala 437:84]
  wire  _T_329 = mtdata1_t_3[6] & mtdata1_t_3[9]; // @[dec_tlu_ctl.scala 532:61]
  wire  _T_332 = mtdata1_t_2[6] & mtdata1_t_2[9]; // @[dec_tlu_ctl.scala 532:121]
  wire  _T_335 = mtdata1_t_1[6] & mtdata1_t_1[9]; // @[dec_tlu_ctl.scala 532:181]
  wire  _T_338 = mtdata1_t_0[6] & mtdata1_t_0[9]; // @[dec_tlu_ctl.scala 532:241]
  wire [3:0] trigger_action = {_T_329,_T_332,_T_335,_T_338}; // @[Cat.scala 29:58]
  wire [3:0] _T_343 = i0_trigger_chain_masked_r & trigger_action; // @[dec_tlu_ctl.scala 538:57]
  wire  i0_trigger_action_r = |_T_343; // @[dec_tlu_ctl.scala 538:75]
  wire  trigger_hit_dmode_r = i0_trigger_hit_raw_r & i0_trigger_action_r; // @[dec_tlu_ctl.scala 540:45]
  wire  _T_180 = trigger_hit_dmode_r | ebreak_to_debug_mode_r; // @[dec_tlu_ctl.scala 444:57]
  wire  _T_182 = request_debug_mode_r_d1 & _T_402; // @[dec_tlu_ctl.scala 444:110]
  reg  request_debug_mode_done_f; // @[dec_tlu_ctl.scala 463:73]
  wire  _T_183 = request_debug_mode_r_d1 | request_debug_mode_done_f; // @[dec_tlu_ctl.scala 446:64]
  reg  _T_190; // @[dec_tlu_ctl.scala 454:81]
  wire  _T_201 = fence_i_r & internal_dbg_halt_mode; // @[dec_tlu_ctl.scala 475:71]
  wire  _T_202 = take_halt | _T_201; // @[dec_tlu_ctl.scala 475:58]
  wire  _T_203 = _T_202 | io_dec_tlu_flush_pause_r; // @[dec_tlu_ctl.scala 475:97]
  wire  _T_204 = i0_trigger_hit_raw_r & trigger_hit_dmode_r; // @[dec_tlu_ctl.scala 475:144]
  wire  _T_205 = _T_203 | _T_204; // @[dec_tlu_ctl.scala 475:124]
  wire  take_ext_int_start = ext_int_ready & _T_704; // @[dec_tlu_ctl.scala 748:45]
  wire  _T_207 = ~interrupt_valid_r; // @[dec_tlu_ctl.scala 480:61]
  wire  _T_208 = dec_tlu_wr_pause_r_d1 & _T_207; // @[dec_tlu_ctl.scala 480:59]
  wire  _T_209 = ~take_ext_int_start; // @[dec_tlu_ctl.scala 480:82]
  wire  _T_231 = io_tlu_exu_dec_tlu_flush_lower_r & dcsr[2]; // @[dec_tlu_ctl.scala 484:82]
  wire  _T_232 = io_dec_tlu_resume_ack | dcsr_single_step_running; // @[dec_tlu_ctl.scala 484:125]
  wire  _T_233 = _T_231 & _T_232; // @[dec_tlu_ctl.scala 484:100]
  wire  _T_234 = ~io_tlu_ifc_dec_tlu_flush_noredir_wb; // @[dec_tlu_ctl.scala 484:155]
  wire [3:0] _T_342 = i0_trigger_hit_raw_r ? 4'hf : 4'h0; // @[Bitwise.scala 72:12]
  wire  _T_345 = ~trigger_hit_dmode_r; // @[dec_tlu_ctl.scala 542:55]
  wire  mepc_trigger_hit_sel_pc_r = i0_trigger_hit_raw_r & _T_345; // @[dec_tlu_ctl.scala 542:53]
  wire  _T_350 = i_cpu_run_req_sync & _T_346; // @[dec_tlu_ctl.scala 570:58]
  wire  _T_351 = _T_350 & pmu_fw_tlu_halted_f; // @[dec_tlu_ctl.scala 570:83]
  wire  i_cpu_run_req_sync_qual = _T_351 & _T_107; // @[dec_tlu_ctl.scala 570:105]
  reg  _T_353; // @[dec_tlu_ctl.scala 574:81]
  reg  _T_354; // @[dec_tlu_ctl.scala 575:81]
  reg  _T_355; // @[dec_tlu_ctl.scala 576:81]
  wire  _T_384 = io_o_cpu_halt_status & _T_375; // @[dec_tlu_ctl.scala 594:89]
  wire  _T_386 = _T_384 & _T_152; // @[dec_tlu_ctl.scala 594:109]
  wire  _T_388 = io_o_cpu_halt_status & i_cpu_run_req_sync_qual; // @[dec_tlu_ctl.scala 595:41]
  wire  _T_389 = io_o_cpu_run_ack & i_cpu_run_req_sync_qual; // @[dec_tlu_ctl.scala 595:88]
  reg  lsu_single_ecc_error_r_d1; // @[dec_tlu_ctl.scala 607:72]
  reg  lsu_i0_exc_r_d1; // @[dec_tlu_ctl.scala 614:73]
  wire  _T_408 = ~io_lsu_error_pkt_r_bits_exc_type; // @[dec_tlu_ctl.scala 615:40]
  wire  lsu_exc_ma_r = lsu_exc_valid_r & _T_408; // @[dec_tlu_ctl.scala 615:38]
  wire  lsu_exc_acc_r = lsu_exc_valid_r & io_lsu_error_pkt_r_bits_exc_type; // @[dec_tlu_ctl.scala 616:38]
  wire  lsu_exc_st_r = lsu_exc_valid_r & io_lsu_error_pkt_r_bits_inst_type; // @[dec_tlu_ctl.scala 617:38]
  wire  _T_424 = rfpc_i0_r | lsu_exc_valid_r; // @[dec_tlu_ctl.scala 627:38]
  wire  _T_425 = _T_424 | inst_acc_r; // @[dec_tlu_ctl.scala 627:53]
  wire  _T_426 = illegal_r & io_dec_tlu_dbg_halted; // @[dec_tlu_ctl.scala 627:79]
  wire  _T_427 = _T_425 | _T_426; // @[dec_tlu_ctl.scala 627:66]
  wire  _T_441 = ~io_tlu_exu_dec_tlu_flush_lower_r; // @[dec_tlu_ctl.scala 636:70]
  wire  _T_442 = iccm_repair_state_d1 & _T_441; // @[dec_tlu_ctl.scala 636:68]
  wire  _T_453 = io_tlu_exu_exu_i0_br_error_r & io_dec_tlu_i0_valid_r; // @[dec_tlu_ctl.scala 645:59]
  wire  _T_455 = io_tlu_exu_exu_i0_br_start_error_r & io_dec_tlu_i0_valid_r; // @[dec_tlu_ctl.scala 646:71]
  wire  _T_457 = io_tlu_exu_exu_i0_br_valid_r & io_dec_tlu_i0_valid_r; // @[dec_tlu_ctl.scala 647:55]
  wire  _T_459 = _T_457 & _T_429; // @[dec_tlu_ctl.scala 647:79]
  wire  _T_460 = ~io_tlu_exu_exu_i0_br_mp_r; // @[dec_tlu_ctl.scala 647:106]
  wire  _T_461 = ~io_tlu_exu_exu_pmu_i0_br_ataken; // @[dec_tlu_ctl.scala 647:135]
  wire  _T_462 = _T_460 | _T_461; // @[dec_tlu_ctl.scala 647:133]
  wire  _T_529 = ~take_nmi; // @[dec_tlu_ctl.scala 695:33]
  wire  _T_530 = take_ext_int & _T_529; // @[dec_tlu_ctl.scala 695:31]
  wire  _T_533 = take_timer_int & _T_529; // @[dec_tlu_ctl.scala 696:25]
  wire  _T_536 = take_soft_int & _T_529; // @[dec_tlu_ctl.scala 697:24]
  wire  _T_539 = take_int_timer0_int & _T_529; // @[dec_tlu_ctl.scala 698:30]
  wire  _T_542 = take_int_timer1_int & _T_529; // @[dec_tlu_ctl.scala 699:30]
  wire  _T_545 = take_ce_int & _T_529; // @[dec_tlu_ctl.scala 700:22]
  wire  _T_548 = illegal_r & _T_529; // @[dec_tlu_ctl.scala 701:20]
  wire  _T_551 = ecall_r & _T_529; // @[dec_tlu_ctl.scala 702:19]
  wire  _T_554 = inst_acc_r & _T_529; // @[dec_tlu_ctl.scala 703:22]
  wire  _T_556 = ebreak_r | i0_trigger_hit_raw_r; // @[dec_tlu_ctl.scala 704:20]
  wire  _T_558 = _T_556 & _T_529; // @[dec_tlu_ctl.scala 704:40]
  wire  _T_560 = ~lsu_exc_st_r; // @[dec_tlu_ctl.scala 705:25]
  wire  _T_561 = lsu_exc_ma_r & _T_560; // @[dec_tlu_ctl.scala 705:23]
  wire  _T_563 = _T_561 & _T_529; // @[dec_tlu_ctl.scala 705:39]
  wire  _T_566 = lsu_exc_acc_r & _T_560; // @[dec_tlu_ctl.scala 706:24]
  wire  _T_568 = _T_566 & _T_529; // @[dec_tlu_ctl.scala 706:40]
  wire  _T_570 = lsu_exc_ma_r & lsu_exc_st_r; // @[dec_tlu_ctl.scala 707:23]
  wire  _T_572 = _T_570 & _T_529; // @[dec_tlu_ctl.scala 707:38]
  wire  _T_574 = lsu_exc_acc_r & lsu_exc_st_r; // @[dec_tlu_ctl.scala 708:24]
  wire  _T_576 = _T_574 & _T_529; // @[dec_tlu_ctl.scala 708:39]
  wire [4:0] _T_578 = _T_530 ? 5'hb : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_579 = _T_533 ? 5'h7 : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_580 = _T_536 ? 5'h3 : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_581 = _T_539 ? 5'h1d : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_582 = _T_542 ? 5'h1c : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_583 = _T_545 ? 5'h1e : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_584 = _T_548 ? 5'h2 : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_585 = _T_551 ? 5'hb : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_586 = _T_554 ? 5'h1 : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_587 = _T_558 ? 5'h3 : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_588 = _T_563 ? 5'h4 : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_589 = _T_568 ? 5'h5 : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_590 = _T_572 ? 5'h6 : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_591 = _T_576 ? 5'h7 : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_592 = _T_578 | _T_579; // @[Mux.scala 27:72]
  wire [4:0] _T_593 = _T_592 | _T_580; // @[Mux.scala 27:72]
  wire [4:0] _T_594 = _T_593 | _T_581; // @[Mux.scala 27:72]
  wire [4:0] _T_595 = _T_594 | _T_582; // @[Mux.scala 27:72]
  wire [4:0] _T_596 = _T_595 | _T_583; // @[Mux.scala 27:72]
  wire [4:0] _T_597 = _T_596 | _T_584; // @[Mux.scala 27:72]
  wire [4:0] _T_598 = _T_597 | _T_585; // @[Mux.scala 27:72]
  wire [4:0] _T_599 = _T_598 | _T_586; // @[Mux.scala 27:72]
  wire [4:0] _T_600 = _T_599 | _T_587; // @[Mux.scala 27:72]
  wire [4:0] _T_601 = _T_600 | _T_588; // @[Mux.scala 27:72]
  wire [4:0] _T_602 = _T_601 | _T_589; // @[Mux.scala 27:72]
  wire [4:0] _T_603 = _T_602 | _T_590; // @[Mux.scala 27:72]
  wire [4:0] exc_cause_r = _T_603 | _T_591; // @[Mux.scala 27:72]
  wire  _T_641 = io_dec_csr_stall_int_ff | synchronous_flush_r; // @[dec_tlu_ctl.scala 733:52]
  wire  _T_642 = _T_641 | exc_or_int_valid_r_d1; // @[dec_tlu_ctl.scala 733:74]
  wire  int_timer_stalled = _T_642 | mret_r; // @[dec_tlu_ctl.scala 733:98]
  wire  _T_643 = pmu_fw_tlu_halted_f | int_timer_stalled; // @[dec_tlu_ctl.scala 735:72]
  wire  _T_644 = int_timer0_int_ready & _T_643; // @[dec_tlu_ctl.scala 735:49]
  wire  _T_645 = int_timer0_int_possible & int_timer0_int_hold_f; // @[dec_tlu_ctl.scala 735:121]
  wire  _T_647 = _T_645 & _T_207; // @[dec_tlu_ctl.scala 735:145]
  wire  _T_649 = _T_647 & _T_209; // @[dec_tlu_ctl.scala 735:166]
  wire  _T_651 = _T_649 & _T_152; // @[dec_tlu_ctl.scala 735:188]
  wire  _T_654 = int_timer1_int_ready & _T_643; // @[dec_tlu_ctl.scala 736:49]
  wire  _T_655 = int_timer1_int_possible & int_timer1_int_hold_f; // @[dec_tlu_ctl.scala 736:121]
  wire  _T_657 = _T_655 & _T_207; // @[dec_tlu_ctl.scala 736:145]
  wire  _T_659 = _T_657 & _T_209; // @[dec_tlu_ctl.scala 736:166]
  wire  _T_661 = _T_659 & _T_152; // @[dec_tlu_ctl.scala 736:188]
  reg  take_ext_int_start_d2; // @[dec_tlu_ctl.scala 745:62]
  wire  _T_681 = take_ext_int_start | take_ext_int_start_d1; // @[dec_tlu_ctl.scala 750:46]
  wire  _T_682 = _T_681 | take_ext_int_start_d2; // @[dec_tlu_ctl.scala 750:70]
  wire  csr_pkt_csr_meicpct = csr_read_io_csr_pkt_csr_meicpct; // @[dec_tlu_ctl.scala 271:41 dec_tlu_ctl.scala 1013:16]
  wire  fast_int_meicpct = csr_pkt_csr_meicpct & io_dec_csr_any_unq_d; // @[dec_tlu_ctl.scala 752:49]
  wire [30:0] mtvec = csr_io_mtvec; // @[dec_tlu_ctl.scala 1008:31]
  wire [30:0] _T_769 = {mtvec[30:1],1'h0}; // @[Cat.scala 29:58]
  wire [30:0] _T_771 = {25'h0,exc_cause_r,1'h0}; // @[Cat.scala 29:58]
  wire [30:0] vectored_path = _T_769 + _T_771; // @[dec_tlu_ctl.scala 780:51]
  wire [30:0] _T_778 = mtvec[0] ? vectored_path : _T_769; // @[dec_tlu_ctl.scala 781:61]
  wire [30:0] interrupt_path = take_nmi ? io_nmi_vec : _T_778; // @[dec_tlu_ctl.scala 781:28]
  wire  _T_779 = lsu_i0_rfnpc_r | fence_i_r; // @[dec_tlu_ctl.scala 782:36]
  wire  _T_780 = _T_779 | iccm_repair_state_rfnpc; // @[dec_tlu_ctl.scala 782:48]
  wire  _T_782 = i_cpu_run_req_d1 & _T_207; // @[dec_tlu_ctl.scala 782:94]
  wire  _T_783 = _T_780 | _T_782; // @[dec_tlu_ctl.scala 782:74]
  wire  _T_785 = rfpc_i0_r & _T_743; // @[dec_tlu_ctl.scala 782:129]
  wire  sel_npc_r = _T_783 | _T_785; // @[dec_tlu_ctl.scala 782:116]
  wire  _T_798 = interrupt_valid_r | mret_r; // @[dec_tlu_ctl.scala 786:43]
  wire  _T_799 = _T_798 | synchronous_flush_r; // @[dec_tlu_ctl.scala 786:52]
  wire  _T_800 = _T_799 | take_halt; // @[dec_tlu_ctl.scala 786:74]
  wire  _T_801 = _T_800 | take_reset; // @[dec_tlu_ctl.scala 786:86]
  wire  _T_807 = _T_529 & sel_npc_r; // @[dec_tlu_ctl.scala 790:73]
  wire  _T_810 = _T_529 & rfpc_i0_r; // @[dec_tlu_ctl.scala 791:73]
  wire  _T_812 = _T_810 & io_dec_tlu_i0_valid_r; // @[dec_tlu_ctl.scala 791:91]
  wire  _T_813 = ~sel_npc_r; // @[dec_tlu_ctl.scala 791:132]
  wire  _T_814 = _T_812 & _T_813; // @[dec_tlu_ctl.scala 791:121]
  wire  _T_816 = ~take_ext_int; // @[dec_tlu_ctl.scala 792:96]
  wire  _T_817 = interrupt_valid_r & _T_816; // @[dec_tlu_ctl.scala 792:82]
  wire  _T_818 = i0_exception_valid_r | lsu_exc_valid_r; // @[dec_tlu_ctl.scala 793:80]
  wire  _T_821 = _T_818 | mepc_trigger_hit_sel_pc_r; // @[dec_tlu_ctl.scala 793:98]
  wire  _T_823 = _T_821 & _T_207; // @[dec_tlu_ctl.scala 793:143]
  wire  _T_825 = _T_823 & _T_816; // @[dec_tlu_ctl.scala 793:164]
  wire  _T_830 = _T_529 & mret_r; // @[dec_tlu_ctl.scala 794:68]
  wire  _T_833 = _T_529 & debug_resume_req_f; // @[dec_tlu_ctl.scala 795:68]
  wire  _T_836 = _T_529 & sel_npc_resume; // @[dec_tlu_ctl.scala 796:68]
  wire [30:0] _T_838 = take_ext_int ? io_lsu_fir_addr : 31'h0; // @[Mux.scala 27:72]
  wire [30:0] npc_r = csr_io_npc_r; // @[dec_tlu_ctl.scala 996:31]
  wire [30:0] _T_839 = _T_807 ? npc_r : 31'h0; // @[Mux.scala 27:72]
  wire [30:0] _T_840 = _T_814 ? io_dec_tlu_i0_pc_r : 31'h0; // @[Mux.scala 27:72]
  wire [30:0] _T_841 = _T_817 ? interrupt_path : 31'h0; // @[Mux.scala 27:72]
  wire [30:0] _T_842 = _T_825 ? _T_769 : 31'h0; // @[Mux.scala 27:72]
  wire [30:0] mepc = csr_io_mepc; // @[dec_tlu_ctl.scala 999:31]
  wire [30:0] _T_843 = _T_830 ? mepc : 31'h0; // @[Mux.scala 27:72]
  wire [30:0] dpc = csr_io_dpc; // @[dec_tlu_ctl.scala 1002:31]
  wire [30:0] _T_844 = _T_833 ? dpc : 31'h0; // @[Mux.scala 27:72]
  wire [30:0] npc_r_d1 = csr_io_npc_r_d1; // @[dec_tlu_ctl.scala 997:31]
  wire [30:0] _T_845 = _T_836 ? npc_r_d1 : 31'h0; // @[Mux.scala 27:72]
  wire [30:0] _T_846 = _T_838 | _T_839; // @[Mux.scala 27:72]
  wire [30:0] _T_847 = _T_846 | _T_840; // @[Mux.scala 27:72]
  wire [30:0] _T_848 = _T_847 | _T_841; // @[Mux.scala 27:72]
  wire [30:0] _T_849 = _T_848 | _T_842; // @[Mux.scala 27:72]
  wire [30:0] _T_850 = _T_849 | _T_843; // @[Mux.scala 27:72]
  wire [30:0] _T_851 = _T_850 | _T_844; // @[Mux.scala 27:72]
  wire [30:0] _T_852 = _T_851 | _T_845; // @[Mux.scala 27:72]
  reg [30:0] tlu_flush_path_r_d1; // @[dec_tlu_ctl.scala 799:64]
  wire  _T_854 = lsu_exc_valid_r | i0_exception_valid_r; // @[dec_tlu_ctl.scala 807:45]
  wire  _T_855 = _T_854 | interrupt_valid_r; // @[dec_tlu_ctl.scala 807:68]
  reg  i0_exception_valid_r_d1; // @[dec_tlu_ctl.scala 810:89]
  reg [4:0] exc_cause_wb; // @[dec_tlu_ctl.scala 812:89]
  wire  _T_860 = ~illegal_r; // @[dec_tlu_ctl.scala 813:119]
  reg  i0_valid_wb; // @[dec_tlu_ctl.scala 813:97]
  reg  trigger_hit_r_d1; // @[dec_tlu_ctl.scala 814:89]
  wire  csr_pkt_presync = csr_read_io_csr_pkt_presync; // @[dec_tlu_ctl.scala 271:41 dec_tlu_ctl.scala 1013:16]
  wire  _T_864 = csr_pkt_presync & io_dec_csr_any_unq_d; // @[dec_tlu_ctl.scala 1015:42]
  wire  _T_865 = ~io_dec_csr_wen_unq_d; // @[dec_tlu_ctl.scala 1015:67]
  wire  csr_pkt_postsync = csr_read_io_csr_pkt_postsync; // @[dec_tlu_ctl.scala 271:41 dec_tlu_ctl.scala 1013:16]
  wire  csr_pkt_csr_dcsr = csr_read_io_csr_pkt_csr_dcsr; // @[dec_tlu_ctl.scala 271:41 dec_tlu_ctl.scala 1013:16]
  wire  csr_pkt_csr_dpc = csr_read_io_csr_pkt_csr_dpc; // @[dec_tlu_ctl.scala 271:41 dec_tlu_ctl.scala 1013:16]
  wire  _T_874 = csr_pkt_csr_dcsr | csr_pkt_csr_dpc; // @[dec_tlu_ctl.scala 1020:55]
  wire  csr_pkt_csr_dmst = csr_read_io_csr_pkt_csr_dmst; // @[dec_tlu_ctl.scala 271:41 dec_tlu_ctl.scala 1013:16]
  wire  _T_875 = _T_874 | csr_pkt_csr_dmst; // @[dec_tlu_ctl.scala 1020:73]
  wire  csr_pkt_csr_dicawics = csr_read_io_csr_pkt_csr_dicawics; // @[dec_tlu_ctl.scala 271:41 dec_tlu_ctl.scala 1013:16]
  wire  _T_876 = _T_875 | csr_pkt_csr_dicawics; // @[dec_tlu_ctl.scala 1020:92]
  wire  csr_pkt_csr_dicad0 = csr_read_io_csr_pkt_csr_dicad0; // @[dec_tlu_ctl.scala 271:41 dec_tlu_ctl.scala 1013:16]
  wire  _T_877 = _T_876 | csr_pkt_csr_dicad0; // @[dec_tlu_ctl.scala 1020:115]
  wire  csr_pkt_csr_dicad0h = csr_read_io_csr_pkt_csr_dicad0h; // @[dec_tlu_ctl.scala 271:41 dec_tlu_ctl.scala 1013:16]
  wire  _T_878 = _T_877 | csr_pkt_csr_dicad0h; // @[dec_tlu_ctl.scala 1020:136]
  wire  csr_pkt_csr_dicad1 = csr_read_io_csr_pkt_csr_dicad1; // @[dec_tlu_ctl.scala 271:41 dec_tlu_ctl.scala 1013:16]
  wire  _T_879 = _T_878 | csr_pkt_csr_dicad1; // @[dec_tlu_ctl.scala 1020:158]
  wire  csr_pkt_csr_dicago = csr_read_io_csr_pkt_csr_dicago; // @[dec_tlu_ctl.scala 271:41 dec_tlu_ctl.scala 1013:16]
  wire  _T_880 = _T_879 | csr_pkt_csr_dicago; // @[dec_tlu_ctl.scala 1020:179]
  wire  _T_881 = ~_T_880; // @[dec_tlu_ctl.scala 1020:36]
  wire  _T_882 = _T_881 | dbg_tlu_halted_f; // @[dec_tlu_ctl.scala 1020:201]
  wire  csr_pkt_legal = csr_read_io_csr_pkt_legal; // @[dec_tlu_ctl.scala 271:41 dec_tlu_ctl.scala 1013:16]
  wire  _T_883 = csr_pkt_legal & _T_882; // @[dec_tlu_ctl.scala 1020:33]
  wire  _T_884 = ~fast_int_meicpct; // @[dec_tlu_ctl.scala 1020:223]
  wire  valid_csr = _T_883 & _T_884; // @[dec_tlu_ctl.scala 1020:221]
  wire  _T_887 = io_dec_csr_any_unq_d & valid_csr; // @[dec_tlu_ctl.scala 1022:46]
  wire  csr_pkt_csr_mvendorid = csr_read_io_csr_pkt_csr_mvendorid; // @[dec_tlu_ctl.scala 271:41 dec_tlu_ctl.scala 1013:16]
  wire  csr_pkt_csr_marchid = csr_read_io_csr_pkt_csr_marchid; // @[dec_tlu_ctl.scala 271:41 dec_tlu_ctl.scala 1013:16]
  wire  _T_888 = csr_pkt_csr_mvendorid | csr_pkt_csr_marchid; // @[dec_tlu_ctl.scala 1022:107]
  wire  csr_pkt_csr_mimpid = csr_read_io_csr_pkt_csr_mimpid; // @[dec_tlu_ctl.scala 271:41 dec_tlu_ctl.scala 1013:16]
  wire  _T_889 = _T_888 | csr_pkt_csr_mimpid; // @[dec_tlu_ctl.scala 1022:129]
  wire  csr_pkt_csr_mhartid = csr_read_io_csr_pkt_csr_mhartid; // @[dec_tlu_ctl.scala 271:41 dec_tlu_ctl.scala 1013:16]
  wire  _T_890 = _T_889 | csr_pkt_csr_mhartid; // @[dec_tlu_ctl.scala 1022:150]
  wire  csr_pkt_csr_mdseac = csr_read_io_csr_pkt_csr_mdseac; // @[dec_tlu_ctl.scala 271:41 dec_tlu_ctl.scala 1013:16]
  wire  _T_891 = _T_890 | csr_pkt_csr_mdseac; // @[dec_tlu_ctl.scala 1022:172]
  wire  csr_pkt_csr_meihap = csr_read_io_csr_pkt_csr_meihap; // @[dec_tlu_ctl.scala 271:41 dec_tlu_ctl.scala 1013:16]
  wire  _T_892 = _T_891 | csr_pkt_csr_meihap; // @[dec_tlu_ctl.scala 1022:193]
  wire  _T_893 = io_dec_csr_wen_unq_d & _T_892; // @[dec_tlu_ctl.scala 1022:82]
  wire  _T_894 = ~_T_893; // @[dec_tlu_ctl.scala 1022:59]
  dec_timer_ctl int_timers ( // @[dec_tlu_ctl.scala 275:30]
    .clock(int_timers_clock),
    .reset(int_timers_reset),
    .io_free_clk(int_timers_io_free_clk),
    .io_scan_mode(int_timers_io_scan_mode),
    .io_dec_csr_wen_r_mod(int_timers_io_dec_csr_wen_r_mod),
    .io_dec_csr_wraddr_r(int_timers_io_dec_csr_wraddr_r),
    .io_dec_csr_wrdata_r(int_timers_io_dec_csr_wrdata_r),
    .io_csr_mitctl0(int_timers_io_csr_mitctl0),
    .io_csr_mitctl1(int_timers_io_csr_mitctl1),
    .io_csr_mitb0(int_timers_io_csr_mitb0),
    .io_csr_mitb1(int_timers_io_csr_mitb1),
    .io_csr_mitcnt0(int_timers_io_csr_mitcnt0),
    .io_csr_mitcnt1(int_timers_io_csr_mitcnt1),
    .io_dec_pause_state(int_timers_io_dec_pause_state),
    .io_dec_tlu_pmu_fw_halted(int_timers_io_dec_tlu_pmu_fw_halted),
    .io_internal_dbg_halt_timers(int_timers_io_internal_dbg_halt_timers),
    .io_dec_timer_rddata_d(int_timers_io_dec_timer_rddata_d),
    .io_dec_timer_read_d(int_timers_io_dec_timer_read_d),
    .io_dec_timer_t0_pulse(int_timers_io_dec_timer_t0_pulse),
    .io_dec_timer_t1_pulse(int_timers_io_dec_timer_t1_pulse)
  );
  rvclkhdr rvclkhdr ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_io_l1clk),
    .io_clk(rvclkhdr_io_clk),
    .io_en(rvclkhdr_io_en),
    .io_scan_mode(rvclkhdr_io_scan_mode)
  );
  rvclkhdr rvclkhdr_1 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_1_io_l1clk),
    .io_clk(rvclkhdr_1_io_clk),
    .io_en(rvclkhdr_1_io_en),
    .io_scan_mode(rvclkhdr_1_io_scan_mode)
  );
  rvclkhdr rvclkhdr_2 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_2_io_l1clk),
    .io_clk(rvclkhdr_2_io_clk),
    .io_en(rvclkhdr_2_io_en),
    .io_scan_mode(rvclkhdr_2_io_scan_mode)
  );
  rvclkhdr rvclkhdr_3 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_3_io_l1clk),
    .io_clk(rvclkhdr_3_io_clk),
    .io_en(rvclkhdr_3_io_en),
    .io_scan_mode(rvclkhdr_3_io_scan_mode)
  );
  csr_tlu csr ( // @[dec_tlu_ctl.scala 818:15]
    .clock(csr_clock),
    .reset(csr_reset),
    .io_free_clk(csr_io_free_clk),
    .io_active_clk(csr_io_active_clk),
    .io_scan_mode(csr_io_scan_mode),
    .io_dec_csr_wrdata_r(csr_io_dec_csr_wrdata_r),
    .io_dec_csr_wraddr_r(csr_io_dec_csr_wraddr_r),
    .io_dec_csr_rdaddr_d(csr_io_dec_csr_rdaddr_d),
    .io_dec_csr_wen_unq_d(csr_io_dec_csr_wen_unq_d),
    .io_dec_i0_decode_d(csr_io_dec_i0_decode_d),
    .io_dec_tlu_ic_diag_pkt_icache_wrdata(csr_io_dec_tlu_ic_diag_pkt_icache_wrdata),
    .io_dec_tlu_ic_diag_pkt_icache_dicawics(csr_io_dec_tlu_ic_diag_pkt_icache_dicawics),
    .io_dec_tlu_ic_diag_pkt_icache_rd_valid(csr_io_dec_tlu_ic_diag_pkt_icache_rd_valid),
    .io_dec_tlu_ic_diag_pkt_icache_wr_valid(csr_io_dec_tlu_ic_diag_pkt_icache_wr_valid),
    .io_ifu_ic_debug_rd_data_valid(csr_io_ifu_ic_debug_rd_data_valid),
    .io_trigger_pkt_any_0_select(csr_io_trigger_pkt_any_0_select),
    .io_trigger_pkt_any_0_match_pkt(csr_io_trigger_pkt_any_0_match_pkt),
    .io_trigger_pkt_any_0_store(csr_io_trigger_pkt_any_0_store),
    .io_trigger_pkt_any_0_load(csr_io_trigger_pkt_any_0_load),
    .io_trigger_pkt_any_0_execute(csr_io_trigger_pkt_any_0_execute),
    .io_trigger_pkt_any_0_m(csr_io_trigger_pkt_any_0_m),
    .io_trigger_pkt_any_0_tdata2(csr_io_trigger_pkt_any_0_tdata2),
    .io_trigger_pkt_any_1_select(csr_io_trigger_pkt_any_1_select),
    .io_trigger_pkt_any_1_match_pkt(csr_io_trigger_pkt_any_1_match_pkt),
    .io_trigger_pkt_any_1_store(csr_io_trigger_pkt_any_1_store),
    .io_trigger_pkt_any_1_load(csr_io_trigger_pkt_any_1_load),
    .io_trigger_pkt_any_1_execute(csr_io_trigger_pkt_any_1_execute),
    .io_trigger_pkt_any_1_m(csr_io_trigger_pkt_any_1_m),
    .io_trigger_pkt_any_1_tdata2(csr_io_trigger_pkt_any_1_tdata2),
    .io_trigger_pkt_any_2_select(csr_io_trigger_pkt_any_2_select),
    .io_trigger_pkt_any_2_match_pkt(csr_io_trigger_pkt_any_2_match_pkt),
    .io_trigger_pkt_any_2_store(csr_io_trigger_pkt_any_2_store),
    .io_trigger_pkt_any_2_load(csr_io_trigger_pkt_any_2_load),
    .io_trigger_pkt_any_2_execute(csr_io_trigger_pkt_any_2_execute),
    .io_trigger_pkt_any_2_m(csr_io_trigger_pkt_any_2_m),
    .io_trigger_pkt_any_2_tdata2(csr_io_trigger_pkt_any_2_tdata2),
    .io_trigger_pkt_any_3_select(csr_io_trigger_pkt_any_3_select),
    .io_trigger_pkt_any_3_match_pkt(csr_io_trigger_pkt_any_3_match_pkt),
    .io_trigger_pkt_any_3_store(csr_io_trigger_pkt_any_3_store),
    .io_trigger_pkt_any_3_load(csr_io_trigger_pkt_any_3_load),
    .io_trigger_pkt_any_3_execute(csr_io_trigger_pkt_any_3_execute),
    .io_trigger_pkt_any_3_m(csr_io_trigger_pkt_any_3_m),
    .io_trigger_pkt_any_3_tdata2(csr_io_trigger_pkt_any_3_tdata2),
    .io_dma_iccm_stall_any(csr_io_dma_iccm_stall_any),
    .io_dma_dccm_stall_any(csr_io_dma_dccm_stall_any),
    .io_lsu_store_stall_any(csr_io_lsu_store_stall_any),
    .io_dec_pmu_presync_stall(csr_io_dec_pmu_presync_stall),
    .io_dec_pmu_postsync_stall(csr_io_dec_pmu_postsync_stall),
    .io_dec_pmu_decode_stall(csr_io_dec_pmu_decode_stall),
    .io_ifu_pmu_fetch_stall(csr_io_ifu_pmu_fetch_stall),
    .io_dec_tlu_packet_r_icaf_type(csr_io_dec_tlu_packet_r_icaf_type),
    .io_dec_tlu_packet_r_pmu_i0_itype(csr_io_dec_tlu_packet_r_pmu_i0_itype),
    .io_dec_tlu_packet_r_pmu_i0_br_unpred(csr_io_dec_tlu_packet_r_pmu_i0_br_unpred),
    .io_dec_tlu_packet_r_pmu_divide(csr_io_dec_tlu_packet_r_pmu_divide),
    .io_dec_tlu_packet_r_pmu_lsu_misaligned(csr_io_dec_tlu_packet_r_pmu_lsu_misaligned),
    .io_exu_pmu_i0_br_ataken(csr_io_exu_pmu_i0_br_ataken),
    .io_exu_pmu_i0_br_misp(csr_io_exu_pmu_i0_br_misp),
    .io_dec_pmu_instr_decoded(csr_io_dec_pmu_instr_decoded),
    .io_ifu_pmu_instr_aligned(csr_io_ifu_pmu_instr_aligned),
    .io_exu_pmu_i0_pc4(csr_io_exu_pmu_i0_pc4),
    .io_ifu_pmu_ic_miss(csr_io_ifu_pmu_ic_miss),
    .io_ifu_pmu_ic_hit(csr_io_ifu_pmu_ic_hit),
    .io_dec_tlu_int_valid_wb1(csr_io_dec_tlu_int_valid_wb1),
    .io_dec_tlu_i0_exc_valid_wb1(csr_io_dec_tlu_i0_exc_valid_wb1),
    .io_dec_tlu_i0_valid_wb1(csr_io_dec_tlu_i0_valid_wb1),
    .io_dec_csr_wen_r(csr_io_dec_csr_wen_r),
    .io_dec_tlu_mtval_wb1(csr_io_dec_tlu_mtval_wb1),
    .io_dec_tlu_exc_cause_wb1(csr_io_dec_tlu_exc_cause_wb1),
    .io_dec_tlu_perfcnt0(csr_io_dec_tlu_perfcnt0),
    .io_dec_tlu_perfcnt1(csr_io_dec_tlu_perfcnt1),
    .io_dec_tlu_perfcnt2(csr_io_dec_tlu_perfcnt2),
    .io_dec_tlu_perfcnt3(csr_io_dec_tlu_perfcnt3),
    .io_dec_tlu_dbg_halted(csr_io_dec_tlu_dbg_halted),
    .io_dma_pmu_dccm_write(csr_io_dma_pmu_dccm_write),
    .io_dma_pmu_dccm_read(csr_io_dma_pmu_dccm_read),
    .io_dma_pmu_any_write(csr_io_dma_pmu_any_write),
    .io_dma_pmu_any_read(csr_io_dma_pmu_any_read),
    .io_lsu_pmu_bus_busy(csr_io_lsu_pmu_bus_busy),
    .io_dec_tlu_i0_pc_r(csr_io_dec_tlu_i0_pc_r),
    .io_dec_tlu_i0_valid_r(csr_io_dec_tlu_i0_valid_r),
    .io_dec_csr_any_unq_d(csr_io_dec_csr_any_unq_d),
    .io_dec_tlu_misc_clk_override(csr_io_dec_tlu_misc_clk_override),
    .io_dec_tlu_dec_clk_override(csr_io_dec_tlu_dec_clk_override),
    .io_dec_tlu_lsu_clk_override(csr_io_dec_tlu_lsu_clk_override),
    .io_dec_tlu_bus_clk_override(csr_io_dec_tlu_bus_clk_override),
    .io_dec_tlu_pic_clk_override(csr_io_dec_tlu_pic_clk_override),
    .io_dec_tlu_dccm_clk_override(csr_io_dec_tlu_dccm_clk_override),
    .io_dec_tlu_icm_clk_override(csr_io_dec_tlu_icm_clk_override),
    .io_dec_csr_rddata_d(csr_io_dec_csr_rddata_d),
    .io_dec_tlu_pipelining_disable(csr_io_dec_tlu_pipelining_disable),
    .io_dec_tlu_wr_pause_r(csr_io_dec_tlu_wr_pause_r),
    .io_ifu_pmu_bus_busy(csr_io_ifu_pmu_bus_busy),
    .io_lsu_pmu_bus_error(csr_io_lsu_pmu_bus_error),
    .io_ifu_pmu_bus_error(csr_io_ifu_pmu_bus_error),
    .io_lsu_pmu_bus_misaligned(csr_io_lsu_pmu_bus_misaligned),
    .io_ifu_ic_debug_rd_data(csr_io_ifu_ic_debug_rd_data),
    .io_dec_tlu_meipt(csr_io_dec_tlu_meipt),
    .io_pic_pl(csr_io_pic_pl),
    .io_dec_tlu_meicurpl(csr_io_dec_tlu_meicurpl),
    .io_dec_tlu_meihap(csr_io_dec_tlu_meihap),
    .io_pic_claimid(csr_io_pic_claimid),
    .io_iccm_dma_sb_error(csr_io_iccm_dma_sb_error),
    .io_lsu_imprecise_error_addr_any(csr_io_lsu_imprecise_error_addr_any),
    .io_lsu_imprecise_error_load_any(csr_io_lsu_imprecise_error_load_any),
    .io_lsu_imprecise_error_store_any(csr_io_lsu_imprecise_error_store_any),
    .io_dec_tlu_mrac_ff(csr_io_dec_tlu_mrac_ff),
    .io_dec_tlu_wb_coalescing_disable(csr_io_dec_tlu_wb_coalescing_disable),
    .io_dec_tlu_bpred_disable(csr_io_dec_tlu_bpred_disable),
    .io_dec_tlu_sideeffect_posted_disable(csr_io_dec_tlu_sideeffect_posted_disable),
    .io_dec_tlu_core_ecc_disable(csr_io_dec_tlu_core_ecc_disable),
    .io_dec_tlu_external_ldfwd_disable(csr_io_dec_tlu_external_ldfwd_disable),
    .io_dec_tlu_dma_qos_prty(csr_io_dec_tlu_dma_qos_prty),
    .io_dec_illegal_inst(csr_io_dec_illegal_inst),
    .io_lsu_error_pkt_r_bits_mscause(csr_io_lsu_error_pkt_r_bits_mscause),
    .io_mexintpend(csr_io_mexintpend),
    .io_exu_npc_r(csr_io_exu_npc_r),
    .io_mpc_reset_run_req(csr_io_mpc_reset_run_req),
    .io_rst_vec(csr_io_rst_vec),
    .io_core_id(csr_io_core_id),
    .io_dec_timer_rddata_d(csr_io_dec_timer_rddata_d),
    .io_dec_timer_read_d(csr_io_dec_timer_read_d),
    .io_dec_csr_wen_r_mod(csr_io_dec_csr_wen_r_mod),
    .io_rfpc_i0_r(csr_io_rfpc_i0_r),
    .io_i0_trigger_hit_r(csr_io_i0_trigger_hit_r),
    .io_fw_halt_req(csr_io_fw_halt_req),
    .io_mstatus(csr_io_mstatus),
    .io_exc_or_int_valid_r(csr_io_exc_or_int_valid_r),
    .io_mret_r(csr_io_mret_r),
    .io_mstatus_mie_ns(csr_io_mstatus_mie_ns),
    .io_dcsr_single_step_running_f(csr_io_dcsr_single_step_running_f),
    .io_dcsr(csr_io_dcsr),
    .io_mtvec(csr_io_mtvec),
    .io_mip(csr_io_mip),
    .io_dec_timer_t0_pulse(csr_io_dec_timer_t0_pulse),
    .io_dec_timer_t1_pulse(csr_io_dec_timer_t1_pulse),
    .io_timer_int_sync(csr_io_timer_int_sync),
    .io_soft_int_sync(csr_io_soft_int_sync),
    .io_mie_ns(csr_io_mie_ns),
    .io_csr_wr_clk(csr_io_csr_wr_clk),
    .io_ebreak_to_debug_mode_r(csr_io_ebreak_to_debug_mode_r),
    .io_dec_tlu_pmu_fw_halted(csr_io_dec_tlu_pmu_fw_halted),
    .io_lsu_fir_error(csr_io_lsu_fir_error),
    .io_npc_r(csr_io_npc_r),
    .io_tlu_flush_lower_r_d1(csr_io_tlu_flush_lower_r_d1),
    .io_dec_tlu_flush_noredir_r_d1(csr_io_dec_tlu_flush_noredir_r_d1),
    .io_tlu_flush_path_r_d1(csr_io_tlu_flush_path_r_d1),
    .io_npc_r_d1(csr_io_npc_r_d1),
    .io_reset_delayed(csr_io_reset_delayed),
    .io_mepc(csr_io_mepc),
    .io_interrupt_valid_r(csr_io_interrupt_valid_r),
    .io_i0_exception_valid_r(csr_io_i0_exception_valid_r),
    .io_lsu_exc_valid_r(csr_io_lsu_exc_valid_r),
    .io_mepc_trigger_hit_sel_pc_r(csr_io_mepc_trigger_hit_sel_pc_r),
    .io_e4e5_int_clk(csr_io_e4e5_int_clk),
    .io_lsu_i0_exc_r(csr_io_lsu_i0_exc_r),
    .io_inst_acc_r(csr_io_inst_acc_r),
    .io_inst_acc_second_r(csr_io_inst_acc_second_r),
    .io_take_nmi(csr_io_take_nmi),
    .io_lsu_error_pkt_addr_r(csr_io_lsu_error_pkt_addr_r),
    .io_exc_cause_r(csr_io_exc_cause_r),
    .io_i0_valid_wb(csr_io_i0_valid_wb),
    .io_exc_or_int_valid_r_d1(csr_io_exc_or_int_valid_r_d1),
    .io_interrupt_valid_r_d1(csr_io_interrupt_valid_r_d1),
    .io_clk_override(csr_io_clk_override),
    .io_i0_exception_valid_r_d1(csr_io_i0_exception_valid_r_d1),
    .io_lsu_i0_exc_r_d1(csr_io_lsu_i0_exc_r_d1),
    .io_exc_cause_wb(csr_io_exc_cause_wb),
    .io_nmi_lsu_store_type(csr_io_nmi_lsu_store_type),
    .io_nmi_lsu_load_type(csr_io_nmi_lsu_load_type),
    .io_tlu_i0_commit_cmt(csr_io_tlu_i0_commit_cmt),
    .io_ebreak_r(csr_io_ebreak_r),
    .io_ecall_r(csr_io_ecall_r),
    .io_illegal_r(csr_io_illegal_r),
    .io_mdseac_locked_ns(csr_io_mdseac_locked_ns),
    .io_mdseac_locked_f(csr_io_mdseac_locked_f),
    .io_nmi_int_detected_f(csr_io_nmi_int_detected_f),
    .io_internal_dbg_halt_mode_f2(csr_io_internal_dbg_halt_mode_f2),
    .io_ext_int_freeze_d1(csr_io_ext_int_freeze_d1),
    .io_ic_perr_r_d1(csr_io_ic_perr_r_d1),
    .io_iccm_sbecc_r_d1(csr_io_iccm_sbecc_r_d1),
    .io_lsu_single_ecc_error_r_d1(csr_io_lsu_single_ecc_error_r_d1),
    .io_ifu_miss_state_idle_f(csr_io_ifu_miss_state_idle_f),
    .io_lsu_idle_any_f(csr_io_lsu_idle_any_f),
    .io_dbg_tlu_halted_f(csr_io_dbg_tlu_halted_f),
    .io_dbg_tlu_halted(csr_io_dbg_tlu_halted),
    .io_debug_halt_req_f(csr_io_debug_halt_req_f),
    .io_force_halt(csr_io_force_halt),
    .io_take_ext_int_start(csr_io_take_ext_int_start),
    .io_trigger_hit_dmode_r_d1(csr_io_trigger_hit_dmode_r_d1),
    .io_trigger_hit_r_d1(csr_io_trigger_hit_r_d1),
    .io_dcsr_single_step_done_f(csr_io_dcsr_single_step_done_f),
    .io_ebreak_to_debug_mode_r_d1(csr_io_ebreak_to_debug_mode_r_d1),
    .io_debug_halt_req(csr_io_debug_halt_req),
    .io_allow_dbg_halt_csr_write(csr_io_allow_dbg_halt_csr_write),
    .io_internal_dbg_halt_mode_f(csr_io_internal_dbg_halt_mode_f),
    .io_enter_debug_halt_req(csr_io_enter_debug_halt_req),
    .io_internal_dbg_halt_mode(csr_io_internal_dbg_halt_mode),
    .io_request_debug_mode_done(csr_io_request_debug_mode_done),
    .io_request_debug_mode_r(csr_io_request_debug_mode_r),
    .io_dpc(csr_io_dpc),
    .io_update_hit_bit_r(csr_io_update_hit_bit_r),
    .io_take_timer_int(csr_io_take_timer_int),
    .io_take_int_timer0_int(csr_io_take_int_timer0_int),
    .io_take_int_timer1_int(csr_io_take_int_timer1_int),
    .io_take_ext_int(csr_io_take_ext_int),
    .io_tlu_flush_lower_r(csr_io_tlu_flush_lower_r),
    .io_dec_tlu_br0_error_r(csr_io_dec_tlu_br0_error_r),
    .io_dec_tlu_br0_start_error_r(csr_io_dec_tlu_br0_start_error_r),
    .io_lsu_pmu_load_external_r(csr_io_lsu_pmu_load_external_r),
    .io_lsu_pmu_store_external_r(csr_io_lsu_pmu_store_external_r),
    .io_csr_pkt_csr_misa(csr_io_csr_pkt_csr_misa),
    .io_csr_pkt_csr_mvendorid(csr_io_csr_pkt_csr_mvendorid),
    .io_csr_pkt_csr_marchid(csr_io_csr_pkt_csr_marchid),
    .io_csr_pkt_csr_mimpid(csr_io_csr_pkt_csr_mimpid),
    .io_csr_pkt_csr_mhartid(csr_io_csr_pkt_csr_mhartid),
    .io_csr_pkt_csr_mstatus(csr_io_csr_pkt_csr_mstatus),
    .io_csr_pkt_csr_mtvec(csr_io_csr_pkt_csr_mtvec),
    .io_csr_pkt_csr_mip(csr_io_csr_pkt_csr_mip),
    .io_csr_pkt_csr_mie(csr_io_csr_pkt_csr_mie),
    .io_csr_pkt_csr_mcyclel(csr_io_csr_pkt_csr_mcyclel),
    .io_csr_pkt_csr_mcycleh(csr_io_csr_pkt_csr_mcycleh),
    .io_csr_pkt_csr_minstretl(csr_io_csr_pkt_csr_minstretl),
    .io_csr_pkt_csr_minstreth(csr_io_csr_pkt_csr_minstreth),
    .io_csr_pkt_csr_mscratch(csr_io_csr_pkt_csr_mscratch),
    .io_csr_pkt_csr_mepc(csr_io_csr_pkt_csr_mepc),
    .io_csr_pkt_csr_mcause(csr_io_csr_pkt_csr_mcause),
    .io_csr_pkt_csr_mscause(csr_io_csr_pkt_csr_mscause),
    .io_csr_pkt_csr_mtval(csr_io_csr_pkt_csr_mtval),
    .io_csr_pkt_csr_mrac(csr_io_csr_pkt_csr_mrac),
    .io_csr_pkt_csr_mdseac(csr_io_csr_pkt_csr_mdseac),
    .io_csr_pkt_csr_meihap(csr_io_csr_pkt_csr_meihap),
    .io_csr_pkt_csr_meivt(csr_io_csr_pkt_csr_meivt),
    .io_csr_pkt_csr_meipt(csr_io_csr_pkt_csr_meipt),
    .io_csr_pkt_csr_meicurpl(csr_io_csr_pkt_csr_meicurpl),
    .io_csr_pkt_csr_meicidpl(csr_io_csr_pkt_csr_meicidpl),
    .io_csr_pkt_csr_dcsr(csr_io_csr_pkt_csr_dcsr),
    .io_csr_pkt_csr_mcgc(csr_io_csr_pkt_csr_mcgc),
    .io_csr_pkt_csr_mfdc(csr_io_csr_pkt_csr_mfdc),
    .io_csr_pkt_csr_dpc(csr_io_csr_pkt_csr_dpc),
    .io_csr_pkt_csr_mtsel(csr_io_csr_pkt_csr_mtsel),
    .io_csr_pkt_csr_mtdata1(csr_io_csr_pkt_csr_mtdata1),
    .io_csr_pkt_csr_mtdata2(csr_io_csr_pkt_csr_mtdata2),
    .io_csr_pkt_csr_mhpmc3(csr_io_csr_pkt_csr_mhpmc3),
    .io_csr_pkt_csr_mhpmc4(csr_io_csr_pkt_csr_mhpmc4),
    .io_csr_pkt_csr_mhpmc5(csr_io_csr_pkt_csr_mhpmc5),
    .io_csr_pkt_csr_mhpmc6(csr_io_csr_pkt_csr_mhpmc6),
    .io_csr_pkt_csr_mhpmc3h(csr_io_csr_pkt_csr_mhpmc3h),
    .io_csr_pkt_csr_mhpmc4h(csr_io_csr_pkt_csr_mhpmc4h),
    .io_csr_pkt_csr_mhpmc5h(csr_io_csr_pkt_csr_mhpmc5h),
    .io_csr_pkt_csr_mhpmc6h(csr_io_csr_pkt_csr_mhpmc6h),
    .io_csr_pkt_csr_mhpme3(csr_io_csr_pkt_csr_mhpme3),
    .io_csr_pkt_csr_mhpme4(csr_io_csr_pkt_csr_mhpme4),
    .io_csr_pkt_csr_mhpme5(csr_io_csr_pkt_csr_mhpme5),
    .io_csr_pkt_csr_mhpme6(csr_io_csr_pkt_csr_mhpme6),
    .io_csr_pkt_csr_mcountinhibit(csr_io_csr_pkt_csr_mcountinhibit),
    .io_csr_pkt_csr_mpmc(csr_io_csr_pkt_csr_mpmc),
    .io_csr_pkt_csr_micect(csr_io_csr_pkt_csr_micect),
    .io_csr_pkt_csr_miccmect(csr_io_csr_pkt_csr_miccmect),
    .io_csr_pkt_csr_mdccmect(csr_io_csr_pkt_csr_mdccmect),
    .io_csr_pkt_csr_mfdht(csr_io_csr_pkt_csr_mfdht),
    .io_csr_pkt_csr_mfdhs(csr_io_csr_pkt_csr_mfdhs),
    .io_csr_pkt_csr_dicawics(csr_io_csr_pkt_csr_dicawics),
    .io_csr_pkt_csr_dicad0h(csr_io_csr_pkt_csr_dicad0h),
    .io_csr_pkt_csr_dicad0(csr_io_csr_pkt_csr_dicad0),
    .io_csr_pkt_csr_dicad1(csr_io_csr_pkt_csr_dicad1),
    .io_mtdata1_t_0(csr_io_mtdata1_t_0),
    .io_mtdata1_t_1(csr_io_mtdata1_t_1),
    .io_mtdata1_t_2(csr_io_mtdata1_t_2),
    .io_mtdata1_t_3(csr_io_mtdata1_t_3)
  );
  dec_decode_csr_read csr_read ( // @[dec_tlu_ctl.scala 1011:22]
    .io_dec_csr_rdaddr_d(csr_read_io_dec_csr_rdaddr_d),
    .io_csr_pkt_csr_misa(csr_read_io_csr_pkt_csr_misa),
    .io_csr_pkt_csr_mvendorid(csr_read_io_csr_pkt_csr_mvendorid),
    .io_csr_pkt_csr_marchid(csr_read_io_csr_pkt_csr_marchid),
    .io_csr_pkt_csr_mimpid(csr_read_io_csr_pkt_csr_mimpid),
    .io_csr_pkt_csr_mhartid(csr_read_io_csr_pkt_csr_mhartid),
    .io_csr_pkt_csr_mstatus(csr_read_io_csr_pkt_csr_mstatus),
    .io_csr_pkt_csr_mtvec(csr_read_io_csr_pkt_csr_mtvec),
    .io_csr_pkt_csr_mip(csr_read_io_csr_pkt_csr_mip),
    .io_csr_pkt_csr_mie(csr_read_io_csr_pkt_csr_mie),
    .io_csr_pkt_csr_mcyclel(csr_read_io_csr_pkt_csr_mcyclel),
    .io_csr_pkt_csr_mcycleh(csr_read_io_csr_pkt_csr_mcycleh),
    .io_csr_pkt_csr_minstretl(csr_read_io_csr_pkt_csr_minstretl),
    .io_csr_pkt_csr_minstreth(csr_read_io_csr_pkt_csr_minstreth),
    .io_csr_pkt_csr_mscratch(csr_read_io_csr_pkt_csr_mscratch),
    .io_csr_pkt_csr_mepc(csr_read_io_csr_pkt_csr_mepc),
    .io_csr_pkt_csr_mcause(csr_read_io_csr_pkt_csr_mcause),
    .io_csr_pkt_csr_mscause(csr_read_io_csr_pkt_csr_mscause),
    .io_csr_pkt_csr_mtval(csr_read_io_csr_pkt_csr_mtval),
    .io_csr_pkt_csr_mrac(csr_read_io_csr_pkt_csr_mrac),
    .io_csr_pkt_csr_dmst(csr_read_io_csr_pkt_csr_dmst),
    .io_csr_pkt_csr_mdseac(csr_read_io_csr_pkt_csr_mdseac),
    .io_csr_pkt_csr_meihap(csr_read_io_csr_pkt_csr_meihap),
    .io_csr_pkt_csr_meivt(csr_read_io_csr_pkt_csr_meivt),
    .io_csr_pkt_csr_meipt(csr_read_io_csr_pkt_csr_meipt),
    .io_csr_pkt_csr_meicurpl(csr_read_io_csr_pkt_csr_meicurpl),
    .io_csr_pkt_csr_meicidpl(csr_read_io_csr_pkt_csr_meicidpl),
    .io_csr_pkt_csr_dcsr(csr_read_io_csr_pkt_csr_dcsr),
    .io_csr_pkt_csr_mcgc(csr_read_io_csr_pkt_csr_mcgc),
    .io_csr_pkt_csr_mfdc(csr_read_io_csr_pkt_csr_mfdc),
    .io_csr_pkt_csr_dpc(csr_read_io_csr_pkt_csr_dpc),
    .io_csr_pkt_csr_mtsel(csr_read_io_csr_pkt_csr_mtsel),
    .io_csr_pkt_csr_mtdata1(csr_read_io_csr_pkt_csr_mtdata1),
    .io_csr_pkt_csr_mtdata2(csr_read_io_csr_pkt_csr_mtdata2),
    .io_csr_pkt_csr_mhpmc3(csr_read_io_csr_pkt_csr_mhpmc3),
    .io_csr_pkt_csr_mhpmc4(csr_read_io_csr_pkt_csr_mhpmc4),
    .io_csr_pkt_csr_mhpmc5(csr_read_io_csr_pkt_csr_mhpmc5),
    .io_csr_pkt_csr_mhpmc6(csr_read_io_csr_pkt_csr_mhpmc6),
    .io_csr_pkt_csr_mhpmc3h(csr_read_io_csr_pkt_csr_mhpmc3h),
    .io_csr_pkt_csr_mhpmc4h(csr_read_io_csr_pkt_csr_mhpmc4h),
    .io_csr_pkt_csr_mhpmc5h(csr_read_io_csr_pkt_csr_mhpmc5h),
    .io_csr_pkt_csr_mhpmc6h(csr_read_io_csr_pkt_csr_mhpmc6h),
    .io_csr_pkt_csr_mhpme3(csr_read_io_csr_pkt_csr_mhpme3),
    .io_csr_pkt_csr_mhpme4(csr_read_io_csr_pkt_csr_mhpme4),
    .io_csr_pkt_csr_mhpme5(csr_read_io_csr_pkt_csr_mhpme5),
    .io_csr_pkt_csr_mhpme6(csr_read_io_csr_pkt_csr_mhpme6),
    .io_csr_pkt_csr_mcountinhibit(csr_read_io_csr_pkt_csr_mcountinhibit),
    .io_csr_pkt_csr_mitctl0(csr_read_io_csr_pkt_csr_mitctl0),
    .io_csr_pkt_csr_mitctl1(csr_read_io_csr_pkt_csr_mitctl1),
    .io_csr_pkt_csr_mitb0(csr_read_io_csr_pkt_csr_mitb0),
    .io_csr_pkt_csr_mitb1(csr_read_io_csr_pkt_csr_mitb1),
    .io_csr_pkt_csr_mitcnt0(csr_read_io_csr_pkt_csr_mitcnt0),
    .io_csr_pkt_csr_mitcnt1(csr_read_io_csr_pkt_csr_mitcnt1),
    .io_csr_pkt_csr_mpmc(csr_read_io_csr_pkt_csr_mpmc),
    .io_csr_pkt_csr_meicpct(csr_read_io_csr_pkt_csr_meicpct),
    .io_csr_pkt_csr_micect(csr_read_io_csr_pkt_csr_micect),
    .io_csr_pkt_csr_miccmect(csr_read_io_csr_pkt_csr_miccmect),
    .io_csr_pkt_csr_mdccmect(csr_read_io_csr_pkt_csr_mdccmect),
    .io_csr_pkt_csr_mfdht(csr_read_io_csr_pkt_csr_mfdht),
    .io_csr_pkt_csr_mfdhs(csr_read_io_csr_pkt_csr_mfdhs),
    .io_csr_pkt_csr_dicawics(csr_read_io_csr_pkt_csr_dicawics),
    .io_csr_pkt_csr_dicad0h(csr_read_io_csr_pkt_csr_dicad0h),
    .io_csr_pkt_csr_dicad0(csr_read_io_csr_pkt_csr_dicad0),
    .io_csr_pkt_csr_dicad1(csr_read_io_csr_pkt_csr_dicad1),
    .io_csr_pkt_csr_dicago(csr_read_io_csr_pkt_csr_dicago),
    .io_csr_pkt_presync(csr_read_io_csr_pkt_presync),
    .io_csr_pkt_postsync(csr_read_io_csr_pkt_postsync),
    .io_csr_pkt_legal(csr_read_io_csr_pkt_legal)
  );
  assign io_tlu_exu_dec_tlu_meihap = csr_io_dec_tlu_meihap; // @[dec_tlu_ctl.scala 877:52]
  assign io_tlu_exu_dec_tlu_flush_lower_r = _T_801 | take_ext_int_start; // @[dec_tlu_ctl.scala 803:49]
  assign io_tlu_exu_dec_tlu_flush_path_r = take_reset ? io_rst_vec : _T_852; // @[dec_tlu_ctl.scala 804:49]
  assign io_tlu_dma_dec_tlu_dma_qos_prty = csr_io_dec_tlu_dma_qos_prty; // @[dec_tlu_ctl.scala 907:48]
  assign io_dec_dbg_cmd_done = io_dec_tlu_i0_valid_r & io_dec_tlu_dbg_halted; // @[dec_tlu_ctl.scala 488:29]
  assign io_dec_dbg_cmd_fail = illegal_r & io_dec_dbg_cmd_done; // @[dec_tlu_ctl.scala 489:29]
  assign io_dec_tlu_dbg_halted = dbg_tlu_halted_f; // @[dec_tlu_ctl.scala 470:41]
  assign io_dec_tlu_debug_mode = debug_mode_status; // @[dec_tlu_ctl.scala 471:41]
  assign io_dec_tlu_resume_ack = _T_190; // @[dec_tlu_ctl.scala 454:49]
  assign io_dec_tlu_debug_stall = debug_halt_req_f; // @[dec_tlu_ctl.scala 469:41]
  assign io_dec_tlu_mpc_halted_only = _T_65; // @[dec_tlu_ctl.scala 369:49]
  assign io_dec_tlu_flush_extint = ext_int_ready & _T_704; // @[dec_tlu_ctl.scala 477:33]
  assign io_trigger_pkt_any_0_select = csr_io_trigger_pkt_any_0_select; // @[dec_tlu_ctl.scala 883:40]
  assign io_trigger_pkt_any_0_match_pkt = csr_io_trigger_pkt_any_0_match_pkt; // @[dec_tlu_ctl.scala 883:40]
  assign io_trigger_pkt_any_0_store = csr_io_trigger_pkt_any_0_store; // @[dec_tlu_ctl.scala 883:40]
  assign io_trigger_pkt_any_0_load = csr_io_trigger_pkt_any_0_load; // @[dec_tlu_ctl.scala 883:40]
  assign io_trigger_pkt_any_0_execute = csr_io_trigger_pkt_any_0_execute; // @[dec_tlu_ctl.scala 883:40]
  assign io_trigger_pkt_any_0_m = csr_io_trigger_pkt_any_0_m; // @[dec_tlu_ctl.scala 883:40]
  assign io_trigger_pkt_any_0_tdata2 = csr_io_trigger_pkt_any_0_tdata2; // @[dec_tlu_ctl.scala 883:40]
  assign io_trigger_pkt_any_1_select = csr_io_trigger_pkt_any_1_select; // @[dec_tlu_ctl.scala 883:40]
  assign io_trigger_pkt_any_1_match_pkt = csr_io_trigger_pkt_any_1_match_pkt; // @[dec_tlu_ctl.scala 883:40]
  assign io_trigger_pkt_any_1_store = csr_io_trigger_pkt_any_1_store; // @[dec_tlu_ctl.scala 883:40]
  assign io_trigger_pkt_any_1_load = csr_io_trigger_pkt_any_1_load; // @[dec_tlu_ctl.scala 883:40]
  assign io_trigger_pkt_any_1_execute = csr_io_trigger_pkt_any_1_execute; // @[dec_tlu_ctl.scala 883:40]
  assign io_trigger_pkt_any_1_m = csr_io_trigger_pkt_any_1_m; // @[dec_tlu_ctl.scala 883:40]
  assign io_trigger_pkt_any_1_tdata2 = csr_io_trigger_pkt_any_1_tdata2; // @[dec_tlu_ctl.scala 883:40]
  assign io_trigger_pkt_any_2_select = csr_io_trigger_pkt_any_2_select; // @[dec_tlu_ctl.scala 883:40]
  assign io_trigger_pkt_any_2_match_pkt = csr_io_trigger_pkt_any_2_match_pkt; // @[dec_tlu_ctl.scala 883:40]
  assign io_trigger_pkt_any_2_store = csr_io_trigger_pkt_any_2_store; // @[dec_tlu_ctl.scala 883:40]
  assign io_trigger_pkt_any_2_load = csr_io_trigger_pkt_any_2_load; // @[dec_tlu_ctl.scala 883:40]
  assign io_trigger_pkt_any_2_execute = csr_io_trigger_pkt_any_2_execute; // @[dec_tlu_ctl.scala 883:40]
  assign io_trigger_pkt_any_2_m = csr_io_trigger_pkt_any_2_m; // @[dec_tlu_ctl.scala 883:40]
  assign io_trigger_pkt_any_2_tdata2 = csr_io_trigger_pkt_any_2_tdata2; // @[dec_tlu_ctl.scala 883:40]
  assign io_trigger_pkt_any_3_select = csr_io_trigger_pkt_any_3_select; // @[dec_tlu_ctl.scala 883:40]
  assign io_trigger_pkt_any_3_match_pkt = csr_io_trigger_pkt_any_3_match_pkt; // @[dec_tlu_ctl.scala 883:40]
  assign io_trigger_pkt_any_3_store = csr_io_trigger_pkt_any_3_store; // @[dec_tlu_ctl.scala 883:40]
  assign io_trigger_pkt_any_3_load = csr_io_trigger_pkt_any_3_load; // @[dec_tlu_ctl.scala 883:40]
  assign io_trigger_pkt_any_3_execute = csr_io_trigger_pkt_any_3_execute; // @[dec_tlu_ctl.scala 883:40]
  assign io_trigger_pkt_any_3_m = csr_io_trigger_pkt_any_3_m; // @[dec_tlu_ctl.scala 883:40]
  assign io_trigger_pkt_any_3_tdata2 = csr_io_trigger_pkt_any_3_tdata2; // @[dec_tlu_ctl.scala 883:40]
  assign io_o_cpu_halt_status = _T_353; // @[dec_tlu_ctl.scala 574:49]
  assign io_o_cpu_halt_ack = _T_354; // @[dec_tlu_ctl.scala 575:49]
  assign io_o_cpu_run_ack = _T_355; // @[dec_tlu_ctl.scala 576:49]
  assign io_o_debug_mode_status = debug_mode_status; // @[dec_tlu_ctl.scala 597:27]
  assign io_mpc_debug_halt_ack = mpc_debug_halt_ack_f; // @[dec_tlu_ctl.scala 394:31]
  assign io_mpc_debug_run_ack = mpc_debug_run_ack_f; // @[dec_tlu_ctl.scala 395:31]
  assign io_debug_brkpt_status = debug_brkpt_status_f; // @[dec_tlu_ctl.scala 396:31]
  assign io_dec_csr_rddata_d = csr_io_dec_csr_rddata_d; // @[dec_tlu_ctl.scala 898:40]
  assign io_dec_csr_legal_d = _T_887 & _T_894; // @[dec_tlu_ctl.scala 1022:20]
  assign io_dec_tlu_i0_kill_writeb_wb = _T_32; // @[dec_tlu_ctl.scala 329:41]
  assign io_dec_tlu_i0_kill_writeb_r = _T_427 | i0_trigger_hit_raw_r; // @[dec_tlu_ctl.scala 335:41]
  assign io_dec_tlu_wr_pause_r = csr_io_dec_tlu_wr_pause_r; // @[dec_tlu_ctl.scala 900:40]
  assign io_dec_tlu_flush_pause_r = _T_208 & _T_209; // @[dec_tlu_ctl.scala 480:34]
  assign io_dec_tlu_presync_d = _T_864 & _T_865; // @[dec_tlu_ctl.scala 1015:23]
  assign io_dec_tlu_postsync_d = csr_pkt_postsync & io_dec_csr_any_unq_d; // @[dec_tlu_ctl.scala 1016:23]
  assign io_dec_tlu_perfcnt0 = csr_io_dec_tlu_perfcnt0; // @[dec_tlu_ctl.scala 886:40]
  assign io_dec_tlu_perfcnt1 = csr_io_dec_tlu_perfcnt1; // @[dec_tlu_ctl.scala 887:40]
  assign io_dec_tlu_perfcnt2 = csr_io_dec_tlu_perfcnt2; // @[dec_tlu_ctl.scala 888:40]
  assign io_dec_tlu_perfcnt3 = csr_io_dec_tlu_perfcnt3; // @[dec_tlu_ctl.scala 889:40]
  assign io_dec_tlu_i0_exc_valid_wb1 = csr_io_dec_tlu_i0_exc_valid_wb1; // @[dec_tlu_ctl.scala 880:44]
  assign io_dec_tlu_i0_valid_wb1 = csr_io_dec_tlu_i0_valid_wb1; // @[dec_tlu_ctl.scala 881:44]
  assign io_dec_tlu_int_valid_wb1 = csr_io_dec_tlu_int_valid_wb1; // @[dec_tlu_ctl.scala 879:44]
  assign io_dec_tlu_exc_cause_wb1 = csr_io_dec_tlu_exc_cause_wb1; // @[dec_tlu_ctl.scala 885:40]
  assign io_dec_tlu_mtval_wb1 = csr_io_dec_tlu_mtval_wb1; // @[dec_tlu_ctl.scala 884:40]
  assign io_dec_tlu_pipelining_disable = csr_io_dec_tlu_pipelining_disable; // @[dec_tlu_ctl.scala 899:40]
  assign io_dec_tlu_misc_clk_override = csr_io_dec_tlu_misc_clk_override; // @[dec_tlu_ctl.scala 890:40]
  assign io_dec_tlu_dec_clk_override = csr_io_dec_tlu_dec_clk_override; // @[dec_tlu_ctl.scala 891:40]
  assign io_dec_tlu_lsu_clk_override = csr_io_dec_tlu_lsu_clk_override; // @[dec_tlu_ctl.scala 893:40]
  assign io_dec_tlu_bus_clk_override = csr_io_dec_tlu_bus_clk_override; // @[dec_tlu_ctl.scala 894:40]
  assign io_dec_tlu_pic_clk_override = csr_io_dec_tlu_pic_clk_override; // @[dec_tlu_ctl.scala 895:40]
  assign io_dec_tlu_dccm_clk_override = csr_io_dec_tlu_dccm_clk_override; // @[dec_tlu_ctl.scala 896:40]
  assign io_dec_tlu_icm_clk_override = csr_io_dec_tlu_icm_clk_override; // @[dec_tlu_ctl.scala 897:40]
  assign io_dec_tlu_flush_lower_wb = tlu_flush_lower_r_d1; // @[dec_tlu_ctl.scala 801:41]
  assign io_tlu_bp_dec_tlu_br0_r_pkt_valid = _T_459 & _T_462; // @[dec_tlu_ctl.scala 653:57]
  assign io_tlu_bp_dec_tlu_br0_r_pkt_bits_hist = io_tlu_exu_exu_i0_br_hist_r; // @[dec_tlu_ctl.scala 650:65]
  assign io_tlu_bp_dec_tlu_br0_r_pkt_bits_br_error = _T_453 & _T_429; // @[dec_tlu_ctl.scala 651:57]
  assign io_tlu_bp_dec_tlu_br0_r_pkt_bits_br_start_error = _T_455 & _T_429; // @[dec_tlu_ctl.scala 652:57]
  assign io_tlu_bp_dec_tlu_br0_r_pkt_bits_way = io_exu_i0_br_way_r; // @[dec_tlu_ctl.scala 654:65]
  assign io_tlu_bp_dec_tlu_br0_r_pkt_bits_middle = io_tlu_exu_exu_i0_br_middle_r; // @[dec_tlu_ctl.scala 655:65]
  assign io_tlu_bp_dec_tlu_flush_leak_one_wb = _T_233 & _T_234; // @[dec_tlu_ctl.scala 484:45]
  assign io_tlu_bp_dec_tlu_bpred_disable = csr_io_dec_tlu_bpred_disable; // @[dec_tlu_ctl.scala 903:47]
  assign io_tlu_ifc_dec_tlu_flush_noredir_wb = _T_205 | take_ext_int_start; // @[dec_tlu_ctl.scala 475:45]
  assign io_tlu_ifc_dec_tlu_mrac_ff = csr_io_dec_tlu_mrac_ff; // @[dec_tlu_ctl.scala 901:48]
  assign io_tlu_mem_dec_tlu_flush_err_wb = io_tlu_exu_dec_tlu_flush_lower_r & _T_433; // @[dec_tlu_ctl.scala 485:41]
  assign io_tlu_mem_dec_tlu_i0_commit_cmt = _T_422 & _T_465; // @[dec_tlu_ctl.scala 628:37]
  assign io_tlu_mem_dec_tlu_force_halt = _T_33; // @[dec_tlu_ctl.scala 331:57]
  assign io_tlu_mem_dec_tlu_fence_i_wb = _T_492 & _T_470; // @[dec_tlu_ctl.scala 673:39]
  assign io_tlu_mem_dec_tlu_ic_diag_pkt_icache_wrdata = csr_io_dec_tlu_ic_diag_pkt_icache_wrdata; // @[dec_tlu_ctl.scala 882:52]
  assign io_tlu_mem_dec_tlu_ic_diag_pkt_icache_dicawics = csr_io_dec_tlu_ic_diag_pkt_icache_dicawics; // @[dec_tlu_ctl.scala 882:52]
  assign io_tlu_mem_dec_tlu_ic_diag_pkt_icache_rd_valid = csr_io_dec_tlu_ic_diag_pkt_icache_rd_valid; // @[dec_tlu_ctl.scala 882:52]
  assign io_tlu_mem_dec_tlu_ic_diag_pkt_icache_wr_valid = csr_io_dec_tlu_ic_diag_pkt_icache_wr_valid; // @[dec_tlu_ctl.scala 882:52]
  assign io_tlu_mem_dec_tlu_core_ecc_disable = csr_io_dec_tlu_core_ecc_disable; // @[dec_tlu_ctl.scala 905:48]
  assign io_tlu_busbuff_dec_tlu_external_ldfwd_disable = csr_io_dec_tlu_external_ldfwd_disable; // @[dec_tlu_ctl.scala 906:52]
  assign io_tlu_busbuff_dec_tlu_wb_coalescing_disable = csr_io_dec_tlu_wb_coalescing_disable; // @[dec_tlu_ctl.scala 902:52]
  assign io_tlu_busbuff_dec_tlu_sideeffect_posted_disable = csr_io_dec_tlu_sideeffect_posted_disable; // @[dec_tlu_ctl.scala 904:52]
  assign io_dec_pic_dec_tlu_meicurpl = csr_io_dec_tlu_meicurpl; // @[dec_tlu_ctl.scala 876:52]
  assign io_dec_pic_dec_tlu_meipt = csr_io_dec_tlu_meipt; // @[dec_tlu_ctl.scala 878:52]
  assign int_timers_clock = clock;
  assign int_timers_reset = reset;
  assign int_timers_io_free_clk = io_free_clk; // @[dec_tlu_ctl.scala 276:57]
  assign int_timers_io_scan_mode = io_scan_mode; // @[dec_tlu_ctl.scala 277:57]
  assign int_timers_io_dec_csr_wen_r_mod = csr_io_dec_csr_wen_r_mod; // @[dec_tlu_ctl.scala 278:49]
  assign int_timers_io_dec_csr_wraddr_r = io_dec_csr_wraddr_r; // @[dec_tlu_ctl.scala 280:49]
  assign int_timers_io_dec_csr_wrdata_r = io_dec_csr_wrdata_r; // @[dec_tlu_ctl.scala 281:49]
  assign int_timers_io_csr_mitctl0 = csr_read_io_csr_pkt_csr_mitctl0; // @[dec_tlu_ctl.scala 282:57]
  assign int_timers_io_csr_mitctl1 = csr_read_io_csr_pkt_csr_mitctl1; // @[dec_tlu_ctl.scala 283:57]
  assign int_timers_io_csr_mitb0 = csr_read_io_csr_pkt_csr_mitb0; // @[dec_tlu_ctl.scala 284:57]
  assign int_timers_io_csr_mitb1 = csr_read_io_csr_pkt_csr_mitb1; // @[dec_tlu_ctl.scala 285:57]
  assign int_timers_io_csr_mitcnt0 = csr_read_io_csr_pkt_csr_mitcnt0; // @[dec_tlu_ctl.scala 286:57]
  assign int_timers_io_csr_mitcnt1 = csr_read_io_csr_pkt_csr_mitcnt1; // @[dec_tlu_ctl.scala 287:57]
  assign int_timers_io_dec_pause_state = io_dec_pause_state; // @[dec_tlu_ctl.scala 288:49]
  assign int_timers_io_dec_tlu_pmu_fw_halted = pmu_fw_tlu_halted_f; // @[dec_tlu_ctl.scala 289:49]
  assign int_timers_io_internal_dbg_halt_timers = debug_mode_status & _T_665; // @[dec_tlu_ctl.scala 290:47]
  assign rvclkhdr_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_io_en = dec_csr_wen_r_mod | io_dec_tlu_dec_clk_override; // @[lib.scala 345:16]
  assign rvclkhdr_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_1_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_1_io_en = _T_11 | io_dec_tlu_dec_clk_override; // @[lib.scala 345:16]
  assign rvclkhdr_1_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_2_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_2_io_en = e4e5_valid | io_dec_tlu_dec_clk_override; // @[lib.scala 345:16]
  assign rvclkhdr_2_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_3_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_3_io_en = e4e5_valid | flush_clkvalid; // @[lib.scala 345:16]
  assign rvclkhdr_3_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign csr_clock = clock;
  assign csr_reset = reset;
  assign csr_io_free_clk = io_free_clk; // @[dec_tlu_ctl.scala 819:44]
  assign csr_io_active_clk = io_active_clk; // @[dec_tlu_ctl.scala 820:44]
  assign csr_io_scan_mode = io_scan_mode; // @[dec_tlu_ctl.scala 821:44]
  assign csr_io_dec_csr_wrdata_r = io_dec_csr_wrdata_r; // @[dec_tlu_ctl.scala 822:44]
  assign csr_io_dec_csr_wraddr_r = io_dec_csr_wraddr_r; // @[dec_tlu_ctl.scala 823:44]
  assign csr_io_dec_csr_rdaddr_d = io_dec_csr_rdaddr_d; // @[dec_tlu_ctl.scala 824:44]
  assign csr_io_dec_csr_wen_unq_d = io_dec_csr_wen_unq_d; // @[dec_tlu_ctl.scala 825:44]
  assign csr_io_dec_i0_decode_d = io_dec_i0_decode_d; // @[dec_tlu_ctl.scala 826:44]
  assign csr_io_ifu_ic_debug_rd_data_valid = io_tlu_mem_ifu_ic_debug_rd_data_valid; // @[dec_tlu_ctl.scala 827:44]
  assign csr_io_dma_iccm_stall_any = io_tlu_dma_dma_iccm_stall_any; // @[dec_tlu_ctl.scala 829:44]
  assign csr_io_dma_dccm_stall_any = io_tlu_dma_dma_dccm_stall_any; // @[dec_tlu_ctl.scala 830:44]
  assign csr_io_lsu_store_stall_any = io_lsu_store_stall_any; // @[dec_tlu_ctl.scala 831:44]
  assign csr_io_dec_pmu_presync_stall = io_dec_pmu_presync_stall; // @[dec_tlu_ctl.scala 832:44]
  assign csr_io_dec_pmu_postsync_stall = io_dec_pmu_postsync_stall; // @[dec_tlu_ctl.scala 833:44]
  assign csr_io_dec_pmu_decode_stall = io_dec_pmu_decode_stall; // @[dec_tlu_ctl.scala 834:44]
  assign csr_io_ifu_pmu_fetch_stall = io_tlu_ifc_ifu_pmu_fetch_stall; // @[dec_tlu_ctl.scala 835:44]
  assign csr_io_dec_tlu_packet_r_icaf_type = io_dec_tlu_packet_r_icaf_type; // @[dec_tlu_ctl.scala 836:44]
  assign csr_io_dec_tlu_packet_r_pmu_i0_itype = io_dec_tlu_packet_r_pmu_i0_itype; // @[dec_tlu_ctl.scala 836:44]
  assign csr_io_dec_tlu_packet_r_pmu_i0_br_unpred = io_dec_tlu_packet_r_pmu_i0_br_unpred; // @[dec_tlu_ctl.scala 836:44]
  assign csr_io_dec_tlu_packet_r_pmu_divide = io_dec_tlu_packet_r_pmu_divide; // @[dec_tlu_ctl.scala 836:44]
  assign csr_io_dec_tlu_packet_r_pmu_lsu_misaligned = io_dec_tlu_packet_r_pmu_lsu_misaligned; // @[dec_tlu_ctl.scala 836:44]
  assign csr_io_exu_pmu_i0_br_ataken = io_tlu_exu_exu_pmu_i0_br_ataken; // @[dec_tlu_ctl.scala 837:44]
  assign csr_io_exu_pmu_i0_br_misp = io_tlu_exu_exu_pmu_i0_br_misp; // @[dec_tlu_ctl.scala 838:44]
  assign csr_io_dec_pmu_instr_decoded = io_dec_pmu_instr_decoded; // @[dec_tlu_ctl.scala 839:44]
  assign csr_io_ifu_pmu_instr_aligned = io_ifu_pmu_instr_aligned; // @[dec_tlu_ctl.scala 840:44]
  assign csr_io_exu_pmu_i0_pc4 = io_tlu_exu_exu_pmu_i0_pc4; // @[dec_tlu_ctl.scala 841:44]
  assign csr_io_ifu_pmu_ic_miss = io_tlu_mem_ifu_pmu_ic_miss; // @[dec_tlu_ctl.scala 842:44]
  assign csr_io_ifu_pmu_ic_hit = io_tlu_mem_ifu_pmu_ic_hit; // @[dec_tlu_ctl.scala 843:44]
  assign csr_io_dec_csr_wen_r = io_dec_csr_wen_r; // @[dec_tlu_ctl.scala 844:44]
  assign csr_io_dec_tlu_dbg_halted = io_dec_tlu_dbg_halted; // @[dec_tlu_ctl.scala 845:44]
  assign csr_io_dma_pmu_dccm_write = io_tlu_dma_dma_pmu_dccm_write; // @[dec_tlu_ctl.scala 846:44]
  assign csr_io_dma_pmu_dccm_read = io_tlu_dma_dma_pmu_dccm_read; // @[dec_tlu_ctl.scala 847:44]
  assign csr_io_dma_pmu_any_write = io_tlu_dma_dma_pmu_any_write; // @[dec_tlu_ctl.scala 848:44]
  assign csr_io_dma_pmu_any_read = io_tlu_dma_dma_pmu_any_read; // @[dec_tlu_ctl.scala 849:44]
  assign csr_io_lsu_pmu_bus_busy = io_tlu_busbuff_lsu_pmu_bus_busy; // @[dec_tlu_ctl.scala 850:44]
  assign csr_io_dec_tlu_i0_pc_r = io_dec_tlu_i0_pc_r; // @[dec_tlu_ctl.scala 851:44]
  assign csr_io_dec_tlu_i0_valid_r = io_dec_tlu_i0_valid_r; // @[dec_tlu_ctl.scala 852:44]
  assign csr_io_dec_csr_any_unq_d = io_dec_csr_any_unq_d; // @[dec_tlu_ctl.scala 854:44]
  assign csr_io_ifu_pmu_bus_busy = io_tlu_mem_ifu_pmu_bus_busy; // @[dec_tlu_ctl.scala 855:44]
  assign csr_io_lsu_pmu_bus_error = io_tlu_busbuff_lsu_pmu_bus_error; // @[dec_tlu_ctl.scala 856:44]
  assign csr_io_ifu_pmu_bus_error = io_tlu_mem_ifu_pmu_bus_error; // @[dec_tlu_ctl.scala 857:44]
  assign csr_io_lsu_pmu_bus_misaligned = io_tlu_busbuff_lsu_pmu_bus_misaligned; // @[dec_tlu_ctl.scala 858:44]
  assign csr_io_ifu_ic_debug_rd_data = io_tlu_mem_ifu_ic_debug_rd_data; // @[dec_tlu_ctl.scala 860:44]
  assign csr_io_pic_pl = io_dec_pic_pic_pl; // @[dec_tlu_ctl.scala 861:44]
  assign csr_io_pic_claimid = io_dec_pic_pic_claimid; // @[dec_tlu_ctl.scala 862:44]
  assign csr_io_iccm_dma_sb_error = io_iccm_dma_sb_error; // @[dec_tlu_ctl.scala 863:44]
  assign csr_io_lsu_imprecise_error_addr_any = io_tlu_busbuff_lsu_imprecise_error_addr_any; // @[dec_tlu_ctl.scala 864:44]
  assign csr_io_lsu_imprecise_error_load_any = io_tlu_busbuff_lsu_imprecise_error_load_any; // @[dec_tlu_ctl.scala 865:44]
  assign csr_io_lsu_imprecise_error_store_any = io_tlu_busbuff_lsu_imprecise_error_store_any; // @[dec_tlu_ctl.scala 866:44]
  assign csr_io_dec_illegal_inst = io_dec_illegal_inst; // @[dec_tlu_ctl.scala 867:44 dec_tlu_ctl.scala 908:44]
  assign csr_io_lsu_error_pkt_r_bits_mscause = io_lsu_error_pkt_r_bits_mscause; // @[dec_tlu_ctl.scala 868:44 dec_tlu_ctl.scala 909:44]
  assign csr_io_mexintpend = io_dec_pic_mexintpend; // @[dec_tlu_ctl.scala 869:44 dec_tlu_ctl.scala 910:44]
  assign csr_io_exu_npc_r = io_tlu_exu_exu_npc_r; // @[dec_tlu_ctl.scala 870:44 dec_tlu_ctl.scala 911:44]
  assign csr_io_mpc_reset_run_req = io_mpc_reset_run_req; // @[dec_tlu_ctl.scala 871:44 dec_tlu_ctl.scala 912:44]
  assign csr_io_rst_vec = io_rst_vec; // @[dec_tlu_ctl.scala 872:44 dec_tlu_ctl.scala 913:44]
  assign csr_io_core_id = io_core_id; // @[dec_tlu_ctl.scala 873:44 dec_tlu_ctl.scala 914:44]
  assign csr_io_dec_timer_rddata_d = int_timers_io_dec_timer_rddata_d; // @[dec_tlu_ctl.scala 874:44 dec_tlu_ctl.scala 915:44]
  assign csr_io_dec_timer_read_d = int_timers_io_dec_timer_read_d; // @[dec_tlu_ctl.scala 875:44 dec_tlu_ctl.scala 916:44]
  assign csr_io_rfpc_i0_r = _T_438 & _T_439; // @[dec_tlu_ctl.scala 919:39]
  assign csr_io_i0_trigger_hit_r = |i0_trigger_chain_masked_r; // @[dec_tlu_ctl.scala 920:39]
  assign csr_io_exc_or_int_valid_r = _T_855 | mepc_trigger_hit_sel_pc_r; // @[dec_tlu_ctl.scala 921:39]
  assign csr_io_mret_r = _T_487 & _T_470; // @[dec_tlu_ctl.scala 922:39]
  assign csr_io_dcsr_single_step_running_f = dcsr_single_step_running_f; // @[dec_tlu_ctl.scala 923:39]
  assign csr_io_dec_timer_t0_pulse = int_timers_io_dec_timer_t0_pulse; // @[dec_tlu_ctl.scala 924:39]
  assign csr_io_dec_timer_t1_pulse = int_timers_io_dec_timer_t1_pulse; // @[dec_tlu_ctl.scala 925:39]
  assign csr_io_timer_int_sync = syncro_ff[5]; // @[dec_tlu_ctl.scala 926:39]
  assign csr_io_soft_int_sync = syncro_ff[4]; // @[dec_tlu_ctl.scala 927:39]
  assign csr_io_csr_wr_clk = rvclkhdr_io_l1clk; // @[dec_tlu_ctl.scala 928:39]
  assign csr_io_ebreak_to_debug_mode_r = _T_519 & _T_470; // @[dec_tlu_ctl.scala 929:39]
  assign csr_io_dec_tlu_pmu_fw_halted = pmu_fw_tlu_halted_f; // @[dec_tlu_ctl.scala 930:39]
  assign csr_io_lsu_fir_error = io_lsu_fir_error; // @[dec_tlu_ctl.scala 931:39]
  assign csr_io_tlu_flush_lower_r_d1 = tlu_flush_lower_r_d1; // @[dec_tlu_ctl.scala 932:39]
  assign csr_io_dec_tlu_flush_noredir_r_d1 = dec_tlu_flush_noredir_r_d1; // @[dec_tlu_ctl.scala 933:39]
  assign csr_io_tlu_flush_path_r_d1 = tlu_flush_path_r_d1; // @[dec_tlu_ctl.scala 934:39]
  assign csr_io_reset_delayed = reset_detect ^ reset_detected; // @[dec_tlu_ctl.scala 935:39]
  assign csr_io_interrupt_valid_r = _T_766 | take_int_timer1_int; // @[dec_tlu_ctl.scala 936:39]
  assign csr_io_i0_exception_valid_r = _T_527 & _T_528; // @[dec_tlu_ctl.scala 937:39]
  assign csr_io_lsu_exc_valid_r = _T_405 & _T_470; // @[dec_tlu_ctl.scala 938:39]
  assign csr_io_mepc_trigger_hit_sel_pc_r = i0_trigger_hit_raw_r & _T_345; // @[dec_tlu_ctl.scala 939:39]
  assign csr_io_e4e5_int_clk = rvclkhdr_3_io_l1clk; // @[dec_tlu_ctl.scala 940:39]
  assign csr_io_lsu_i0_exc_r = _T_405 & _T_470; // @[dec_tlu_ctl.scala 941:39]
  assign csr_io_inst_acc_r = _T_511 & _T_465; // @[dec_tlu_ctl.scala 942:39]
  assign csr_io_inst_acc_second_r = io_dec_tlu_packet_r_icaf_f1; // @[dec_tlu_ctl.scala 943:39]
  assign csr_io_take_nmi = _T_756 & _T_760; // @[dec_tlu_ctl.scala 944:39]
  assign csr_io_lsu_error_pkt_addr_r = io_lsu_error_pkt_r_bits_addr; // @[dec_tlu_ctl.scala 945:39]
  assign csr_io_exc_cause_r = _T_603 | _T_591; // @[dec_tlu_ctl.scala 946:39]
  assign csr_io_i0_valid_wb = i0_valid_wb; // @[dec_tlu_ctl.scala 947:39]
  assign csr_io_exc_or_int_valid_r_d1 = exc_or_int_valid_r_d1; // @[dec_tlu_ctl.scala 948:39]
  assign csr_io_interrupt_valid_r_d1 = interrupt_valid_r_d1; // @[dec_tlu_ctl.scala 949:39]
  assign csr_io_clk_override = io_dec_tlu_dec_clk_override; // @[dec_tlu_ctl.scala 950:39]
  assign csr_io_i0_exception_valid_r_d1 = i0_exception_valid_r_d1; // @[dec_tlu_ctl.scala 951:39]
  assign csr_io_lsu_i0_exc_r_d1 = lsu_i0_exc_r_d1; // @[dec_tlu_ctl.scala 952:39]
  assign csr_io_exc_cause_wb = exc_cause_wb; // @[dec_tlu_ctl.scala 953:39]
  assign csr_io_nmi_lsu_store_type = _T_58 | _T_60; // @[dec_tlu_ctl.scala 954:39]
  assign csr_io_nmi_lsu_load_type = _T_50 | _T_52; // @[dec_tlu_ctl.scala 955:39]
  assign csr_io_tlu_i0_commit_cmt = _T_422 & _T_465; // @[dec_tlu_ctl.scala 956:39]
  assign csr_io_ebreak_r = _T_469 & _T_470; // @[dec_tlu_ctl.scala 957:39]
  assign csr_io_ecall_r = _T_475 & _T_470; // @[dec_tlu_ctl.scala 958:39]
  assign csr_io_illegal_r = _T_481 & _T_470; // @[dec_tlu_ctl.scala 959:39]
  assign csr_io_mdseac_locked_f = mdseac_locked_f; // @[dec_tlu_ctl.scala 960:39]
  assign csr_io_nmi_int_detected_f = nmi_int_detected_f; // @[dec_tlu_ctl.scala 961:39]
  assign csr_io_internal_dbg_halt_mode_f2 = internal_dbg_halt_mode_f2; // @[dec_tlu_ctl.scala 962:39]
  assign csr_io_ext_int_freeze_d1 = ext_int_freeze_d1; // @[dec_tlu_ctl.scala 963:39]
  assign csr_io_ic_perr_r_d1 = ic_perr_r_d1; // @[dec_tlu_ctl.scala 964:39]
  assign csr_io_iccm_sbecc_r_d1 = iccm_sbecc_r_d1; // @[dec_tlu_ctl.scala 965:39]
  assign csr_io_lsu_single_ecc_error_r_d1 = lsu_single_ecc_error_r_d1; // @[dec_tlu_ctl.scala 966:39]
  assign csr_io_ifu_miss_state_idle_f = ifu_miss_state_idle_f; // @[dec_tlu_ctl.scala 967:39]
  assign csr_io_lsu_idle_any_f = lsu_idle_any_f; // @[dec_tlu_ctl.scala 968:39]
  assign csr_io_dbg_tlu_halted_f = dbg_tlu_halted_f; // @[dec_tlu_ctl.scala 969:39]
  assign csr_io_dbg_tlu_halted = _T_164 | _T_166; // @[dec_tlu_ctl.scala 970:39]
  assign csr_io_debug_halt_req_f = debug_halt_req_f; // @[dec_tlu_ctl.scala 971:51]
  assign csr_io_take_ext_int_start = ext_int_ready & _T_704; // @[dec_tlu_ctl.scala 972:47]
  assign csr_io_trigger_hit_dmode_r_d1 = trigger_hit_dmode_r_d1; // @[dec_tlu_ctl.scala 973:43]
  assign csr_io_trigger_hit_r_d1 = trigger_hit_r_d1; // @[dec_tlu_ctl.scala 974:43]
  assign csr_io_dcsr_single_step_done_f = dcsr_single_step_done_f; // @[dec_tlu_ctl.scala 975:43]
  assign csr_io_ebreak_to_debug_mode_r_d1 = ebreak_to_debug_mode_r_d1; // @[dec_tlu_ctl.scala 976:39]
  assign csr_io_debug_halt_req = _T_114 & _T_107; // @[dec_tlu_ctl.scala 977:51]
  assign csr_io_allow_dbg_halt_csr_write = debug_mode_status & _T_77; // @[dec_tlu_ctl.scala 978:39]
  assign csr_io_internal_dbg_halt_mode_f = debug_mode_status; // @[dec_tlu_ctl.scala 979:39]
  assign csr_io_enter_debug_halt_req = _T_155 | ebreak_to_debug_mode_r_d1; // @[dec_tlu_ctl.scala 980:39]
  assign csr_io_internal_dbg_halt_mode = debug_halt_req_ns | _T_160; // @[dec_tlu_ctl.scala 981:39]
  assign csr_io_request_debug_mode_done = _T_183 & _T_136; // @[dec_tlu_ctl.scala 982:39]
  assign csr_io_request_debug_mode_r = _T_180 | _T_182; // @[dec_tlu_ctl.scala 983:39]
  assign csr_io_update_hit_bit_r = _T_342 & i0_trigger_chain_masked_r; // @[dec_tlu_ctl.scala 984:39]
  assign csr_io_take_timer_int = _T_703 & _T_704; // @[dec_tlu_ctl.scala 985:39]
  assign csr_io_take_int_timer0_int = _T_717 & _T_704; // @[dec_tlu_ctl.scala 986:39]
  assign csr_io_take_int_timer1_int = _T_734 & _T_704; // @[dec_tlu_ctl.scala 987:39]
  assign csr_io_take_ext_int = take_ext_int_start_d3 & _T_685; // @[dec_tlu_ctl.scala 988:39]
  assign csr_io_tlu_flush_lower_r = _T_801 | take_ext_int_start; // @[dec_tlu_ctl.scala 989:39]
  assign csr_io_dec_tlu_br0_error_r = _T_453 & _T_429; // @[dec_tlu_ctl.scala 990:39]
  assign csr_io_dec_tlu_br0_start_error_r = _T_455 & _T_429; // @[dec_tlu_ctl.scala 991:39]
  assign csr_io_lsu_pmu_load_external_r = lsu_pmu_load_external_r; // @[dec_tlu_ctl.scala 992:39]
  assign csr_io_lsu_pmu_store_external_r = lsu_pmu_store_external_r; // @[dec_tlu_ctl.scala 993:39]
  assign csr_io_csr_pkt_csr_misa = csr_read_io_csr_pkt_csr_misa; // @[dec_tlu_ctl.scala 994:39]
  assign csr_io_csr_pkt_csr_mvendorid = csr_read_io_csr_pkt_csr_mvendorid; // @[dec_tlu_ctl.scala 994:39]
  assign csr_io_csr_pkt_csr_marchid = csr_read_io_csr_pkt_csr_marchid; // @[dec_tlu_ctl.scala 994:39]
  assign csr_io_csr_pkt_csr_mimpid = csr_read_io_csr_pkt_csr_mimpid; // @[dec_tlu_ctl.scala 994:39]
  assign csr_io_csr_pkt_csr_mhartid = csr_read_io_csr_pkt_csr_mhartid; // @[dec_tlu_ctl.scala 994:39]
  assign csr_io_csr_pkt_csr_mstatus = csr_read_io_csr_pkt_csr_mstatus; // @[dec_tlu_ctl.scala 994:39]
  assign csr_io_csr_pkt_csr_mtvec = csr_read_io_csr_pkt_csr_mtvec; // @[dec_tlu_ctl.scala 994:39]
  assign csr_io_csr_pkt_csr_mip = csr_read_io_csr_pkt_csr_mip; // @[dec_tlu_ctl.scala 994:39]
  assign csr_io_csr_pkt_csr_mie = csr_read_io_csr_pkt_csr_mie; // @[dec_tlu_ctl.scala 994:39]
  assign csr_io_csr_pkt_csr_mcyclel = csr_read_io_csr_pkt_csr_mcyclel; // @[dec_tlu_ctl.scala 994:39]
  assign csr_io_csr_pkt_csr_mcycleh = csr_read_io_csr_pkt_csr_mcycleh; // @[dec_tlu_ctl.scala 994:39]
  assign csr_io_csr_pkt_csr_minstretl = csr_read_io_csr_pkt_csr_minstretl; // @[dec_tlu_ctl.scala 994:39]
  assign csr_io_csr_pkt_csr_minstreth = csr_read_io_csr_pkt_csr_minstreth; // @[dec_tlu_ctl.scala 994:39]
  assign csr_io_csr_pkt_csr_mscratch = csr_read_io_csr_pkt_csr_mscratch; // @[dec_tlu_ctl.scala 994:39]
  assign csr_io_csr_pkt_csr_mepc = csr_read_io_csr_pkt_csr_mepc; // @[dec_tlu_ctl.scala 994:39]
  assign csr_io_csr_pkt_csr_mcause = csr_read_io_csr_pkt_csr_mcause; // @[dec_tlu_ctl.scala 994:39]
  assign csr_io_csr_pkt_csr_mscause = csr_read_io_csr_pkt_csr_mscause; // @[dec_tlu_ctl.scala 994:39]
  assign csr_io_csr_pkt_csr_mtval = csr_read_io_csr_pkt_csr_mtval; // @[dec_tlu_ctl.scala 994:39]
  assign csr_io_csr_pkt_csr_mrac = csr_read_io_csr_pkt_csr_mrac; // @[dec_tlu_ctl.scala 994:39]
  assign csr_io_csr_pkt_csr_mdseac = csr_read_io_csr_pkt_csr_mdseac; // @[dec_tlu_ctl.scala 994:39]
  assign csr_io_csr_pkt_csr_meihap = csr_read_io_csr_pkt_csr_meihap; // @[dec_tlu_ctl.scala 994:39]
  assign csr_io_csr_pkt_csr_meivt = csr_read_io_csr_pkt_csr_meivt; // @[dec_tlu_ctl.scala 994:39]
  assign csr_io_csr_pkt_csr_meipt = csr_read_io_csr_pkt_csr_meipt; // @[dec_tlu_ctl.scala 994:39]
  assign csr_io_csr_pkt_csr_meicurpl = csr_read_io_csr_pkt_csr_meicurpl; // @[dec_tlu_ctl.scala 994:39]
  assign csr_io_csr_pkt_csr_meicidpl = csr_read_io_csr_pkt_csr_meicidpl; // @[dec_tlu_ctl.scala 994:39]
  assign csr_io_csr_pkt_csr_dcsr = csr_read_io_csr_pkt_csr_dcsr; // @[dec_tlu_ctl.scala 994:39]
  assign csr_io_csr_pkt_csr_mcgc = csr_read_io_csr_pkt_csr_mcgc; // @[dec_tlu_ctl.scala 994:39]
  assign csr_io_csr_pkt_csr_mfdc = csr_read_io_csr_pkt_csr_mfdc; // @[dec_tlu_ctl.scala 994:39]
  assign csr_io_csr_pkt_csr_dpc = csr_read_io_csr_pkt_csr_dpc; // @[dec_tlu_ctl.scala 994:39]
  assign csr_io_csr_pkt_csr_mtsel = csr_read_io_csr_pkt_csr_mtsel; // @[dec_tlu_ctl.scala 994:39]
  assign csr_io_csr_pkt_csr_mtdata1 = csr_read_io_csr_pkt_csr_mtdata1; // @[dec_tlu_ctl.scala 994:39]
  assign csr_io_csr_pkt_csr_mtdata2 = csr_read_io_csr_pkt_csr_mtdata2; // @[dec_tlu_ctl.scala 994:39]
  assign csr_io_csr_pkt_csr_mhpmc3 = csr_read_io_csr_pkt_csr_mhpmc3; // @[dec_tlu_ctl.scala 994:39]
  assign csr_io_csr_pkt_csr_mhpmc4 = csr_read_io_csr_pkt_csr_mhpmc4; // @[dec_tlu_ctl.scala 994:39]
  assign csr_io_csr_pkt_csr_mhpmc5 = csr_read_io_csr_pkt_csr_mhpmc5; // @[dec_tlu_ctl.scala 994:39]
  assign csr_io_csr_pkt_csr_mhpmc6 = csr_read_io_csr_pkt_csr_mhpmc6; // @[dec_tlu_ctl.scala 994:39]
  assign csr_io_csr_pkt_csr_mhpmc3h = csr_read_io_csr_pkt_csr_mhpmc3h; // @[dec_tlu_ctl.scala 994:39]
  assign csr_io_csr_pkt_csr_mhpmc4h = csr_read_io_csr_pkt_csr_mhpmc4h; // @[dec_tlu_ctl.scala 994:39]
  assign csr_io_csr_pkt_csr_mhpmc5h = csr_read_io_csr_pkt_csr_mhpmc5h; // @[dec_tlu_ctl.scala 994:39]
  assign csr_io_csr_pkt_csr_mhpmc6h = csr_read_io_csr_pkt_csr_mhpmc6h; // @[dec_tlu_ctl.scala 994:39]
  assign csr_io_csr_pkt_csr_mhpme3 = csr_read_io_csr_pkt_csr_mhpme3; // @[dec_tlu_ctl.scala 994:39]
  assign csr_io_csr_pkt_csr_mhpme4 = csr_read_io_csr_pkt_csr_mhpme4; // @[dec_tlu_ctl.scala 994:39]
  assign csr_io_csr_pkt_csr_mhpme5 = csr_read_io_csr_pkt_csr_mhpme5; // @[dec_tlu_ctl.scala 994:39]
  assign csr_io_csr_pkt_csr_mhpme6 = csr_read_io_csr_pkt_csr_mhpme6; // @[dec_tlu_ctl.scala 994:39]
  assign csr_io_csr_pkt_csr_mcountinhibit = csr_read_io_csr_pkt_csr_mcountinhibit; // @[dec_tlu_ctl.scala 994:39]
  assign csr_io_csr_pkt_csr_mpmc = csr_read_io_csr_pkt_csr_mpmc; // @[dec_tlu_ctl.scala 994:39]
  assign csr_io_csr_pkt_csr_micect = csr_read_io_csr_pkt_csr_micect; // @[dec_tlu_ctl.scala 994:39]
  assign csr_io_csr_pkt_csr_miccmect = csr_read_io_csr_pkt_csr_miccmect; // @[dec_tlu_ctl.scala 994:39]
  assign csr_io_csr_pkt_csr_mdccmect = csr_read_io_csr_pkt_csr_mdccmect; // @[dec_tlu_ctl.scala 994:39]
  assign csr_io_csr_pkt_csr_mfdht = csr_read_io_csr_pkt_csr_mfdht; // @[dec_tlu_ctl.scala 994:39]
  assign csr_io_csr_pkt_csr_mfdhs = csr_read_io_csr_pkt_csr_mfdhs; // @[dec_tlu_ctl.scala 994:39]
  assign csr_io_csr_pkt_csr_dicawics = csr_read_io_csr_pkt_csr_dicawics; // @[dec_tlu_ctl.scala 994:39]
  assign csr_io_csr_pkt_csr_dicad0h = csr_read_io_csr_pkt_csr_dicad0h; // @[dec_tlu_ctl.scala 994:39]
  assign csr_io_csr_pkt_csr_dicad0 = csr_read_io_csr_pkt_csr_dicad0; // @[dec_tlu_ctl.scala 994:39]
  assign csr_io_csr_pkt_csr_dicad1 = csr_read_io_csr_pkt_csr_dicad1; // @[dec_tlu_ctl.scala 994:39]
  assign csr_read_io_dec_csr_rdaddr_d = io_dec_csr_rdaddr_d; // @[dec_tlu_ctl.scala 1012:37]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  dbg_halt_state_f = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  mpc_halt_state_f = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  _T_8 = _RAND_2[6:0];
  _RAND_3 = {1{`RANDOM}};
  syncro_ff = _RAND_3[6:0];
  _RAND_4 = {1{`RANDOM}};
  lsu_exc_valid_r_d1 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  e5_valid = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  debug_mode_status = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  i_cpu_run_req_d1_raw = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  nmi_int_delayed = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  mdseac_locked_f = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  nmi_int_detected_f = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  take_nmi_r_d1 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  take_ext_int_start_d3 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  int_timer0_int_hold_f = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  int_timer1_int_hold_f = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  i_cpu_halt_req_d1 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  dbg_halt_req_held = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  ext_int_freeze_d1 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  reset_detect = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  reset_detected = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  dcsr_single_step_done_f = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  trigger_hit_dmode_r_d1 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  ebreak_to_debug_mode_r_d1 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  debug_halt_req_f = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  lsu_idle_any_f = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  ifu_miss_state_idle_f = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  debug_halt_req_d1 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  dec_tlu_flush_noredir_r_d1 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  dec_tlu_flush_pause_r_d1 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  take_ext_int_start_d1 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  halt_taken_f = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  dbg_tlu_halted_f = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  pmu_fw_tlu_halted_f = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  interrupt_valid_r_d1 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  debug_resume_req_f = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  dcsr_single_step_running_f = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  pmu_fw_halt_req_f = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  internal_pmu_fw_halt_mode_f = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  tlu_flush_lower_r_d1 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  ic_perr_r_d1 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  iccm_sbecc_r_d1 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  request_debug_mode_r_d1 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  iccm_repair_state_d1 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  dec_pause_state_f = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  dec_tlu_wr_pause_r_d1 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  exc_or_int_valid_r_d1 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  pause_expired_wb = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  lsu_pmu_load_external_r = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  lsu_pmu_store_external_r = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  _T_32 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  internal_dbg_halt_mode_f2 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  _T_33 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  nmi_lsu_load_type_f = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  nmi_lsu_store_type_f = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  mpc_debug_halt_req_sync_f = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  mpc_debug_run_req_sync_f = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  mpc_run_state_f = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  debug_brkpt_status_f = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  mpc_debug_halt_ack_f = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  mpc_debug_run_ack_f = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  dbg_run_state_f = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  _T_65 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  request_debug_mode_done_f = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  _T_190 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  _T_353 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  _T_354 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  _T_355 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  lsu_single_ecc_error_r_d1 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  lsu_i0_exc_r_d1 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  take_ext_int_start_d2 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  tlu_flush_path_r_d1 = _RAND_70[30:0];
  _RAND_71 = {1{`RANDOM}};
  i0_exception_valid_r_d1 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  exc_cause_wb = _RAND_72[4:0];
  _RAND_73 = {1{`RANDOM}};
  i0_valid_wb = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  trigger_hit_r_d1 = _RAND_74[0:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    dbg_halt_state_f = 1'h0;
  end
  if (reset) begin
    mpc_halt_state_f = 1'h0;
  end
  if (reset) begin
    _T_8 = 7'h0;
  end
  if (reset) begin
    syncro_ff = 7'h0;
  end
  if (reset) begin
    lsu_exc_valid_r_d1 = 1'h0;
  end
  if (reset) begin
    e5_valid = 1'h0;
  end
  if (reset) begin
    debug_mode_status = 1'h0;
  end
  if (reset) begin
    i_cpu_run_req_d1_raw = 1'h0;
  end
  if (reset) begin
    nmi_int_delayed = 1'h0;
  end
  if (reset) begin
    mdseac_locked_f = 1'h0;
  end
  if (reset) begin
    nmi_int_detected_f = 1'h0;
  end
  if (reset) begin
    take_nmi_r_d1 = 1'h0;
  end
  if (reset) begin
    take_ext_int_start_d3 = 1'h0;
  end
  if (reset) begin
    int_timer0_int_hold_f = 1'h0;
  end
  if (reset) begin
    int_timer1_int_hold_f = 1'h0;
  end
  if (reset) begin
    i_cpu_halt_req_d1 = 1'h0;
  end
  if (reset) begin
    dbg_halt_req_held = 1'h0;
  end
  if (reset) begin
    ext_int_freeze_d1 = 1'h0;
  end
  if (reset) begin
    reset_detect = 1'h0;
  end
  if (reset) begin
    reset_detected = 1'h0;
  end
  if (reset) begin
    dcsr_single_step_done_f = 1'h0;
  end
  if (reset) begin
    trigger_hit_dmode_r_d1 = 1'h0;
  end
  if (reset) begin
    ebreak_to_debug_mode_r_d1 = 1'h0;
  end
  if (reset) begin
    debug_halt_req_f = 1'h0;
  end
  if (reset) begin
    lsu_idle_any_f = 1'h0;
  end
  if (reset) begin
    ifu_miss_state_idle_f = 1'h0;
  end
  if (reset) begin
    debug_halt_req_d1 = 1'h0;
  end
  if (reset) begin
    dec_tlu_flush_noredir_r_d1 = 1'h0;
  end
  if (reset) begin
    dec_tlu_flush_pause_r_d1 = 1'h0;
  end
  if (reset) begin
    take_ext_int_start_d1 = 1'h0;
  end
  if (reset) begin
    halt_taken_f = 1'h0;
  end
  if (reset) begin
    dbg_tlu_halted_f = 1'h0;
  end
  if (reset) begin
    pmu_fw_tlu_halted_f = 1'h0;
  end
  if (reset) begin
    interrupt_valid_r_d1 = 1'h0;
  end
  if (reset) begin
    debug_resume_req_f = 1'h0;
  end
  if (reset) begin
    dcsr_single_step_running_f = 1'h0;
  end
  if (reset) begin
    pmu_fw_halt_req_f = 1'h0;
  end
  if (reset) begin
    internal_pmu_fw_halt_mode_f = 1'h0;
  end
  if (reset) begin
    tlu_flush_lower_r_d1 = 1'h0;
  end
  if (reset) begin
    ic_perr_r_d1 = 1'h0;
  end
  if (reset) begin
    iccm_sbecc_r_d1 = 1'h0;
  end
  if (reset) begin
    request_debug_mode_r_d1 = 1'h0;
  end
  if (reset) begin
    iccm_repair_state_d1 = 1'h0;
  end
  if (reset) begin
    dec_pause_state_f = 1'h0;
  end
  if (reset) begin
    dec_tlu_wr_pause_r_d1 = 1'h0;
  end
  if (reset) begin
    exc_or_int_valid_r_d1 = 1'h0;
  end
  if (reset) begin
    pause_expired_wb = 1'h0;
  end
  if (reset) begin
    lsu_pmu_load_external_r = 1'h0;
  end
  if (reset) begin
    lsu_pmu_store_external_r = 1'h0;
  end
  if (reset) begin
    _T_32 = 1'h0;
  end
  if (reset) begin
    internal_dbg_halt_mode_f2 = 1'h0;
  end
  if (reset) begin
    _T_33 = 1'h0;
  end
  if (reset) begin
    nmi_lsu_load_type_f = 1'h0;
  end
  if (reset) begin
    nmi_lsu_store_type_f = 1'h0;
  end
  if (reset) begin
    mpc_debug_halt_req_sync_f = 1'h0;
  end
  if (reset) begin
    mpc_debug_run_req_sync_f = 1'h0;
  end
  if (reset) begin
    mpc_run_state_f = 1'h0;
  end
  if (reset) begin
    debug_brkpt_status_f = 1'h0;
  end
  if (reset) begin
    mpc_debug_halt_ack_f = 1'h0;
  end
  if (reset) begin
    mpc_debug_run_ack_f = 1'h0;
  end
  if (reset) begin
    dbg_run_state_f = 1'h0;
  end
  if (reset) begin
    _T_65 = 1'h0;
  end
  if (reset) begin
    request_debug_mode_done_f = 1'h0;
  end
  if (reset) begin
    _T_190 = 1'h0;
  end
  if (reset) begin
    _T_353 = 1'h0;
  end
  if (reset) begin
    _T_354 = 1'h0;
  end
  if (reset) begin
    _T_355 = 1'h0;
  end
  if (reset) begin
    lsu_single_ecc_error_r_d1 = 1'h0;
  end
  if (reset) begin
    lsu_i0_exc_r_d1 = 1'h0;
  end
  if (reset) begin
    take_ext_int_start_d2 = 1'h0;
  end
  if (reset) begin
    tlu_flush_path_r_d1 = 31'h0;
  end
  if (reset) begin
    i0_exception_valid_r_d1 = 1'h0;
  end
  if (reset) begin
    exc_cause_wb = 5'h0;
  end
  if (reset) begin
    i0_valid_wb = 1'h0;
  end
  if (reset) begin
    trigger_hit_r_d1 = 1'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      dbg_halt_state_f <= 1'h0;
    end else begin
      dbg_halt_state_f <= _T_83 & _T_84;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      mpc_halt_state_f <= 1'h0;
    end else begin
      mpc_halt_state_f <= _T_71 & _T_72;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      _T_8 <= 7'h0;
    end else begin
      _T_8 <= {_T_6,_T_3};
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      syncro_ff <= 7'h0;
    end else begin
      syncro_ff <= _T_8;
    end
  end
  always @(posedge rvclkhdr_1_io_l1clk or posedge reset) begin
    if (reset) begin
      lsu_exc_valid_r_d1 <= 1'h0;
    end else begin
      lsu_exc_valid_r_d1 <= _T_405 & _T_470;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      e5_valid <= 1'h0;
    end else begin
      e5_valid <= io_dec_tlu_i0_valid_r;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      debug_mode_status <= 1'h0;
    end else begin
      debug_mode_status <= debug_halt_req_ns | _T_160;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      i_cpu_run_req_d1_raw <= 1'h0;
    end else begin
      i_cpu_run_req_d1_raw <= _T_351 & _T_107;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      nmi_int_delayed <= 1'h0;
    end else begin
      nmi_int_delayed <= syncro_ff[6];
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      mdseac_locked_f <= 1'h0;
    end else begin
      mdseac_locked_f <= csr_io_mdseac_locked_ns;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      nmi_int_detected_f <= 1'h0;
    end else begin
      nmi_int_detected_f <= _T_42 | _T_44;
    end
  end
  always @(posedge rvclkhdr_3_io_l1clk or posedge reset) begin
    if (reset) begin
      take_nmi_r_d1 <= 1'h0;
    end else begin
      take_nmi_r_d1 <= _T_756 & _T_760;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      take_ext_int_start_d3 <= 1'h0;
    end else begin
      take_ext_int_start_d3 <= take_ext_int_start_d2;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      int_timer0_int_hold_f <= 1'h0;
    end else begin
      int_timer0_int_hold_f <= _T_644 | _T_651;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      int_timer1_int_hold_f <= 1'h0;
    end else begin
      int_timer1_int_hold_f <= _T_654 | _T_661;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      i_cpu_halt_req_d1 <= 1'h0;
    end else begin
      i_cpu_halt_req_d1 <= _T_347 & _T_107;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      dbg_halt_req_held <= 1'h0;
    end else begin
      dbg_halt_req_held <= _T_106 & ext_int_freeze_d1;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      ext_int_freeze_d1 <= 1'h0;
    end else begin
      ext_int_freeze_d1 <= _T_682 | take_ext_int_start_d3;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      reset_detect <= 1'h0;
    end else begin
      reset_detect <= 1'h1;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      reset_detected <= 1'h0;
    end else begin
      reset_detected <= reset_detect;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      dcsr_single_step_done_f <= 1'h0;
    end else begin
      dcsr_single_step_done_f <= _T_174 & _T_470;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      trigger_hit_dmode_r_d1 <= 1'h0;
    end else begin
      trigger_hit_dmode_r_d1 <= i0_trigger_hit_raw_r & i0_trigger_action_r;
    end
  end
  always @(posedge rvclkhdr_2_io_l1clk or posedge reset) begin
    if (reset) begin
      ebreak_to_debug_mode_r_d1 <= 1'h0;
    end else begin
      ebreak_to_debug_mode_r_d1 <= _T_519 & _T_470;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      debug_halt_req_f <= 1'h0;
    end else begin
      debug_halt_req_f <= enter_debug_halt_req | _T_168;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      lsu_idle_any_f <= 1'h0;
    end else begin
      lsu_idle_any_f <= io_lsu_idle_any;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      ifu_miss_state_idle_f <= 1'h0;
    end else begin
      ifu_miss_state_idle_f <= io_tlu_mem_ifu_miss_state_idle;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      debug_halt_req_d1 <= 1'h0;
    end else begin
      debug_halt_req_d1 <= _T_114 & _T_107;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      dec_tlu_flush_noredir_r_d1 <= 1'h0;
    end else begin
      dec_tlu_flush_noredir_r_d1 <= io_tlu_ifc_dec_tlu_flush_noredir_wb;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      dec_tlu_flush_pause_r_d1 <= 1'h0;
    end else begin
      dec_tlu_flush_pause_r_d1 <= io_dec_tlu_flush_pause_r;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      take_ext_int_start_d1 <= 1'h0;
    end else begin
      take_ext_int_start_d1 <= ext_int_ready & _T_704;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      halt_taken_f <= 1'h0;
    end else begin
      halt_taken_f <= _T_135 | _T_141;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      dbg_tlu_halted_f <= 1'h0;
    end else begin
      dbg_tlu_halted_f <= _T_164 | _T_166;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      pmu_fw_tlu_halted_f <= 1'h0;
    end else begin
      pmu_fw_tlu_halted_f <= _T_377 & _T_378;
    end
  end
  always @(posedge rvclkhdr_3_io_l1clk or posedge reset) begin
    if (reset) begin
      interrupt_valid_r_d1 <= 1'h0;
    end else begin
      interrupt_valid_r_d1 <= _T_766 | take_int_timer1_int;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      debug_resume_req_f <= 1'h0;
    end else begin
      debug_resume_req_f <= _T_165 & _T_121;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      dcsr_single_step_running_f <= 1'h0;
    end else begin
      dcsr_single_step_running_f <= _T_177 | _T_179;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      pmu_fw_halt_req_f <= 1'h0;
    end else begin
      pmu_fw_halt_req_f <= _T_363 & _T_378;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      internal_pmu_fw_halt_mode_f <= 1'h0;
    end else begin
      internal_pmu_fw_halt_mode_f <= pmu_fw_halt_req_ns | _T_369;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      tlu_flush_lower_r_d1 <= 1'h0;
    end else begin
      tlu_flush_lower_r_d1 <= _T_801 | take_ext_int_start;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      ic_perr_r_d1 <= 1'h0;
    end else begin
      ic_perr_r_d1 <= _T_499 & _T_500;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      iccm_sbecc_r_d1 <= 1'h0;
    end else begin
      iccm_sbecc_r_d1 <= _T_506 & _T_500;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      request_debug_mode_r_d1 <= 1'h0;
    end else begin
      request_debug_mode_r_d1 <= _T_180 | _T_182;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      iccm_repair_state_d1 <= 1'h0;
    end else begin
      iccm_repair_state_d1 <= iccm_sbecc_r_d1 | _T_442;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      dec_pause_state_f <= 1'h0;
    end else begin
      dec_pause_state_f <= io_dec_pause_state;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      dec_tlu_wr_pause_r_d1 <= 1'h0;
    end else begin
      dec_tlu_wr_pause_r_d1 <= io_dec_tlu_wr_pause_r;
    end
  end
  always @(posedge rvclkhdr_3_io_l1clk or posedge reset) begin
    if (reset) begin
      exc_or_int_valid_r_d1 <= 1'h0;
    end else begin
      exc_or_int_valid_r_d1 <= _T_855 | mepc_trigger_hit_sel_pc_r;
    end
  end
  always @(posedge rvclkhdr_3_io_l1clk or posedge reset) begin
    if (reset) begin
      pause_expired_wb <= 1'h0;
    end else begin
      pause_expired_wb <= _T_227 & _T_228;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      lsu_pmu_load_external_r <= 1'h0;
    end else begin
      lsu_pmu_load_external_r <= io_lsu_tlu_lsu_pmu_load_external_m;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      lsu_pmu_store_external_r <= 1'h0;
    end else begin
      lsu_pmu_store_external_r <= io_lsu_tlu_lsu_pmu_store_external_m;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      _T_32 <= 1'h0;
    end else begin
      _T_32 <= _T_427 | i0_trigger_hit_raw_r;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      internal_dbg_halt_mode_f2 <= 1'h0;
    end else begin
      internal_dbg_halt_mode_f2 <= debug_mode_status;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      _T_33 <= 1'h0;
    end else begin
      _T_33 <= csr_io_force_halt;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      nmi_lsu_load_type_f <= 1'h0;
    end else begin
      nmi_lsu_load_type_f <= _T_50 | _T_52;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      nmi_lsu_store_type_f <= 1'h0;
    end else begin
      nmi_lsu_store_type_f <= _T_58 | _T_60;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      mpc_debug_halt_req_sync_f <= 1'h0;
    end else begin
      mpc_debug_halt_req_sync_f <= mpc_debug_halt_req_sync_raw & _T_107;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      mpc_debug_run_req_sync_f <= 1'h0;
    end else begin
      mpc_debug_run_req_sync_f <= syncro_ff[0];
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      mpc_run_state_f <= 1'h0;
    end else begin
      mpc_run_state_f <= _T_76 & _T_78;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      debug_brkpt_status_f <= 1'h0;
    end else begin
      debug_brkpt_status_f <= _T_92 & _T_94;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      mpc_debug_halt_ack_f <= 1'h0;
    end else begin
      mpc_debug_halt_ack_f <= _T_97 & core_empty;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      mpc_debug_run_ack_f <= 1'h0;
    end else begin
      mpc_debug_run_ack_f <= _T_102 | _T_103;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      dbg_run_state_f <= 1'h0;
    end else begin
      dbg_run_state_f <= _T_86 & _T_78;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      _T_65 <= 1'h0;
    end else begin
      _T_65 <= _T & mpc_halt_state_f;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      request_debug_mode_done_f <= 1'h0;
    end else begin
      request_debug_mode_done_f <= _T_183 & _T_136;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      _T_190 <= 1'h0;
    end else begin
      _T_190 <= _T_170 & dbg_run_state_ns;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      _T_353 <= 1'h0;
    end else begin
      _T_353 <= _T_376 | _T_386;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      _T_354 <= 1'h0;
    end else begin
      _T_354 <= i_cpu_halt_req_d1 & pmu_fw_tlu_halted_f;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      _T_355 <= 1'h0;
    end else begin
      _T_355 <= _T_388 | _T_389;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      lsu_single_ecc_error_r_d1 <= 1'h0;
    end else begin
      lsu_single_ecc_error_r_d1 <= io_lsu_single_ecc_error_incr;
    end
  end
  always @(posedge rvclkhdr_1_io_l1clk or posedge reset) begin
    if (reset) begin
      lsu_i0_exc_r_d1 <= 1'h0;
    end else begin
      lsu_i0_exc_r_d1 <= _T_405 & _T_470;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      take_ext_int_start_d2 <= 1'h0;
    end else begin
      take_ext_int_start_d2 <= take_ext_int_start_d1;
    end
  end
  always @(posedge rvclkhdr_3_io_l1clk or posedge reset) begin
    if (reset) begin
      tlu_flush_path_r_d1 <= 31'h0;
    end else if (take_reset) begin
      tlu_flush_path_r_d1 <= io_rst_vec;
    end else begin
      tlu_flush_path_r_d1 <= _T_852;
    end
  end
  always @(posedge rvclkhdr_3_io_l1clk or posedge reset) begin
    if (reset) begin
      i0_exception_valid_r_d1 <= 1'h0;
    end else begin
      i0_exception_valid_r_d1 <= _T_527 & _T_528;
    end
  end
  always @(posedge rvclkhdr_3_io_l1clk or posedge reset) begin
    if (reset) begin
      exc_cause_wb <= 5'h0;
    end else begin
      exc_cause_wb <= _T_603 | _T_591;
    end
  end
  always @(posedge rvclkhdr_3_io_l1clk or posedge reset) begin
    if (reset) begin
      i0_valid_wb <= 1'h0;
    end else begin
      i0_valid_wb <= tlu_i0_commit_cmt & _T_860;
    end
  end
  always @(posedge rvclkhdr_3_io_l1clk or posedge reset) begin
    if (reset) begin
      trigger_hit_r_d1 <= 1'h0;
    end else begin
      trigger_hit_r_d1 <= |i0_trigger_chain_masked_r;
    end
  end
endmodule
module dec_trigger(
  input         io_trigger_pkt_any_0_select,
  input         io_trigger_pkt_any_0_match_pkt,
  input         io_trigger_pkt_any_0_execute,
  input         io_trigger_pkt_any_0_m,
  input  [31:0] io_trigger_pkt_any_0_tdata2,
  input         io_trigger_pkt_any_1_select,
  input         io_trigger_pkt_any_1_match_pkt,
  input         io_trigger_pkt_any_1_execute,
  input         io_trigger_pkt_any_1_m,
  input  [31:0] io_trigger_pkt_any_1_tdata2,
  input         io_trigger_pkt_any_2_select,
  input         io_trigger_pkt_any_2_match_pkt,
  input         io_trigger_pkt_any_2_execute,
  input         io_trigger_pkt_any_2_m,
  input  [31:0] io_trigger_pkt_any_2_tdata2,
  input         io_trigger_pkt_any_3_select,
  input         io_trigger_pkt_any_3_match_pkt,
  input         io_trigger_pkt_any_3_execute,
  input         io_trigger_pkt_any_3_m,
  input  [31:0] io_trigger_pkt_any_3_tdata2,
  input  [30:0] io_dec_i0_pc_d,
  output [3:0]  io_dec_i0_trigger_match_d
);
  wire  _T = ~io_trigger_pkt_any_0_select; // @[dec_trigger.scala 14:63]
  wire  _T_1 = _T & io_trigger_pkt_any_0_execute; // @[dec_trigger.scala 14:93]
  wire [9:0] _T_11 = {_T_1,_T_1,_T_1,_T_1,_T_1,_T_1,_T_1,_T_1,_T_1,_T_1}; // @[Cat.scala 29:58]
  wire [18:0] _T_20 = {_T_11,_T_1,_T_1,_T_1,_T_1,_T_1,_T_1,_T_1,_T_1,_T_1}; // @[Cat.scala 29:58]
  wire [27:0] _T_29 = {_T_20,_T_1,_T_1,_T_1,_T_1,_T_1,_T_1,_T_1,_T_1,_T_1}; // @[Cat.scala 29:58]
  wire [31:0] _T_33 = {_T_29,_T_1,_T_1,_T_1,_T_1}; // @[Cat.scala 29:58]
  wire [31:0] _T_35 = {io_dec_i0_pc_d,io_trigger_pkt_any_0_tdata2[0]}; // @[Cat.scala 29:58]
  wire [31:0] dec_i0_match_data_0 = _T_33 & _T_35; // @[dec_trigger.scala 14:127]
  wire  _T_37 = ~io_trigger_pkt_any_1_select; // @[dec_trigger.scala 14:63]
  wire  _T_38 = _T_37 & io_trigger_pkt_any_1_execute; // @[dec_trigger.scala 14:93]
  wire [9:0] _T_48 = {_T_38,_T_38,_T_38,_T_38,_T_38,_T_38,_T_38,_T_38,_T_38,_T_38}; // @[Cat.scala 29:58]
  wire [18:0] _T_57 = {_T_48,_T_38,_T_38,_T_38,_T_38,_T_38,_T_38,_T_38,_T_38,_T_38}; // @[Cat.scala 29:58]
  wire [27:0] _T_66 = {_T_57,_T_38,_T_38,_T_38,_T_38,_T_38,_T_38,_T_38,_T_38,_T_38}; // @[Cat.scala 29:58]
  wire [31:0] _T_70 = {_T_66,_T_38,_T_38,_T_38,_T_38}; // @[Cat.scala 29:58]
  wire [31:0] _T_72 = {io_dec_i0_pc_d,io_trigger_pkt_any_1_tdata2[0]}; // @[Cat.scala 29:58]
  wire [31:0] dec_i0_match_data_1 = _T_70 & _T_72; // @[dec_trigger.scala 14:127]
  wire  _T_74 = ~io_trigger_pkt_any_2_select; // @[dec_trigger.scala 14:63]
  wire  _T_75 = _T_74 & io_trigger_pkt_any_2_execute; // @[dec_trigger.scala 14:93]
  wire [9:0] _T_85 = {_T_75,_T_75,_T_75,_T_75,_T_75,_T_75,_T_75,_T_75,_T_75,_T_75}; // @[Cat.scala 29:58]
  wire [18:0] _T_94 = {_T_85,_T_75,_T_75,_T_75,_T_75,_T_75,_T_75,_T_75,_T_75,_T_75}; // @[Cat.scala 29:58]
  wire [27:0] _T_103 = {_T_94,_T_75,_T_75,_T_75,_T_75,_T_75,_T_75,_T_75,_T_75,_T_75}; // @[Cat.scala 29:58]
  wire [31:0] _T_107 = {_T_103,_T_75,_T_75,_T_75,_T_75}; // @[Cat.scala 29:58]
  wire [31:0] _T_109 = {io_dec_i0_pc_d,io_trigger_pkt_any_2_tdata2[0]}; // @[Cat.scala 29:58]
  wire [31:0] dec_i0_match_data_2 = _T_107 & _T_109; // @[dec_trigger.scala 14:127]
  wire  _T_111 = ~io_trigger_pkt_any_3_select; // @[dec_trigger.scala 14:63]
  wire  _T_112 = _T_111 & io_trigger_pkt_any_3_execute; // @[dec_trigger.scala 14:93]
  wire [9:0] _T_122 = {_T_112,_T_112,_T_112,_T_112,_T_112,_T_112,_T_112,_T_112,_T_112,_T_112}; // @[Cat.scala 29:58]
  wire [18:0] _T_131 = {_T_122,_T_112,_T_112,_T_112,_T_112,_T_112,_T_112,_T_112,_T_112,_T_112}; // @[Cat.scala 29:58]
  wire [27:0] _T_140 = {_T_131,_T_112,_T_112,_T_112,_T_112,_T_112,_T_112,_T_112,_T_112,_T_112}; // @[Cat.scala 29:58]
  wire [31:0] _T_144 = {_T_140,_T_112,_T_112,_T_112,_T_112}; // @[Cat.scala 29:58]
  wire [31:0] _T_146 = {io_dec_i0_pc_d,io_trigger_pkt_any_3_tdata2[0]}; // @[Cat.scala 29:58]
  wire [31:0] dec_i0_match_data_3 = _T_144 & _T_146; // @[dec_trigger.scala 14:127]
  wire  _T_148 = io_trigger_pkt_any_0_execute & io_trigger_pkt_any_0_m; // @[dec_trigger.scala 15:83]
  wire  _T_151 = &io_trigger_pkt_any_0_tdata2; // @[lib.scala 101:45]
  wire  _T_152 = ~_T_151; // @[lib.scala 101:39]
  wire  _T_153 = io_trigger_pkt_any_0_match_pkt & _T_152; // @[lib.scala 101:37]
  wire  _T_156 = io_trigger_pkt_any_0_tdata2[0] == dec_i0_match_data_0[0]; // @[lib.scala 102:52]
  wire  _T_157 = _T_153 | _T_156; // @[lib.scala 102:41]
  wire  _T_159 = &io_trigger_pkt_any_0_tdata2[0]; // @[lib.scala 104:36]
  wire  _T_160 = _T_159 & _T_153; // @[lib.scala 104:41]
  wire  _T_163 = io_trigger_pkt_any_0_tdata2[1] == dec_i0_match_data_0[1]; // @[lib.scala 104:78]
  wire  _T_164 = _T_160 | _T_163; // @[lib.scala 104:23]
  wire  _T_166 = &io_trigger_pkt_any_0_tdata2[1:0]; // @[lib.scala 104:36]
  wire  _T_167 = _T_166 & _T_153; // @[lib.scala 104:41]
  wire  _T_170 = io_trigger_pkt_any_0_tdata2[2] == dec_i0_match_data_0[2]; // @[lib.scala 104:78]
  wire  _T_171 = _T_167 | _T_170; // @[lib.scala 104:23]
  wire  _T_173 = &io_trigger_pkt_any_0_tdata2[2:0]; // @[lib.scala 104:36]
  wire  _T_174 = _T_173 & _T_153; // @[lib.scala 104:41]
  wire  _T_177 = io_trigger_pkt_any_0_tdata2[3] == dec_i0_match_data_0[3]; // @[lib.scala 104:78]
  wire  _T_178 = _T_174 | _T_177; // @[lib.scala 104:23]
  wire  _T_180 = &io_trigger_pkt_any_0_tdata2[3:0]; // @[lib.scala 104:36]
  wire  _T_181 = _T_180 & _T_153; // @[lib.scala 104:41]
  wire  _T_184 = io_trigger_pkt_any_0_tdata2[4] == dec_i0_match_data_0[4]; // @[lib.scala 104:78]
  wire  _T_185 = _T_181 | _T_184; // @[lib.scala 104:23]
  wire  _T_187 = &io_trigger_pkt_any_0_tdata2[4:0]; // @[lib.scala 104:36]
  wire  _T_188 = _T_187 & _T_153; // @[lib.scala 104:41]
  wire  _T_191 = io_trigger_pkt_any_0_tdata2[5] == dec_i0_match_data_0[5]; // @[lib.scala 104:78]
  wire  _T_192 = _T_188 | _T_191; // @[lib.scala 104:23]
  wire  _T_194 = &io_trigger_pkt_any_0_tdata2[5:0]; // @[lib.scala 104:36]
  wire  _T_195 = _T_194 & _T_153; // @[lib.scala 104:41]
  wire  _T_198 = io_trigger_pkt_any_0_tdata2[6] == dec_i0_match_data_0[6]; // @[lib.scala 104:78]
  wire  _T_199 = _T_195 | _T_198; // @[lib.scala 104:23]
  wire  _T_201 = &io_trigger_pkt_any_0_tdata2[6:0]; // @[lib.scala 104:36]
  wire  _T_202 = _T_201 & _T_153; // @[lib.scala 104:41]
  wire  _T_205 = io_trigger_pkt_any_0_tdata2[7] == dec_i0_match_data_0[7]; // @[lib.scala 104:78]
  wire  _T_206 = _T_202 | _T_205; // @[lib.scala 104:23]
  wire  _T_208 = &io_trigger_pkt_any_0_tdata2[7:0]; // @[lib.scala 104:36]
  wire  _T_209 = _T_208 & _T_153; // @[lib.scala 104:41]
  wire  _T_212 = io_trigger_pkt_any_0_tdata2[8] == dec_i0_match_data_0[8]; // @[lib.scala 104:78]
  wire  _T_213 = _T_209 | _T_212; // @[lib.scala 104:23]
  wire  _T_215 = &io_trigger_pkt_any_0_tdata2[8:0]; // @[lib.scala 104:36]
  wire  _T_216 = _T_215 & _T_153; // @[lib.scala 104:41]
  wire  _T_219 = io_trigger_pkt_any_0_tdata2[9] == dec_i0_match_data_0[9]; // @[lib.scala 104:78]
  wire  _T_220 = _T_216 | _T_219; // @[lib.scala 104:23]
  wire  _T_222 = &io_trigger_pkt_any_0_tdata2[9:0]; // @[lib.scala 104:36]
  wire  _T_223 = _T_222 & _T_153; // @[lib.scala 104:41]
  wire  _T_226 = io_trigger_pkt_any_0_tdata2[10] == dec_i0_match_data_0[10]; // @[lib.scala 104:78]
  wire  _T_227 = _T_223 | _T_226; // @[lib.scala 104:23]
  wire  _T_229 = &io_trigger_pkt_any_0_tdata2[10:0]; // @[lib.scala 104:36]
  wire  _T_230 = _T_229 & _T_153; // @[lib.scala 104:41]
  wire  _T_233 = io_trigger_pkt_any_0_tdata2[11] == dec_i0_match_data_0[11]; // @[lib.scala 104:78]
  wire  _T_234 = _T_230 | _T_233; // @[lib.scala 104:23]
  wire  _T_236 = &io_trigger_pkt_any_0_tdata2[11:0]; // @[lib.scala 104:36]
  wire  _T_237 = _T_236 & _T_153; // @[lib.scala 104:41]
  wire  _T_240 = io_trigger_pkt_any_0_tdata2[12] == dec_i0_match_data_0[12]; // @[lib.scala 104:78]
  wire  _T_241 = _T_237 | _T_240; // @[lib.scala 104:23]
  wire  _T_243 = &io_trigger_pkt_any_0_tdata2[12:0]; // @[lib.scala 104:36]
  wire  _T_244 = _T_243 & _T_153; // @[lib.scala 104:41]
  wire  _T_247 = io_trigger_pkt_any_0_tdata2[13] == dec_i0_match_data_0[13]; // @[lib.scala 104:78]
  wire  _T_248 = _T_244 | _T_247; // @[lib.scala 104:23]
  wire  _T_250 = &io_trigger_pkt_any_0_tdata2[13:0]; // @[lib.scala 104:36]
  wire  _T_251 = _T_250 & _T_153; // @[lib.scala 104:41]
  wire  _T_254 = io_trigger_pkt_any_0_tdata2[14] == dec_i0_match_data_0[14]; // @[lib.scala 104:78]
  wire  _T_255 = _T_251 | _T_254; // @[lib.scala 104:23]
  wire  _T_257 = &io_trigger_pkt_any_0_tdata2[14:0]; // @[lib.scala 104:36]
  wire  _T_258 = _T_257 & _T_153; // @[lib.scala 104:41]
  wire  _T_261 = io_trigger_pkt_any_0_tdata2[15] == dec_i0_match_data_0[15]; // @[lib.scala 104:78]
  wire  _T_262 = _T_258 | _T_261; // @[lib.scala 104:23]
  wire  _T_264 = &io_trigger_pkt_any_0_tdata2[15:0]; // @[lib.scala 104:36]
  wire  _T_265 = _T_264 & _T_153; // @[lib.scala 104:41]
  wire  _T_268 = io_trigger_pkt_any_0_tdata2[16] == dec_i0_match_data_0[16]; // @[lib.scala 104:78]
  wire  _T_269 = _T_265 | _T_268; // @[lib.scala 104:23]
  wire  _T_271 = &io_trigger_pkt_any_0_tdata2[16:0]; // @[lib.scala 104:36]
  wire  _T_272 = _T_271 & _T_153; // @[lib.scala 104:41]
  wire  _T_275 = io_trigger_pkt_any_0_tdata2[17] == dec_i0_match_data_0[17]; // @[lib.scala 104:78]
  wire  _T_276 = _T_272 | _T_275; // @[lib.scala 104:23]
  wire  _T_278 = &io_trigger_pkt_any_0_tdata2[17:0]; // @[lib.scala 104:36]
  wire  _T_279 = _T_278 & _T_153; // @[lib.scala 104:41]
  wire  _T_282 = io_trigger_pkt_any_0_tdata2[18] == dec_i0_match_data_0[18]; // @[lib.scala 104:78]
  wire  _T_283 = _T_279 | _T_282; // @[lib.scala 104:23]
  wire  _T_285 = &io_trigger_pkt_any_0_tdata2[18:0]; // @[lib.scala 104:36]
  wire  _T_286 = _T_285 & _T_153; // @[lib.scala 104:41]
  wire  _T_289 = io_trigger_pkt_any_0_tdata2[19] == dec_i0_match_data_0[19]; // @[lib.scala 104:78]
  wire  _T_290 = _T_286 | _T_289; // @[lib.scala 104:23]
  wire  _T_292 = &io_trigger_pkt_any_0_tdata2[19:0]; // @[lib.scala 104:36]
  wire  _T_293 = _T_292 & _T_153; // @[lib.scala 104:41]
  wire  _T_296 = io_trigger_pkt_any_0_tdata2[20] == dec_i0_match_data_0[20]; // @[lib.scala 104:78]
  wire  _T_297 = _T_293 | _T_296; // @[lib.scala 104:23]
  wire  _T_299 = &io_trigger_pkt_any_0_tdata2[20:0]; // @[lib.scala 104:36]
  wire  _T_300 = _T_299 & _T_153; // @[lib.scala 104:41]
  wire  _T_303 = io_trigger_pkt_any_0_tdata2[21] == dec_i0_match_data_0[21]; // @[lib.scala 104:78]
  wire  _T_304 = _T_300 | _T_303; // @[lib.scala 104:23]
  wire  _T_306 = &io_trigger_pkt_any_0_tdata2[21:0]; // @[lib.scala 104:36]
  wire  _T_307 = _T_306 & _T_153; // @[lib.scala 104:41]
  wire  _T_310 = io_trigger_pkt_any_0_tdata2[22] == dec_i0_match_data_0[22]; // @[lib.scala 104:78]
  wire  _T_311 = _T_307 | _T_310; // @[lib.scala 104:23]
  wire  _T_313 = &io_trigger_pkt_any_0_tdata2[22:0]; // @[lib.scala 104:36]
  wire  _T_314 = _T_313 & _T_153; // @[lib.scala 104:41]
  wire  _T_317 = io_trigger_pkt_any_0_tdata2[23] == dec_i0_match_data_0[23]; // @[lib.scala 104:78]
  wire  _T_318 = _T_314 | _T_317; // @[lib.scala 104:23]
  wire  _T_320 = &io_trigger_pkt_any_0_tdata2[23:0]; // @[lib.scala 104:36]
  wire  _T_321 = _T_320 & _T_153; // @[lib.scala 104:41]
  wire  _T_324 = io_trigger_pkt_any_0_tdata2[24] == dec_i0_match_data_0[24]; // @[lib.scala 104:78]
  wire  _T_325 = _T_321 | _T_324; // @[lib.scala 104:23]
  wire  _T_327 = &io_trigger_pkt_any_0_tdata2[24:0]; // @[lib.scala 104:36]
  wire  _T_328 = _T_327 & _T_153; // @[lib.scala 104:41]
  wire  _T_331 = io_trigger_pkt_any_0_tdata2[25] == dec_i0_match_data_0[25]; // @[lib.scala 104:78]
  wire  _T_332 = _T_328 | _T_331; // @[lib.scala 104:23]
  wire  _T_334 = &io_trigger_pkt_any_0_tdata2[25:0]; // @[lib.scala 104:36]
  wire  _T_335 = _T_334 & _T_153; // @[lib.scala 104:41]
  wire  _T_338 = io_trigger_pkt_any_0_tdata2[26] == dec_i0_match_data_0[26]; // @[lib.scala 104:78]
  wire  _T_339 = _T_335 | _T_338; // @[lib.scala 104:23]
  wire  _T_341 = &io_trigger_pkt_any_0_tdata2[26:0]; // @[lib.scala 104:36]
  wire  _T_342 = _T_341 & _T_153; // @[lib.scala 104:41]
  wire  _T_345 = io_trigger_pkt_any_0_tdata2[27] == dec_i0_match_data_0[27]; // @[lib.scala 104:78]
  wire  _T_346 = _T_342 | _T_345; // @[lib.scala 104:23]
  wire  _T_348 = &io_trigger_pkt_any_0_tdata2[27:0]; // @[lib.scala 104:36]
  wire  _T_349 = _T_348 & _T_153; // @[lib.scala 104:41]
  wire  _T_352 = io_trigger_pkt_any_0_tdata2[28] == dec_i0_match_data_0[28]; // @[lib.scala 104:78]
  wire  _T_353 = _T_349 | _T_352; // @[lib.scala 104:23]
  wire  _T_355 = &io_trigger_pkt_any_0_tdata2[28:0]; // @[lib.scala 104:36]
  wire  _T_356 = _T_355 & _T_153; // @[lib.scala 104:41]
  wire  _T_359 = io_trigger_pkt_any_0_tdata2[29] == dec_i0_match_data_0[29]; // @[lib.scala 104:78]
  wire  _T_360 = _T_356 | _T_359; // @[lib.scala 104:23]
  wire  _T_362 = &io_trigger_pkt_any_0_tdata2[29:0]; // @[lib.scala 104:36]
  wire  _T_363 = _T_362 & _T_153; // @[lib.scala 104:41]
  wire  _T_366 = io_trigger_pkt_any_0_tdata2[30] == dec_i0_match_data_0[30]; // @[lib.scala 104:78]
  wire  _T_367 = _T_363 | _T_366; // @[lib.scala 104:23]
  wire  _T_369 = &io_trigger_pkt_any_0_tdata2[30:0]; // @[lib.scala 104:36]
  wire  _T_370 = _T_369 & _T_153; // @[lib.scala 104:41]
  wire  _T_373 = io_trigger_pkt_any_0_tdata2[31] == dec_i0_match_data_0[31]; // @[lib.scala 104:78]
  wire  _T_374 = _T_370 | _T_373; // @[lib.scala 104:23]
  wire [7:0] _T_381 = {_T_206,_T_199,_T_192,_T_185,_T_178,_T_171,_T_164,_T_157}; // @[lib.scala 105:14]
  wire [15:0] _T_389 = {_T_262,_T_255,_T_248,_T_241,_T_234,_T_227,_T_220,_T_213,_T_381}; // @[lib.scala 105:14]
  wire [7:0] _T_396 = {_T_318,_T_311,_T_304,_T_297,_T_290,_T_283,_T_276,_T_269}; // @[lib.scala 105:14]
  wire [31:0] _T_405 = {_T_374,_T_367,_T_360,_T_353,_T_346,_T_339,_T_332,_T_325,_T_396,_T_389}; // @[lib.scala 105:14]
  wire  _T_406 = &_T_405; // @[lib.scala 105:25]
  wire  _T_407 = _T_148 & _T_406; // @[dec_trigger.scala 15:109]
  wire  _T_408 = io_trigger_pkt_any_1_execute & io_trigger_pkt_any_1_m; // @[dec_trigger.scala 15:83]
  wire  _T_411 = &io_trigger_pkt_any_1_tdata2; // @[lib.scala 101:45]
  wire  _T_412 = ~_T_411; // @[lib.scala 101:39]
  wire  _T_413 = io_trigger_pkt_any_1_match_pkt & _T_412; // @[lib.scala 101:37]
  wire  _T_416 = io_trigger_pkt_any_1_tdata2[0] == dec_i0_match_data_1[0]; // @[lib.scala 102:52]
  wire  _T_417 = _T_413 | _T_416; // @[lib.scala 102:41]
  wire  _T_419 = &io_trigger_pkt_any_1_tdata2[0]; // @[lib.scala 104:36]
  wire  _T_420 = _T_419 & _T_413; // @[lib.scala 104:41]
  wire  _T_423 = io_trigger_pkt_any_1_tdata2[1] == dec_i0_match_data_1[1]; // @[lib.scala 104:78]
  wire  _T_424 = _T_420 | _T_423; // @[lib.scala 104:23]
  wire  _T_426 = &io_trigger_pkt_any_1_tdata2[1:0]; // @[lib.scala 104:36]
  wire  _T_427 = _T_426 & _T_413; // @[lib.scala 104:41]
  wire  _T_430 = io_trigger_pkt_any_1_tdata2[2] == dec_i0_match_data_1[2]; // @[lib.scala 104:78]
  wire  _T_431 = _T_427 | _T_430; // @[lib.scala 104:23]
  wire  _T_433 = &io_trigger_pkt_any_1_tdata2[2:0]; // @[lib.scala 104:36]
  wire  _T_434 = _T_433 & _T_413; // @[lib.scala 104:41]
  wire  _T_437 = io_trigger_pkt_any_1_tdata2[3] == dec_i0_match_data_1[3]; // @[lib.scala 104:78]
  wire  _T_438 = _T_434 | _T_437; // @[lib.scala 104:23]
  wire  _T_440 = &io_trigger_pkt_any_1_tdata2[3:0]; // @[lib.scala 104:36]
  wire  _T_441 = _T_440 & _T_413; // @[lib.scala 104:41]
  wire  _T_444 = io_trigger_pkt_any_1_tdata2[4] == dec_i0_match_data_1[4]; // @[lib.scala 104:78]
  wire  _T_445 = _T_441 | _T_444; // @[lib.scala 104:23]
  wire  _T_447 = &io_trigger_pkt_any_1_tdata2[4:0]; // @[lib.scala 104:36]
  wire  _T_448 = _T_447 & _T_413; // @[lib.scala 104:41]
  wire  _T_451 = io_trigger_pkt_any_1_tdata2[5] == dec_i0_match_data_1[5]; // @[lib.scala 104:78]
  wire  _T_452 = _T_448 | _T_451; // @[lib.scala 104:23]
  wire  _T_454 = &io_trigger_pkt_any_1_tdata2[5:0]; // @[lib.scala 104:36]
  wire  _T_455 = _T_454 & _T_413; // @[lib.scala 104:41]
  wire  _T_458 = io_trigger_pkt_any_1_tdata2[6] == dec_i0_match_data_1[6]; // @[lib.scala 104:78]
  wire  _T_459 = _T_455 | _T_458; // @[lib.scala 104:23]
  wire  _T_461 = &io_trigger_pkt_any_1_tdata2[6:0]; // @[lib.scala 104:36]
  wire  _T_462 = _T_461 & _T_413; // @[lib.scala 104:41]
  wire  _T_465 = io_trigger_pkt_any_1_tdata2[7] == dec_i0_match_data_1[7]; // @[lib.scala 104:78]
  wire  _T_466 = _T_462 | _T_465; // @[lib.scala 104:23]
  wire  _T_468 = &io_trigger_pkt_any_1_tdata2[7:0]; // @[lib.scala 104:36]
  wire  _T_469 = _T_468 & _T_413; // @[lib.scala 104:41]
  wire  _T_472 = io_trigger_pkt_any_1_tdata2[8] == dec_i0_match_data_1[8]; // @[lib.scala 104:78]
  wire  _T_473 = _T_469 | _T_472; // @[lib.scala 104:23]
  wire  _T_475 = &io_trigger_pkt_any_1_tdata2[8:0]; // @[lib.scala 104:36]
  wire  _T_476 = _T_475 & _T_413; // @[lib.scala 104:41]
  wire  _T_479 = io_trigger_pkt_any_1_tdata2[9] == dec_i0_match_data_1[9]; // @[lib.scala 104:78]
  wire  _T_480 = _T_476 | _T_479; // @[lib.scala 104:23]
  wire  _T_482 = &io_trigger_pkt_any_1_tdata2[9:0]; // @[lib.scala 104:36]
  wire  _T_483 = _T_482 & _T_413; // @[lib.scala 104:41]
  wire  _T_486 = io_trigger_pkt_any_1_tdata2[10] == dec_i0_match_data_1[10]; // @[lib.scala 104:78]
  wire  _T_487 = _T_483 | _T_486; // @[lib.scala 104:23]
  wire  _T_489 = &io_trigger_pkt_any_1_tdata2[10:0]; // @[lib.scala 104:36]
  wire  _T_490 = _T_489 & _T_413; // @[lib.scala 104:41]
  wire  _T_493 = io_trigger_pkt_any_1_tdata2[11] == dec_i0_match_data_1[11]; // @[lib.scala 104:78]
  wire  _T_494 = _T_490 | _T_493; // @[lib.scala 104:23]
  wire  _T_496 = &io_trigger_pkt_any_1_tdata2[11:0]; // @[lib.scala 104:36]
  wire  _T_497 = _T_496 & _T_413; // @[lib.scala 104:41]
  wire  _T_500 = io_trigger_pkt_any_1_tdata2[12] == dec_i0_match_data_1[12]; // @[lib.scala 104:78]
  wire  _T_501 = _T_497 | _T_500; // @[lib.scala 104:23]
  wire  _T_503 = &io_trigger_pkt_any_1_tdata2[12:0]; // @[lib.scala 104:36]
  wire  _T_504 = _T_503 & _T_413; // @[lib.scala 104:41]
  wire  _T_507 = io_trigger_pkt_any_1_tdata2[13] == dec_i0_match_data_1[13]; // @[lib.scala 104:78]
  wire  _T_508 = _T_504 | _T_507; // @[lib.scala 104:23]
  wire  _T_510 = &io_trigger_pkt_any_1_tdata2[13:0]; // @[lib.scala 104:36]
  wire  _T_511 = _T_510 & _T_413; // @[lib.scala 104:41]
  wire  _T_514 = io_trigger_pkt_any_1_tdata2[14] == dec_i0_match_data_1[14]; // @[lib.scala 104:78]
  wire  _T_515 = _T_511 | _T_514; // @[lib.scala 104:23]
  wire  _T_517 = &io_trigger_pkt_any_1_tdata2[14:0]; // @[lib.scala 104:36]
  wire  _T_518 = _T_517 & _T_413; // @[lib.scala 104:41]
  wire  _T_521 = io_trigger_pkt_any_1_tdata2[15] == dec_i0_match_data_1[15]; // @[lib.scala 104:78]
  wire  _T_522 = _T_518 | _T_521; // @[lib.scala 104:23]
  wire  _T_524 = &io_trigger_pkt_any_1_tdata2[15:0]; // @[lib.scala 104:36]
  wire  _T_525 = _T_524 & _T_413; // @[lib.scala 104:41]
  wire  _T_528 = io_trigger_pkt_any_1_tdata2[16] == dec_i0_match_data_1[16]; // @[lib.scala 104:78]
  wire  _T_529 = _T_525 | _T_528; // @[lib.scala 104:23]
  wire  _T_531 = &io_trigger_pkt_any_1_tdata2[16:0]; // @[lib.scala 104:36]
  wire  _T_532 = _T_531 & _T_413; // @[lib.scala 104:41]
  wire  _T_535 = io_trigger_pkt_any_1_tdata2[17] == dec_i0_match_data_1[17]; // @[lib.scala 104:78]
  wire  _T_536 = _T_532 | _T_535; // @[lib.scala 104:23]
  wire  _T_538 = &io_trigger_pkt_any_1_tdata2[17:0]; // @[lib.scala 104:36]
  wire  _T_539 = _T_538 & _T_413; // @[lib.scala 104:41]
  wire  _T_542 = io_trigger_pkt_any_1_tdata2[18] == dec_i0_match_data_1[18]; // @[lib.scala 104:78]
  wire  _T_543 = _T_539 | _T_542; // @[lib.scala 104:23]
  wire  _T_545 = &io_trigger_pkt_any_1_tdata2[18:0]; // @[lib.scala 104:36]
  wire  _T_546 = _T_545 & _T_413; // @[lib.scala 104:41]
  wire  _T_549 = io_trigger_pkt_any_1_tdata2[19] == dec_i0_match_data_1[19]; // @[lib.scala 104:78]
  wire  _T_550 = _T_546 | _T_549; // @[lib.scala 104:23]
  wire  _T_552 = &io_trigger_pkt_any_1_tdata2[19:0]; // @[lib.scala 104:36]
  wire  _T_553 = _T_552 & _T_413; // @[lib.scala 104:41]
  wire  _T_556 = io_trigger_pkt_any_1_tdata2[20] == dec_i0_match_data_1[20]; // @[lib.scala 104:78]
  wire  _T_557 = _T_553 | _T_556; // @[lib.scala 104:23]
  wire  _T_559 = &io_trigger_pkt_any_1_tdata2[20:0]; // @[lib.scala 104:36]
  wire  _T_560 = _T_559 & _T_413; // @[lib.scala 104:41]
  wire  _T_563 = io_trigger_pkt_any_1_tdata2[21] == dec_i0_match_data_1[21]; // @[lib.scala 104:78]
  wire  _T_564 = _T_560 | _T_563; // @[lib.scala 104:23]
  wire  _T_566 = &io_trigger_pkt_any_1_tdata2[21:0]; // @[lib.scala 104:36]
  wire  _T_567 = _T_566 & _T_413; // @[lib.scala 104:41]
  wire  _T_570 = io_trigger_pkt_any_1_tdata2[22] == dec_i0_match_data_1[22]; // @[lib.scala 104:78]
  wire  _T_571 = _T_567 | _T_570; // @[lib.scala 104:23]
  wire  _T_573 = &io_trigger_pkt_any_1_tdata2[22:0]; // @[lib.scala 104:36]
  wire  _T_574 = _T_573 & _T_413; // @[lib.scala 104:41]
  wire  _T_577 = io_trigger_pkt_any_1_tdata2[23] == dec_i0_match_data_1[23]; // @[lib.scala 104:78]
  wire  _T_578 = _T_574 | _T_577; // @[lib.scala 104:23]
  wire  _T_580 = &io_trigger_pkt_any_1_tdata2[23:0]; // @[lib.scala 104:36]
  wire  _T_581 = _T_580 & _T_413; // @[lib.scala 104:41]
  wire  _T_584 = io_trigger_pkt_any_1_tdata2[24] == dec_i0_match_data_1[24]; // @[lib.scala 104:78]
  wire  _T_585 = _T_581 | _T_584; // @[lib.scala 104:23]
  wire  _T_587 = &io_trigger_pkt_any_1_tdata2[24:0]; // @[lib.scala 104:36]
  wire  _T_588 = _T_587 & _T_413; // @[lib.scala 104:41]
  wire  _T_591 = io_trigger_pkt_any_1_tdata2[25] == dec_i0_match_data_1[25]; // @[lib.scala 104:78]
  wire  _T_592 = _T_588 | _T_591; // @[lib.scala 104:23]
  wire  _T_594 = &io_trigger_pkt_any_1_tdata2[25:0]; // @[lib.scala 104:36]
  wire  _T_595 = _T_594 & _T_413; // @[lib.scala 104:41]
  wire  _T_598 = io_trigger_pkt_any_1_tdata2[26] == dec_i0_match_data_1[26]; // @[lib.scala 104:78]
  wire  _T_599 = _T_595 | _T_598; // @[lib.scala 104:23]
  wire  _T_601 = &io_trigger_pkt_any_1_tdata2[26:0]; // @[lib.scala 104:36]
  wire  _T_602 = _T_601 & _T_413; // @[lib.scala 104:41]
  wire  _T_605 = io_trigger_pkt_any_1_tdata2[27] == dec_i0_match_data_1[27]; // @[lib.scala 104:78]
  wire  _T_606 = _T_602 | _T_605; // @[lib.scala 104:23]
  wire  _T_608 = &io_trigger_pkt_any_1_tdata2[27:0]; // @[lib.scala 104:36]
  wire  _T_609 = _T_608 & _T_413; // @[lib.scala 104:41]
  wire  _T_612 = io_trigger_pkt_any_1_tdata2[28] == dec_i0_match_data_1[28]; // @[lib.scala 104:78]
  wire  _T_613 = _T_609 | _T_612; // @[lib.scala 104:23]
  wire  _T_615 = &io_trigger_pkt_any_1_tdata2[28:0]; // @[lib.scala 104:36]
  wire  _T_616 = _T_615 & _T_413; // @[lib.scala 104:41]
  wire  _T_619 = io_trigger_pkt_any_1_tdata2[29] == dec_i0_match_data_1[29]; // @[lib.scala 104:78]
  wire  _T_620 = _T_616 | _T_619; // @[lib.scala 104:23]
  wire  _T_622 = &io_trigger_pkt_any_1_tdata2[29:0]; // @[lib.scala 104:36]
  wire  _T_623 = _T_622 & _T_413; // @[lib.scala 104:41]
  wire  _T_626 = io_trigger_pkt_any_1_tdata2[30] == dec_i0_match_data_1[30]; // @[lib.scala 104:78]
  wire  _T_627 = _T_623 | _T_626; // @[lib.scala 104:23]
  wire  _T_629 = &io_trigger_pkt_any_1_tdata2[30:0]; // @[lib.scala 104:36]
  wire  _T_630 = _T_629 & _T_413; // @[lib.scala 104:41]
  wire  _T_633 = io_trigger_pkt_any_1_tdata2[31] == dec_i0_match_data_1[31]; // @[lib.scala 104:78]
  wire  _T_634 = _T_630 | _T_633; // @[lib.scala 104:23]
  wire [7:0] _T_641 = {_T_466,_T_459,_T_452,_T_445,_T_438,_T_431,_T_424,_T_417}; // @[lib.scala 105:14]
  wire [15:0] _T_649 = {_T_522,_T_515,_T_508,_T_501,_T_494,_T_487,_T_480,_T_473,_T_641}; // @[lib.scala 105:14]
  wire [7:0] _T_656 = {_T_578,_T_571,_T_564,_T_557,_T_550,_T_543,_T_536,_T_529}; // @[lib.scala 105:14]
  wire [31:0] _T_665 = {_T_634,_T_627,_T_620,_T_613,_T_606,_T_599,_T_592,_T_585,_T_656,_T_649}; // @[lib.scala 105:14]
  wire  _T_666 = &_T_665; // @[lib.scala 105:25]
  wire  _T_667 = _T_408 & _T_666; // @[dec_trigger.scala 15:109]
  wire  _T_668 = io_trigger_pkt_any_2_execute & io_trigger_pkt_any_2_m; // @[dec_trigger.scala 15:83]
  wire  _T_671 = &io_trigger_pkt_any_2_tdata2; // @[lib.scala 101:45]
  wire  _T_672 = ~_T_671; // @[lib.scala 101:39]
  wire  _T_673 = io_trigger_pkt_any_2_match_pkt & _T_672; // @[lib.scala 101:37]
  wire  _T_676 = io_trigger_pkt_any_2_tdata2[0] == dec_i0_match_data_2[0]; // @[lib.scala 102:52]
  wire  _T_677 = _T_673 | _T_676; // @[lib.scala 102:41]
  wire  _T_679 = &io_trigger_pkt_any_2_tdata2[0]; // @[lib.scala 104:36]
  wire  _T_680 = _T_679 & _T_673; // @[lib.scala 104:41]
  wire  _T_683 = io_trigger_pkt_any_2_tdata2[1] == dec_i0_match_data_2[1]; // @[lib.scala 104:78]
  wire  _T_684 = _T_680 | _T_683; // @[lib.scala 104:23]
  wire  _T_686 = &io_trigger_pkt_any_2_tdata2[1:0]; // @[lib.scala 104:36]
  wire  _T_687 = _T_686 & _T_673; // @[lib.scala 104:41]
  wire  _T_690 = io_trigger_pkt_any_2_tdata2[2] == dec_i0_match_data_2[2]; // @[lib.scala 104:78]
  wire  _T_691 = _T_687 | _T_690; // @[lib.scala 104:23]
  wire  _T_693 = &io_trigger_pkt_any_2_tdata2[2:0]; // @[lib.scala 104:36]
  wire  _T_694 = _T_693 & _T_673; // @[lib.scala 104:41]
  wire  _T_697 = io_trigger_pkt_any_2_tdata2[3] == dec_i0_match_data_2[3]; // @[lib.scala 104:78]
  wire  _T_698 = _T_694 | _T_697; // @[lib.scala 104:23]
  wire  _T_700 = &io_trigger_pkt_any_2_tdata2[3:0]; // @[lib.scala 104:36]
  wire  _T_701 = _T_700 & _T_673; // @[lib.scala 104:41]
  wire  _T_704 = io_trigger_pkt_any_2_tdata2[4] == dec_i0_match_data_2[4]; // @[lib.scala 104:78]
  wire  _T_705 = _T_701 | _T_704; // @[lib.scala 104:23]
  wire  _T_707 = &io_trigger_pkt_any_2_tdata2[4:0]; // @[lib.scala 104:36]
  wire  _T_708 = _T_707 & _T_673; // @[lib.scala 104:41]
  wire  _T_711 = io_trigger_pkt_any_2_tdata2[5] == dec_i0_match_data_2[5]; // @[lib.scala 104:78]
  wire  _T_712 = _T_708 | _T_711; // @[lib.scala 104:23]
  wire  _T_714 = &io_trigger_pkt_any_2_tdata2[5:0]; // @[lib.scala 104:36]
  wire  _T_715 = _T_714 & _T_673; // @[lib.scala 104:41]
  wire  _T_718 = io_trigger_pkt_any_2_tdata2[6] == dec_i0_match_data_2[6]; // @[lib.scala 104:78]
  wire  _T_719 = _T_715 | _T_718; // @[lib.scala 104:23]
  wire  _T_721 = &io_trigger_pkt_any_2_tdata2[6:0]; // @[lib.scala 104:36]
  wire  _T_722 = _T_721 & _T_673; // @[lib.scala 104:41]
  wire  _T_725 = io_trigger_pkt_any_2_tdata2[7] == dec_i0_match_data_2[7]; // @[lib.scala 104:78]
  wire  _T_726 = _T_722 | _T_725; // @[lib.scala 104:23]
  wire  _T_728 = &io_trigger_pkt_any_2_tdata2[7:0]; // @[lib.scala 104:36]
  wire  _T_729 = _T_728 & _T_673; // @[lib.scala 104:41]
  wire  _T_732 = io_trigger_pkt_any_2_tdata2[8] == dec_i0_match_data_2[8]; // @[lib.scala 104:78]
  wire  _T_733 = _T_729 | _T_732; // @[lib.scala 104:23]
  wire  _T_735 = &io_trigger_pkt_any_2_tdata2[8:0]; // @[lib.scala 104:36]
  wire  _T_736 = _T_735 & _T_673; // @[lib.scala 104:41]
  wire  _T_739 = io_trigger_pkt_any_2_tdata2[9] == dec_i0_match_data_2[9]; // @[lib.scala 104:78]
  wire  _T_740 = _T_736 | _T_739; // @[lib.scala 104:23]
  wire  _T_742 = &io_trigger_pkt_any_2_tdata2[9:0]; // @[lib.scala 104:36]
  wire  _T_743 = _T_742 & _T_673; // @[lib.scala 104:41]
  wire  _T_746 = io_trigger_pkt_any_2_tdata2[10] == dec_i0_match_data_2[10]; // @[lib.scala 104:78]
  wire  _T_747 = _T_743 | _T_746; // @[lib.scala 104:23]
  wire  _T_749 = &io_trigger_pkt_any_2_tdata2[10:0]; // @[lib.scala 104:36]
  wire  _T_750 = _T_749 & _T_673; // @[lib.scala 104:41]
  wire  _T_753 = io_trigger_pkt_any_2_tdata2[11] == dec_i0_match_data_2[11]; // @[lib.scala 104:78]
  wire  _T_754 = _T_750 | _T_753; // @[lib.scala 104:23]
  wire  _T_756 = &io_trigger_pkt_any_2_tdata2[11:0]; // @[lib.scala 104:36]
  wire  _T_757 = _T_756 & _T_673; // @[lib.scala 104:41]
  wire  _T_760 = io_trigger_pkt_any_2_tdata2[12] == dec_i0_match_data_2[12]; // @[lib.scala 104:78]
  wire  _T_761 = _T_757 | _T_760; // @[lib.scala 104:23]
  wire  _T_763 = &io_trigger_pkt_any_2_tdata2[12:0]; // @[lib.scala 104:36]
  wire  _T_764 = _T_763 & _T_673; // @[lib.scala 104:41]
  wire  _T_767 = io_trigger_pkt_any_2_tdata2[13] == dec_i0_match_data_2[13]; // @[lib.scala 104:78]
  wire  _T_768 = _T_764 | _T_767; // @[lib.scala 104:23]
  wire  _T_770 = &io_trigger_pkt_any_2_tdata2[13:0]; // @[lib.scala 104:36]
  wire  _T_771 = _T_770 & _T_673; // @[lib.scala 104:41]
  wire  _T_774 = io_trigger_pkt_any_2_tdata2[14] == dec_i0_match_data_2[14]; // @[lib.scala 104:78]
  wire  _T_775 = _T_771 | _T_774; // @[lib.scala 104:23]
  wire  _T_777 = &io_trigger_pkt_any_2_tdata2[14:0]; // @[lib.scala 104:36]
  wire  _T_778 = _T_777 & _T_673; // @[lib.scala 104:41]
  wire  _T_781 = io_trigger_pkt_any_2_tdata2[15] == dec_i0_match_data_2[15]; // @[lib.scala 104:78]
  wire  _T_782 = _T_778 | _T_781; // @[lib.scala 104:23]
  wire  _T_784 = &io_trigger_pkt_any_2_tdata2[15:0]; // @[lib.scala 104:36]
  wire  _T_785 = _T_784 & _T_673; // @[lib.scala 104:41]
  wire  _T_788 = io_trigger_pkt_any_2_tdata2[16] == dec_i0_match_data_2[16]; // @[lib.scala 104:78]
  wire  _T_789 = _T_785 | _T_788; // @[lib.scala 104:23]
  wire  _T_791 = &io_trigger_pkt_any_2_tdata2[16:0]; // @[lib.scala 104:36]
  wire  _T_792 = _T_791 & _T_673; // @[lib.scala 104:41]
  wire  _T_795 = io_trigger_pkt_any_2_tdata2[17] == dec_i0_match_data_2[17]; // @[lib.scala 104:78]
  wire  _T_796 = _T_792 | _T_795; // @[lib.scala 104:23]
  wire  _T_798 = &io_trigger_pkt_any_2_tdata2[17:0]; // @[lib.scala 104:36]
  wire  _T_799 = _T_798 & _T_673; // @[lib.scala 104:41]
  wire  _T_802 = io_trigger_pkt_any_2_tdata2[18] == dec_i0_match_data_2[18]; // @[lib.scala 104:78]
  wire  _T_803 = _T_799 | _T_802; // @[lib.scala 104:23]
  wire  _T_805 = &io_trigger_pkt_any_2_tdata2[18:0]; // @[lib.scala 104:36]
  wire  _T_806 = _T_805 & _T_673; // @[lib.scala 104:41]
  wire  _T_809 = io_trigger_pkt_any_2_tdata2[19] == dec_i0_match_data_2[19]; // @[lib.scala 104:78]
  wire  _T_810 = _T_806 | _T_809; // @[lib.scala 104:23]
  wire  _T_812 = &io_trigger_pkt_any_2_tdata2[19:0]; // @[lib.scala 104:36]
  wire  _T_813 = _T_812 & _T_673; // @[lib.scala 104:41]
  wire  _T_816 = io_trigger_pkt_any_2_tdata2[20] == dec_i0_match_data_2[20]; // @[lib.scala 104:78]
  wire  _T_817 = _T_813 | _T_816; // @[lib.scala 104:23]
  wire  _T_819 = &io_trigger_pkt_any_2_tdata2[20:0]; // @[lib.scala 104:36]
  wire  _T_820 = _T_819 & _T_673; // @[lib.scala 104:41]
  wire  _T_823 = io_trigger_pkt_any_2_tdata2[21] == dec_i0_match_data_2[21]; // @[lib.scala 104:78]
  wire  _T_824 = _T_820 | _T_823; // @[lib.scala 104:23]
  wire  _T_826 = &io_trigger_pkt_any_2_tdata2[21:0]; // @[lib.scala 104:36]
  wire  _T_827 = _T_826 & _T_673; // @[lib.scala 104:41]
  wire  _T_830 = io_trigger_pkt_any_2_tdata2[22] == dec_i0_match_data_2[22]; // @[lib.scala 104:78]
  wire  _T_831 = _T_827 | _T_830; // @[lib.scala 104:23]
  wire  _T_833 = &io_trigger_pkt_any_2_tdata2[22:0]; // @[lib.scala 104:36]
  wire  _T_834 = _T_833 & _T_673; // @[lib.scala 104:41]
  wire  _T_837 = io_trigger_pkt_any_2_tdata2[23] == dec_i0_match_data_2[23]; // @[lib.scala 104:78]
  wire  _T_838 = _T_834 | _T_837; // @[lib.scala 104:23]
  wire  _T_840 = &io_trigger_pkt_any_2_tdata2[23:0]; // @[lib.scala 104:36]
  wire  _T_841 = _T_840 & _T_673; // @[lib.scala 104:41]
  wire  _T_844 = io_trigger_pkt_any_2_tdata2[24] == dec_i0_match_data_2[24]; // @[lib.scala 104:78]
  wire  _T_845 = _T_841 | _T_844; // @[lib.scala 104:23]
  wire  _T_847 = &io_trigger_pkt_any_2_tdata2[24:0]; // @[lib.scala 104:36]
  wire  _T_848 = _T_847 & _T_673; // @[lib.scala 104:41]
  wire  _T_851 = io_trigger_pkt_any_2_tdata2[25] == dec_i0_match_data_2[25]; // @[lib.scala 104:78]
  wire  _T_852 = _T_848 | _T_851; // @[lib.scala 104:23]
  wire  _T_854 = &io_trigger_pkt_any_2_tdata2[25:0]; // @[lib.scala 104:36]
  wire  _T_855 = _T_854 & _T_673; // @[lib.scala 104:41]
  wire  _T_858 = io_trigger_pkt_any_2_tdata2[26] == dec_i0_match_data_2[26]; // @[lib.scala 104:78]
  wire  _T_859 = _T_855 | _T_858; // @[lib.scala 104:23]
  wire  _T_861 = &io_trigger_pkt_any_2_tdata2[26:0]; // @[lib.scala 104:36]
  wire  _T_862 = _T_861 & _T_673; // @[lib.scala 104:41]
  wire  _T_865 = io_trigger_pkt_any_2_tdata2[27] == dec_i0_match_data_2[27]; // @[lib.scala 104:78]
  wire  _T_866 = _T_862 | _T_865; // @[lib.scala 104:23]
  wire  _T_868 = &io_trigger_pkt_any_2_tdata2[27:0]; // @[lib.scala 104:36]
  wire  _T_869 = _T_868 & _T_673; // @[lib.scala 104:41]
  wire  _T_872 = io_trigger_pkt_any_2_tdata2[28] == dec_i0_match_data_2[28]; // @[lib.scala 104:78]
  wire  _T_873 = _T_869 | _T_872; // @[lib.scala 104:23]
  wire  _T_875 = &io_trigger_pkt_any_2_tdata2[28:0]; // @[lib.scala 104:36]
  wire  _T_876 = _T_875 & _T_673; // @[lib.scala 104:41]
  wire  _T_879 = io_trigger_pkt_any_2_tdata2[29] == dec_i0_match_data_2[29]; // @[lib.scala 104:78]
  wire  _T_880 = _T_876 | _T_879; // @[lib.scala 104:23]
  wire  _T_882 = &io_trigger_pkt_any_2_tdata2[29:0]; // @[lib.scala 104:36]
  wire  _T_883 = _T_882 & _T_673; // @[lib.scala 104:41]
  wire  _T_886 = io_trigger_pkt_any_2_tdata2[30] == dec_i0_match_data_2[30]; // @[lib.scala 104:78]
  wire  _T_887 = _T_883 | _T_886; // @[lib.scala 104:23]
  wire  _T_889 = &io_trigger_pkt_any_2_tdata2[30:0]; // @[lib.scala 104:36]
  wire  _T_890 = _T_889 & _T_673; // @[lib.scala 104:41]
  wire  _T_893 = io_trigger_pkt_any_2_tdata2[31] == dec_i0_match_data_2[31]; // @[lib.scala 104:78]
  wire  _T_894 = _T_890 | _T_893; // @[lib.scala 104:23]
  wire [7:0] _T_901 = {_T_726,_T_719,_T_712,_T_705,_T_698,_T_691,_T_684,_T_677}; // @[lib.scala 105:14]
  wire [15:0] _T_909 = {_T_782,_T_775,_T_768,_T_761,_T_754,_T_747,_T_740,_T_733,_T_901}; // @[lib.scala 105:14]
  wire [7:0] _T_916 = {_T_838,_T_831,_T_824,_T_817,_T_810,_T_803,_T_796,_T_789}; // @[lib.scala 105:14]
  wire [31:0] _T_925 = {_T_894,_T_887,_T_880,_T_873,_T_866,_T_859,_T_852,_T_845,_T_916,_T_909}; // @[lib.scala 105:14]
  wire  _T_926 = &_T_925; // @[lib.scala 105:25]
  wire  _T_927 = _T_668 & _T_926; // @[dec_trigger.scala 15:109]
  wire  _T_928 = io_trigger_pkt_any_3_execute & io_trigger_pkt_any_3_m; // @[dec_trigger.scala 15:83]
  wire  _T_931 = &io_trigger_pkt_any_3_tdata2; // @[lib.scala 101:45]
  wire  _T_932 = ~_T_931; // @[lib.scala 101:39]
  wire  _T_933 = io_trigger_pkt_any_3_match_pkt & _T_932; // @[lib.scala 101:37]
  wire  _T_936 = io_trigger_pkt_any_3_tdata2[0] == dec_i0_match_data_3[0]; // @[lib.scala 102:52]
  wire  _T_937 = _T_933 | _T_936; // @[lib.scala 102:41]
  wire  _T_939 = &io_trigger_pkt_any_3_tdata2[0]; // @[lib.scala 104:36]
  wire  _T_940 = _T_939 & _T_933; // @[lib.scala 104:41]
  wire  _T_943 = io_trigger_pkt_any_3_tdata2[1] == dec_i0_match_data_3[1]; // @[lib.scala 104:78]
  wire  _T_944 = _T_940 | _T_943; // @[lib.scala 104:23]
  wire  _T_946 = &io_trigger_pkt_any_3_tdata2[1:0]; // @[lib.scala 104:36]
  wire  _T_947 = _T_946 & _T_933; // @[lib.scala 104:41]
  wire  _T_950 = io_trigger_pkt_any_3_tdata2[2] == dec_i0_match_data_3[2]; // @[lib.scala 104:78]
  wire  _T_951 = _T_947 | _T_950; // @[lib.scala 104:23]
  wire  _T_953 = &io_trigger_pkt_any_3_tdata2[2:0]; // @[lib.scala 104:36]
  wire  _T_954 = _T_953 & _T_933; // @[lib.scala 104:41]
  wire  _T_957 = io_trigger_pkt_any_3_tdata2[3] == dec_i0_match_data_3[3]; // @[lib.scala 104:78]
  wire  _T_958 = _T_954 | _T_957; // @[lib.scala 104:23]
  wire  _T_960 = &io_trigger_pkt_any_3_tdata2[3:0]; // @[lib.scala 104:36]
  wire  _T_961 = _T_960 & _T_933; // @[lib.scala 104:41]
  wire  _T_964 = io_trigger_pkt_any_3_tdata2[4] == dec_i0_match_data_3[4]; // @[lib.scala 104:78]
  wire  _T_965 = _T_961 | _T_964; // @[lib.scala 104:23]
  wire  _T_967 = &io_trigger_pkt_any_3_tdata2[4:0]; // @[lib.scala 104:36]
  wire  _T_968 = _T_967 & _T_933; // @[lib.scala 104:41]
  wire  _T_971 = io_trigger_pkt_any_3_tdata2[5] == dec_i0_match_data_3[5]; // @[lib.scala 104:78]
  wire  _T_972 = _T_968 | _T_971; // @[lib.scala 104:23]
  wire  _T_974 = &io_trigger_pkt_any_3_tdata2[5:0]; // @[lib.scala 104:36]
  wire  _T_975 = _T_974 & _T_933; // @[lib.scala 104:41]
  wire  _T_978 = io_trigger_pkt_any_3_tdata2[6] == dec_i0_match_data_3[6]; // @[lib.scala 104:78]
  wire  _T_979 = _T_975 | _T_978; // @[lib.scala 104:23]
  wire  _T_981 = &io_trigger_pkt_any_3_tdata2[6:0]; // @[lib.scala 104:36]
  wire  _T_982 = _T_981 & _T_933; // @[lib.scala 104:41]
  wire  _T_985 = io_trigger_pkt_any_3_tdata2[7] == dec_i0_match_data_3[7]; // @[lib.scala 104:78]
  wire  _T_986 = _T_982 | _T_985; // @[lib.scala 104:23]
  wire  _T_988 = &io_trigger_pkt_any_3_tdata2[7:0]; // @[lib.scala 104:36]
  wire  _T_989 = _T_988 & _T_933; // @[lib.scala 104:41]
  wire  _T_992 = io_trigger_pkt_any_3_tdata2[8] == dec_i0_match_data_3[8]; // @[lib.scala 104:78]
  wire  _T_993 = _T_989 | _T_992; // @[lib.scala 104:23]
  wire  _T_995 = &io_trigger_pkt_any_3_tdata2[8:0]; // @[lib.scala 104:36]
  wire  _T_996 = _T_995 & _T_933; // @[lib.scala 104:41]
  wire  _T_999 = io_trigger_pkt_any_3_tdata2[9] == dec_i0_match_data_3[9]; // @[lib.scala 104:78]
  wire  _T_1000 = _T_996 | _T_999; // @[lib.scala 104:23]
  wire  _T_1002 = &io_trigger_pkt_any_3_tdata2[9:0]; // @[lib.scala 104:36]
  wire  _T_1003 = _T_1002 & _T_933; // @[lib.scala 104:41]
  wire  _T_1006 = io_trigger_pkt_any_3_tdata2[10] == dec_i0_match_data_3[10]; // @[lib.scala 104:78]
  wire  _T_1007 = _T_1003 | _T_1006; // @[lib.scala 104:23]
  wire  _T_1009 = &io_trigger_pkt_any_3_tdata2[10:0]; // @[lib.scala 104:36]
  wire  _T_1010 = _T_1009 & _T_933; // @[lib.scala 104:41]
  wire  _T_1013 = io_trigger_pkt_any_3_tdata2[11] == dec_i0_match_data_3[11]; // @[lib.scala 104:78]
  wire  _T_1014 = _T_1010 | _T_1013; // @[lib.scala 104:23]
  wire  _T_1016 = &io_trigger_pkt_any_3_tdata2[11:0]; // @[lib.scala 104:36]
  wire  _T_1017 = _T_1016 & _T_933; // @[lib.scala 104:41]
  wire  _T_1020 = io_trigger_pkt_any_3_tdata2[12] == dec_i0_match_data_3[12]; // @[lib.scala 104:78]
  wire  _T_1021 = _T_1017 | _T_1020; // @[lib.scala 104:23]
  wire  _T_1023 = &io_trigger_pkt_any_3_tdata2[12:0]; // @[lib.scala 104:36]
  wire  _T_1024 = _T_1023 & _T_933; // @[lib.scala 104:41]
  wire  _T_1027 = io_trigger_pkt_any_3_tdata2[13] == dec_i0_match_data_3[13]; // @[lib.scala 104:78]
  wire  _T_1028 = _T_1024 | _T_1027; // @[lib.scala 104:23]
  wire  _T_1030 = &io_trigger_pkt_any_3_tdata2[13:0]; // @[lib.scala 104:36]
  wire  _T_1031 = _T_1030 & _T_933; // @[lib.scala 104:41]
  wire  _T_1034 = io_trigger_pkt_any_3_tdata2[14] == dec_i0_match_data_3[14]; // @[lib.scala 104:78]
  wire  _T_1035 = _T_1031 | _T_1034; // @[lib.scala 104:23]
  wire  _T_1037 = &io_trigger_pkt_any_3_tdata2[14:0]; // @[lib.scala 104:36]
  wire  _T_1038 = _T_1037 & _T_933; // @[lib.scala 104:41]
  wire  _T_1041 = io_trigger_pkt_any_3_tdata2[15] == dec_i0_match_data_3[15]; // @[lib.scala 104:78]
  wire  _T_1042 = _T_1038 | _T_1041; // @[lib.scala 104:23]
  wire  _T_1044 = &io_trigger_pkt_any_3_tdata2[15:0]; // @[lib.scala 104:36]
  wire  _T_1045 = _T_1044 & _T_933; // @[lib.scala 104:41]
  wire  _T_1048 = io_trigger_pkt_any_3_tdata2[16] == dec_i0_match_data_3[16]; // @[lib.scala 104:78]
  wire  _T_1049 = _T_1045 | _T_1048; // @[lib.scala 104:23]
  wire  _T_1051 = &io_trigger_pkt_any_3_tdata2[16:0]; // @[lib.scala 104:36]
  wire  _T_1052 = _T_1051 & _T_933; // @[lib.scala 104:41]
  wire  _T_1055 = io_trigger_pkt_any_3_tdata2[17] == dec_i0_match_data_3[17]; // @[lib.scala 104:78]
  wire  _T_1056 = _T_1052 | _T_1055; // @[lib.scala 104:23]
  wire  _T_1058 = &io_trigger_pkt_any_3_tdata2[17:0]; // @[lib.scala 104:36]
  wire  _T_1059 = _T_1058 & _T_933; // @[lib.scala 104:41]
  wire  _T_1062 = io_trigger_pkt_any_3_tdata2[18] == dec_i0_match_data_3[18]; // @[lib.scala 104:78]
  wire  _T_1063 = _T_1059 | _T_1062; // @[lib.scala 104:23]
  wire  _T_1065 = &io_trigger_pkt_any_3_tdata2[18:0]; // @[lib.scala 104:36]
  wire  _T_1066 = _T_1065 & _T_933; // @[lib.scala 104:41]
  wire  _T_1069 = io_trigger_pkt_any_3_tdata2[19] == dec_i0_match_data_3[19]; // @[lib.scala 104:78]
  wire  _T_1070 = _T_1066 | _T_1069; // @[lib.scala 104:23]
  wire  _T_1072 = &io_trigger_pkt_any_3_tdata2[19:0]; // @[lib.scala 104:36]
  wire  _T_1073 = _T_1072 & _T_933; // @[lib.scala 104:41]
  wire  _T_1076 = io_trigger_pkt_any_3_tdata2[20] == dec_i0_match_data_3[20]; // @[lib.scala 104:78]
  wire  _T_1077 = _T_1073 | _T_1076; // @[lib.scala 104:23]
  wire  _T_1079 = &io_trigger_pkt_any_3_tdata2[20:0]; // @[lib.scala 104:36]
  wire  _T_1080 = _T_1079 & _T_933; // @[lib.scala 104:41]
  wire  _T_1083 = io_trigger_pkt_any_3_tdata2[21] == dec_i0_match_data_3[21]; // @[lib.scala 104:78]
  wire  _T_1084 = _T_1080 | _T_1083; // @[lib.scala 104:23]
  wire  _T_1086 = &io_trigger_pkt_any_3_tdata2[21:0]; // @[lib.scala 104:36]
  wire  _T_1087 = _T_1086 & _T_933; // @[lib.scala 104:41]
  wire  _T_1090 = io_trigger_pkt_any_3_tdata2[22] == dec_i0_match_data_3[22]; // @[lib.scala 104:78]
  wire  _T_1091 = _T_1087 | _T_1090; // @[lib.scala 104:23]
  wire  _T_1093 = &io_trigger_pkt_any_3_tdata2[22:0]; // @[lib.scala 104:36]
  wire  _T_1094 = _T_1093 & _T_933; // @[lib.scala 104:41]
  wire  _T_1097 = io_trigger_pkt_any_3_tdata2[23] == dec_i0_match_data_3[23]; // @[lib.scala 104:78]
  wire  _T_1098 = _T_1094 | _T_1097; // @[lib.scala 104:23]
  wire  _T_1100 = &io_trigger_pkt_any_3_tdata2[23:0]; // @[lib.scala 104:36]
  wire  _T_1101 = _T_1100 & _T_933; // @[lib.scala 104:41]
  wire  _T_1104 = io_trigger_pkt_any_3_tdata2[24] == dec_i0_match_data_3[24]; // @[lib.scala 104:78]
  wire  _T_1105 = _T_1101 | _T_1104; // @[lib.scala 104:23]
  wire  _T_1107 = &io_trigger_pkt_any_3_tdata2[24:0]; // @[lib.scala 104:36]
  wire  _T_1108 = _T_1107 & _T_933; // @[lib.scala 104:41]
  wire  _T_1111 = io_trigger_pkt_any_3_tdata2[25] == dec_i0_match_data_3[25]; // @[lib.scala 104:78]
  wire  _T_1112 = _T_1108 | _T_1111; // @[lib.scala 104:23]
  wire  _T_1114 = &io_trigger_pkt_any_3_tdata2[25:0]; // @[lib.scala 104:36]
  wire  _T_1115 = _T_1114 & _T_933; // @[lib.scala 104:41]
  wire  _T_1118 = io_trigger_pkt_any_3_tdata2[26] == dec_i0_match_data_3[26]; // @[lib.scala 104:78]
  wire  _T_1119 = _T_1115 | _T_1118; // @[lib.scala 104:23]
  wire  _T_1121 = &io_trigger_pkt_any_3_tdata2[26:0]; // @[lib.scala 104:36]
  wire  _T_1122 = _T_1121 & _T_933; // @[lib.scala 104:41]
  wire  _T_1125 = io_trigger_pkt_any_3_tdata2[27] == dec_i0_match_data_3[27]; // @[lib.scala 104:78]
  wire  _T_1126 = _T_1122 | _T_1125; // @[lib.scala 104:23]
  wire  _T_1128 = &io_trigger_pkt_any_3_tdata2[27:0]; // @[lib.scala 104:36]
  wire  _T_1129 = _T_1128 & _T_933; // @[lib.scala 104:41]
  wire  _T_1132 = io_trigger_pkt_any_3_tdata2[28] == dec_i0_match_data_3[28]; // @[lib.scala 104:78]
  wire  _T_1133 = _T_1129 | _T_1132; // @[lib.scala 104:23]
  wire  _T_1135 = &io_trigger_pkt_any_3_tdata2[28:0]; // @[lib.scala 104:36]
  wire  _T_1136 = _T_1135 & _T_933; // @[lib.scala 104:41]
  wire  _T_1139 = io_trigger_pkt_any_3_tdata2[29] == dec_i0_match_data_3[29]; // @[lib.scala 104:78]
  wire  _T_1140 = _T_1136 | _T_1139; // @[lib.scala 104:23]
  wire  _T_1142 = &io_trigger_pkt_any_3_tdata2[29:0]; // @[lib.scala 104:36]
  wire  _T_1143 = _T_1142 & _T_933; // @[lib.scala 104:41]
  wire  _T_1146 = io_trigger_pkt_any_3_tdata2[30] == dec_i0_match_data_3[30]; // @[lib.scala 104:78]
  wire  _T_1147 = _T_1143 | _T_1146; // @[lib.scala 104:23]
  wire  _T_1149 = &io_trigger_pkt_any_3_tdata2[30:0]; // @[lib.scala 104:36]
  wire  _T_1150 = _T_1149 & _T_933; // @[lib.scala 104:41]
  wire  _T_1153 = io_trigger_pkt_any_3_tdata2[31] == dec_i0_match_data_3[31]; // @[lib.scala 104:78]
  wire  _T_1154 = _T_1150 | _T_1153; // @[lib.scala 104:23]
  wire [7:0] _T_1161 = {_T_986,_T_979,_T_972,_T_965,_T_958,_T_951,_T_944,_T_937}; // @[lib.scala 105:14]
  wire [15:0] _T_1169 = {_T_1042,_T_1035,_T_1028,_T_1021,_T_1014,_T_1007,_T_1000,_T_993,_T_1161}; // @[lib.scala 105:14]
  wire [7:0] _T_1176 = {_T_1098,_T_1091,_T_1084,_T_1077,_T_1070,_T_1063,_T_1056,_T_1049}; // @[lib.scala 105:14]
  wire [31:0] _T_1185 = {_T_1154,_T_1147,_T_1140,_T_1133,_T_1126,_T_1119,_T_1112,_T_1105,_T_1176,_T_1169}; // @[lib.scala 105:14]
  wire  _T_1186 = &_T_1185; // @[lib.scala 105:25]
  wire  _T_1187 = _T_928 & _T_1186; // @[dec_trigger.scala 15:109]
  wire [2:0] _T_1189 = {_T_1187,_T_927,_T_667}; // @[Cat.scala 29:58]
  assign io_dec_i0_trigger_match_d = {_T_1189,_T_407}; // @[dec_trigger.scala 15:29]
endmodule
module dec(
  input         clock,
  input         reset,
  input         io_free_clk,
  input         io_active_clk,
  input         io_lsu_fastint_stall_any,
  output        io_dec_pause_state_cg,
  input  [30:0] io_rst_vec,
  input         io_nmi_int,
  input  [30:0] io_nmi_vec,
  input         io_i_cpu_halt_req,
  input         io_i_cpu_run_req,
  output        io_o_cpu_halt_status,
  output        io_o_cpu_halt_ack,
  output        io_o_cpu_run_ack,
  output        io_o_debug_mode_status,
  input  [27:0] io_core_id,
  input         io_mpc_debug_halt_req,
  input         io_mpc_debug_run_req,
  input         io_mpc_reset_run_req,
  output        io_mpc_debug_halt_ack,
  output        io_mpc_debug_run_ack,
  output        io_debug_brkpt_status,
  input         io_lsu_pmu_misaligned_m,
  input  [30:0] io_lsu_fir_addr,
  input  [1:0]  io_lsu_fir_error,
  input  [3:0]  io_lsu_trigger_match_m,
  input         io_lsu_idle_any,
  input         io_lsu_error_pkt_r_valid,
  input         io_lsu_error_pkt_r_bits_single_ecc_error,
  input         io_lsu_error_pkt_r_bits_inst_type,
  input         io_lsu_error_pkt_r_bits_exc_type,
  input  [3:0]  io_lsu_error_pkt_r_bits_mscause,
  input  [31:0] io_lsu_error_pkt_r_bits_addr,
  input         io_lsu_single_ecc_error_incr,
  input  [31:0] io_exu_div_result,
  input         io_exu_div_wren,
  input  [31:0] io_lsu_result_m,
  input  [31:0] io_lsu_result_corr_r,
  input         io_lsu_load_stall_any,
  input         io_lsu_store_stall_any,
  input         io_iccm_dma_sb_error,
  input         io_exu_flush_final,
  input         io_timer_int,
  input         io_soft_int,
  input         io_dbg_halt_req,
  input         io_dbg_resume_req,
  output        io_dec_tlu_dbg_halted,
  output        io_dec_tlu_debug_mode,
  output        io_dec_tlu_resume_ack,
  output        io_dec_tlu_mpc_halted_only,
  output [31:0] io_dec_dbg_rddata,
  output        io_dec_dbg_cmd_done,
  output        io_dec_dbg_cmd_fail,
  output        io_trigger_pkt_any_0_select,
  output        io_trigger_pkt_any_0_match_pkt,
  output        io_trigger_pkt_any_0_store,
  output        io_trigger_pkt_any_0_load,
  output [31:0] io_trigger_pkt_any_0_tdata2,
  output        io_trigger_pkt_any_1_select,
  output        io_trigger_pkt_any_1_match_pkt,
  output        io_trigger_pkt_any_1_store,
  output        io_trigger_pkt_any_1_load,
  output [31:0] io_trigger_pkt_any_1_tdata2,
  output        io_trigger_pkt_any_2_select,
  output        io_trigger_pkt_any_2_match_pkt,
  output        io_trigger_pkt_any_2_store,
  output        io_trigger_pkt_any_2_load,
  output [31:0] io_trigger_pkt_any_2_tdata2,
  output        io_trigger_pkt_any_3_select,
  output        io_trigger_pkt_any_3_match_pkt,
  output        io_trigger_pkt_any_3_store,
  output        io_trigger_pkt_any_3_load,
  output [31:0] io_trigger_pkt_any_3_tdata2,
  input         io_exu_i0_br_way_r,
  output        io_lsu_p_valid,
  output        io_lsu_p_bits_fast_int,
  output        io_lsu_p_bits_by,
  output        io_lsu_p_bits_half,
  output        io_lsu_p_bits_word,
  output        io_lsu_p_bits_load,
  output        io_lsu_p_bits_store,
  output        io_lsu_p_bits_unsign,
  output        io_lsu_p_bits_store_data_bypass_d,
  output        io_lsu_p_bits_load_ldst_bypass_d,
  output [11:0] io_dec_lsu_offset_d,
  output        io_dec_tlu_i0_kill_writeb_r,
  output        io_dec_tlu_perfcnt0,
  output        io_dec_tlu_perfcnt1,
  output        io_dec_tlu_perfcnt2,
  output        io_dec_tlu_perfcnt3,
  output        io_dec_lsu_valid_raw_d,
  output [1:0]  io_rv_trace_pkt_rv_i_valid_ip,
  output [31:0] io_rv_trace_pkt_rv_i_insn_ip,
  output [31:0] io_rv_trace_pkt_rv_i_address_ip,
  output [1:0]  io_rv_trace_pkt_rv_i_exception_ip,
  output [4:0]  io_rv_trace_pkt_rv_i_ecause_ip,
  output [1:0]  io_rv_trace_pkt_rv_i_interrupt_ip,
  output [31:0] io_rv_trace_pkt_rv_i_tval_ip,
  output        io_dec_tlu_misc_clk_override,
  output        io_dec_tlu_lsu_clk_override,
  output        io_dec_tlu_bus_clk_override,
  output        io_dec_tlu_pic_clk_override,
  output        io_dec_tlu_dccm_clk_override,
  output        io_dec_tlu_icm_clk_override,
  input         io_scan_mode,
  output        io_ifu_dec_dec_aln_aln_dec_dec_i0_decode_d,
  input  [15:0] io_ifu_dec_dec_aln_aln_dec_ifu_i0_cinst,
  input         io_ifu_dec_dec_aln_aln_ib_ifu_i0_icaf,
  input  [1:0]  io_ifu_dec_dec_aln_aln_ib_ifu_i0_icaf_type,
  input         io_ifu_dec_dec_aln_aln_ib_ifu_i0_icaf_f1,
  input         io_ifu_dec_dec_aln_aln_ib_ifu_i0_dbecc,
  input  [7:0]  io_ifu_dec_dec_aln_aln_ib_ifu_i0_bp_index,
  input  [7:0]  io_ifu_dec_dec_aln_aln_ib_ifu_i0_bp_fghr,
  input  [4:0]  io_ifu_dec_dec_aln_aln_ib_ifu_i0_bp_btag,
  input         io_ifu_dec_dec_aln_aln_ib_ifu_i0_valid,
  input  [31:0] io_ifu_dec_dec_aln_aln_ib_ifu_i0_instr,
  input  [30:0] io_ifu_dec_dec_aln_aln_ib_ifu_i0_pc,
  input         io_ifu_dec_dec_aln_aln_ib_ifu_i0_pc4,
  input         io_ifu_dec_dec_aln_aln_ib_i0_brp_valid,
  input  [11:0] io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_toffset,
  input  [1:0]  io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_hist,
  input         io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_br_error,
  input         io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_br_start_error,
  input  [30:0] io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_prett,
  input         io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_way,
  input         io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_ret,
  input         io_ifu_dec_dec_aln_ifu_pmu_instr_aligned,
  output        io_ifu_dec_dec_mem_ctrl_dec_tlu_flush_err_wb,
  output        io_ifu_dec_dec_mem_ctrl_dec_tlu_i0_commit_cmt,
  output        io_ifu_dec_dec_mem_ctrl_dec_tlu_force_halt,
  output        io_ifu_dec_dec_mem_ctrl_dec_tlu_fence_i_wb,
  output [70:0] io_ifu_dec_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_wrdata,
  output [16:0] io_ifu_dec_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_dicawics,
  output        io_ifu_dec_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_rd_valid,
  output        io_ifu_dec_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_wr_valid,
  output        io_ifu_dec_dec_mem_ctrl_dec_tlu_core_ecc_disable,
  input         io_ifu_dec_dec_mem_ctrl_ifu_pmu_ic_miss,
  input         io_ifu_dec_dec_mem_ctrl_ifu_pmu_ic_hit,
  input         io_ifu_dec_dec_mem_ctrl_ifu_pmu_bus_error,
  input         io_ifu_dec_dec_mem_ctrl_ifu_pmu_bus_busy,
  input         io_ifu_dec_dec_mem_ctrl_ifu_ic_error_start,
  input         io_ifu_dec_dec_mem_ctrl_ifu_iccm_rd_ecc_single_err,
  input  [70:0] io_ifu_dec_dec_mem_ctrl_ifu_ic_debug_rd_data,
  input         io_ifu_dec_dec_mem_ctrl_ifu_ic_debug_rd_data_valid,
  input         io_ifu_dec_dec_mem_ctrl_ifu_miss_state_idle,
  output        io_ifu_dec_dec_ifc_dec_tlu_flush_noredir_wb,
  output [31:0] io_ifu_dec_dec_ifc_dec_tlu_mrac_ff,
  input         io_ifu_dec_dec_ifc_ifu_pmu_fetch_stall,
  output        io_ifu_dec_dec_bp_dec_tlu_br0_r_pkt_valid,
  output [1:0]  io_ifu_dec_dec_bp_dec_tlu_br0_r_pkt_bits_hist,
  output        io_ifu_dec_dec_bp_dec_tlu_br0_r_pkt_bits_br_error,
  output        io_ifu_dec_dec_bp_dec_tlu_br0_r_pkt_bits_br_start_error,
  output        io_ifu_dec_dec_bp_dec_tlu_br0_r_pkt_bits_way,
  output        io_ifu_dec_dec_bp_dec_tlu_br0_r_pkt_bits_middle,
  output        io_ifu_dec_dec_bp_dec_tlu_flush_leak_one_wb,
  output        io_ifu_dec_dec_bp_dec_tlu_bpred_disable,
  output        io_dec_exu_dec_alu_dec_i0_alu_decode_d,
  output        io_dec_exu_dec_alu_dec_csr_ren_d,
  output [11:0] io_dec_exu_dec_alu_dec_i0_br_immed_d,
  input  [30:0] io_dec_exu_dec_alu_exu_i0_pc_x,
  output        io_dec_exu_dec_div_div_p_valid,
  output        io_dec_exu_dec_div_div_p_bits_unsign,
  output        io_dec_exu_dec_div_div_p_bits_rem,
  output        io_dec_exu_dec_div_dec_div_cancel,
  output [1:0]  io_dec_exu_decode_exu_dec_data_en,
  output [1:0]  io_dec_exu_decode_exu_dec_ctl_en,
  output        io_dec_exu_decode_exu_i0_ap_land,
  output        io_dec_exu_decode_exu_i0_ap_lor,
  output        io_dec_exu_decode_exu_i0_ap_lxor,
  output        io_dec_exu_decode_exu_i0_ap_sll,
  output        io_dec_exu_decode_exu_i0_ap_srl,
  output        io_dec_exu_decode_exu_i0_ap_sra,
  output        io_dec_exu_decode_exu_i0_ap_beq,
  output        io_dec_exu_decode_exu_i0_ap_bne,
  output        io_dec_exu_decode_exu_i0_ap_blt,
  output        io_dec_exu_decode_exu_i0_ap_bge,
  output        io_dec_exu_decode_exu_i0_ap_add,
  output        io_dec_exu_decode_exu_i0_ap_sub,
  output        io_dec_exu_decode_exu_i0_ap_slt,
  output        io_dec_exu_decode_exu_i0_ap_unsign,
  output        io_dec_exu_decode_exu_i0_ap_jal,
  output        io_dec_exu_decode_exu_i0_ap_predict_t,
  output        io_dec_exu_decode_exu_i0_ap_predict_nt,
  output        io_dec_exu_decode_exu_i0_ap_csr_write,
  output        io_dec_exu_decode_exu_i0_ap_csr_imm,
  output        io_dec_exu_decode_exu_dec_i0_predict_p_d_valid,
  output        io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_pc4,
  output [1:0]  io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_hist,
  output [11:0] io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_toffset,
  output        io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_br_error,
  output        io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_br_start_error,
  output [30:0] io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_prett,
  output        io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_pcall,
  output        io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_pret,
  output        io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_pja,
  output        io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_way,
  output [7:0]  io_dec_exu_decode_exu_i0_predict_fghr_d,
  output [7:0]  io_dec_exu_decode_exu_i0_predict_index_d,
  output [4:0]  io_dec_exu_decode_exu_i0_predict_btag_d,
  output        io_dec_exu_decode_exu_dec_i0_rs1_en_d,
  output        io_dec_exu_decode_exu_dec_i0_rs2_en_d,
  output [31:0] io_dec_exu_decode_exu_dec_i0_immed_d,
  output [31:0] io_dec_exu_decode_exu_dec_i0_rs1_bypass_data_d,
  output [31:0] io_dec_exu_decode_exu_dec_i0_rs2_bypass_data_d,
  output        io_dec_exu_decode_exu_dec_i0_select_pc_d,
  output [1:0]  io_dec_exu_decode_exu_dec_i0_rs1_bypass_en_d,
  output [1:0]  io_dec_exu_decode_exu_dec_i0_rs2_bypass_en_d,
  output        io_dec_exu_decode_exu_mul_p_valid,
  output        io_dec_exu_decode_exu_mul_p_bits_rs1_sign,
  output        io_dec_exu_decode_exu_mul_p_bits_rs2_sign,
  output        io_dec_exu_decode_exu_mul_p_bits_low,
  output [30:0] io_dec_exu_decode_exu_pred_correct_npc_x,
  output        io_dec_exu_decode_exu_dec_extint_stall,
  input  [31:0] io_dec_exu_decode_exu_exu_i0_result_x,
  input  [31:0] io_dec_exu_decode_exu_exu_csr_rs1_x,
  output [29:0] io_dec_exu_tlu_exu_dec_tlu_meihap,
  output        io_dec_exu_tlu_exu_dec_tlu_flush_lower_r,
  output [30:0] io_dec_exu_tlu_exu_dec_tlu_flush_path_r,
  input  [1:0]  io_dec_exu_tlu_exu_exu_i0_br_hist_r,
  input         io_dec_exu_tlu_exu_exu_i0_br_error_r,
  input         io_dec_exu_tlu_exu_exu_i0_br_start_error_r,
  input         io_dec_exu_tlu_exu_exu_i0_br_valid_r,
  input         io_dec_exu_tlu_exu_exu_i0_br_mp_r,
  input         io_dec_exu_tlu_exu_exu_i0_br_middle_r,
  input         io_dec_exu_tlu_exu_exu_pmu_i0_br_misp,
  input         io_dec_exu_tlu_exu_exu_pmu_i0_br_ataken,
  input         io_dec_exu_tlu_exu_exu_pmu_i0_pc4,
  input  [30:0] io_dec_exu_tlu_exu_exu_npc_r,
  output [30:0] io_dec_exu_ib_exu_dec_i0_pc_d,
  output        io_dec_exu_ib_exu_dec_debug_wdata_rs1_d,
  output [31:0] io_dec_exu_gpr_exu_gpr_i0_rs1_d,
  output [31:0] io_dec_exu_gpr_exu_gpr_i0_rs2_d,
  input         io_lsu_dec_tlu_busbuff_lsu_pmu_bus_misaligned,
  input         io_lsu_dec_tlu_busbuff_lsu_pmu_bus_error,
  input         io_lsu_dec_tlu_busbuff_lsu_pmu_bus_busy,
  output        io_lsu_dec_tlu_busbuff_dec_tlu_external_ldfwd_disable,
  output        io_lsu_dec_tlu_busbuff_dec_tlu_wb_coalescing_disable,
  output        io_lsu_dec_tlu_busbuff_dec_tlu_sideeffect_posted_disable,
  input         io_lsu_dec_tlu_busbuff_lsu_imprecise_error_load_any,
  input         io_lsu_dec_tlu_busbuff_lsu_imprecise_error_store_any,
  input  [31:0] io_lsu_dec_tlu_busbuff_lsu_imprecise_error_addr_any,
  input         io_lsu_dec_dctl_busbuff_lsu_nonblock_load_valid_m,
  input  [1:0]  io_lsu_dec_dctl_busbuff_lsu_nonblock_load_tag_m,
  input         io_lsu_dec_dctl_busbuff_lsu_nonblock_load_inv_r,
  input  [1:0]  io_lsu_dec_dctl_busbuff_lsu_nonblock_load_inv_tag_r,
  input         io_lsu_dec_dctl_busbuff_lsu_nonblock_load_data_valid,
  input         io_lsu_dec_dctl_busbuff_lsu_nonblock_load_data_error,
  input  [1:0]  io_lsu_dec_dctl_busbuff_lsu_nonblock_load_data_tag,
  input  [31:0] io_lsu_dec_dctl_busbuff_lsu_nonblock_load_data,
  input         io_lsu_tlu_lsu_pmu_load_external_m,
  input         io_lsu_tlu_lsu_pmu_store_external_m,
  input         io_dec_dbg_dbg_ib_dbg_cmd_valid,
  input         io_dec_dbg_dbg_ib_dbg_cmd_write,
  input  [1:0]  io_dec_dbg_dbg_ib_dbg_cmd_type,
  input  [31:0] io_dec_dbg_dbg_ib_dbg_cmd_addr,
  input  [31:0] io_dec_dbg_dbg_dctl_dbg_cmd_wrdata,
  input         io_dec_dma_dctl_dma_dma_dccm_stall_any,
  input         io_dec_dma_tlu_dma_dma_pmu_dccm_read,
  input         io_dec_dma_tlu_dma_dma_pmu_dccm_write,
  input         io_dec_dma_tlu_dma_dma_pmu_any_read,
  input         io_dec_dma_tlu_dma_dma_pmu_any_write,
  output [2:0]  io_dec_dma_tlu_dma_dec_tlu_dma_qos_prty,
  input         io_dec_dma_tlu_dma_dma_dccm_stall_any,
  input         io_dec_dma_tlu_dma_dma_iccm_stall_any,
  input  [7:0]  io_dec_pic_pic_claimid,
  input  [3:0]  io_dec_pic_pic_pl,
  input         io_dec_pic_mhwakeup,
  output [3:0]  io_dec_pic_dec_tlu_meicurpl,
  output [3:0]  io_dec_pic_dec_tlu_meipt,
  input         io_dec_pic_mexintpend
);
  wire  instbuff_io_ifu_ib_ifu_i0_icaf; // @[dec.scala 117:24]
  wire [1:0] instbuff_io_ifu_ib_ifu_i0_icaf_type; // @[dec.scala 117:24]
  wire  instbuff_io_ifu_ib_ifu_i0_icaf_f1; // @[dec.scala 117:24]
  wire  instbuff_io_ifu_ib_ifu_i0_dbecc; // @[dec.scala 117:24]
  wire [7:0] instbuff_io_ifu_ib_ifu_i0_bp_index; // @[dec.scala 117:24]
  wire [7:0] instbuff_io_ifu_ib_ifu_i0_bp_fghr; // @[dec.scala 117:24]
  wire [4:0] instbuff_io_ifu_ib_ifu_i0_bp_btag; // @[dec.scala 117:24]
  wire  instbuff_io_ifu_ib_ifu_i0_valid; // @[dec.scala 117:24]
  wire [31:0] instbuff_io_ifu_ib_ifu_i0_instr; // @[dec.scala 117:24]
  wire [30:0] instbuff_io_ifu_ib_ifu_i0_pc; // @[dec.scala 117:24]
  wire  instbuff_io_ifu_ib_ifu_i0_pc4; // @[dec.scala 117:24]
  wire  instbuff_io_ifu_ib_i0_brp_valid; // @[dec.scala 117:24]
  wire [11:0] instbuff_io_ifu_ib_i0_brp_bits_toffset; // @[dec.scala 117:24]
  wire [1:0] instbuff_io_ifu_ib_i0_brp_bits_hist; // @[dec.scala 117:24]
  wire  instbuff_io_ifu_ib_i0_brp_bits_br_error; // @[dec.scala 117:24]
  wire  instbuff_io_ifu_ib_i0_brp_bits_br_start_error; // @[dec.scala 117:24]
  wire [30:0] instbuff_io_ifu_ib_i0_brp_bits_prett; // @[dec.scala 117:24]
  wire  instbuff_io_ifu_ib_i0_brp_bits_way; // @[dec.scala 117:24]
  wire  instbuff_io_ifu_ib_i0_brp_bits_ret; // @[dec.scala 117:24]
  wire [30:0] instbuff_io_ib_exu_dec_i0_pc_d; // @[dec.scala 117:24]
  wire  instbuff_io_ib_exu_dec_debug_wdata_rs1_d; // @[dec.scala 117:24]
  wire  instbuff_io_dbg_ib_dbg_cmd_valid; // @[dec.scala 117:24]
  wire  instbuff_io_dbg_ib_dbg_cmd_write; // @[dec.scala 117:24]
  wire [1:0] instbuff_io_dbg_ib_dbg_cmd_type; // @[dec.scala 117:24]
  wire [31:0] instbuff_io_dbg_ib_dbg_cmd_addr; // @[dec.scala 117:24]
  wire  instbuff_io_dec_ib0_valid_d; // @[dec.scala 117:24]
  wire [1:0] instbuff_io_dec_i0_icaf_type_d; // @[dec.scala 117:24]
  wire [31:0] instbuff_io_dec_i0_instr_d; // @[dec.scala 117:24]
  wire  instbuff_io_dec_i0_pc4_d; // @[dec.scala 117:24]
  wire  instbuff_io_dec_i0_brp_valid; // @[dec.scala 117:24]
  wire [11:0] instbuff_io_dec_i0_brp_bits_toffset; // @[dec.scala 117:24]
  wire [1:0] instbuff_io_dec_i0_brp_bits_hist; // @[dec.scala 117:24]
  wire  instbuff_io_dec_i0_brp_bits_br_error; // @[dec.scala 117:24]
  wire  instbuff_io_dec_i0_brp_bits_br_start_error; // @[dec.scala 117:24]
  wire [30:0] instbuff_io_dec_i0_brp_bits_prett; // @[dec.scala 117:24]
  wire  instbuff_io_dec_i0_brp_bits_way; // @[dec.scala 117:24]
  wire  instbuff_io_dec_i0_brp_bits_ret; // @[dec.scala 117:24]
  wire [7:0] instbuff_io_dec_i0_bp_index; // @[dec.scala 117:24]
  wire [7:0] instbuff_io_dec_i0_bp_fghr; // @[dec.scala 117:24]
  wire [4:0] instbuff_io_dec_i0_bp_btag; // @[dec.scala 117:24]
  wire  instbuff_io_dec_i0_icaf_d; // @[dec.scala 117:24]
  wire  instbuff_io_dec_i0_icaf_f1_d; // @[dec.scala 117:24]
  wire  instbuff_io_dec_i0_dbecc_d; // @[dec.scala 117:24]
  wire  instbuff_io_dec_debug_fence_d; // @[dec.scala 117:24]
  wire  decode_clock; // @[dec.scala 118:22]
  wire  decode_reset; // @[dec.scala 118:22]
  wire [1:0] decode_io_decode_exu_dec_data_en; // @[dec.scala 118:22]
  wire [1:0] decode_io_decode_exu_dec_ctl_en; // @[dec.scala 118:22]
  wire  decode_io_decode_exu_i0_ap_land; // @[dec.scala 118:22]
  wire  decode_io_decode_exu_i0_ap_lor; // @[dec.scala 118:22]
  wire  decode_io_decode_exu_i0_ap_lxor; // @[dec.scala 118:22]
  wire  decode_io_decode_exu_i0_ap_sll; // @[dec.scala 118:22]
  wire  decode_io_decode_exu_i0_ap_srl; // @[dec.scala 118:22]
  wire  decode_io_decode_exu_i0_ap_sra; // @[dec.scala 118:22]
  wire  decode_io_decode_exu_i0_ap_beq; // @[dec.scala 118:22]
  wire  decode_io_decode_exu_i0_ap_bne; // @[dec.scala 118:22]
  wire  decode_io_decode_exu_i0_ap_blt; // @[dec.scala 118:22]
  wire  decode_io_decode_exu_i0_ap_bge; // @[dec.scala 118:22]
  wire  decode_io_decode_exu_i0_ap_add; // @[dec.scala 118:22]
  wire  decode_io_decode_exu_i0_ap_sub; // @[dec.scala 118:22]
  wire  decode_io_decode_exu_i0_ap_slt; // @[dec.scala 118:22]
  wire  decode_io_decode_exu_i0_ap_unsign; // @[dec.scala 118:22]
  wire  decode_io_decode_exu_i0_ap_jal; // @[dec.scala 118:22]
  wire  decode_io_decode_exu_i0_ap_predict_t; // @[dec.scala 118:22]
  wire  decode_io_decode_exu_i0_ap_predict_nt; // @[dec.scala 118:22]
  wire  decode_io_decode_exu_i0_ap_csr_write; // @[dec.scala 118:22]
  wire  decode_io_decode_exu_i0_ap_csr_imm; // @[dec.scala 118:22]
  wire  decode_io_decode_exu_dec_i0_predict_p_d_valid; // @[dec.scala 118:22]
  wire  decode_io_decode_exu_dec_i0_predict_p_d_bits_pc4; // @[dec.scala 118:22]
  wire [1:0] decode_io_decode_exu_dec_i0_predict_p_d_bits_hist; // @[dec.scala 118:22]
  wire [11:0] decode_io_decode_exu_dec_i0_predict_p_d_bits_toffset; // @[dec.scala 118:22]
  wire  decode_io_decode_exu_dec_i0_predict_p_d_bits_br_error; // @[dec.scala 118:22]
  wire  decode_io_decode_exu_dec_i0_predict_p_d_bits_br_start_error; // @[dec.scala 118:22]
  wire [30:0] decode_io_decode_exu_dec_i0_predict_p_d_bits_prett; // @[dec.scala 118:22]
  wire  decode_io_decode_exu_dec_i0_predict_p_d_bits_pcall; // @[dec.scala 118:22]
  wire  decode_io_decode_exu_dec_i0_predict_p_d_bits_pret; // @[dec.scala 118:22]
  wire  decode_io_decode_exu_dec_i0_predict_p_d_bits_pja; // @[dec.scala 118:22]
  wire  decode_io_decode_exu_dec_i0_predict_p_d_bits_way; // @[dec.scala 118:22]
  wire [7:0] decode_io_decode_exu_i0_predict_fghr_d; // @[dec.scala 118:22]
  wire [7:0] decode_io_decode_exu_i0_predict_index_d; // @[dec.scala 118:22]
  wire [4:0] decode_io_decode_exu_i0_predict_btag_d; // @[dec.scala 118:22]
  wire  decode_io_decode_exu_dec_i0_rs1_en_d; // @[dec.scala 118:22]
  wire  decode_io_decode_exu_dec_i0_rs2_en_d; // @[dec.scala 118:22]
  wire [31:0] decode_io_decode_exu_dec_i0_immed_d; // @[dec.scala 118:22]
  wire [31:0] decode_io_decode_exu_dec_i0_rs1_bypass_data_d; // @[dec.scala 118:22]
  wire [31:0] decode_io_decode_exu_dec_i0_rs2_bypass_data_d; // @[dec.scala 118:22]
  wire  decode_io_decode_exu_dec_i0_select_pc_d; // @[dec.scala 118:22]
  wire [1:0] decode_io_decode_exu_dec_i0_rs1_bypass_en_d; // @[dec.scala 118:22]
  wire [1:0] decode_io_decode_exu_dec_i0_rs2_bypass_en_d; // @[dec.scala 118:22]
  wire  decode_io_decode_exu_mul_p_valid; // @[dec.scala 118:22]
  wire  decode_io_decode_exu_mul_p_bits_rs1_sign; // @[dec.scala 118:22]
  wire  decode_io_decode_exu_mul_p_bits_rs2_sign; // @[dec.scala 118:22]
  wire  decode_io_decode_exu_mul_p_bits_low; // @[dec.scala 118:22]
  wire [30:0] decode_io_decode_exu_pred_correct_npc_x; // @[dec.scala 118:22]
  wire  decode_io_decode_exu_dec_extint_stall; // @[dec.scala 118:22]
  wire [31:0] decode_io_decode_exu_exu_i0_result_x; // @[dec.scala 118:22]
  wire [31:0] decode_io_decode_exu_exu_csr_rs1_x; // @[dec.scala 118:22]
  wire  decode_io_dec_alu_dec_i0_alu_decode_d; // @[dec.scala 118:22]
  wire  decode_io_dec_alu_dec_csr_ren_d; // @[dec.scala 118:22]
  wire [11:0] decode_io_dec_alu_dec_i0_br_immed_d; // @[dec.scala 118:22]
  wire [30:0] decode_io_dec_alu_exu_i0_pc_x; // @[dec.scala 118:22]
  wire  decode_io_dec_div_div_p_valid; // @[dec.scala 118:22]
  wire  decode_io_dec_div_div_p_bits_unsign; // @[dec.scala 118:22]
  wire  decode_io_dec_div_div_p_bits_rem; // @[dec.scala 118:22]
  wire  decode_io_dec_div_dec_div_cancel; // @[dec.scala 118:22]
  wire  decode_io_dctl_busbuff_lsu_nonblock_load_valid_m; // @[dec.scala 118:22]
  wire [1:0] decode_io_dctl_busbuff_lsu_nonblock_load_tag_m; // @[dec.scala 118:22]
  wire  decode_io_dctl_busbuff_lsu_nonblock_load_inv_r; // @[dec.scala 118:22]
  wire [1:0] decode_io_dctl_busbuff_lsu_nonblock_load_inv_tag_r; // @[dec.scala 118:22]
  wire  decode_io_dctl_busbuff_lsu_nonblock_load_data_valid; // @[dec.scala 118:22]
  wire  decode_io_dctl_busbuff_lsu_nonblock_load_data_error; // @[dec.scala 118:22]
  wire [1:0] decode_io_dctl_busbuff_lsu_nonblock_load_data_tag; // @[dec.scala 118:22]
  wire [31:0] decode_io_dctl_busbuff_lsu_nonblock_load_data; // @[dec.scala 118:22]
  wire  decode_io_dctl_dma_dma_dccm_stall_any; // @[dec.scala 118:22]
  wire  decode_io_dec_aln_dec_i0_decode_d; // @[dec.scala 118:22]
  wire [15:0] decode_io_dec_aln_ifu_i0_cinst; // @[dec.scala 118:22]
  wire [31:0] decode_io_dbg_dctl_dbg_cmd_wrdata; // @[dec.scala 118:22]
  wire  decode_io_dec_tlu_flush_extint; // @[dec.scala 118:22]
  wire  decode_io_dec_tlu_force_halt; // @[dec.scala 118:22]
  wire [31:0] decode_io_dec_i0_inst_wb1; // @[dec.scala 118:22]
  wire [30:0] decode_io_dec_i0_pc_wb1; // @[dec.scala 118:22]
  wire [3:0] decode_io_dec_i0_trigger_match_d; // @[dec.scala 118:22]
  wire  decode_io_dec_tlu_wr_pause_r; // @[dec.scala 118:22]
  wire  decode_io_dec_tlu_pipelining_disable; // @[dec.scala 118:22]
  wire [3:0] decode_io_lsu_trigger_match_m; // @[dec.scala 118:22]
  wire  decode_io_lsu_pmu_misaligned_m; // @[dec.scala 118:22]
  wire  decode_io_dec_tlu_debug_stall; // @[dec.scala 118:22]
  wire  decode_io_dec_tlu_flush_leak_one_r; // @[dec.scala 118:22]
  wire  decode_io_dec_debug_fence_d; // @[dec.scala 118:22]
  wire  decode_io_dec_i0_icaf_d; // @[dec.scala 118:22]
  wire  decode_io_dec_i0_icaf_f1_d; // @[dec.scala 118:22]
  wire [1:0] decode_io_dec_i0_icaf_type_d; // @[dec.scala 118:22]
  wire  decode_io_dec_i0_dbecc_d; // @[dec.scala 118:22]
  wire  decode_io_dec_i0_brp_valid; // @[dec.scala 118:22]
  wire [11:0] decode_io_dec_i0_brp_bits_toffset; // @[dec.scala 118:22]
  wire [1:0] decode_io_dec_i0_brp_bits_hist; // @[dec.scala 118:22]
  wire  decode_io_dec_i0_brp_bits_br_error; // @[dec.scala 118:22]
  wire  decode_io_dec_i0_brp_bits_br_start_error; // @[dec.scala 118:22]
  wire [30:0] decode_io_dec_i0_brp_bits_prett; // @[dec.scala 118:22]
  wire  decode_io_dec_i0_brp_bits_way; // @[dec.scala 118:22]
  wire  decode_io_dec_i0_brp_bits_ret; // @[dec.scala 118:22]
  wire [7:0] decode_io_dec_i0_bp_index; // @[dec.scala 118:22]
  wire [7:0] decode_io_dec_i0_bp_fghr; // @[dec.scala 118:22]
  wire [4:0] decode_io_dec_i0_bp_btag; // @[dec.scala 118:22]
  wire  decode_io_lsu_idle_any; // @[dec.scala 118:22]
  wire  decode_io_lsu_load_stall_any; // @[dec.scala 118:22]
  wire  decode_io_lsu_store_stall_any; // @[dec.scala 118:22]
  wire  decode_io_exu_div_wren; // @[dec.scala 118:22]
  wire  decode_io_dec_tlu_i0_kill_writeb_wb; // @[dec.scala 118:22]
  wire  decode_io_dec_tlu_flush_lower_wb; // @[dec.scala 118:22]
  wire  decode_io_dec_tlu_i0_kill_writeb_r; // @[dec.scala 118:22]
  wire  decode_io_dec_tlu_flush_lower_r; // @[dec.scala 118:22]
  wire  decode_io_dec_tlu_flush_pause_r; // @[dec.scala 118:22]
  wire  decode_io_dec_tlu_presync_d; // @[dec.scala 118:22]
  wire  decode_io_dec_tlu_postsync_d; // @[dec.scala 118:22]
  wire  decode_io_dec_i0_pc4_d; // @[dec.scala 118:22]
  wire [31:0] decode_io_dec_csr_rddata_d; // @[dec.scala 118:22]
  wire  decode_io_dec_csr_legal_d; // @[dec.scala 118:22]
  wire [31:0] decode_io_lsu_result_m; // @[dec.scala 118:22]
  wire [31:0] decode_io_lsu_result_corr_r; // @[dec.scala 118:22]
  wire  decode_io_exu_flush_final; // @[dec.scala 118:22]
  wire [31:0] decode_io_dec_i0_instr_d; // @[dec.scala 118:22]
  wire  decode_io_dec_ib0_valid_d; // @[dec.scala 118:22]
  wire  decode_io_free_clk; // @[dec.scala 118:22]
  wire  decode_io_active_clk; // @[dec.scala 118:22]
  wire  decode_io_clk_override; // @[dec.scala 118:22]
  wire [4:0] decode_io_dec_i0_rs1_d; // @[dec.scala 118:22]
  wire [4:0] decode_io_dec_i0_rs2_d; // @[dec.scala 118:22]
  wire [4:0] decode_io_dec_i0_waddr_r; // @[dec.scala 118:22]
  wire  decode_io_dec_i0_wen_r; // @[dec.scala 118:22]
  wire [31:0] decode_io_dec_i0_wdata_r; // @[dec.scala 118:22]
  wire  decode_io_lsu_p_valid; // @[dec.scala 118:22]
  wire  decode_io_lsu_p_bits_fast_int; // @[dec.scala 118:22]
  wire  decode_io_lsu_p_bits_by; // @[dec.scala 118:22]
  wire  decode_io_lsu_p_bits_half; // @[dec.scala 118:22]
  wire  decode_io_lsu_p_bits_word; // @[dec.scala 118:22]
  wire  decode_io_lsu_p_bits_load; // @[dec.scala 118:22]
  wire  decode_io_lsu_p_bits_store; // @[dec.scala 118:22]
  wire  decode_io_lsu_p_bits_unsign; // @[dec.scala 118:22]
  wire  decode_io_lsu_p_bits_store_data_bypass_d; // @[dec.scala 118:22]
  wire  decode_io_lsu_p_bits_load_ldst_bypass_d; // @[dec.scala 118:22]
  wire [4:0] decode_io_div_waddr_wb; // @[dec.scala 118:22]
  wire  decode_io_dec_lsu_valid_raw_d; // @[dec.scala 118:22]
  wire [11:0] decode_io_dec_lsu_offset_d; // @[dec.scala 118:22]
  wire  decode_io_dec_csr_wen_unq_d; // @[dec.scala 118:22]
  wire  decode_io_dec_csr_any_unq_d; // @[dec.scala 118:22]
  wire [11:0] decode_io_dec_csr_rdaddr_d; // @[dec.scala 118:22]
  wire  decode_io_dec_csr_wen_r; // @[dec.scala 118:22]
  wire [11:0] decode_io_dec_csr_wraddr_r; // @[dec.scala 118:22]
  wire [31:0] decode_io_dec_csr_wrdata_r; // @[dec.scala 118:22]
  wire  decode_io_dec_csr_stall_int_ff; // @[dec.scala 118:22]
  wire  decode_io_dec_tlu_i0_valid_r; // @[dec.scala 118:22]
  wire  decode_io_dec_tlu_packet_r_legal; // @[dec.scala 118:22]
  wire  decode_io_dec_tlu_packet_r_icaf; // @[dec.scala 118:22]
  wire  decode_io_dec_tlu_packet_r_icaf_f1; // @[dec.scala 118:22]
  wire [1:0] decode_io_dec_tlu_packet_r_icaf_type; // @[dec.scala 118:22]
  wire  decode_io_dec_tlu_packet_r_fence_i; // @[dec.scala 118:22]
  wire [3:0] decode_io_dec_tlu_packet_r_i0trigger; // @[dec.scala 118:22]
  wire [3:0] decode_io_dec_tlu_packet_r_pmu_i0_itype; // @[dec.scala 118:22]
  wire  decode_io_dec_tlu_packet_r_pmu_i0_br_unpred; // @[dec.scala 118:22]
  wire  decode_io_dec_tlu_packet_r_pmu_divide; // @[dec.scala 118:22]
  wire  decode_io_dec_tlu_packet_r_pmu_lsu_misaligned; // @[dec.scala 118:22]
  wire [30:0] decode_io_dec_tlu_i0_pc_r; // @[dec.scala 118:22]
  wire [31:0] decode_io_dec_illegal_inst; // @[dec.scala 118:22]
  wire  decode_io_dec_pmu_instr_decoded; // @[dec.scala 118:22]
  wire  decode_io_dec_pmu_decode_stall; // @[dec.scala 118:22]
  wire  decode_io_dec_pmu_presync_stall; // @[dec.scala 118:22]
  wire  decode_io_dec_pmu_postsync_stall; // @[dec.scala 118:22]
  wire  decode_io_dec_nonblock_load_wen; // @[dec.scala 118:22]
  wire [4:0] decode_io_dec_nonblock_load_waddr; // @[dec.scala 118:22]
  wire  decode_io_dec_pause_state; // @[dec.scala 118:22]
  wire  decode_io_dec_pause_state_cg; // @[dec.scala 118:22]
  wire  decode_io_dec_div_active; // @[dec.scala 118:22]
  wire  decode_io_scan_mode; // @[dec.scala 118:22]
  wire  gpr_clock; // @[dec.scala 119:19]
  wire  gpr_reset; // @[dec.scala 119:19]
  wire [4:0] gpr_io_raddr0; // @[dec.scala 119:19]
  wire [4:0] gpr_io_raddr1; // @[dec.scala 119:19]
  wire  gpr_io_wen0; // @[dec.scala 119:19]
  wire [4:0] gpr_io_waddr0; // @[dec.scala 119:19]
  wire [31:0] gpr_io_wd0; // @[dec.scala 119:19]
  wire  gpr_io_wen1; // @[dec.scala 119:19]
  wire [4:0] gpr_io_waddr1; // @[dec.scala 119:19]
  wire [31:0] gpr_io_wd1; // @[dec.scala 119:19]
  wire  gpr_io_wen2; // @[dec.scala 119:19]
  wire [4:0] gpr_io_waddr2; // @[dec.scala 119:19]
  wire [31:0] gpr_io_wd2; // @[dec.scala 119:19]
  wire  gpr_io_scan_mode; // @[dec.scala 119:19]
  wire [31:0] gpr_io_gpr_exu_gpr_i0_rs1_d; // @[dec.scala 119:19]
  wire [31:0] gpr_io_gpr_exu_gpr_i0_rs2_d; // @[dec.scala 119:19]
  wire  tlu_clock; // @[dec.scala 120:19]
  wire  tlu_reset; // @[dec.scala 120:19]
  wire [29:0] tlu_io_tlu_exu_dec_tlu_meihap; // @[dec.scala 120:19]
  wire  tlu_io_tlu_exu_dec_tlu_flush_lower_r; // @[dec.scala 120:19]
  wire [30:0] tlu_io_tlu_exu_dec_tlu_flush_path_r; // @[dec.scala 120:19]
  wire [1:0] tlu_io_tlu_exu_exu_i0_br_hist_r; // @[dec.scala 120:19]
  wire  tlu_io_tlu_exu_exu_i0_br_error_r; // @[dec.scala 120:19]
  wire  tlu_io_tlu_exu_exu_i0_br_start_error_r; // @[dec.scala 120:19]
  wire  tlu_io_tlu_exu_exu_i0_br_valid_r; // @[dec.scala 120:19]
  wire  tlu_io_tlu_exu_exu_i0_br_mp_r; // @[dec.scala 120:19]
  wire  tlu_io_tlu_exu_exu_i0_br_middle_r; // @[dec.scala 120:19]
  wire  tlu_io_tlu_exu_exu_pmu_i0_br_misp; // @[dec.scala 120:19]
  wire  tlu_io_tlu_exu_exu_pmu_i0_br_ataken; // @[dec.scala 120:19]
  wire  tlu_io_tlu_exu_exu_pmu_i0_pc4; // @[dec.scala 120:19]
  wire [30:0] tlu_io_tlu_exu_exu_npc_r; // @[dec.scala 120:19]
  wire  tlu_io_tlu_dma_dma_pmu_dccm_read; // @[dec.scala 120:19]
  wire  tlu_io_tlu_dma_dma_pmu_dccm_write; // @[dec.scala 120:19]
  wire  tlu_io_tlu_dma_dma_pmu_any_read; // @[dec.scala 120:19]
  wire  tlu_io_tlu_dma_dma_pmu_any_write; // @[dec.scala 120:19]
  wire [2:0] tlu_io_tlu_dma_dec_tlu_dma_qos_prty; // @[dec.scala 120:19]
  wire  tlu_io_tlu_dma_dma_dccm_stall_any; // @[dec.scala 120:19]
  wire  tlu_io_tlu_dma_dma_iccm_stall_any; // @[dec.scala 120:19]
  wire  tlu_io_active_clk; // @[dec.scala 120:19]
  wire  tlu_io_free_clk; // @[dec.scala 120:19]
  wire  tlu_io_scan_mode; // @[dec.scala 120:19]
  wire [30:0] tlu_io_rst_vec; // @[dec.scala 120:19]
  wire  tlu_io_nmi_int; // @[dec.scala 120:19]
  wire [30:0] tlu_io_nmi_vec; // @[dec.scala 120:19]
  wire  tlu_io_i_cpu_halt_req; // @[dec.scala 120:19]
  wire  tlu_io_i_cpu_run_req; // @[dec.scala 120:19]
  wire  tlu_io_lsu_fastint_stall_any; // @[dec.scala 120:19]
  wire  tlu_io_lsu_idle_any; // @[dec.scala 120:19]
  wire  tlu_io_dec_pmu_instr_decoded; // @[dec.scala 120:19]
  wire  tlu_io_dec_pmu_decode_stall; // @[dec.scala 120:19]
  wire  tlu_io_dec_pmu_presync_stall; // @[dec.scala 120:19]
  wire  tlu_io_dec_pmu_postsync_stall; // @[dec.scala 120:19]
  wire  tlu_io_lsu_store_stall_any; // @[dec.scala 120:19]
  wire [30:0] tlu_io_lsu_fir_addr; // @[dec.scala 120:19]
  wire [1:0] tlu_io_lsu_fir_error; // @[dec.scala 120:19]
  wire  tlu_io_iccm_dma_sb_error; // @[dec.scala 120:19]
  wire  tlu_io_lsu_error_pkt_r_valid; // @[dec.scala 120:19]
  wire  tlu_io_lsu_error_pkt_r_bits_single_ecc_error; // @[dec.scala 120:19]
  wire  tlu_io_lsu_error_pkt_r_bits_inst_type; // @[dec.scala 120:19]
  wire  tlu_io_lsu_error_pkt_r_bits_exc_type; // @[dec.scala 120:19]
  wire [3:0] tlu_io_lsu_error_pkt_r_bits_mscause; // @[dec.scala 120:19]
  wire [31:0] tlu_io_lsu_error_pkt_r_bits_addr; // @[dec.scala 120:19]
  wire  tlu_io_lsu_single_ecc_error_incr; // @[dec.scala 120:19]
  wire  tlu_io_dec_pause_state; // @[dec.scala 120:19]
  wire  tlu_io_dec_csr_wen_unq_d; // @[dec.scala 120:19]
  wire  tlu_io_dec_csr_any_unq_d; // @[dec.scala 120:19]
  wire [11:0] tlu_io_dec_csr_rdaddr_d; // @[dec.scala 120:19]
  wire  tlu_io_dec_csr_wen_r; // @[dec.scala 120:19]
  wire [11:0] tlu_io_dec_csr_wraddr_r; // @[dec.scala 120:19]
  wire [31:0] tlu_io_dec_csr_wrdata_r; // @[dec.scala 120:19]
  wire  tlu_io_dec_csr_stall_int_ff; // @[dec.scala 120:19]
  wire  tlu_io_dec_tlu_i0_valid_r; // @[dec.scala 120:19]
  wire [30:0] tlu_io_dec_tlu_i0_pc_r; // @[dec.scala 120:19]
  wire  tlu_io_dec_tlu_packet_r_legal; // @[dec.scala 120:19]
  wire  tlu_io_dec_tlu_packet_r_icaf; // @[dec.scala 120:19]
  wire  tlu_io_dec_tlu_packet_r_icaf_f1; // @[dec.scala 120:19]
  wire [1:0] tlu_io_dec_tlu_packet_r_icaf_type; // @[dec.scala 120:19]
  wire  tlu_io_dec_tlu_packet_r_fence_i; // @[dec.scala 120:19]
  wire [3:0] tlu_io_dec_tlu_packet_r_i0trigger; // @[dec.scala 120:19]
  wire [3:0] tlu_io_dec_tlu_packet_r_pmu_i0_itype; // @[dec.scala 120:19]
  wire  tlu_io_dec_tlu_packet_r_pmu_i0_br_unpred; // @[dec.scala 120:19]
  wire  tlu_io_dec_tlu_packet_r_pmu_divide; // @[dec.scala 120:19]
  wire  tlu_io_dec_tlu_packet_r_pmu_lsu_misaligned; // @[dec.scala 120:19]
  wire [31:0] tlu_io_dec_illegal_inst; // @[dec.scala 120:19]
  wire  tlu_io_dec_i0_decode_d; // @[dec.scala 120:19]
  wire  tlu_io_exu_i0_br_way_r; // @[dec.scala 120:19]
  wire  tlu_io_dec_dbg_cmd_done; // @[dec.scala 120:19]
  wire  tlu_io_dec_dbg_cmd_fail; // @[dec.scala 120:19]
  wire  tlu_io_dec_tlu_dbg_halted; // @[dec.scala 120:19]
  wire  tlu_io_dec_tlu_debug_mode; // @[dec.scala 120:19]
  wire  tlu_io_dec_tlu_resume_ack; // @[dec.scala 120:19]
  wire  tlu_io_dec_tlu_debug_stall; // @[dec.scala 120:19]
  wire  tlu_io_dec_tlu_mpc_halted_only; // @[dec.scala 120:19]
  wire  tlu_io_dec_tlu_flush_extint; // @[dec.scala 120:19]
  wire  tlu_io_dbg_halt_req; // @[dec.scala 120:19]
  wire  tlu_io_dbg_resume_req; // @[dec.scala 120:19]
  wire  tlu_io_dec_div_active; // @[dec.scala 120:19]
  wire  tlu_io_trigger_pkt_any_0_select; // @[dec.scala 120:19]
  wire  tlu_io_trigger_pkt_any_0_match_pkt; // @[dec.scala 120:19]
  wire  tlu_io_trigger_pkt_any_0_store; // @[dec.scala 120:19]
  wire  tlu_io_trigger_pkt_any_0_load; // @[dec.scala 120:19]
  wire  tlu_io_trigger_pkt_any_0_execute; // @[dec.scala 120:19]
  wire  tlu_io_trigger_pkt_any_0_m; // @[dec.scala 120:19]
  wire [31:0] tlu_io_trigger_pkt_any_0_tdata2; // @[dec.scala 120:19]
  wire  tlu_io_trigger_pkt_any_1_select; // @[dec.scala 120:19]
  wire  tlu_io_trigger_pkt_any_1_match_pkt; // @[dec.scala 120:19]
  wire  tlu_io_trigger_pkt_any_1_store; // @[dec.scala 120:19]
  wire  tlu_io_trigger_pkt_any_1_load; // @[dec.scala 120:19]
  wire  tlu_io_trigger_pkt_any_1_execute; // @[dec.scala 120:19]
  wire  tlu_io_trigger_pkt_any_1_m; // @[dec.scala 120:19]
  wire [31:0] tlu_io_trigger_pkt_any_1_tdata2; // @[dec.scala 120:19]
  wire  tlu_io_trigger_pkt_any_2_select; // @[dec.scala 120:19]
  wire  tlu_io_trigger_pkt_any_2_match_pkt; // @[dec.scala 120:19]
  wire  tlu_io_trigger_pkt_any_2_store; // @[dec.scala 120:19]
  wire  tlu_io_trigger_pkt_any_2_load; // @[dec.scala 120:19]
  wire  tlu_io_trigger_pkt_any_2_execute; // @[dec.scala 120:19]
  wire  tlu_io_trigger_pkt_any_2_m; // @[dec.scala 120:19]
  wire [31:0] tlu_io_trigger_pkt_any_2_tdata2; // @[dec.scala 120:19]
  wire  tlu_io_trigger_pkt_any_3_select; // @[dec.scala 120:19]
  wire  tlu_io_trigger_pkt_any_3_match_pkt; // @[dec.scala 120:19]
  wire  tlu_io_trigger_pkt_any_3_store; // @[dec.scala 120:19]
  wire  tlu_io_trigger_pkt_any_3_load; // @[dec.scala 120:19]
  wire  tlu_io_trigger_pkt_any_3_execute; // @[dec.scala 120:19]
  wire  tlu_io_trigger_pkt_any_3_m; // @[dec.scala 120:19]
  wire [31:0] tlu_io_trigger_pkt_any_3_tdata2; // @[dec.scala 120:19]
  wire  tlu_io_timer_int; // @[dec.scala 120:19]
  wire  tlu_io_soft_int; // @[dec.scala 120:19]
  wire  tlu_io_o_cpu_halt_status; // @[dec.scala 120:19]
  wire  tlu_io_o_cpu_halt_ack; // @[dec.scala 120:19]
  wire  tlu_io_o_cpu_run_ack; // @[dec.scala 120:19]
  wire  tlu_io_o_debug_mode_status; // @[dec.scala 120:19]
  wire [27:0] tlu_io_core_id; // @[dec.scala 120:19]
  wire  tlu_io_mpc_debug_halt_req; // @[dec.scala 120:19]
  wire  tlu_io_mpc_debug_run_req; // @[dec.scala 120:19]
  wire  tlu_io_mpc_reset_run_req; // @[dec.scala 120:19]
  wire  tlu_io_mpc_debug_halt_ack; // @[dec.scala 120:19]
  wire  tlu_io_mpc_debug_run_ack; // @[dec.scala 120:19]
  wire  tlu_io_debug_brkpt_status; // @[dec.scala 120:19]
  wire [31:0] tlu_io_dec_csr_rddata_d; // @[dec.scala 120:19]
  wire  tlu_io_dec_csr_legal_d; // @[dec.scala 120:19]
  wire  tlu_io_dec_tlu_i0_kill_writeb_wb; // @[dec.scala 120:19]
  wire  tlu_io_dec_tlu_i0_kill_writeb_r; // @[dec.scala 120:19]
  wire  tlu_io_dec_tlu_wr_pause_r; // @[dec.scala 120:19]
  wire  tlu_io_dec_tlu_flush_pause_r; // @[dec.scala 120:19]
  wire  tlu_io_dec_tlu_presync_d; // @[dec.scala 120:19]
  wire  tlu_io_dec_tlu_postsync_d; // @[dec.scala 120:19]
  wire  tlu_io_dec_tlu_perfcnt0; // @[dec.scala 120:19]
  wire  tlu_io_dec_tlu_perfcnt1; // @[dec.scala 120:19]
  wire  tlu_io_dec_tlu_perfcnt2; // @[dec.scala 120:19]
  wire  tlu_io_dec_tlu_perfcnt3; // @[dec.scala 120:19]
  wire  tlu_io_dec_tlu_i0_exc_valid_wb1; // @[dec.scala 120:19]
  wire  tlu_io_dec_tlu_i0_valid_wb1; // @[dec.scala 120:19]
  wire  tlu_io_dec_tlu_int_valid_wb1; // @[dec.scala 120:19]
  wire [4:0] tlu_io_dec_tlu_exc_cause_wb1; // @[dec.scala 120:19]
  wire [31:0] tlu_io_dec_tlu_mtval_wb1; // @[dec.scala 120:19]
  wire  tlu_io_dec_tlu_pipelining_disable; // @[dec.scala 120:19]
  wire  tlu_io_dec_tlu_misc_clk_override; // @[dec.scala 120:19]
  wire  tlu_io_dec_tlu_dec_clk_override; // @[dec.scala 120:19]
  wire  tlu_io_dec_tlu_lsu_clk_override; // @[dec.scala 120:19]
  wire  tlu_io_dec_tlu_bus_clk_override; // @[dec.scala 120:19]
  wire  tlu_io_dec_tlu_pic_clk_override; // @[dec.scala 120:19]
  wire  tlu_io_dec_tlu_dccm_clk_override; // @[dec.scala 120:19]
  wire  tlu_io_dec_tlu_icm_clk_override; // @[dec.scala 120:19]
  wire  tlu_io_dec_tlu_flush_lower_wb; // @[dec.scala 120:19]
  wire  tlu_io_ifu_pmu_instr_aligned; // @[dec.scala 120:19]
  wire  tlu_io_tlu_bp_dec_tlu_br0_r_pkt_valid; // @[dec.scala 120:19]
  wire [1:0] tlu_io_tlu_bp_dec_tlu_br0_r_pkt_bits_hist; // @[dec.scala 120:19]
  wire  tlu_io_tlu_bp_dec_tlu_br0_r_pkt_bits_br_error; // @[dec.scala 120:19]
  wire  tlu_io_tlu_bp_dec_tlu_br0_r_pkt_bits_br_start_error; // @[dec.scala 120:19]
  wire  tlu_io_tlu_bp_dec_tlu_br0_r_pkt_bits_way; // @[dec.scala 120:19]
  wire  tlu_io_tlu_bp_dec_tlu_br0_r_pkt_bits_middle; // @[dec.scala 120:19]
  wire  tlu_io_tlu_bp_dec_tlu_flush_leak_one_wb; // @[dec.scala 120:19]
  wire  tlu_io_tlu_bp_dec_tlu_bpred_disable; // @[dec.scala 120:19]
  wire  tlu_io_tlu_ifc_dec_tlu_flush_noredir_wb; // @[dec.scala 120:19]
  wire [31:0] tlu_io_tlu_ifc_dec_tlu_mrac_ff; // @[dec.scala 120:19]
  wire  tlu_io_tlu_ifc_ifu_pmu_fetch_stall; // @[dec.scala 120:19]
  wire  tlu_io_tlu_mem_dec_tlu_flush_err_wb; // @[dec.scala 120:19]
  wire  tlu_io_tlu_mem_dec_tlu_i0_commit_cmt; // @[dec.scala 120:19]
  wire  tlu_io_tlu_mem_dec_tlu_force_halt; // @[dec.scala 120:19]
  wire  tlu_io_tlu_mem_dec_tlu_fence_i_wb; // @[dec.scala 120:19]
  wire [70:0] tlu_io_tlu_mem_dec_tlu_ic_diag_pkt_icache_wrdata; // @[dec.scala 120:19]
  wire [16:0] tlu_io_tlu_mem_dec_tlu_ic_diag_pkt_icache_dicawics; // @[dec.scala 120:19]
  wire  tlu_io_tlu_mem_dec_tlu_ic_diag_pkt_icache_rd_valid; // @[dec.scala 120:19]
  wire  tlu_io_tlu_mem_dec_tlu_ic_diag_pkt_icache_wr_valid; // @[dec.scala 120:19]
  wire  tlu_io_tlu_mem_dec_tlu_core_ecc_disable; // @[dec.scala 120:19]
  wire  tlu_io_tlu_mem_ifu_pmu_ic_miss; // @[dec.scala 120:19]
  wire  tlu_io_tlu_mem_ifu_pmu_ic_hit; // @[dec.scala 120:19]
  wire  tlu_io_tlu_mem_ifu_pmu_bus_error; // @[dec.scala 120:19]
  wire  tlu_io_tlu_mem_ifu_pmu_bus_busy; // @[dec.scala 120:19]
  wire  tlu_io_tlu_mem_ifu_ic_error_start; // @[dec.scala 120:19]
  wire  tlu_io_tlu_mem_ifu_iccm_rd_ecc_single_err; // @[dec.scala 120:19]
  wire [70:0] tlu_io_tlu_mem_ifu_ic_debug_rd_data; // @[dec.scala 120:19]
  wire  tlu_io_tlu_mem_ifu_ic_debug_rd_data_valid; // @[dec.scala 120:19]
  wire  tlu_io_tlu_mem_ifu_miss_state_idle; // @[dec.scala 120:19]
  wire  tlu_io_tlu_busbuff_lsu_pmu_bus_misaligned; // @[dec.scala 120:19]
  wire  tlu_io_tlu_busbuff_lsu_pmu_bus_error; // @[dec.scala 120:19]
  wire  tlu_io_tlu_busbuff_lsu_pmu_bus_busy; // @[dec.scala 120:19]
  wire  tlu_io_tlu_busbuff_dec_tlu_external_ldfwd_disable; // @[dec.scala 120:19]
  wire  tlu_io_tlu_busbuff_dec_tlu_wb_coalescing_disable; // @[dec.scala 120:19]
  wire  tlu_io_tlu_busbuff_dec_tlu_sideeffect_posted_disable; // @[dec.scala 120:19]
  wire  tlu_io_tlu_busbuff_lsu_imprecise_error_load_any; // @[dec.scala 120:19]
  wire  tlu_io_tlu_busbuff_lsu_imprecise_error_store_any; // @[dec.scala 120:19]
  wire [31:0] tlu_io_tlu_busbuff_lsu_imprecise_error_addr_any; // @[dec.scala 120:19]
  wire  tlu_io_lsu_tlu_lsu_pmu_load_external_m; // @[dec.scala 120:19]
  wire  tlu_io_lsu_tlu_lsu_pmu_store_external_m; // @[dec.scala 120:19]
  wire [7:0] tlu_io_dec_pic_pic_claimid; // @[dec.scala 120:19]
  wire [3:0] tlu_io_dec_pic_pic_pl; // @[dec.scala 120:19]
  wire  tlu_io_dec_pic_mhwakeup; // @[dec.scala 120:19]
  wire [3:0] tlu_io_dec_pic_dec_tlu_meicurpl; // @[dec.scala 120:19]
  wire [3:0] tlu_io_dec_pic_dec_tlu_meipt; // @[dec.scala 120:19]
  wire  tlu_io_dec_pic_mexintpend; // @[dec.scala 120:19]
  wire  dec_trigger_io_trigger_pkt_any_0_select; // @[dec.scala 121:27]
  wire  dec_trigger_io_trigger_pkt_any_0_match_pkt; // @[dec.scala 121:27]
  wire  dec_trigger_io_trigger_pkt_any_0_execute; // @[dec.scala 121:27]
  wire  dec_trigger_io_trigger_pkt_any_0_m; // @[dec.scala 121:27]
  wire [31:0] dec_trigger_io_trigger_pkt_any_0_tdata2; // @[dec.scala 121:27]
  wire  dec_trigger_io_trigger_pkt_any_1_select; // @[dec.scala 121:27]
  wire  dec_trigger_io_trigger_pkt_any_1_match_pkt; // @[dec.scala 121:27]
  wire  dec_trigger_io_trigger_pkt_any_1_execute; // @[dec.scala 121:27]
  wire  dec_trigger_io_trigger_pkt_any_1_m; // @[dec.scala 121:27]
  wire [31:0] dec_trigger_io_trigger_pkt_any_1_tdata2; // @[dec.scala 121:27]
  wire  dec_trigger_io_trigger_pkt_any_2_select; // @[dec.scala 121:27]
  wire  dec_trigger_io_trigger_pkt_any_2_match_pkt; // @[dec.scala 121:27]
  wire  dec_trigger_io_trigger_pkt_any_2_execute; // @[dec.scala 121:27]
  wire  dec_trigger_io_trigger_pkt_any_2_m; // @[dec.scala 121:27]
  wire [31:0] dec_trigger_io_trigger_pkt_any_2_tdata2; // @[dec.scala 121:27]
  wire  dec_trigger_io_trigger_pkt_any_3_select; // @[dec.scala 121:27]
  wire  dec_trigger_io_trigger_pkt_any_3_match_pkt; // @[dec.scala 121:27]
  wire  dec_trigger_io_trigger_pkt_any_3_execute; // @[dec.scala 121:27]
  wire  dec_trigger_io_trigger_pkt_any_3_m; // @[dec.scala 121:27]
  wire [31:0] dec_trigger_io_trigger_pkt_any_3_tdata2; // @[dec.scala 121:27]
  wire [30:0] dec_trigger_io_dec_i0_pc_d; // @[dec.scala 121:27]
  wire [3:0] dec_trigger_io_dec_i0_trigger_match_d; // @[dec.scala 121:27]
  wire  _T_1 = tlu_io_dec_tlu_i0_valid_wb1 | tlu_io_dec_tlu_i0_exc_valid_wb1; // @[dec.scala 296:98]
  dec_ib_ctl instbuff ( // @[dec.scala 117:24]
    .io_ifu_ib_ifu_i0_icaf(instbuff_io_ifu_ib_ifu_i0_icaf),
    .io_ifu_ib_ifu_i0_icaf_type(instbuff_io_ifu_ib_ifu_i0_icaf_type),
    .io_ifu_ib_ifu_i0_icaf_f1(instbuff_io_ifu_ib_ifu_i0_icaf_f1),
    .io_ifu_ib_ifu_i0_dbecc(instbuff_io_ifu_ib_ifu_i0_dbecc),
    .io_ifu_ib_ifu_i0_bp_index(instbuff_io_ifu_ib_ifu_i0_bp_index),
    .io_ifu_ib_ifu_i0_bp_fghr(instbuff_io_ifu_ib_ifu_i0_bp_fghr),
    .io_ifu_ib_ifu_i0_bp_btag(instbuff_io_ifu_ib_ifu_i0_bp_btag),
    .io_ifu_ib_ifu_i0_valid(instbuff_io_ifu_ib_ifu_i0_valid),
    .io_ifu_ib_ifu_i0_instr(instbuff_io_ifu_ib_ifu_i0_instr),
    .io_ifu_ib_ifu_i0_pc(instbuff_io_ifu_ib_ifu_i0_pc),
    .io_ifu_ib_ifu_i0_pc4(instbuff_io_ifu_ib_ifu_i0_pc4),
    .io_ifu_ib_i0_brp_valid(instbuff_io_ifu_ib_i0_brp_valid),
    .io_ifu_ib_i0_brp_bits_toffset(instbuff_io_ifu_ib_i0_brp_bits_toffset),
    .io_ifu_ib_i0_brp_bits_hist(instbuff_io_ifu_ib_i0_brp_bits_hist),
    .io_ifu_ib_i0_brp_bits_br_error(instbuff_io_ifu_ib_i0_brp_bits_br_error),
    .io_ifu_ib_i0_brp_bits_br_start_error(instbuff_io_ifu_ib_i0_brp_bits_br_start_error),
    .io_ifu_ib_i0_brp_bits_prett(instbuff_io_ifu_ib_i0_brp_bits_prett),
    .io_ifu_ib_i0_brp_bits_way(instbuff_io_ifu_ib_i0_brp_bits_way),
    .io_ifu_ib_i0_brp_bits_ret(instbuff_io_ifu_ib_i0_brp_bits_ret),
    .io_ib_exu_dec_i0_pc_d(instbuff_io_ib_exu_dec_i0_pc_d),
    .io_ib_exu_dec_debug_wdata_rs1_d(instbuff_io_ib_exu_dec_debug_wdata_rs1_d),
    .io_dbg_ib_dbg_cmd_valid(instbuff_io_dbg_ib_dbg_cmd_valid),
    .io_dbg_ib_dbg_cmd_write(instbuff_io_dbg_ib_dbg_cmd_write),
    .io_dbg_ib_dbg_cmd_type(instbuff_io_dbg_ib_dbg_cmd_type),
    .io_dbg_ib_dbg_cmd_addr(instbuff_io_dbg_ib_dbg_cmd_addr),
    .io_dec_ib0_valid_d(instbuff_io_dec_ib0_valid_d),
    .io_dec_i0_icaf_type_d(instbuff_io_dec_i0_icaf_type_d),
    .io_dec_i0_instr_d(instbuff_io_dec_i0_instr_d),
    .io_dec_i0_pc4_d(instbuff_io_dec_i0_pc4_d),
    .io_dec_i0_brp_valid(instbuff_io_dec_i0_brp_valid),
    .io_dec_i0_brp_bits_toffset(instbuff_io_dec_i0_brp_bits_toffset),
    .io_dec_i0_brp_bits_hist(instbuff_io_dec_i0_brp_bits_hist),
    .io_dec_i0_brp_bits_br_error(instbuff_io_dec_i0_brp_bits_br_error),
    .io_dec_i0_brp_bits_br_start_error(instbuff_io_dec_i0_brp_bits_br_start_error),
    .io_dec_i0_brp_bits_prett(instbuff_io_dec_i0_brp_bits_prett),
    .io_dec_i0_brp_bits_way(instbuff_io_dec_i0_brp_bits_way),
    .io_dec_i0_brp_bits_ret(instbuff_io_dec_i0_brp_bits_ret),
    .io_dec_i0_bp_index(instbuff_io_dec_i0_bp_index),
    .io_dec_i0_bp_fghr(instbuff_io_dec_i0_bp_fghr),
    .io_dec_i0_bp_btag(instbuff_io_dec_i0_bp_btag),
    .io_dec_i0_icaf_d(instbuff_io_dec_i0_icaf_d),
    .io_dec_i0_icaf_f1_d(instbuff_io_dec_i0_icaf_f1_d),
    .io_dec_i0_dbecc_d(instbuff_io_dec_i0_dbecc_d),
    .io_dec_debug_fence_d(instbuff_io_dec_debug_fence_d)
  );
  dec_decode_ctl decode ( // @[dec.scala 118:22]
    .clock(decode_clock),
    .reset(decode_reset),
    .io_decode_exu_dec_data_en(decode_io_decode_exu_dec_data_en),
    .io_decode_exu_dec_ctl_en(decode_io_decode_exu_dec_ctl_en),
    .io_decode_exu_i0_ap_land(decode_io_decode_exu_i0_ap_land),
    .io_decode_exu_i0_ap_lor(decode_io_decode_exu_i0_ap_lor),
    .io_decode_exu_i0_ap_lxor(decode_io_decode_exu_i0_ap_lxor),
    .io_decode_exu_i0_ap_sll(decode_io_decode_exu_i0_ap_sll),
    .io_decode_exu_i0_ap_srl(decode_io_decode_exu_i0_ap_srl),
    .io_decode_exu_i0_ap_sra(decode_io_decode_exu_i0_ap_sra),
    .io_decode_exu_i0_ap_beq(decode_io_decode_exu_i0_ap_beq),
    .io_decode_exu_i0_ap_bne(decode_io_decode_exu_i0_ap_bne),
    .io_decode_exu_i0_ap_blt(decode_io_decode_exu_i0_ap_blt),
    .io_decode_exu_i0_ap_bge(decode_io_decode_exu_i0_ap_bge),
    .io_decode_exu_i0_ap_add(decode_io_decode_exu_i0_ap_add),
    .io_decode_exu_i0_ap_sub(decode_io_decode_exu_i0_ap_sub),
    .io_decode_exu_i0_ap_slt(decode_io_decode_exu_i0_ap_slt),
    .io_decode_exu_i0_ap_unsign(decode_io_decode_exu_i0_ap_unsign),
    .io_decode_exu_i0_ap_jal(decode_io_decode_exu_i0_ap_jal),
    .io_decode_exu_i0_ap_predict_t(decode_io_decode_exu_i0_ap_predict_t),
    .io_decode_exu_i0_ap_predict_nt(decode_io_decode_exu_i0_ap_predict_nt),
    .io_decode_exu_i0_ap_csr_write(decode_io_decode_exu_i0_ap_csr_write),
    .io_decode_exu_i0_ap_csr_imm(decode_io_decode_exu_i0_ap_csr_imm),
    .io_decode_exu_dec_i0_predict_p_d_valid(decode_io_decode_exu_dec_i0_predict_p_d_valid),
    .io_decode_exu_dec_i0_predict_p_d_bits_pc4(decode_io_decode_exu_dec_i0_predict_p_d_bits_pc4),
    .io_decode_exu_dec_i0_predict_p_d_bits_hist(decode_io_decode_exu_dec_i0_predict_p_d_bits_hist),
    .io_decode_exu_dec_i0_predict_p_d_bits_toffset(decode_io_decode_exu_dec_i0_predict_p_d_bits_toffset),
    .io_decode_exu_dec_i0_predict_p_d_bits_br_error(decode_io_decode_exu_dec_i0_predict_p_d_bits_br_error),
    .io_decode_exu_dec_i0_predict_p_d_bits_br_start_error(decode_io_decode_exu_dec_i0_predict_p_d_bits_br_start_error),
    .io_decode_exu_dec_i0_predict_p_d_bits_prett(decode_io_decode_exu_dec_i0_predict_p_d_bits_prett),
    .io_decode_exu_dec_i0_predict_p_d_bits_pcall(decode_io_decode_exu_dec_i0_predict_p_d_bits_pcall),
    .io_decode_exu_dec_i0_predict_p_d_bits_pret(decode_io_decode_exu_dec_i0_predict_p_d_bits_pret),
    .io_decode_exu_dec_i0_predict_p_d_bits_pja(decode_io_decode_exu_dec_i0_predict_p_d_bits_pja),
    .io_decode_exu_dec_i0_predict_p_d_bits_way(decode_io_decode_exu_dec_i0_predict_p_d_bits_way),
    .io_decode_exu_i0_predict_fghr_d(decode_io_decode_exu_i0_predict_fghr_d),
    .io_decode_exu_i0_predict_index_d(decode_io_decode_exu_i0_predict_index_d),
    .io_decode_exu_i0_predict_btag_d(decode_io_decode_exu_i0_predict_btag_d),
    .io_decode_exu_dec_i0_rs1_en_d(decode_io_decode_exu_dec_i0_rs1_en_d),
    .io_decode_exu_dec_i0_rs2_en_d(decode_io_decode_exu_dec_i0_rs2_en_d),
    .io_decode_exu_dec_i0_immed_d(decode_io_decode_exu_dec_i0_immed_d),
    .io_decode_exu_dec_i0_rs1_bypass_data_d(decode_io_decode_exu_dec_i0_rs1_bypass_data_d),
    .io_decode_exu_dec_i0_rs2_bypass_data_d(decode_io_decode_exu_dec_i0_rs2_bypass_data_d),
    .io_decode_exu_dec_i0_select_pc_d(decode_io_decode_exu_dec_i0_select_pc_d),
    .io_decode_exu_dec_i0_rs1_bypass_en_d(decode_io_decode_exu_dec_i0_rs1_bypass_en_d),
    .io_decode_exu_dec_i0_rs2_bypass_en_d(decode_io_decode_exu_dec_i0_rs2_bypass_en_d),
    .io_decode_exu_mul_p_valid(decode_io_decode_exu_mul_p_valid),
    .io_decode_exu_mul_p_bits_rs1_sign(decode_io_decode_exu_mul_p_bits_rs1_sign),
    .io_decode_exu_mul_p_bits_rs2_sign(decode_io_decode_exu_mul_p_bits_rs2_sign),
    .io_decode_exu_mul_p_bits_low(decode_io_decode_exu_mul_p_bits_low),
    .io_decode_exu_pred_correct_npc_x(decode_io_decode_exu_pred_correct_npc_x),
    .io_decode_exu_dec_extint_stall(decode_io_decode_exu_dec_extint_stall),
    .io_decode_exu_exu_i0_result_x(decode_io_decode_exu_exu_i0_result_x),
    .io_decode_exu_exu_csr_rs1_x(decode_io_decode_exu_exu_csr_rs1_x),
    .io_dec_alu_dec_i0_alu_decode_d(decode_io_dec_alu_dec_i0_alu_decode_d),
    .io_dec_alu_dec_csr_ren_d(decode_io_dec_alu_dec_csr_ren_d),
    .io_dec_alu_dec_i0_br_immed_d(decode_io_dec_alu_dec_i0_br_immed_d),
    .io_dec_alu_exu_i0_pc_x(decode_io_dec_alu_exu_i0_pc_x),
    .io_dec_div_div_p_valid(decode_io_dec_div_div_p_valid),
    .io_dec_div_div_p_bits_unsign(decode_io_dec_div_div_p_bits_unsign),
    .io_dec_div_div_p_bits_rem(decode_io_dec_div_div_p_bits_rem),
    .io_dec_div_dec_div_cancel(decode_io_dec_div_dec_div_cancel),
    .io_dctl_busbuff_lsu_nonblock_load_valid_m(decode_io_dctl_busbuff_lsu_nonblock_load_valid_m),
    .io_dctl_busbuff_lsu_nonblock_load_tag_m(decode_io_dctl_busbuff_lsu_nonblock_load_tag_m),
    .io_dctl_busbuff_lsu_nonblock_load_inv_r(decode_io_dctl_busbuff_lsu_nonblock_load_inv_r),
    .io_dctl_busbuff_lsu_nonblock_load_inv_tag_r(decode_io_dctl_busbuff_lsu_nonblock_load_inv_tag_r),
    .io_dctl_busbuff_lsu_nonblock_load_data_valid(decode_io_dctl_busbuff_lsu_nonblock_load_data_valid),
    .io_dctl_busbuff_lsu_nonblock_load_data_error(decode_io_dctl_busbuff_lsu_nonblock_load_data_error),
    .io_dctl_busbuff_lsu_nonblock_load_data_tag(decode_io_dctl_busbuff_lsu_nonblock_load_data_tag),
    .io_dctl_busbuff_lsu_nonblock_load_data(decode_io_dctl_busbuff_lsu_nonblock_load_data),
    .io_dctl_dma_dma_dccm_stall_any(decode_io_dctl_dma_dma_dccm_stall_any),
    .io_dec_aln_dec_i0_decode_d(decode_io_dec_aln_dec_i0_decode_d),
    .io_dec_aln_ifu_i0_cinst(decode_io_dec_aln_ifu_i0_cinst),
    .io_dbg_dctl_dbg_cmd_wrdata(decode_io_dbg_dctl_dbg_cmd_wrdata),
    .io_dec_tlu_flush_extint(decode_io_dec_tlu_flush_extint),
    .io_dec_tlu_force_halt(decode_io_dec_tlu_force_halt),
    .io_dec_i0_inst_wb1(decode_io_dec_i0_inst_wb1),
    .io_dec_i0_pc_wb1(decode_io_dec_i0_pc_wb1),
    .io_dec_i0_trigger_match_d(decode_io_dec_i0_trigger_match_d),
    .io_dec_tlu_wr_pause_r(decode_io_dec_tlu_wr_pause_r),
    .io_dec_tlu_pipelining_disable(decode_io_dec_tlu_pipelining_disable),
    .io_lsu_trigger_match_m(decode_io_lsu_trigger_match_m),
    .io_lsu_pmu_misaligned_m(decode_io_lsu_pmu_misaligned_m),
    .io_dec_tlu_debug_stall(decode_io_dec_tlu_debug_stall),
    .io_dec_tlu_flush_leak_one_r(decode_io_dec_tlu_flush_leak_one_r),
    .io_dec_debug_fence_d(decode_io_dec_debug_fence_d),
    .io_dec_i0_icaf_d(decode_io_dec_i0_icaf_d),
    .io_dec_i0_icaf_f1_d(decode_io_dec_i0_icaf_f1_d),
    .io_dec_i0_icaf_type_d(decode_io_dec_i0_icaf_type_d),
    .io_dec_i0_dbecc_d(decode_io_dec_i0_dbecc_d),
    .io_dec_i0_brp_valid(decode_io_dec_i0_brp_valid),
    .io_dec_i0_brp_bits_toffset(decode_io_dec_i0_brp_bits_toffset),
    .io_dec_i0_brp_bits_hist(decode_io_dec_i0_brp_bits_hist),
    .io_dec_i0_brp_bits_br_error(decode_io_dec_i0_brp_bits_br_error),
    .io_dec_i0_brp_bits_br_start_error(decode_io_dec_i0_brp_bits_br_start_error),
    .io_dec_i0_brp_bits_prett(decode_io_dec_i0_brp_bits_prett),
    .io_dec_i0_brp_bits_way(decode_io_dec_i0_brp_bits_way),
    .io_dec_i0_brp_bits_ret(decode_io_dec_i0_brp_bits_ret),
    .io_dec_i0_bp_index(decode_io_dec_i0_bp_index),
    .io_dec_i0_bp_fghr(decode_io_dec_i0_bp_fghr),
    .io_dec_i0_bp_btag(decode_io_dec_i0_bp_btag),
    .io_lsu_idle_any(decode_io_lsu_idle_any),
    .io_lsu_load_stall_any(decode_io_lsu_load_stall_any),
    .io_lsu_store_stall_any(decode_io_lsu_store_stall_any),
    .io_exu_div_wren(decode_io_exu_div_wren),
    .io_dec_tlu_i0_kill_writeb_wb(decode_io_dec_tlu_i0_kill_writeb_wb),
    .io_dec_tlu_flush_lower_wb(decode_io_dec_tlu_flush_lower_wb),
    .io_dec_tlu_i0_kill_writeb_r(decode_io_dec_tlu_i0_kill_writeb_r),
    .io_dec_tlu_flush_lower_r(decode_io_dec_tlu_flush_lower_r),
    .io_dec_tlu_flush_pause_r(decode_io_dec_tlu_flush_pause_r),
    .io_dec_tlu_presync_d(decode_io_dec_tlu_presync_d),
    .io_dec_tlu_postsync_d(decode_io_dec_tlu_postsync_d),
    .io_dec_i0_pc4_d(decode_io_dec_i0_pc4_d),
    .io_dec_csr_rddata_d(decode_io_dec_csr_rddata_d),
    .io_dec_csr_legal_d(decode_io_dec_csr_legal_d),
    .io_lsu_result_m(decode_io_lsu_result_m),
    .io_lsu_result_corr_r(decode_io_lsu_result_corr_r),
    .io_exu_flush_final(decode_io_exu_flush_final),
    .io_dec_i0_instr_d(decode_io_dec_i0_instr_d),
    .io_dec_ib0_valid_d(decode_io_dec_ib0_valid_d),
    .io_free_clk(decode_io_free_clk),
    .io_active_clk(decode_io_active_clk),
    .io_clk_override(decode_io_clk_override),
    .io_dec_i0_rs1_d(decode_io_dec_i0_rs1_d),
    .io_dec_i0_rs2_d(decode_io_dec_i0_rs2_d),
    .io_dec_i0_waddr_r(decode_io_dec_i0_waddr_r),
    .io_dec_i0_wen_r(decode_io_dec_i0_wen_r),
    .io_dec_i0_wdata_r(decode_io_dec_i0_wdata_r),
    .io_lsu_p_valid(decode_io_lsu_p_valid),
    .io_lsu_p_bits_fast_int(decode_io_lsu_p_bits_fast_int),
    .io_lsu_p_bits_by(decode_io_lsu_p_bits_by),
    .io_lsu_p_bits_half(decode_io_lsu_p_bits_half),
    .io_lsu_p_bits_word(decode_io_lsu_p_bits_word),
    .io_lsu_p_bits_load(decode_io_lsu_p_bits_load),
    .io_lsu_p_bits_store(decode_io_lsu_p_bits_store),
    .io_lsu_p_bits_unsign(decode_io_lsu_p_bits_unsign),
    .io_lsu_p_bits_store_data_bypass_d(decode_io_lsu_p_bits_store_data_bypass_d),
    .io_lsu_p_bits_load_ldst_bypass_d(decode_io_lsu_p_bits_load_ldst_bypass_d),
    .io_div_waddr_wb(decode_io_div_waddr_wb),
    .io_dec_lsu_valid_raw_d(decode_io_dec_lsu_valid_raw_d),
    .io_dec_lsu_offset_d(decode_io_dec_lsu_offset_d),
    .io_dec_csr_wen_unq_d(decode_io_dec_csr_wen_unq_d),
    .io_dec_csr_any_unq_d(decode_io_dec_csr_any_unq_d),
    .io_dec_csr_rdaddr_d(decode_io_dec_csr_rdaddr_d),
    .io_dec_csr_wen_r(decode_io_dec_csr_wen_r),
    .io_dec_csr_wraddr_r(decode_io_dec_csr_wraddr_r),
    .io_dec_csr_wrdata_r(decode_io_dec_csr_wrdata_r),
    .io_dec_csr_stall_int_ff(decode_io_dec_csr_stall_int_ff),
    .io_dec_tlu_i0_valid_r(decode_io_dec_tlu_i0_valid_r),
    .io_dec_tlu_packet_r_legal(decode_io_dec_tlu_packet_r_legal),
    .io_dec_tlu_packet_r_icaf(decode_io_dec_tlu_packet_r_icaf),
    .io_dec_tlu_packet_r_icaf_f1(decode_io_dec_tlu_packet_r_icaf_f1),
    .io_dec_tlu_packet_r_icaf_type(decode_io_dec_tlu_packet_r_icaf_type),
    .io_dec_tlu_packet_r_fence_i(decode_io_dec_tlu_packet_r_fence_i),
    .io_dec_tlu_packet_r_i0trigger(decode_io_dec_tlu_packet_r_i0trigger),
    .io_dec_tlu_packet_r_pmu_i0_itype(decode_io_dec_tlu_packet_r_pmu_i0_itype),
    .io_dec_tlu_packet_r_pmu_i0_br_unpred(decode_io_dec_tlu_packet_r_pmu_i0_br_unpred),
    .io_dec_tlu_packet_r_pmu_divide(decode_io_dec_tlu_packet_r_pmu_divide),
    .io_dec_tlu_packet_r_pmu_lsu_misaligned(decode_io_dec_tlu_packet_r_pmu_lsu_misaligned),
    .io_dec_tlu_i0_pc_r(decode_io_dec_tlu_i0_pc_r),
    .io_dec_illegal_inst(decode_io_dec_illegal_inst),
    .io_dec_pmu_instr_decoded(decode_io_dec_pmu_instr_decoded),
    .io_dec_pmu_decode_stall(decode_io_dec_pmu_decode_stall),
    .io_dec_pmu_presync_stall(decode_io_dec_pmu_presync_stall),
    .io_dec_pmu_postsync_stall(decode_io_dec_pmu_postsync_stall),
    .io_dec_nonblock_load_wen(decode_io_dec_nonblock_load_wen),
    .io_dec_nonblock_load_waddr(decode_io_dec_nonblock_load_waddr),
    .io_dec_pause_state(decode_io_dec_pause_state),
    .io_dec_pause_state_cg(decode_io_dec_pause_state_cg),
    .io_dec_div_active(decode_io_dec_div_active),
    .io_scan_mode(decode_io_scan_mode)
  );
  dec_gpr_ctl gpr ( // @[dec.scala 119:19]
    .clock(gpr_clock),
    .reset(gpr_reset),
    .io_raddr0(gpr_io_raddr0),
    .io_raddr1(gpr_io_raddr1),
    .io_wen0(gpr_io_wen0),
    .io_waddr0(gpr_io_waddr0),
    .io_wd0(gpr_io_wd0),
    .io_wen1(gpr_io_wen1),
    .io_waddr1(gpr_io_waddr1),
    .io_wd1(gpr_io_wd1),
    .io_wen2(gpr_io_wen2),
    .io_waddr2(gpr_io_waddr2),
    .io_wd2(gpr_io_wd2),
    .io_scan_mode(gpr_io_scan_mode),
    .io_gpr_exu_gpr_i0_rs1_d(gpr_io_gpr_exu_gpr_i0_rs1_d),
    .io_gpr_exu_gpr_i0_rs2_d(gpr_io_gpr_exu_gpr_i0_rs2_d)
  );
  dec_tlu_ctl tlu ( // @[dec.scala 120:19]
    .clock(tlu_clock),
    .reset(tlu_reset),
    .io_tlu_exu_dec_tlu_meihap(tlu_io_tlu_exu_dec_tlu_meihap),
    .io_tlu_exu_dec_tlu_flush_lower_r(tlu_io_tlu_exu_dec_tlu_flush_lower_r),
    .io_tlu_exu_dec_tlu_flush_path_r(tlu_io_tlu_exu_dec_tlu_flush_path_r),
    .io_tlu_exu_exu_i0_br_hist_r(tlu_io_tlu_exu_exu_i0_br_hist_r),
    .io_tlu_exu_exu_i0_br_error_r(tlu_io_tlu_exu_exu_i0_br_error_r),
    .io_tlu_exu_exu_i0_br_start_error_r(tlu_io_tlu_exu_exu_i0_br_start_error_r),
    .io_tlu_exu_exu_i0_br_valid_r(tlu_io_tlu_exu_exu_i0_br_valid_r),
    .io_tlu_exu_exu_i0_br_mp_r(tlu_io_tlu_exu_exu_i0_br_mp_r),
    .io_tlu_exu_exu_i0_br_middle_r(tlu_io_tlu_exu_exu_i0_br_middle_r),
    .io_tlu_exu_exu_pmu_i0_br_misp(tlu_io_tlu_exu_exu_pmu_i0_br_misp),
    .io_tlu_exu_exu_pmu_i0_br_ataken(tlu_io_tlu_exu_exu_pmu_i0_br_ataken),
    .io_tlu_exu_exu_pmu_i0_pc4(tlu_io_tlu_exu_exu_pmu_i0_pc4),
    .io_tlu_exu_exu_npc_r(tlu_io_tlu_exu_exu_npc_r),
    .io_tlu_dma_dma_pmu_dccm_read(tlu_io_tlu_dma_dma_pmu_dccm_read),
    .io_tlu_dma_dma_pmu_dccm_write(tlu_io_tlu_dma_dma_pmu_dccm_write),
    .io_tlu_dma_dma_pmu_any_read(tlu_io_tlu_dma_dma_pmu_any_read),
    .io_tlu_dma_dma_pmu_any_write(tlu_io_tlu_dma_dma_pmu_any_write),
    .io_tlu_dma_dec_tlu_dma_qos_prty(tlu_io_tlu_dma_dec_tlu_dma_qos_prty),
    .io_tlu_dma_dma_dccm_stall_any(tlu_io_tlu_dma_dma_dccm_stall_any),
    .io_tlu_dma_dma_iccm_stall_any(tlu_io_tlu_dma_dma_iccm_stall_any),
    .io_active_clk(tlu_io_active_clk),
    .io_free_clk(tlu_io_free_clk),
    .io_scan_mode(tlu_io_scan_mode),
    .io_rst_vec(tlu_io_rst_vec),
    .io_nmi_int(tlu_io_nmi_int),
    .io_nmi_vec(tlu_io_nmi_vec),
    .io_i_cpu_halt_req(tlu_io_i_cpu_halt_req),
    .io_i_cpu_run_req(tlu_io_i_cpu_run_req),
    .io_lsu_fastint_stall_any(tlu_io_lsu_fastint_stall_any),
    .io_lsu_idle_any(tlu_io_lsu_idle_any),
    .io_dec_pmu_instr_decoded(tlu_io_dec_pmu_instr_decoded),
    .io_dec_pmu_decode_stall(tlu_io_dec_pmu_decode_stall),
    .io_dec_pmu_presync_stall(tlu_io_dec_pmu_presync_stall),
    .io_dec_pmu_postsync_stall(tlu_io_dec_pmu_postsync_stall),
    .io_lsu_store_stall_any(tlu_io_lsu_store_stall_any),
    .io_lsu_fir_addr(tlu_io_lsu_fir_addr),
    .io_lsu_fir_error(tlu_io_lsu_fir_error),
    .io_iccm_dma_sb_error(tlu_io_iccm_dma_sb_error),
    .io_lsu_error_pkt_r_valid(tlu_io_lsu_error_pkt_r_valid),
    .io_lsu_error_pkt_r_bits_single_ecc_error(tlu_io_lsu_error_pkt_r_bits_single_ecc_error),
    .io_lsu_error_pkt_r_bits_inst_type(tlu_io_lsu_error_pkt_r_bits_inst_type),
    .io_lsu_error_pkt_r_bits_exc_type(tlu_io_lsu_error_pkt_r_bits_exc_type),
    .io_lsu_error_pkt_r_bits_mscause(tlu_io_lsu_error_pkt_r_bits_mscause),
    .io_lsu_error_pkt_r_bits_addr(tlu_io_lsu_error_pkt_r_bits_addr),
    .io_lsu_single_ecc_error_incr(tlu_io_lsu_single_ecc_error_incr),
    .io_dec_pause_state(tlu_io_dec_pause_state),
    .io_dec_csr_wen_unq_d(tlu_io_dec_csr_wen_unq_d),
    .io_dec_csr_any_unq_d(tlu_io_dec_csr_any_unq_d),
    .io_dec_csr_rdaddr_d(tlu_io_dec_csr_rdaddr_d),
    .io_dec_csr_wen_r(tlu_io_dec_csr_wen_r),
    .io_dec_csr_wraddr_r(tlu_io_dec_csr_wraddr_r),
    .io_dec_csr_wrdata_r(tlu_io_dec_csr_wrdata_r),
    .io_dec_csr_stall_int_ff(tlu_io_dec_csr_stall_int_ff),
    .io_dec_tlu_i0_valid_r(tlu_io_dec_tlu_i0_valid_r),
    .io_dec_tlu_i0_pc_r(tlu_io_dec_tlu_i0_pc_r),
    .io_dec_tlu_packet_r_legal(tlu_io_dec_tlu_packet_r_legal),
    .io_dec_tlu_packet_r_icaf(tlu_io_dec_tlu_packet_r_icaf),
    .io_dec_tlu_packet_r_icaf_f1(tlu_io_dec_tlu_packet_r_icaf_f1),
    .io_dec_tlu_packet_r_icaf_type(tlu_io_dec_tlu_packet_r_icaf_type),
    .io_dec_tlu_packet_r_fence_i(tlu_io_dec_tlu_packet_r_fence_i),
    .io_dec_tlu_packet_r_i0trigger(tlu_io_dec_tlu_packet_r_i0trigger),
    .io_dec_tlu_packet_r_pmu_i0_itype(tlu_io_dec_tlu_packet_r_pmu_i0_itype),
    .io_dec_tlu_packet_r_pmu_i0_br_unpred(tlu_io_dec_tlu_packet_r_pmu_i0_br_unpred),
    .io_dec_tlu_packet_r_pmu_divide(tlu_io_dec_tlu_packet_r_pmu_divide),
    .io_dec_tlu_packet_r_pmu_lsu_misaligned(tlu_io_dec_tlu_packet_r_pmu_lsu_misaligned),
    .io_dec_illegal_inst(tlu_io_dec_illegal_inst),
    .io_dec_i0_decode_d(tlu_io_dec_i0_decode_d),
    .io_exu_i0_br_way_r(tlu_io_exu_i0_br_way_r),
    .io_dec_dbg_cmd_done(tlu_io_dec_dbg_cmd_done),
    .io_dec_dbg_cmd_fail(tlu_io_dec_dbg_cmd_fail),
    .io_dec_tlu_dbg_halted(tlu_io_dec_tlu_dbg_halted),
    .io_dec_tlu_debug_mode(tlu_io_dec_tlu_debug_mode),
    .io_dec_tlu_resume_ack(tlu_io_dec_tlu_resume_ack),
    .io_dec_tlu_debug_stall(tlu_io_dec_tlu_debug_stall),
    .io_dec_tlu_mpc_halted_only(tlu_io_dec_tlu_mpc_halted_only),
    .io_dec_tlu_flush_extint(tlu_io_dec_tlu_flush_extint),
    .io_dbg_halt_req(tlu_io_dbg_halt_req),
    .io_dbg_resume_req(tlu_io_dbg_resume_req),
    .io_dec_div_active(tlu_io_dec_div_active),
    .io_trigger_pkt_any_0_select(tlu_io_trigger_pkt_any_0_select),
    .io_trigger_pkt_any_0_match_pkt(tlu_io_trigger_pkt_any_0_match_pkt),
    .io_trigger_pkt_any_0_store(tlu_io_trigger_pkt_any_0_store),
    .io_trigger_pkt_any_0_load(tlu_io_trigger_pkt_any_0_load),
    .io_trigger_pkt_any_0_execute(tlu_io_trigger_pkt_any_0_execute),
    .io_trigger_pkt_any_0_m(tlu_io_trigger_pkt_any_0_m),
    .io_trigger_pkt_any_0_tdata2(tlu_io_trigger_pkt_any_0_tdata2),
    .io_trigger_pkt_any_1_select(tlu_io_trigger_pkt_any_1_select),
    .io_trigger_pkt_any_1_match_pkt(tlu_io_trigger_pkt_any_1_match_pkt),
    .io_trigger_pkt_any_1_store(tlu_io_trigger_pkt_any_1_store),
    .io_trigger_pkt_any_1_load(tlu_io_trigger_pkt_any_1_load),
    .io_trigger_pkt_any_1_execute(tlu_io_trigger_pkt_any_1_execute),
    .io_trigger_pkt_any_1_m(tlu_io_trigger_pkt_any_1_m),
    .io_trigger_pkt_any_1_tdata2(tlu_io_trigger_pkt_any_1_tdata2),
    .io_trigger_pkt_any_2_select(tlu_io_trigger_pkt_any_2_select),
    .io_trigger_pkt_any_2_match_pkt(tlu_io_trigger_pkt_any_2_match_pkt),
    .io_trigger_pkt_any_2_store(tlu_io_trigger_pkt_any_2_store),
    .io_trigger_pkt_any_2_load(tlu_io_trigger_pkt_any_2_load),
    .io_trigger_pkt_any_2_execute(tlu_io_trigger_pkt_any_2_execute),
    .io_trigger_pkt_any_2_m(tlu_io_trigger_pkt_any_2_m),
    .io_trigger_pkt_any_2_tdata2(tlu_io_trigger_pkt_any_2_tdata2),
    .io_trigger_pkt_any_3_select(tlu_io_trigger_pkt_any_3_select),
    .io_trigger_pkt_any_3_match_pkt(tlu_io_trigger_pkt_any_3_match_pkt),
    .io_trigger_pkt_any_3_store(tlu_io_trigger_pkt_any_3_store),
    .io_trigger_pkt_any_3_load(tlu_io_trigger_pkt_any_3_load),
    .io_trigger_pkt_any_3_execute(tlu_io_trigger_pkt_any_3_execute),
    .io_trigger_pkt_any_3_m(tlu_io_trigger_pkt_any_3_m),
    .io_trigger_pkt_any_3_tdata2(tlu_io_trigger_pkt_any_3_tdata2),
    .io_timer_int(tlu_io_timer_int),
    .io_soft_int(tlu_io_soft_int),
    .io_o_cpu_halt_status(tlu_io_o_cpu_halt_status),
    .io_o_cpu_halt_ack(tlu_io_o_cpu_halt_ack),
    .io_o_cpu_run_ack(tlu_io_o_cpu_run_ack),
    .io_o_debug_mode_status(tlu_io_o_debug_mode_status),
    .io_core_id(tlu_io_core_id),
    .io_mpc_debug_halt_req(tlu_io_mpc_debug_halt_req),
    .io_mpc_debug_run_req(tlu_io_mpc_debug_run_req),
    .io_mpc_reset_run_req(tlu_io_mpc_reset_run_req),
    .io_mpc_debug_halt_ack(tlu_io_mpc_debug_halt_ack),
    .io_mpc_debug_run_ack(tlu_io_mpc_debug_run_ack),
    .io_debug_brkpt_status(tlu_io_debug_brkpt_status),
    .io_dec_csr_rddata_d(tlu_io_dec_csr_rddata_d),
    .io_dec_csr_legal_d(tlu_io_dec_csr_legal_d),
    .io_dec_tlu_i0_kill_writeb_wb(tlu_io_dec_tlu_i0_kill_writeb_wb),
    .io_dec_tlu_i0_kill_writeb_r(tlu_io_dec_tlu_i0_kill_writeb_r),
    .io_dec_tlu_wr_pause_r(tlu_io_dec_tlu_wr_pause_r),
    .io_dec_tlu_flush_pause_r(tlu_io_dec_tlu_flush_pause_r),
    .io_dec_tlu_presync_d(tlu_io_dec_tlu_presync_d),
    .io_dec_tlu_postsync_d(tlu_io_dec_tlu_postsync_d),
    .io_dec_tlu_perfcnt0(tlu_io_dec_tlu_perfcnt0),
    .io_dec_tlu_perfcnt1(tlu_io_dec_tlu_perfcnt1),
    .io_dec_tlu_perfcnt2(tlu_io_dec_tlu_perfcnt2),
    .io_dec_tlu_perfcnt3(tlu_io_dec_tlu_perfcnt3),
    .io_dec_tlu_i0_exc_valid_wb1(tlu_io_dec_tlu_i0_exc_valid_wb1),
    .io_dec_tlu_i0_valid_wb1(tlu_io_dec_tlu_i0_valid_wb1),
    .io_dec_tlu_int_valid_wb1(tlu_io_dec_tlu_int_valid_wb1),
    .io_dec_tlu_exc_cause_wb1(tlu_io_dec_tlu_exc_cause_wb1),
    .io_dec_tlu_mtval_wb1(tlu_io_dec_tlu_mtval_wb1),
    .io_dec_tlu_pipelining_disable(tlu_io_dec_tlu_pipelining_disable),
    .io_dec_tlu_misc_clk_override(tlu_io_dec_tlu_misc_clk_override),
    .io_dec_tlu_dec_clk_override(tlu_io_dec_tlu_dec_clk_override),
    .io_dec_tlu_lsu_clk_override(tlu_io_dec_tlu_lsu_clk_override),
    .io_dec_tlu_bus_clk_override(tlu_io_dec_tlu_bus_clk_override),
    .io_dec_tlu_pic_clk_override(tlu_io_dec_tlu_pic_clk_override),
    .io_dec_tlu_dccm_clk_override(tlu_io_dec_tlu_dccm_clk_override),
    .io_dec_tlu_icm_clk_override(tlu_io_dec_tlu_icm_clk_override),
    .io_dec_tlu_flush_lower_wb(tlu_io_dec_tlu_flush_lower_wb),
    .io_ifu_pmu_instr_aligned(tlu_io_ifu_pmu_instr_aligned),
    .io_tlu_bp_dec_tlu_br0_r_pkt_valid(tlu_io_tlu_bp_dec_tlu_br0_r_pkt_valid),
    .io_tlu_bp_dec_tlu_br0_r_pkt_bits_hist(tlu_io_tlu_bp_dec_tlu_br0_r_pkt_bits_hist),
    .io_tlu_bp_dec_tlu_br0_r_pkt_bits_br_error(tlu_io_tlu_bp_dec_tlu_br0_r_pkt_bits_br_error),
    .io_tlu_bp_dec_tlu_br0_r_pkt_bits_br_start_error(tlu_io_tlu_bp_dec_tlu_br0_r_pkt_bits_br_start_error),
    .io_tlu_bp_dec_tlu_br0_r_pkt_bits_way(tlu_io_tlu_bp_dec_tlu_br0_r_pkt_bits_way),
    .io_tlu_bp_dec_tlu_br0_r_pkt_bits_middle(tlu_io_tlu_bp_dec_tlu_br0_r_pkt_bits_middle),
    .io_tlu_bp_dec_tlu_flush_leak_one_wb(tlu_io_tlu_bp_dec_tlu_flush_leak_one_wb),
    .io_tlu_bp_dec_tlu_bpred_disable(tlu_io_tlu_bp_dec_tlu_bpred_disable),
    .io_tlu_ifc_dec_tlu_flush_noredir_wb(tlu_io_tlu_ifc_dec_tlu_flush_noredir_wb),
    .io_tlu_ifc_dec_tlu_mrac_ff(tlu_io_tlu_ifc_dec_tlu_mrac_ff),
    .io_tlu_ifc_ifu_pmu_fetch_stall(tlu_io_tlu_ifc_ifu_pmu_fetch_stall),
    .io_tlu_mem_dec_tlu_flush_err_wb(tlu_io_tlu_mem_dec_tlu_flush_err_wb),
    .io_tlu_mem_dec_tlu_i0_commit_cmt(tlu_io_tlu_mem_dec_tlu_i0_commit_cmt),
    .io_tlu_mem_dec_tlu_force_halt(tlu_io_tlu_mem_dec_tlu_force_halt),
    .io_tlu_mem_dec_tlu_fence_i_wb(tlu_io_tlu_mem_dec_tlu_fence_i_wb),
    .io_tlu_mem_dec_tlu_ic_diag_pkt_icache_wrdata(tlu_io_tlu_mem_dec_tlu_ic_diag_pkt_icache_wrdata),
    .io_tlu_mem_dec_tlu_ic_diag_pkt_icache_dicawics(tlu_io_tlu_mem_dec_tlu_ic_diag_pkt_icache_dicawics),
    .io_tlu_mem_dec_tlu_ic_diag_pkt_icache_rd_valid(tlu_io_tlu_mem_dec_tlu_ic_diag_pkt_icache_rd_valid),
    .io_tlu_mem_dec_tlu_ic_diag_pkt_icache_wr_valid(tlu_io_tlu_mem_dec_tlu_ic_diag_pkt_icache_wr_valid),
    .io_tlu_mem_dec_tlu_core_ecc_disable(tlu_io_tlu_mem_dec_tlu_core_ecc_disable),
    .io_tlu_mem_ifu_pmu_ic_miss(tlu_io_tlu_mem_ifu_pmu_ic_miss),
    .io_tlu_mem_ifu_pmu_ic_hit(tlu_io_tlu_mem_ifu_pmu_ic_hit),
    .io_tlu_mem_ifu_pmu_bus_error(tlu_io_tlu_mem_ifu_pmu_bus_error),
    .io_tlu_mem_ifu_pmu_bus_busy(tlu_io_tlu_mem_ifu_pmu_bus_busy),
    .io_tlu_mem_ifu_ic_error_start(tlu_io_tlu_mem_ifu_ic_error_start),
    .io_tlu_mem_ifu_iccm_rd_ecc_single_err(tlu_io_tlu_mem_ifu_iccm_rd_ecc_single_err),
    .io_tlu_mem_ifu_ic_debug_rd_data(tlu_io_tlu_mem_ifu_ic_debug_rd_data),
    .io_tlu_mem_ifu_ic_debug_rd_data_valid(tlu_io_tlu_mem_ifu_ic_debug_rd_data_valid),
    .io_tlu_mem_ifu_miss_state_idle(tlu_io_tlu_mem_ifu_miss_state_idle),
    .io_tlu_busbuff_lsu_pmu_bus_misaligned(tlu_io_tlu_busbuff_lsu_pmu_bus_misaligned),
    .io_tlu_busbuff_lsu_pmu_bus_error(tlu_io_tlu_busbuff_lsu_pmu_bus_error),
    .io_tlu_busbuff_lsu_pmu_bus_busy(tlu_io_tlu_busbuff_lsu_pmu_bus_busy),
    .io_tlu_busbuff_dec_tlu_external_ldfwd_disable(tlu_io_tlu_busbuff_dec_tlu_external_ldfwd_disable),
    .io_tlu_busbuff_dec_tlu_wb_coalescing_disable(tlu_io_tlu_busbuff_dec_tlu_wb_coalescing_disable),
    .io_tlu_busbuff_dec_tlu_sideeffect_posted_disable(tlu_io_tlu_busbuff_dec_tlu_sideeffect_posted_disable),
    .io_tlu_busbuff_lsu_imprecise_error_load_any(tlu_io_tlu_busbuff_lsu_imprecise_error_load_any),
    .io_tlu_busbuff_lsu_imprecise_error_store_any(tlu_io_tlu_busbuff_lsu_imprecise_error_store_any),
    .io_tlu_busbuff_lsu_imprecise_error_addr_any(tlu_io_tlu_busbuff_lsu_imprecise_error_addr_any),
    .io_lsu_tlu_lsu_pmu_load_external_m(tlu_io_lsu_tlu_lsu_pmu_load_external_m),
    .io_lsu_tlu_lsu_pmu_store_external_m(tlu_io_lsu_tlu_lsu_pmu_store_external_m),
    .io_dec_pic_pic_claimid(tlu_io_dec_pic_pic_claimid),
    .io_dec_pic_pic_pl(tlu_io_dec_pic_pic_pl),
    .io_dec_pic_mhwakeup(tlu_io_dec_pic_mhwakeup),
    .io_dec_pic_dec_tlu_meicurpl(tlu_io_dec_pic_dec_tlu_meicurpl),
    .io_dec_pic_dec_tlu_meipt(tlu_io_dec_pic_dec_tlu_meipt),
    .io_dec_pic_mexintpend(tlu_io_dec_pic_mexintpend)
  );
  dec_trigger dec_trigger ( // @[dec.scala 121:27]
    .io_trigger_pkt_any_0_select(dec_trigger_io_trigger_pkt_any_0_select),
    .io_trigger_pkt_any_0_match_pkt(dec_trigger_io_trigger_pkt_any_0_match_pkt),
    .io_trigger_pkt_any_0_execute(dec_trigger_io_trigger_pkt_any_0_execute),
    .io_trigger_pkt_any_0_m(dec_trigger_io_trigger_pkt_any_0_m),
    .io_trigger_pkt_any_0_tdata2(dec_trigger_io_trigger_pkt_any_0_tdata2),
    .io_trigger_pkt_any_1_select(dec_trigger_io_trigger_pkt_any_1_select),
    .io_trigger_pkt_any_1_match_pkt(dec_trigger_io_trigger_pkt_any_1_match_pkt),
    .io_trigger_pkt_any_1_execute(dec_trigger_io_trigger_pkt_any_1_execute),
    .io_trigger_pkt_any_1_m(dec_trigger_io_trigger_pkt_any_1_m),
    .io_trigger_pkt_any_1_tdata2(dec_trigger_io_trigger_pkt_any_1_tdata2),
    .io_trigger_pkt_any_2_select(dec_trigger_io_trigger_pkt_any_2_select),
    .io_trigger_pkt_any_2_match_pkt(dec_trigger_io_trigger_pkt_any_2_match_pkt),
    .io_trigger_pkt_any_2_execute(dec_trigger_io_trigger_pkt_any_2_execute),
    .io_trigger_pkt_any_2_m(dec_trigger_io_trigger_pkt_any_2_m),
    .io_trigger_pkt_any_2_tdata2(dec_trigger_io_trigger_pkt_any_2_tdata2),
    .io_trigger_pkt_any_3_select(dec_trigger_io_trigger_pkt_any_3_select),
    .io_trigger_pkt_any_3_match_pkt(dec_trigger_io_trigger_pkt_any_3_match_pkt),
    .io_trigger_pkt_any_3_execute(dec_trigger_io_trigger_pkt_any_3_execute),
    .io_trigger_pkt_any_3_m(dec_trigger_io_trigger_pkt_any_3_m),
    .io_trigger_pkt_any_3_tdata2(dec_trigger_io_trigger_pkt_any_3_tdata2),
    .io_dec_i0_pc_d(dec_trigger_io_dec_i0_pc_d),
    .io_dec_i0_trigger_match_d(dec_trigger_io_dec_i0_trigger_match_d)
  );
  assign io_dec_pause_state_cg = decode_io_dec_pause_state_cg; // @[dec.scala 188:40]
  assign io_o_cpu_halt_status = tlu_io_o_cpu_halt_status; // @[dec.scala 265:29]
  assign io_o_cpu_halt_ack = tlu_io_o_cpu_halt_ack; // @[dec.scala 266:29]
  assign io_o_cpu_run_ack = tlu_io_o_cpu_run_ack; // @[dec.scala 267:29]
  assign io_o_debug_mode_status = tlu_io_o_debug_mode_status; // @[dec.scala 268:29]
  assign io_mpc_debug_halt_ack = tlu_io_mpc_debug_halt_ack; // @[dec.scala 269:29]
  assign io_mpc_debug_run_ack = tlu_io_mpc_debug_run_ack; // @[dec.scala 270:29]
  assign io_debug_brkpt_status = tlu_io_debug_brkpt_status; // @[dec.scala 271:29]
  assign io_dec_tlu_dbg_halted = tlu_io_dec_tlu_dbg_halted; // @[dec.scala 260:28]
  assign io_dec_tlu_debug_mode = tlu_io_dec_tlu_debug_mode; // @[dec.scala 261:28]
  assign io_dec_tlu_resume_ack = tlu_io_dec_tlu_resume_ack; // @[dec.scala 262:28]
  assign io_dec_tlu_mpc_halted_only = tlu_io_dec_tlu_mpc_halted_only; // @[dec.scala 263:51]
  assign io_dec_dbg_rddata = decode_io_dec_i0_wdata_r; // @[dec.scala 304:21]
  assign io_dec_dbg_cmd_done = tlu_io_dec_dbg_cmd_done; // @[dec.scala 258:28]
  assign io_dec_dbg_cmd_fail = tlu_io_dec_dbg_cmd_fail; // @[dec.scala 259:28]
  assign io_trigger_pkt_any_0_select = tlu_io_trigger_pkt_any_0_select; // @[dec.scala 264:29]
  assign io_trigger_pkt_any_0_match_pkt = tlu_io_trigger_pkt_any_0_match_pkt; // @[dec.scala 264:29]
  assign io_trigger_pkt_any_0_store = tlu_io_trigger_pkt_any_0_store; // @[dec.scala 264:29]
  assign io_trigger_pkt_any_0_load = tlu_io_trigger_pkt_any_0_load; // @[dec.scala 264:29]
  assign io_trigger_pkt_any_0_tdata2 = tlu_io_trigger_pkt_any_0_tdata2; // @[dec.scala 264:29]
  assign io_trigger_pkt_any_1_select = tlu_io_trigger_pkt_any_1_select; // @[dec.scala 264:29]
  assign io_trigger_pkt_any_1_match_pkt = tlu_io_trigger_pkt_any_1_match_pkt; // @[dec.scala 264:29]
  assign io_trigger_pkt_any_1_store = tlu_io_trigger_pkt_any_1_store; // @[dec.scala 264:29]
  assign io_trigger_pkt_any_1_load = tlu_io_trigger_pkt_any_1_load; // @[dec.scala 264:29]
  assign io_trigger_pkt_any_1_tdata2 = tlu_io_trigger_pkt_any_1_tdata2; // @[dec.scala 264:29]
  assign io_trigger_pkt_any_2_select = tlu_io_trigger_pkt_any_2_select; // @[dec.scala 264:29]
  assign io_trigger_pkt_any_2_match_pkt = tlu_io_trigger_pkt_any_2_match_pkt; // @[dec.scala 264:29]
  assign io_trigger_pkt_any_2_store = tlu_io_trigger_pkt_any_2_store; // @[dec.scala 264:29]
  assign io_trigger_pkt_any_2_load = tlu_io_trigger_pkt_any_2_load; // @[dec.scala 264:29]
  assign io_trigger_pkt_any_2_tdata2 = tlu_io_trigger_pkt_any_2_tdata2; // @[dec.scala 264:29]
  assign io_trigger_pkt_any_3_select = tlu_io_trigger_pkt_any_3_select; // @[dec.scala 264:29]
  assign io_trigger_pkt_any_3_match_pkt = tlu_io_trigger_pkt_any_3_match_pkt; // @[dec.scala 264:29]
  assign io_trigger_pkt_any_3_store = tlu_io_trigger_pkt_any_3_store; // @[dec.scala 264:29]
  assign io_trigger_pkt_any_3_load = tlu_io_trigger_pkt_any_3_load; // @[dec.scala 264:29]
  assign io_trigger_pkt_any_3_tdata2 = tlu_io_trigger_pkt_any_3_tdata2; // @[dec.scala 264:29]
  assign io_lsu_p_valid = decode_io_lsu_p_valid; // @[dec.scala 185:40]
  assign io_lsu_p_bits_fast_int = decode_io_lsu_p_bits_fast_int; // @[dec.scala 185:40]
  assign io_lsu_p_bits_by = decode_io_lsu_p_bits_by; // @[dec.scala 185:40]
  assign io_lsu_p_bits_half = decode_io_lsu_p_bits_half; // @[dec.scala 185:40]
  assign io_lsu_p_bits_word = decode_io_lsu_p_bits_word; // @[dec.scala 185:40]
  assign io_lsu_p_bits_load = decode_io_lsu_p_bits_load; // @[dec.scala 185:40]
  assign io_lsu_p_bits_store = decode_io_lsu_p_bits_store; // @[dec.scala 185:40]
  assign io_lsu_p_bits_unsign = decode_io_lsu_p_bits_unsign; // @[dec.scala 185:40]
  assign io_lsu_p_bits_store_data_bypass_d = decode_io_lsu_p_bits_store_data_bypass_d; // @[dec.scala 185:40]
  assign io_lsu_p_bits_load_ldst_bypass_d = decode_io_lsu_p_bits_load_ldst_bypass_d; // @[dec.scala 185:40]
  assign io_dec_lsu_offset_d = decode_io_dec_lsu_offset_d; // @[dec.scala 187:40]
  assign io_dec_tlu_i0_kill_writeb_r = tlu_io_dec_tlu_i0_kill_writeb_r; // @[dec.scala 274:34]
  assign io_dec_tlu_perfcnt0 = tlu_io_dec_tlu_perfcnt0; // @[dec.scala 275:29]
  assign io_dec_tlu_perfcnt1 = tlu_io_dec_tlu_perfcnt1; // @[dec.scala 276:29]
  assign io_dec_tlu_perfcnt2 = tlu_io_dec_tlu_perfcnt2; // @[dec.scala 277:29]
  assign io_dec_tlu_perfcnt3 = tlu_io_dec_tlu_perfcnt3; // @[dec.scala 278:29]
  assign io_dec_lsu_valid_raw_d = decode_io_dec_lsu_valid_raw_d; // @[dec.scala 186:40]
  assign io_rv_trace_pkt_rv_i_valid_ip = {tlu_io_dec_tlu_int_valid_wb1,_T_1}; // @[dec.scala 296:33]
  assign io_rv_trace_pkt_rv_i_insn_ip = decode_io_dec_i0_inst_wb1; // @[dec.scala 294:32]
  assign io_rv_trace_pkt_rv_i_address_ip = {decode_io_dec_i0_pc_wb1,1'h0}; // @[dec.scala 295:35]
  assign io_rv_trace_pkt_rv_i_exception_ip = {tlu_io_dec_tlu_int_valid_wb1,tlu_io_dec_tlu_i0_exc_valid_wb1}; // @[dec.scala 297:37]
  assign io_rv_trace_pkt_rv_i_ecause_ip = tlu_io_dec_tlu_exc_cause_wb1; // @[dec.scala 298:34]
  assign io_rv_trace_pkt_rv_i_interrupt_ip = {tlu_io_dec_tlu_int_valid_wb1,1'h0}; // @[dec.scala 299:37]
  assign io_rv_trace_pkt_rv_i_tval_ip = tlu_io_dec_tlu_mtval_wb1; // @[dec.scala 300:32]
  assign io_dec_tlu_misc_clk_override = tlu_io_dec_tlu_misc_clk_override; // @[dec.scala 284:35]
  assign io_dec_tlu_lsu_clk_override = tlu_io_dec_tlu_lsu_clk_override; // @[dec.scala 286:36]
  assign io_dec_tlu_bus_clk_override = tlu_io_dec_tlu_bus_clk_override; // @[dec.scala 287:36]
  assign io_dec_tlu_pic_clk_override = tlu_io_dec_tlu_pic_clk_override; // @[dec.scala 288:36]
  assign io_dec_tlu_dccm_clk_override = tlu_io_dec_tlu_dccm_clk_override; // @[dec.scala 289:36]
  assign io_dec_tlu_icm_clk_override = tlu_io_dec_tlu_icm_clk_override; // @[dec.scala 290:36]
  assign io_ifu_dec_dec_aln_aln_dec_dec_i0_decode_d = decode_io_dec_aln_dec_i0_decode_d; // @[dec.scala 133:21]
  assign io_ifu_dec_dec_mem_ctrl_dec_tlu_flush_err_wb = tlu_io_tlu_mem_dec_tlu_flush_err_wb; // @[dec.scala 202:18]
  assign io_ifu_dec_dec_mem_ctrl_dec_tlu_i0_commit_cmt = tlu_io_tlu_mem_dec_tlu_i0_commit_cmt; // @[dec.scala 202:18]
  assign io_ifu_dec_dec_mem_ctrl_dec_tlu_force_halt = tlu_io_tlu_mem_dec_tlu_force_halt; // @[dec.scala 202:18]
  assign io_ifu_dec_dec_mem_ctrl_dec_tlu_fence_i_wb = tlu_io_tlu_mem_dec_tlu_fence_i_wb; // @[dec.scala 202:18]
  assign io_ifu_dec_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_wrdata = tlu_io_tlu_mem_dec_tlu_ic_diag_pkt_icache_wrdata; // @[dec.scala 202:18]
  assign io_ifu_dec_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_dicawics = tlu_io_tlu_mem_dec_tlu_ic_diag_pkt_icache_dicawics; // @[dec.scala 202:18]
  assign io_ifu_dec_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_rd_valid = tlu_io_tlu_mem_dec_tlu_ic_diag_pkt_icache_rd_valid; // @[dec.scala 202:18]
  assign io_ifu_dec_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_wr_valid = tlu_io_tlu_mem_dec_tlu_ic_diag_pkt_icache_wr_valid; // @[dec.scala 202:18]
  assign io_ifu_dec_dec_mem_ctrl_dec_tlu_core_ecc_disable = tlu_io_tlu_mem_dec_tlu_core_ecc_disable; // @[dec.scala 202:18]
  assign io_ifu_dec_dec_ifc_dec_tlu_flush_noredir_wb = tlu_io_tlu_ifc_dec_tlu_flush_noredir_wb; // @[dec.scala 203:18]
  assign io_ifu_dec_dec_ifc_dec_tlu_mrac_ff = tlu_io_tlu_ifc_dec_tlu_mrac_ff; // @[dec.scala 203:18]
  assign io_ifu_dec_dec_bp_dec_tlu_br0_r_pkt_valid = tlu_io_tlu_bp_dec_tlu_br0_r_pkt_valid; // @[dec.scala 204:18]
  assign io_ifu_dec_dec_bp_dec_tlu_br0_r_pkt_bits_hist = tlu_io_tlu_bp_dec_tlu_br0_r_pkt_bits_hist; // @[dec.scala 204:18]
  assign io_ifu_dec_dec_bp_dec_tlu_br0_r_pkt_bits_br_error = tlu_io_tlu_bp_dec_tlu_br0_r_pkt_bits_br_error; // @[dec.scala 204:18]
  assign io_ifu_dec_dec_bp_dec_tlu_br0_r_pkt_bits_br_start_error = tlu_io_tlu_bp_dec_tlu_br0_r_pkt_bits_br_start_error; // @[dec.scala 204:18]
  assign io_ifu_dec_dec_bp_dec_tlu_br0_r_pkt_bits_way = tlu_io_tlu_bp_dec_tlu_br0_r_pkt_bits_way; // @[dec.scala 204:18]
  assign io_ifu_dec_dec_bp_dec_tlu_br0_r_pkt_bits_middle = tlu_io_tlu_bp_dec_tlu_br0_r_pkt_bits_middle; // @[dec.scala 204:18]
  assign io_ifu_dec_dec_bp_dec_tlu_flush_leak_one_wb = tlu_io_tlu_bp_dec_tlu_flush_leak_one_wb; // @[dec.scala 204:18]
  assign io_ifu_dec_dec_bp_dec_tlu_bpred_disable = tlu_io_tlu_bp_dec_tlu_bpred_disable; // @[dec.scala 204:18]
  assign io_dec_exu_dec_alu_dec_i0_alu_decode_d = decode_io_dec_alu_dec_i0_alu_decode_d; // @[dec.scala 136:20]
  assign io_dec_exu_dec_alu_dec_csr_ren_d = decode_io_dec_alu_dec_csr_ren_d; // @[dec.scala 136:20]
  assign io_dec_exu_dec_alu_dec_i0_br_immed_d = decode_io_dec_alu_dec_i0_br_immed_d; // @[dec.scala 136:20]
  assign io_dec_exu_dec_div_div_p_valid = decode_io_dec_div_div_p_valid; // @[dec.scala 137:20]
  assign io_dec_exu_dec_div_div_p_bits_unsign = decode_io_dec_div_div_p_bits_unsign; // @[dec.scala 137:20]
  assign io_dec_exu_dec_div_div_p_bits_rem = decode_io_dec_div_div_p_bits_rem; // @[dec.scala 137:20]
  assign io_dec_exu_dec_div_dec_div_cancel = decode_io_dec_div_dec_div_cancel; // @[dec.scala 137:20]
  assign io_dec_exu_decode_exu_dec_data_en = decode_io_decode_exu_dec_data_en; // @[dec.scala 135:23]
  assign io_dec_exu_decode_exu_dec_ctl_en = decode_io_decode_exu_dec_ctl_en; // @[dec.scala 135:23]
  assign io_dec_exu_decode_exu_i0_ap_land = decode_io_decode_exu_i0_ap_land; // @[dec.scala 135:23]
  assign io_dec_exu_decode_exu_i0_ap_lor = decode_io_decode_exu_i0_ap_lor; // @[dec.scala 135:23]
  assign io_dec_exu_decode_exu_i0_ap_lxor = decode_io_decode_exu_i0_ap_lxor; // @[dec.scala 135:23]
  assign io_dec_exu_decode_exu_i0_ap_sll = decode_io_decode_exu_i0_ap_sll; // @[dec.scala 135:23]
  assign io_dec_exu_decode_exu_i0_ap_srl = decode_io_decode_exu_i0_ap_srl; // @[dec.scala 135:23]
  assign io_dec_exu_decode_exu_i0_ap_sra = decode_io_decode_exu_i0_ap_sra; // @[dec.scala 135:23]
  assign io_dec_exu_decode_exu_i0_ap_beq = decode_io_decode_exu_i0_ap_beq; // @[dec.scala 135:23]
  assign io_dec_exu_decode_exu_i0_ap_bne = decode_io_decode_exu_i0_ap_bne; // @[dec.scala 135:23]
  assign io_dec_exu_decode_exu_i0_ap_blt = decode_io_decode_exu_i0_ap_blt; // @[dec.scala 135:23]
  assign io_dec_exu_decode_exu_i0_ap_bge = decode_io_decode_exu_i0_ap_bge; // @[dec.scala 135:23]
  assign io_dec_exu_decode_exu_i0_ap_add = decode_io_decode_exu_i0_ap_add; // @[dec.scala 135:23]
  assign io_dec_exu_decode_exu_i0_ap_sub = decode_io_decode_exu_i0_ap_sub; // @[dec.scala 135:23]
  assign io_dec_exu_decode_exu_i0_ap_slt = decode_io_decode_exu_i0_ap_slt; // @[dec.scala 135:23]
  assign io_dec_exu_decode_exu_i0_ap_unsign = decode_io_decode_exu_i0_ap_unsign; // @[dec.scala 135:23]
  assign io_dec_exu_decode_exu_i0_ap_jal = decode_io_decode_exu_i0_ap_jal; // @[dec.scala 135:23]
  assign io_dec_exu_decode_exu_i0_ap_predict_t = decode_io_decode_exu_i0_ap_predict_t; // @[dec.scala 135:23]
  assign io_dec_exu_decode_exu_i0_ap_predict_nt = decode_io_decode_exu_i0_ap_predict_nt; // @[dec.scala 135:23]
  assign io_dec_exu_decode_exu_i0_ap_csr_write = decode_io_decode_exu_i0_ap_csr_write; // @[dec.scala 135:23]
  assign io_dec_exu_decode_exu_i0_ap_csr_imm = decode_io_decode_exu_i0_ap_csr_imm; // @[dec.scala 135:23]
  assign io_dec_exu_decode_exu_dec_i0_predict_p_d_valid = decode_io_decode_exu_dec_i0_predict_p_d_valid; // @[dec.scala 135:23]
  assign io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_pc4 = decode_io_decode_exu_dec_i0_predict_p_d_bits_pc4; // @[dec.scala 135:23]
  assign io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_hist = decode_io_decode_exu_dec_i0_predict_p_d_bits_hist; // @[dec.scala 135:23]
  assign io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_toffset = decode_io_decode_exu_dec_i0_predict_p_d_bits_toffset; // @[dec.scala 135:23]
  assign io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_br_error = decode_io_decode_exu_dec_i0_predict_p_d_bits_br_error; // @[dec.scala 135:23]
  assign io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_br_start_error = decode_io_decode_exu_dec_i0_predict_p_d_bits_br_start_error; // @[dec.scala 135:23]
  assign io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_prett = decode_io_decode_exu_dec_i0_predict_p_d_bits_prett; // @[dec.scala 135:23]
  assign io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_pcall = decode_io_decode_exu_dec_i0_predict_p_d_bits_pcall; // @[dec.scala 135:23]
  assign io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_pret = decode_io_decode_exu_dec_i0_predict_p_d_bits_pret; // @[dec.scala 135:23]
  assign io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_pja = decode_io_decode_exu_dec_i0_predict_p_d_bits_pja; // @[dec.scala 135:23]
  assign io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_way = decode_io_decode_exu_dec_i0_predict_p_d_bits_way; // @[dec.scala 135:23]
  assign io_dec_exu_decode_exu_i0_predict_fghr_d = decode_io_decode_exu_i0_predict_fghr_d; // @[dec.scala 135:23]
  assign io_dec_exu_decode_exu_i0_predict_index_d = decode_io_decode_exu_i0_predict_index_d; // @[dec.scala 135:23]
  assign io_dec_exu_decode_exu_i0_predict_btag_d = decode_io_decode_exu_i0_predict_btag_d; // @[dec.scala 135:23]
  assign io_dec_exu_decode_exu_dec_i0_rs1_en_d = decode_io_decode_exu_dec_i0_rs1_en_d; // @[dec.scala 135:23]
  assign io_dec_exu_decode_exu_dec_i0_rs2_en_d = decode_io_decode_exu_dec_i0_rs2_en_d; // @[dec.scala 135:23]
  assign io_dec_exu_decode_exu_dec_i0_immed_d = decode_io_decode_exu_dec_i0_immed_d; // @[dec.scala 135:23]
  assign io_dec_exu_decode_exu_dec_i0_rs1_bypass_data_d = decode_io_decode_exu_dec_i0_rs1_bypass_data_d; // @[dec.scala 135:23]
  assign io_dec_exu_decode_exu_dec_i0_rs2_bypass_data_d = decode_io_decode_exu_dec_i0_rs2_bypass_data_d; // @[dec.scala 135:23]
  assign io_dec_exu_decode_exu_dec_i0_select_pc_d = decode_io_decode_exu_dec_i0_select_pc_d; // @[dec.scala 135:23]
  assign io_dec_exu_decode_exu_dec_i0_rs1_bypass_en_d = decode_io_decode_exu_dec_i0_rs1_bypass_en_d; // @[dec.scala 135:23]
  assign io_dec_exu_decode_exu_dec_i0_rs2_bypass_en_d = decode_io_decode_exu_dec_i0_rs2_bypass_en_d; // @[dec.scala 135:23]
  assign io_dec_exu_decode_exu_mul_p_valid = decode_io_decode_exu_mul_p_valid; // @[dec.scala 135:23]
  assign io_dec_exu_decode_exu_mul_p_bits_rs1_sign = decode_io_decode_exu_mul_p_bits_rs1_sign; // @[dec.scala 135:23]
  assign io_dec_exu_decode_exu_mul_p_bits_rs2_sign = decode_io_decode_exu_mul_p_bits_rs2_sign; // @[dec.scala 135:23]
  assign io_dec_exu_decode_exu_mul_p_bits_low = decode_io_decode_exu_mul_p_bits_low; // @[dec.scala 135:23]
  assign io_dec_exu_decode_exu_pred_correct_npc_x = decode_io_decode_exu_pred_correct_npc_x; // @[dec.scala 135:23]
  assign io_dec_exu_decode_exu_dec_extint_stall = decode_io_decode_exu_dec_extint_stall; // @[dec.scala 135:23]
  assign io_dec_exu_tlu_exu_dec_tlu_meihap = tlu_io_tlu_exu_dec_tlu_meihap; // @[dec.scala 205:18]
  assign io_dec_exu_tlu_exu_dec_tlu_flush_lower_r = tlu_io_tlu_exu_dec_tlu_flush_lower_r; // @[dec.scala 205:18]
  assign io_dec_exu_tlu_exu_dec_tlu_flush_path_r = tlu_io_tlu_exu_dec_tlu_flush_path_r; // @[dec.scala 205:18]
  assign io_dec_exu_ib_exu_dec_i0_pc_d = instbuff_io_ib_exu_dec_i0_pc_d; // @[dec.scala 126:22]
  assign io_dec_exu_ib_exu_dec_debug_wdata_rs1_d = instbuff_io_ib_exu_dec_debug_wdata_rs1_d; // @[dec.scala 126:22]
  assign io_dec_exu_gpr_exu_gpr_i0_rs1_d = gpr_io_gpr_exu_gpr_i0_rs1_d; // @[dec.scala 201:22]
  assign io_dec_exu_gpr_exu_gpr_i0_rs2_d = gpr_io_gpr_exu_gpr_i0_rs2_d; // @[dec.scala 201:22]
  assign io_lsu_dec_tlu_busbuff_dec_tlu_external_ldfwd_disable = tlu_io_tlu_busbuff_dec_tlu_external_ldfwd_disable; // @[dec.scala 222:26]
  assign io_lsu_dec_tlu_busbuff_dec_tlu_wb_coalescing_disable = tlu_io_tlu_busbuff_dec_tlu_wb_coalescing_disable; // @[dec.scala 222:26]
  assign io_lsu_dec_tlu_busbuff_dec_tlu_sideeffect_posted_disable = tlu_io_tlu_busbuff_dec_tlu_sideeffect_posted_disable; // @[dec.scala 222:26]
  assign io_dec_dma_tlu_dma_dec_tlu_dma_qos_prty = tlu_io_tlu_dma_dec_tlu_dma_qos_prty; // @[dec.scala 206:18]
  assign io_dec_pic_dec_tlu_meicurpl = tlu_io_dec_pic_dec_tlu_meicurpl; // @[dec.scala 224:14]
  assign io_dec_pic_dec_tlu_meipt = tlu_io_dec_pic_dec_tlu_meipt; // @[dec.scala 224:14]
  assign instbuff_io_ifu_ib_ifu_i0_icaf = io_ifu_dec_dec_aln_aln_ib_ifu_i0_icaf; // @[dec.scala 125:22]
  assign instbuff_io_ifu_ib_ifu_i0_icaf_type = io_ifu_dec_dec_aln_aln_ib_ifu_i0_icaf_type; // @[dec.scala 125:22]
  assign instbuff_io_ifu_ib_ifu_i0_icaf_f1 = io_ifu_dec_dec_aln_aln_ib_ifu_i0_icaf_f1; // @[dec.scala 125:22]
  assign instbuff_io_ifu_ib_ifu_i0_dbecc = io_ifu_dec_dec_aln_aln_ib_ifu_i0_dbecc; // @[dec.scala 125:22]
  assign instbuff_io_ifu_ib_ifu_i0_bp_index = io_ifu_dec_dec_aln_aln_ib_ifu_i0_bp_index; // @[dec.scala 125:22]
  assign instbuff_io_ifu_ib_ifu_i0_bp_fghr = io_ifu_dec_dec_aln_aln_ib_ifu_i0_bp_fghr; // @[dec.scala 125:22]
  assign instbuff_io_ifu_ib_ifu_i0_bp_btag = io_ifu_dec_dec_aln_aln_ib_ifu_i0_bp_btag; // @[dec.scala 125:22]
  assign instbuff_io_ifu_ib_ifu_i0_valid = io_ifu_dec_dec_aln_aln_ib_ifu_i0_valid; // @[dec.scala 125:22]
  assign instbuff_io_ifu_ib_ifu_i0_instr = io_ifu_dec_dec_aln_aln_ib_ifu_i0_instr; // @[dec.scala 125:22]
  assign instbuff_io_ifu_ib_ifu_i0_pc = io_ifu_dec_dec_aln_aln_ib_ifu_i0_pc; // @[dec.scala 125:22]
  assign instbuff_io_ifu_ib_ifu_i0_pc4 = io_ifu_dec_dec_aln_aln_ib_ifu_i0_pc4; // @[dec.scala 125:22]
  assign instbuff_io_ifu_ib_i0_brp_valid = io_ifu_dec_dec_aln_aln_ib_i0_brp_valid; // @[dec.scala 125:22]
  assign instbuff_io_ifu_ib_i0_brp_bits_toffset = io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_toffset; // @[dec.scala 125:22]
  assign instbuff_io_ifu_ib_i0_brp_bits_hist = io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_hist; // @[dec.scala 125:22]
  assign instbuff_io_ifu_ib_i0_brp_bits_br_error = io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_br_error; // @[dec.scala 125:22]
  assign instbuff_io_ifu_ib_i0_brp_bits_br_start_error = io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_br_start_error; // @[dec.scala 125:22]
  assign instbuff_io_ifu_ib_i0_brp_bits_prett = io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_prett; // @[dec.scala 125:22]
  assign instbuff_io_ifu_ib_i0_brp_bits_way = io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_way; // @[dec.scala 125:22]
  assign instbuff_io_ifu_ib_i0_brp_bits_ret = io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_ret; // @[dec.scala 125:22]
  assign instbuff_io_dbg_ib_dbg_cmd_valid = io_dec_dbg_dbg_ib_dbg_cmd_valid; // @[dec.scala 127:22]
  assign instbuff_io_dbg_ib_dbg_cmd_write = io_dec_dbg_dbg_ib_dbg_cmd_write; // @[dec.scala 127:22]
  assign instbuff_io_dbg_ib_dbg_cmd_type = io_dec_dbg_dbg_ib_dbg_cmd_type; // @[dec.scala 127:22]
  assign instbuff_io_dbg_ib_dbg_cmd_addr = io_dec_dbg_dbg_ib_dbg_cmd_addr; // @[dec.scala 127:22]
  assign decode_clock = clock;
  assign decode_reset = reset;
  assign decode_io_decode_exu_exu_i0_result_x = io_dec_exu_decode_exu_exu_i0_result_x; // @[dec.scala 135:23]
  assign decode_io_decode_exu_exu_csr_rs1_x = io_dec_exu_decode_exu_exu_csr_rs1_x; // @[dec.scala 135:23]
  assign decode_io_dec_alu_exu_i0_pc_x = io_dec_exu_dec_alu_exu_i0_pc_x; // @[dec.scala 136:20]
  assign decode_io_dctl_busbuff_lsu_nonblock_load_valid_m = io_lsu_dec_dctl_busbuff_lsu_nonblock_load_valid_m; // @[dec.scala 141:26]
  assign decode_io_dctl_busbuff_lsu_nonblock_load_tag_m = io_lsu_dec_dctl_busbuff_lsu_nonblock_load_tag_m; // @[dec.scala 141:26]
  assign decode_io_dctl_busbuff_lsu_nonblock_load_inv_r = io_lsu_dec_dctl_busbuff_lsu_nonblock_load_inv_r; // @[dec.scala 141:26]
  assign decode_io_dctl_busbuff_lsu_nonblock_load_inv_tag_r = io_lsu_dec_dctl_busbuff_lsu_nonblock_load_inv_tag_r; // @[dec.scala 141:26]
  assign decode_io_dctl_busbuff_lsu_nonblock_load_data_valid = io_lsu_dec_dctl_busbuff_lsu_nonblock_load_data_valid; // @[dec.scala 141:26]
  assign decode_io_dctl_busbuff_lsu_nonblock_load_data_error = io_lsu_dec_dctl_busbuff_lsu_nonblock_load_data_error; // @[dec.scala 141:26]
  assign decode_io_dctl_busbuff_lsu_nonblock_load_data_tag = io_lsu_dec_dctl_busbuff_lsu_nonblock_load_data_tag; // @[dec.scala 141:26]
  assign decode_io_dctl_busbuff_lsu_nonblock_load_data = io_lsu_dec_dctl_busbuff_lsu_nonblock_load_data; // @[dec.scala 141:26]
  assign decode_io_dctl_dma_dma_dccm_stall_any = io_dec_dma_dctl_dma_dma_dccm_stall_any; // @[dec.scala 138:22]
  assign decode_io_dec_aln_ifu_i0_cinst = io_ifu_dec_dec_aln_aln_dec_ifu_i0_cinst; // @[dec.scala 133:21]
  assign decode_io_dbg_dctl_dbg_cmd_wrdata = io_dec_dbg_dbg_dctl_dbg_cmd_wrdata; // @[dec.scala 150:22]
  assign decode_io_dec_tlu_flush_extint = tlu_io_dec_tlu_flush_extint; // @[dec.scala 139:48]
  assign decode_io_dec_tlu_force_halt = tlu_io_tlu_mem_dec_tlu_force_halt; // @[dec.scala 140:48]
  assign decode_io_dec_i0_trigger_match_d = dec_trigger_io_dec_i0_trigger_match_d; // @[dec.scala 142:48]
  assign decode_io_dec_tlu_wr_pause_r = tlu_io_dec_tlu_wr_pause_r; // @[dec.scala 143:48]
  assign decode_io_dec_tlu_pipelining_disable = tlu_io_dec_tlu_pipelining_disable; // @[dec.scala 144:48]
  assign decode_io_lsu_trigger_match_m = io_lsu_trigger_match_m; // @[dec.scala 145:48]
  assign decode_io_lsu_pmu_misaligned_m = io_lsu_pmu_misaligned_m; // @[dec.scala 146:48]
  assign decode_io_dec_tlu_debug_stall = tlu_io_dec_tlu_debug_stall; // @[dec.scala 147:48]
  assign decode_io_dec_tlu_flush_leak_one_r = tlu_io_tlu_bp_dec_tlu_flush_leak_one_wb; // @[dec.scala 148:48]
  assign decode_io_dec_debug_fence_d = instbuff_io_dec_debug_fence_d; // @[dec.scala 149:48]
  assign decode_io_dec_i0_icaf_d = instbuff_io_dec_i0_icaf_d; // @[dec.scala 151:48]
  assign decode_io_dec_i0_icaf_f1_d = instbuff_io_dec_i0_icaf_f1_d; // @[dec.scala 152:48]
  assign decode_io_dec_i0_icaf_type_d = instbuff_io_dec_i0_icaf_type_d; // @[dec.scala 153:48]
  assign decode_io_dec_i0_dbecc_d = instbuff_io_dec_i0_dbecc_d; // @[dec.scala 154:48]
  assign decode_io_dec_i0_brp_valid = instbuff_io_dec_i0_brp_valid; // @[dec.scala 155:48]
  assign decode_io_dec_i0_brp_bits_toffset = instbuff_io_dec_i0_brp_bits_toffset; // @[dec.scala 155:48]
  assign decode_io_dec_i0_brp_bits_hist = instbuff_io_dec_i0_brp_bits_hist; // @[dec.scala 155:48]
  assign decode_io_dec_i0_brp_bits_br_error = instbuff_io_dec_i0_brp_bits_br_error; // @[dec.scala 155:48]
  assign decode_io_dec_i0_brp_bits_br_start_error = instbuff_io_dec_i0_brp_bits_br_start_error; // @[dec.scala 155:48]
  assign decode_io_dec_i0_brp_bits_prett = instbuff_io_dec_i0_brp_bits_prett; // @[dec.scala 155:48]
  assign decode_io_dec_i0_brp_bits_way = instbuff_io_dec_i0_brp_bits_way; // @[dec.scala 155:48]
  assign decode_io_dec_i0_brp_bits_ret = instbuff_io_dec_i0_brp_bits_ret; // @[dec.scala 155:48]
  assign decode_io_dec_i0_bp_index = instbuff_io_dec_i0_bp_index; // @[dec.scala 156:48]
  assign decode_io_dec_i0_bp_fghr = instbuff_io_dec_i0_bp_fghr; // @[dec.scala 157:48]
  assign decode_io_dec_i0_bp_btag = instbuff_io_dec_i0_bp_btag; // @[dec.scala 158:48]
  assign decode_io_lsu_idle_any = io_lsu_idle_any; // @[dec.scala 160:48]
  assign decode_io_lsu_load_stall_any = io_lsu_load_stall_any; // @[dec.scala 161:48]
  assign decode_io_lsu_store_stall_any = io_lsu_store_stall_any; // @[dec.scala 162:48]
  assign decode_io_exu_div_wren = io_exu_div_wren; // @[dec.scala 163:48]
  assign decode_io_dec_tlu_i0_kill_writeb_wb = tlu_io_dec_tlu_i0_kill_writeb_wb; // @[dec.scala 164:48]
  assign decode_io_dec_tlu_flush_lower_wb = tlu_io_dec_tlu_flush_lower_wb; // @[dec.scala 165:48]
  assign decode_io_dec_tlu_i0_kill_writeb_r = tlu_io_dec_tlu_i0_kill_writeb_r; // @[dec.scala 166:48]
  assign decode_io_dec_tlu_flush_lower_r = tlu_io_tlu_exu_dec_tlu_flush_lower_r; // @[dec.scala 167:48]
  assign decode_io_dec_tlu_flush_pause_r = tlu_io_dec_tlu_flush_pause_r; // @[dec.scala 168:48]
  assign decode_io_dec_tlu_presync_d = tlu_io_dec_tlu_presync_d; // @[dec.scala 169:48]
  assign decode_io_dec_tlu_postsync_d = tlu_io_dec_tlu_postsync_d; // @[dec.scala 170:48]
  assign decode_io_dec_i0_pc4_d = instbuff_io_dec_i0_pc4_d; // @[dec.scala 171:48]
  assign decode_io_dec_csr_rddata_d = tlu_io_dec_csr_rddata_d; // @[dec.scala 172:48]
  assign decode_io_dec_csr_legal_d = tlu_io_dec_csr_legal_d; // @[dec.scala 173:48]
  assign decode_io_lsu_result_m = io_lsu_result_m; // @[dec.scala 174:48]
  assign decode_io_lsu_result_corr_r = io_lsu_result_corr_r; // @[dec.scala 175:48]
  assign decode_io_exu_flush_final = io_exu_flush_final; // @[dec.scala 176:48]
  assign decode_io_dec_i0_instr_d = instbuff_io_dec_i0_instr_d; // @[dec.scala 177:48]
  assign decode_io_dec_ib0_valid_d = instbuff_io_dec_ib0_valid_d; // @[dec.scala 178:48]
  assign decode_io_free_clk = io_free_clk; // @[dec.scala 179:48]
  assign decode_io_active_clk = io_active_clk; // @[dec.scala 180:48]
  assign decode_io_clk_override = tlu_io_dec_tlu_dec_clk_override; // @[dec.scala 181:48]
  assign decode_io_scan_mode = io_scan_mode; // @[dec.scala 182:48]
  assign gpr_clock = clock;
  assign gpr_reset = reset;
  assign gpr_io_raddr0 = decode_io_dec_i0_rs1_d; // @[dec.scala 189:23]
  assign gpr_io_raddr1 = decode_io_dec_i0_rs2_d; // @[dec.scala 190:23]
  assign gpr_io_wen0 = decode_io_dec_i0_wen_r; // @[dec.scala 191:23]
  assign gpr_io_waddr0 = decode_io_dec_i0_waddr_r; // @[dec.scala 192:23]
  assign gpr_io_wd0 = decode_io_dec_i0_wdata_r; // @[dec.scala 193:23]
  assign gpr_io_wen1 = decode_io_dec_nonblock_load_wen; // @[dec.scala 194:23]
  assign gpr_io_waddr1 = decode_io_dec_nonblock_load_waddr; // @[dec.scala 195:23]
  assign gpr_io_wd1 = io_lsu_dec_dctl_busbuff_lsu_nonblock_load_data; // @[dec.scala 196:23]
  assign gpr_io_wen2 = io_exu_div_wren; // @[dec.scala 197:23]
  assign gpr_io_waddr2 = decode_io_div_waddr_wb; // @[dec.scala 198:23]
  assign gpr_io_wd2 = io_exu_div_result; // @[dec.scala 199:23]
  assign gpr_io_scan_mode = io_scan_mode; // @[dec.scala 200:23]
  assign tlu_clock = clock;
  assign tlu_reset = reset;
  assign tlu_io_tlu_exu_exu_i0_br_hist_r = io_dec_exu_tlu_exu_exu_i0_br_hist_r; // @[dec.scala 205:18]
  assign tlu_io_tlu_exu_exu_i0_br_error_r = io_dec_exu_tlu_exu_exu_i0_br_error_r; // @[dec.scala 205:18]
  assign tlu_io_tlu_exu_exu_i0_br_start_error_r = io_dec_exu_tlu_exu_exu_i0_br_start_error_r; // @[dec.scala 205:18]
  assign tlu_io_tlu_exu_exu_i0_br_valid_r = io_dec_exu_tlu_exu_exu_i0_br_valid_r; // @[dec.scala 205:18]
  assign tlu_io_tlu_exu_exu_i0_br_mp_r = io_dec_exu_tlu_exu_exu_i0_br_mp_r; // @[dec.scala 205:18]
  assign tlu_io_tlu_exu_exu_i0_br_middle_r = io_dec_exu_tlu_exu_exu_i0_br_middle_r; // @[dec.scala 205:18]
  assign tlu_io_tlu_exu_exu_pmu_i0_br_misp = io_dec_exu_tlu_exu_exu_pmu_i0_br_misp; // @[dec.scala 205:18]
  assign tlu_io_tlu_exu_exu_pmu_i0_br_ataken = io_dec_exu_tlu_exu_exu_pmu_i0_br_ataken; // @[dec.scala 205:18]
  assign tlu_io_tlu_exu_exu_pmu_i0_pc4 = io_dec_exu_tlu_exu_exu_pmu_i0_pc4; // @[dec.scala 205:18]
  assign tlu_io_tlu_exu_exu_npc_r = io_dec_exu_tlu_exu_exu_npc_r; // @[dec.scala 205:18]
  assign tlu_io_tlu_dma_dma_pmu_dccm_read = io_dec_dma_tlu_dma_dma_pmu_dccm_read; // @[dec.scala 206:18]
  assign tlu_io_tlu_dma_dma_pmu_dccm_write = io_dec_dma_tlu_dma_dma_pmu_dccm_write; // @[dec.scala 206:18]
  assign tlu_io_tlu_dma_dma_pmu_any_read = io_dec_dma_tlu_dma_dma_pmu_any_read; // @[dec.scala 206:18]
  assign tlu_io_tlu_dma_dma_pmu_any_write = io_dec_dma_tlu_dma_dma_pmu_any_write; // @[dec.scala 206:18]
  assign tlu_io_tlu_dma_dma_dccm_stall_any = io_dec_dma_tlu_dma_dma_dccm_stall_any; // @[dec.scala 206:18]
  assign tlu_io_tlu_dma_dma_iccm_stall_any = io_dec_dma_tlu_dma_dma_iccm_stall_any; // @[dec.scala 206:18]
  assign tlu_io_active_clk = io_active_clk; // @[dec.scala 207:45]
  assign tlu_io_free_clk = io_free_clk; // @[dec.scala 208:45]
  assign tlu_io_scan_mode = io_scan_mode; // @[dec.scala 209:45]
  assign tlu_io_rst_vec = io_rst_vec; // @[dec.scala 210:45]
  assign tlu_io_nmi_int = io_nmi_int; // @[dec.scala 211:45]
  assign tlu_io_nmi_vec = io_nmi_vec; // @[dec.scala 212:45]
  assign tlu_io_i_cpu_halt_req = io_i_cpu_halt_req; // @[dec.scala 213:45]
  assign tlu_io_i_cpu_run_req = io_i_cpu_run_req; // @[dec.scala 214:45]
  assign tlu_io_lsu_fastint_stall_any = io_lsu_fastint_stall_any; // @[dec.scala 215:45]
  assign tlu_io_lsu_idle_any = io_lsu_idle_any; // @[dec.scala 246:45]
  assign tlu_io_dec_pmu_instr_decoded = decode_io_dec_pmu_instr_decoded; // @[dec.scala 217:45]
  assign tlu_io_dec_pmu_decode_stall = decode_io_dec_pmu_decode_stall; // @[dec.scala 218:45]
  assign tlu_io_dec_pmu_presync_stall = decode_io_dec_pmu_presync_stall; // @[dec.scala 219:45]
  assign tlu_io_dec_pmu_postsync_stall = decode_io_dec_pmu_postsync_stall; // @[dec.scala 220:45]
  assign tlu_io_lsu_store_stall_any = io_lsu_store_stall_any; // @[dec.scala 221:45]
  assign tlu_io_lsu_fir_addr = io_lsu_fir_addr; // @[dec.scala 225:45]
  assign tlu_io_lsu_fir_error = io_lsu_fir_error; // @[dec.scala 226:45]
  assign tlu_io_iccm_dma_sb_error = io_iccm_dma_sb_error; // @[dec.scala 227:45]
  assign tlu_io_lsu_error_pkt_r_valid = io_lsu_error_pkt_r_valid; // @[dec.scala 228:45]
  assign tlu_io_lsu_error_pkt_r_bits_single_ecc_error = io_lsu_error_pkt_r_bits_single_ecc_error; // @[dec.scala 228:45]
  assign tlu_io_lsu_error_pkt_r_bits_inst_type = io_lsu_error_pkt_r_bits_inst_type; // @[dec.scala 228:45]
  assign tlu_io_lsu_error_pkt_r_bits_exc_type = io_lsu_error_pkt_r_bits_exc_type; // @[dec.scala 228:45]
  assign tlu_io_lsu_error_pkt_r_bits_mscause = io_lsu_error_pkt_r_bits_mscause; // @[dec.scala 228:45]
  assign tlu_io_lsu_error_pkt_r_bits_addr = io_lsu_error_pkt_r_bits_addr; // @[dec.scala 228:45]
  assign tlu_io_lsu_single_ecc_error_incr = io_lsu_single_ecc_error_incr; // @[dec.scala 229:45]
  assign tlu_io_dec_pause_state = decode_io_dec_pause_state; // @[dec.scala 230:45]
  assign tlu_io_dec_csr_wen_unq_d = decode_io_dec_csr_wen_unq_d; // @[dec.scala 231:45]
  assign tlu_io_dec_csr_any_unq_d = decode_io_dec_csr_any_unq_d; // @[dec.scala 232:45]
  assign tlu_io_dec_csr_rdaddr_d = decode_io_dec_csr_rdaddr_d; // @[dec.scala 233:45]
  assign tlu_io_dec_csr_wen_r = decode_io_dec_csr_wen_r; // @[dec.scala 234:45]
  assign tlu_io_dec_csr_wraddr_r = decode_io_dec_csr_wraddr_r; // @[dec.scala 235:45]
  assign tlu_io_dec_csr_wrdata_r = decode_io_dec_csr_wrdata_r; // @[dec.scala 236:45]
  assign tlu_io_dec_csr_stall_int_ff = decode_io_dec_csr_stall_int_ff; // @[dec.scala 237:45]
  assign tlu_io_dec_tlu_i0_valid_r = decode_io_dec_tlu_i0_valid_r; // @[dec.scala 238:45]
  assign tlu_io_dec_tlu_i0_pc_r = decode_io_dec_tlu_i0_pc_r; // @[dec.scala 239:45]
  assign tlu_io_dec_tlu_packet_r_legal = decode_io_dec_tlu_packet_r_legal; // @[dec.scala 240:45]
  assign tlu_io_dec_tlu_packet_r_icaf = decode_io_dec_tlu_packet_r_icaf; // @[dec.scala 240:45]
  assign tlu_io_dec_tlu_packet_r_icaf_f1 = decode_io_dec_tlu_packet_r_icaf_f1; // @[dec.scala 240:45]
  assign tlu_io_dec_tlu_packet_r_icaf_type = decode_io_dec_tlu_packet_r_icaf_type; // @[dec.scala 240:45]
  assign tlu_io_dec_tlu_packet_r_fence_i = decode_io_dec_tlu_packet_r_fence_i; // @[dec.scala 240:45]
  assign tlu_io_dec_tlu_packet_r_i0trigger = decode_io_dec_tlu_packet_r_i0trigger; // @[dec.scala 240:45]
  assign tlu_io_dec_tlu_packet_r_pmu_i0_itype = decode_io_dec_tlu_packet_r_pmu_i0_itype; // @[dec.scala 240:45]
  assign tlu_io_dec_tlu_packet_r_pmu_i0_br_unpred = decode_io_dec_tlu_packet_r_pmu_i0_br_unpred; // @[dec.scala 240:45]
  assign tlu_io_dec_tlu_packet_r_pmu_divide = decode_io_dec_tlu_packet_r_pmu_divide; // @[dec.scala 240:45]
  assign tlu_io_dec_tlu_packet_r_pmu_lsu_misaligned = decode_io_dec_tlu_packet_r_pmu_lsu_misaligned; // @[dec.scala 240:45]
  assign tlu_io_dec_illegal_inst = decode_io_dec_illegal_inst; // @[dec.scala 241:45]
  assign tlu_io_dec_i0_decode_d = decode_io_dec_aln_dec_i0_decode_d; // @[dec.scala 242:45]
  assign tlu_io_exu_i0_br_way_r = io_exu_i0_br_way_r; // @[dec.scala 243:45]
  assign tlu_io_dbg_halt_req = io_dbg_halt_req; // @[dec.scala 244:45]
  assign tlu_io_dbg_resume_req = io_dbg_resume_req; // @[dec.scala 245:45]
  assign tlu_io_dec_div_active = decode_io_dec_div_active; // @[dec.scala 247:45]
  assign tlu_io_timer_int = io_timer_int; // @[dec.scala 252:45]
  assign tlu_io_soft_int = io_soft_int; // @[dec.scala 253:45]
  assign tlu_io_core_id = io_core_id; // @[dec.scala 254:45]
  assign tlu_io_mpc_debug_halt_req = io_mpc_debug_halt_req; // @[dec.scala 255:45]
  assign tlu_io_mpc_debug_run_req = io_mpc_debug_run_req; // @[dec.scala 256:45]
  assign tlu_io_mpc_reset_run_req = io_mpc_reset_run_req; // @[dec.scala 257:45]
  assign tlu_io_ifu_pmu_instr_aligned = io_ifu_dec_dec_aln_ifu_pmu_instr_aligned; // @[dec.scala 216:45]
  assign tlu_io_tlu_ifc_ifu_pmu_fetch_stall = io_ifu_dec_dec_ifc_ifu_pmu_fetch_stall; // @[dec.scala 203:18]
  assign tlu_io_tlu_mem_ifu_pmu_ic_miss = io_ifu_dec_dec_mem_ctrl_ifu_pmu_ic_miss; // @[dec.scala 202:18]
  assign tlu_io_tlu_mem_ifu_pmu_ic_hit = io_ifu_dec_dec_mem_ctrl_ifu_pmu_ic_hit; // @[dec.scala 202:18]
  assign tlu_io_tlu_mem_ifu_pmu_bus_error = io_ifu_dec_dec_mem_ctrl_ifu_pmu_bus_error; // @[dec.scala 202:18]
  assign tlu_io_tlu_mem_ifu_pmu_bus_busy = io_ifu_dec_dec_mem_ctrl_ifu_pmu_bus_busy; // @[dec.scala 202:18]
  assign tlu_io_tlu_mem_ifu_ic_error_start = io_ifu_dec_dec_mem_ctrl_ifu_ic_error_start; // @[dec.scala 202:18]
  assign tlu_io_tlu_mem_ifu_iccm_rd_ecc_single_err = io_ifu_dec_dec_mem_ctrl_ifu_iccm_rd_ecc_single_err; // @[dec.scala 202:18]
  assign tlu_io_tlu_mem_ifu_ic_debug_rd_data = io_ifu_dec_dec_mem_ctrl_ifu_ic_debug_rd_data; // @[dec.scala 202:18]
  assign tlu_io_tlu_mem_ifu_ic_debug_rd_data_valid = io_ifu_dec_dec_mem_ctrl_ifu_ic_debug_rd_data_valid; // @[dec.scala 202:18]
  assign tlu_io_tlu_mem_ifu_miss_state_idle = io_ifu_dec_dec_mem_ctrl_ifu_miss_state_idle; // @[dec.scala 202:18]
  assign tlu_io_tlu_busbuff_lsu_pmu_bus_misaligned = io_lsu_dec_tlu_busbuff_lsu_pmu_bus_misaligned; // @[dec.scala 222:26]
  assign tlu_io_tlu_busbuff_lsu_pmu_bus_error = io_lsu_dec_tlu_busbuff_lsu_pmu_bus_error; // @[dec.scala 222:26]
  assign tlu_io_tlu_busbuff_lsu_pmu_bus_busy = io_lsu_dec_tlu_busbuff_lsu_pmu_bus_busy; // @[dec.scala 222:26]
  assign tlu_io_tlu_busbuff_lsu_imprecise_error_load_any = io_lsu_dec_tlu_busbuff_lsu_imprecise_error_load_any; // @[dec.scala 222:26]
  assign tlu_io_tlu_busbuff_lsu_imprecise_error_store_any = io_lsu_dec_tlu_busbuff_lsu_imprecise_error_store_any; // @[dec.scala 222:26]
  assign tlu_io_tlu_busbuff_lsu_imprecise_error_addr_any = io_lsu_dec_tlu_busbuff_lsu_imprecise_error_addr_any; // @[dec.scala 222:26]
  assign tlu_io_lsu_tlu_lsu_pmu_load_external_m = io_lsu_tlu_lsu_pmu_load_external_m; // @[dec.scala 223:14]
  assign tlu_io_lsu_tlu_lsu_pmu_store_external_m = io_lsu_tlu_lsu_pmu_store_external_m; // @[dec.scala 223:14]
  assign tlu_io_dec_pic_pic_claimid = io_dec_pic_pic_claimid; // @[dec.scala 224:14]
  assign tlu_io_dec_pic_pic_pl = io_dec_pic_pic_pl; // @[dec.scala 224:14]
  assign tlu_io_dec_pic_mhwakeup = io_dec_pic_mhwakeup; // @[dec.scala 224:14]
  assign tlu_io_dec_pic_mexintpend = io_dec_pic_mexintpend; // @[dec.scala 224:14]
  assign dec_trigger_io_trigger_pkt_any_0_select = tlu_io_trigger_pkt_any_0_select; // @[dec.scala 129:34]
  assign dec_trigger_io_trigger_pkt_any_0_match_pkt = tlu_io_trigger_pkt_any_0_match_pkt; // @[dec.scala 129:34]
  assign dec_trigger_io_trigger_pkt_any_0_execute = tlu_io_trigger_pkt_any_0_execute; // @[dec.scala 129:34]
  assign dec_trigger_io_trigger_pkt_any_0_m = tlu_io_trigger_pkt_any_0_m; // @[dec.scala 129:34]
  assign dec_trigger_io_trigger_pkt_any_0_tdata2 = tlu_io_trigger_pkt_any_0_tdata2; // @[dec.scala 129:34]
  assign dec_trigger_io_trigger_pkt_any_1_select = tlu_io_trigger_pkt_any_1_select; // @[dec.scala 129:34]
  assign dec_trigger_io_trigger_pkt_any_1_match_pkt = tlu_io_trigger_pkt_any_1_match_pkt; // @[dec.scala 129:34]
  assign dec_trigger_io_trigger_pkt_any_1_execute = tlu_io_trigger_pkt_any_1_execute; // @[dec.scala 129:34]
  assign dec_trigger_io_trigger_pkt_any_1_m = tlu_io_trigger_pkt_any_1_m; // @[dec.scala 129:34]
  assign dec_trigger_io_trigger_pkt_any_1_tdata2 = tlu_io_trigger_pkt_any_1_tdata2; // @[dec.scala 129:34]
  assign dec_trigger_io_trigger_pkt_any_2_select = tlu_io_trigger_pkt_any_2_select; // @[dec.scala 129:34]
  assign dec_trigger_io_trigger_pkt_any_2_match_pkt = tlu_io_trigger_pkt_any_2_match_pkt; // @[dec.scala 129:34]
  assign dec_trigger_io_trigger_pkt_any_2_execute = tlu_io_trigger_pkt_any_2_execute; // @[dec.scala 129:34]
  assign dec_trigger_io_trigger_pkt_any_2_m = tlu_io_trigger_pkt_any_2_m; // @[dec.scala 129:34]
  assign dec_trigger_io_trigger_pkt_any_2_tdata2 = tlu_io_trigger_pkt_any_2_tdata2; // @[dec.scala 129:34]
  assign dec_trigger_io_trigger_pkt_any_3_select = tlu_io_trigger_pkt_any_3_select; // @[dec.scala 129:34]
  assign dec_trigger_io_trigger_pkt_any_3_match_pkt = tlu_io_trigger_pkt_any_3_match_pkt; // @[dec.scala 129:34]
  assign dec_trigger_io_trigger_pkt_any_3_execute = tlu_io_trigger_pkt_any_3_execute; // @[dec.scala 129:34]
  assign dec_trigger_io_trigger_pkt_any_3_m = tlu_io_trigger_pkt_any_3_m; // @[dec.scala 129:34]
  assign dec_trigger_io_trigger_pkt_any_3_tdata2 = tlu_io_trigger_pkt_any_3_tdata2; // @[dec.scala 129:34]
  assign dec_trigger_io_dec_i0_pc_d = instbuff_io_ib_exu_dec_i0_pc_d; // @[dec.scala 128:30]
endmodule
module dbg(
  input         clock,
  input         reset,
  output [1:0]  io_dbg_cmd_size,
  output        io_dbg_core_rst_l,
  input  [31:0] io_core_dbg_rddata,
  input         io_core_dbg_cmd_done,
  input         io_core_dbg_cmd_fail,
  output        io_dbg_halt_req,
  output        io_dbg_resume_req,
  input         io_dec_tlu_debug_mode,
  input         io_dec_tlu_dbg_halted,
  input         io_dec_tlu_mpc_halted_only,
  input         io_dec_tlu_resume_ack,
  input         io_dmi_reg_en,
  input  [6:0]  io_dmi_reg_addr,
  input         io_dmi_reg_wr_en,
  input  [31:0] io_dmi_reg_wdata,
  output        io_sb_axi_aw_valid,
  output [31:0] io_sb_axi_aw_bits_addr,
  output [2:0]  io_sb_axi_aw_bits_size,
  output        io_sb_axi_w_valid,
  output [7:0]  io_sb_axi_w_bits_strb,
  output        io_sb_axi_ar_valid,
  output [31:0] io_sb_axi_ar_bits_addr,
  output [2:0]  io_sb_axi_ar_bits_size,
  output        io_dbg_dec_dbg_ib_dbg_cmd_valid,
  output        io_dbg_dec_dbg_ib_dbg_cmd_write,
  output [1:0]  io_dbg_dec_dbg_ib_dbg_cmd_type,
  output [31:0] io_dbg_dec_dbg_ib_dbg_cmd_addr,
  output [31:0] io_dbg_dec_dbg_dctl_dbg_cmd_wrdata,
  output        io_dbg_dma_dbg_ib_dbg_cmd_valid,
  output        io_dbg_dma_dbg_ib_dbg_cmd_write,
  output [1:0]  io_dbg_dma_dbg_ib_dbg_cmd_type,
  output [31:0] io_dbg_dma_dbg_ib_dbg_cmd_addr,
  output [31:0] io_dbg_dma_dbg_dctl_dbg_cmd_wrdata,
  output        io_dbg_dma_io_dbg_dma_bubble,
  input         io_dbg_dma_io_dma_dbg_ready,
  input         io_dbg_bus_clk_en,
  input         io_dbg_rst_l,
  input         io_clk_override,
  input         io_scan_mode
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
`endif // RANDOMIZE_REG_INIT
  wire [2:0] dbg_state;
  wire  dbg_state_en;
  wire [3:0] sb_state;
  wire  sb_state_en;
  wire [31:0] dmcontrol_reg;
  wire [31:0] sbaddress0_reg;
  wire  sbcs_sbbusy_wren;
  wire  sbcs_sberror_wren;
  wire  sbaddress0_reg_wren1;
  wire [31:0] dmstatus_reg;
  wire  dmstatus_havereset;
  wire  dmstatus_resumeack;
  wire  dmstatus_unavail;
  wire  dmstatus_running;
  wire  dmstatus_halted;
  wire  abstractcs_busy_wren;
  wire  sbcs_sbbusy_din;
  wire [31:0] data1_reg;
  wire [31:0] sbcs_reg;
  wire  _T = dbg_state != 3'h0; // @[dbg.scala 95:51]
  wire  _T_1 = io_dmi_reg_en | _T; // @[dbg.scala 95:38]
  wire  _T_2 = _T_1 | dbg_state_en; // @[dbg.scala 95:69]
  wire  _T_3 = _T_2 | io_dec_tlu_dbg_halted; // @[dbg.scala 95:84]
  wire  _T_4 = io_dmi_reg_en | sb_state_en; // @[dbg.scala 96:37]
  wire  _T_5 = sb_state != 4'h0; // @[dbg.scala 96:63]
  wire  _T_6 = _T_4 | _T_5; // @[dbg.scala 96:51]
  wire  rvclkhdr_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_1_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_1_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_1_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_1_io_scan_mode; // @[lib.scala 343:22]
  wire  _T_9 = dmcontrol_reg[0] | io_scan_mode; // @[dbg.scala 100:65]
  wire  dbg_dm_rst_l = io_dbg_rst_l & _T_9; // @[dbg.scala 100:94]
  wire  _T_11 = io_dbg_rst_l & _T_9; // @[dbg.scala 102:38]
  wire  rst_temp = _T_11 & reset; // @[dbg.scala 102:71]
  wire  rst_not = ~_T_11; // @[dbg.scala 104:52]
  wire  _T_17 = ~dmcontrol_reg[1]; // @[dbg.scala 107:25]
  wire  _T_19 = io_dmi_reg_addr == 7'h38; // @[dbg.scala 108:36]
  wire  _T_20 = _T_19 & io_dmi_reg_en; // @[dbg.scala 108:49]
  wire  _T_21 = _T_20 & io_dmi_reg_wr_en; // @[dbg.scala 108:65]
  wire  _T_22 = sb_state == 4'h0; // @[dbg.scala 108:96]
  wire  sbcs_wren = _T_21 & _T_22; // @[dbg.scala 108:84]
  wire  _T_24 = sbcs_wren & io_dmi_reg_wdata[22]; // @[dbg.scala 109:42]
  wire  _T_26 = _T_5 & io_dmi_reg_en; // @[dbg.scala 109:102]
  wire  _T_27 = io_dmi_reg_addr == 7'h39; // @[dbg.scala 110:23]
  wire  _T_28 = io_dmi_reg_addr == 7'h3c; // @[dbg.scala 110:55]
  wire  _T_29 = _T_27 | _T_28; // @[dbg.scala 110:36]
  wire  _T_30 = io_dmi_reg_addr == 7'h3d; // @[dbg.scala 110:87]
  wire  _T_31 = _T_29 | _T_30; // @[dbg.scala 110:68]
  wire  _T_32 = _T_26 & _T_31; // @[dbg.scala 109:118]
  wire  sbcs_sbbusyerror_wren = _T_24 | _T_32; // @[dbg.scala 109:66]
  wire  sbcs_sbbusyerror_din = ~_T_24; // @[dbg.scala 112:31]
  reg  temp_sbcs_22; // @[Reg.scala 27:20]
  reg  temp_sbcs_21; // @[Reg.scala 27:20]
  reg  temp_sbcs_20; // @[Reg.scala 27:20]
  reg [4:0] temp_sbcs_19_15; // @[Reg.scala 27:20]
  reg [2:0] temp_sbcs_14_12; // @[Reg.scala 27:20]
  wire [19:0] _T_40 = {temp_sbcs_19_15,temp_sbcs_14_12,12'h40f}; // @[Cat.scala 29:58]
  wire [11:0] _T_44 = {9'h40,temp_sbcs_22,temp_sbcs_21,temp_sbcs_20}; // @[Cat.scala 29:58]
  wire  _T_47 = sbcs_reg[19:17] == 3'h1; // @[dbg.scala 134:42]
  wire  _T_49 = _T_47 & sbaddress0_reg[0]; // @[dbg.scala 134:61]
  wire  _T_51 = sbcs_reg[19:17] == 3'h2; // @[dbg.scala 135:23]
  wire  _T_53 = |sbaddress0_reg[1:0]; // @[dbg.scala 135:65]
  wire  _T_54 = _T_51 & _T_53; // @[dbg.scala 135:42]
  wire  _T_55 = _T_49 | _T_54; // @[dbg.scala 134:81]
  wire  _T_57 = sbcs_reg[19:17] == 3'h3; // @[dbg.scala 136:23]
  wire  _T_59 = |sbaddress0_reg[2:0]; // @[dbg.scala 136:65]
  wire  _T_60 = _T_57 & _T_59; // @[dbg.scala 136:42]
  wire  sbcs_unaligned = _T_55 | _T_60; // @[dbg.scala 135:69]
  wire  sbcs_illegal_size = sbcs_reg[19]; // @[dbg.scala 138:35]
  wire  _T_62 = sbcs_reg[19:17] == 3'h0; // @[dbg.scala 139:51]
  wire [3:0] _T_64 = _T_62 ? 4'hf : 4'h0; // @[Bitwise.scala 72:12]
  wire [3:0] _T_65 = _T_64 & 4'h1; // @[dbg.scala 139:64]
  wire [3:0] _T_69 = _T_47 ? 4'hf : 4'h0; // @[Bitwise.scala 72:12]
  wire [3:0] _T_70 = _T_69 & 4'h2; // @[dbg.scala 139:122]
  wire [3:0] _T_71 = _T_65 | _T_70; // @[dbg.scala 139:81]
  wire [3:0] _T_75 = _T_51 ? 4'hf : 4'h0; // @[Bitwise.scala 72:12]
  wire [3:0] _T_76 = _T_75 & 4'h4; // @[dbg.scala 140:44]
  wire [3:0] _T_77 = _T_71 | _T_76; // @[dbg.scala 139:139]
  wire [3:0] _T_81 = _T_57 ? 4'hf : 4'h0; // @[Bitwise.scala 72:12]
  wire [3:0] _T_82 = _T_81 & 4'h8; // @[dbg.scala 140:102]
  wire [3:0] sbaddress0_incr = _T_77 | _T_82; // @[dbg.scala 140:61]
  wire  _T_83 = io_dmi_reg_en & io_dmi_reg_wr_en; // @[dbg.scala 142:41]
  wire  sbdata0_reg_wren0 = _T_83 & _T_28; // @[dbg.scala 142:60]
  wire  _T_85 = sb_state == 4'h7; // @[dbg.scala 143:37]
  wire  _T_86 = _T_85 & sb_state_en; // @[dbg.scala 143:60]
  wire  _T_87 = ~sbcs_sberror_wren; // @[dbg.scala 143:76]
  wire  sbdata0_reg_wren1 = _T_86 & _T_87; // @[dbg.scala 143:74]
  wire  sbdata1_reg_wren0 = _T_83 & _T_30; // @[dbg.scala 145:60]
  wire  rvclkhdr_2_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_2_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_2_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_2_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_3_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_3_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_3_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_3_io_scan_mode; // @[lib.scala 368:23]
  wire  sbaddress0_reg_wren0 = _T_83 & _T_27; // @[dbg.scala 162:63]
  wire [31:0] _T_110 = sbaddress0_reg_wren0 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_111 = _T_110 & io_dmi_reg_wdata; // @[dbg.scala 164:59]
  wire [31:0] _T_113 = sbaddress0_reg_wren1 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_114 = {28'h0,sbaddress0_incr}; // @[Cat.scala 29:58]
  wire [31:0] _T_116 = sbaddress0_reg + _T_114; // @[dbg.scala 165:54]
  wire [31:0] _T_117 = _T_113 & _T_116; // @[dbg.scala 165:36]
  wire  rvclkhdr_4_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_4_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_4_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_4_io_scan_mode; // @[lib.scala 368:23]
  reg [31:0] _T_118; // @[lib.scala 374:16]
  wire  sbreadonaddr_access = sbaddress0_reg_wren0 & sbcs_reg[20]; // @[dbg.scala 170:94]
  wire  _T_123 = ~io_dmi_reg_wr_en; // @[dbg.scala 171:45]
  wire  _T_124 = io_dmi_reg_en & _T_123; // @[dbg.scala 171:43]
  wire  _T_126 = _T_124 & _T_28; // @[dbg.scala 171:63]
  wire  sbreadondata_access = _T_126 & sbcs_reg[15]; // @[dbg.scala 171:95]
  wire  _T_130 = io_dmi_reg_addr == 7'h10; // @[dbg.scala 173:41]
  wire  _T_131 = _T_130 & io_dmi_reg_en; // @[dbg.scala 173:54]
  wire  dmcontrol_wren = _T_131 & io_dmi_reg_wr_en; // @[dbg.scala 173:70]
  wire [3:0] _T_136 = {io_dmi_reg_wdata[31:30],io_dmi_reg_wdata[28],io_dmi_reg_wdata[1]}; // @[Cat.scala 29:58]
  reg [3:0] dm_temp; // @[Reg.scala 27:20]
  reg  dm_temp_0; // @[Reg.scala 27:20]
  wire [27:0] _T_143 = {26'h0,dm_temp[0],dm_temp_0}; // @[Cat.scala 29:58]
  wire [3:0] _T_145 = {dm_temp[3:2],1'h0,dm_temp[1]}; // @[Cat.scala 29:58]
  reg  dmcontrol_wren_Q; // @[dbg.scala 188:12]
  wire [1:0] _T_147 = dmstatus_havereset ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [1:0] _T_149 = dmstatus_resumeack ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [1:0] _T_151 = dmstatus_unavail ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [1:0] _T_153 = dmstatus_running ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [1:0] _T_155 = dmstatus_halted ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [11:0] _T_159 = {_T_153,_T_155,1'h1,7'h2}; // @[Cat.scala 29:58]
  wire [19:0] _T_163 = {12'h0,_T_147,_T_149,2'h0,_T_151}; // @[Cat.scala 29:58]
  wire  _T_165 = dbg_state == 3'h6; // @[dbg.scala 193:44]
  wire  _T_166 = _T_165 & io_dec_tlu_resume_ack; // @[dbg.scala 193:66]
  wire  _T_168 = ~dmcontrol_reg[30]; // @[dbg.scala 193:113]
  wire  _T_169 = dmstatus_resumeack & _T_168; // @[dbg.scala 193:111]
  wire  dmstatus_resumeack_wren = _T_166 | _T_169; // @[dbg.scala 193:90]
  wire  _T_173 = _T_130 & io_dmi_reg_wdata[1]; // @[dbg.scala 195:63]
  wire  _T_174 = _T_173 & io_dmi_reg_en; // @[dbg.scala 195:85]
  wire  dmstatus_havereset_wren = _T_174 & io_dmi_reg_wr_en; // @[dbg.scala 195:101]
  wire  _T_177 = _T_130 & io_dmi_reg_wdata[28]; // @[dbg.scala 196:62]
  wire  _T_178 = _T_177 & io_dmi_reg_en; // @[dbg.scala 196:85]
  wire  dmstatus_havereset_rst = _T_178 & io_dmi_reg_wr_en; // @[dbg.scala 196:101]
  wire  _T_180 = ~reset; // @[dbg.scala 198:43]
  wire  _T_183 = dmstatus_unavail | dmstatus_halted; // @[dbg.scala 199:42]
  reg  _T_185; // @[Reg.scala 27:20]
  wire  _T_186 = ~io_dec_tlu_mpc_halted_only; // @[dbg.scala 205:37]
  reg  _T_188; // @[dbg.scala 205:12]
  wire  _T_189 = dmstatus_havereset_wren | dmstatus_havereset; // @[dbg.scala 209:16]
  wire  _T_190 = ~dmstatus_havereset_rst; // @[dbg.scala 209:72]
  reg  _T_192; // @[dbg.scala 209:12]
  wire [31:0] abstractcs_reg;
  wire  _T_194 = abstractcs_reg[12] & io_dmi_reg_en; // @[dbg.scala 215:50]
  wire  _T_195 = io_dmi_reg_addr == 7'h16; // @[dbg.scala 215:106]
  wire  _T_196 = io_dmi_reg_addr == 7'h17; // @[dbg.scala 215:138]
  wire  _T_197 = _T_195 | _T_196; // @[dbg.scala 215:119]
  wire  _T_198 = io_dmi_reg_wr_en & _T_197; // @[dbg.scala 215:86]
  wire  _T_199 = io_dmi_reg_addr == 7'h4; // @[dbg.scala 215:171]
  wire  _T_200 = _T_198 | _T_199; // @[dbg.scala 215:152]
  wire  abstractcs_error_sel0 = _T_194 & _T_200; // @[dbg.scala 215:66]
  wire  _T_203 = _T_83 & _T_196; // @[dbg.scala 216:64]
  wire  _T_205 = io_dmi_reg_wdata[31:24] == 8'h0; // @[dbg.scala 216:126]
  wire  _T_207 = io_dmi_reg_wdata[31:24] == 8'h2; // @[dbg.scala 216:163]
  wire  _T_208 = _T_205 | _T_207; // @[dbg.scala 216:135]
  wire  _T_209 = ~_T_208; // @[dbg.scala 216:98]
  wire  abstractcs_error_sel1 = _T_203 & _T_209; // @[dbg.scala 216:96]
  wire  abstractcs_error_sel2 = io_core_dbg_cmd_done & io_core_dbg_cmd_fail; // @[dbg.scala 217:52]
  wire  _T_214 = ~dmstatus_reg[9]; // @[dbg.scala 218:98]
  wire  abstractcs_error_sel3 = _T_203 & _T_214; // @[dbg.scala 218:96]
  wire  _T_216 = _T_196 & io_dmi_reg_en; // @[dbg.scala 219:61]
  wire  _T_217 = _T_216 & io_dmi_reg_wr_en; // @[dbg.scala 219:77]
  wire  _T_219 = io_dmi_reg_wdata[22:20] != 3'h2; // @[dbg.scala 220:32]
  wire  _T_223 = |data1_reg[1:0]; // @[dbg.scala 220:111]
  wire  _T_224 = _T_207 & _T_223; // @[dbg.scala 220:92]
  wire  _T_225 = _T_219 | _T_224; // @[dbg.scala 220:51]
  wire  abstractcs_error_sel4 = _T_217 & _T_225; // @[dbg.scala 219:96]
  wire  _T_227 = _T_195 & io_dmi_reg_en; // @[dbg.scala 222:61]
  wire  abstractcs_error_sel5 = _T_227 & io_dmi_reg_wr_en; // @[dbg.scala 222:77]
  wire  _T_228 = abstractcs_error_sel0 | abstractcs_error_sel1; // @[dbg.scala 223:54]
  wire  _T_229 = _T_228 | abstractcs_error_sel2; // @[dbg.scala 223:78]
  wire  _T_230 = _T_229 | abstractcs_error_sel3; // @[dbg.scala 223:102]
  wire  _T_231 = _T_230 | abstractcs_error_sel4; // @[dbg.scala 223:126]
  wire  abstractcs_error_selor = _T_231 | abstractcs_error_sel5; // @[dbg.scala 223:150]
  wire [2:0] _T_233 = abstractcs_error_sel0 ? 3'h7 : 3'h0; // @[Bitwise.scala 72:12]
  wire [2:0] _T_234 = _T_233 & 3'h1; // @[dbg.scala 224:62]
  wire [2:0] _T_236 = abstractcs_error_sel1 ? 3'h7 : 3'h0; // @[Bitwise.scala 72:12]
  wire [2:0] _T_237 = _T_236 & 3'h2; // @[dbg.scala 225:37]
  wire [2:0] _T_238 = _T_234 | _T_237; // @[dbg.scala 224:79]
  wire [2:0] _T_240 = abstractcs_error_sel2 ? 3'h7 : 3'h0; // @[Bitwise.scala 72:12]
  wire [2:0] _T_241 = _T_240 & 3'h3; // @[dbg.scala 226:37]
  wire [2:0] _T_242 = _T_238 | _T_241; // @[dbg.scala 225:54]
  wire [2:0] _T_244 = abstractcs_error_sel3 ? 3'h7 : 3'h0; // @[Bitwise.scala 72:12]
  wire [2:0] _T_245 = _T_244 & 3'h4; // @[dbg.scala 227:37]
  wire [2:0] _T_246 = _T_242 | _T_245; // @[dbg.scala 226:54]
  wire [2:0] _T_248 = abstractcs_error_sel4 ? 3'h7 : 3'h0; // @[Bitwise.scala 72:12]
  wire [2:0] _T_250 = _T_246 | _T_248; // @[dbg.scala 227:54]
  wire [2:0] _T_252 = abstractcs_error_sel5 ? 3'h7 : 3'h0; // @[Bitwise.scala 72:12]
  wire [2:0] _T_254 = ~io_dmi_reg_wdata[10:8]; // @[dbg.scala 229:40]
  wire [2:0] _T_255 = _T_252 & _T_254; // @[dbg.scala 229:37]
  wire [2:0] _T_257 = _T_255 & abstractcs_reg[10:8]; // @[dbg.scala 229:75]
  wire [2:0] _T_258 = _T_250 | _T_257; // @[dbg.scala 228:54]
  wire  _T_259 = ~abstractcs_error_selor; // @[dbg.scala 230:15]
  wire [2:0] _T_261 = _T_259 ? 3'h7 : 3'h0; // @[Bitwise.scala 72:12]
  wire [2:0] _T_263 = _T_261 & abstractcs_reg[10:8]; // @[dbg.scala 230:50]
  reg  abs_temp_12; // @[Reg.scala 27:20]
  reg [2:0] abs_temp_10_8; // @[dbg.scala 237:12]
  wire [10:0] _T_265 = {abs_temp_10_8,8'h2}; // @[Cat.scala 29:58]
  wire [20:0] _T_267 = {19'h0,abs_temp_12,1'h0}; // @[Cat.scala 29:58]
  wire  _T_272 = dbg_state == 3'h2; // @[dbg.scala 242:100]
  wire  command_wren = _T_217 & _T_272; // @[dbg.scala 242:87]
  wire [19:0] _T_276 = {3'h0,io_dmi_reg_wdata[16:0]}; // @[Cat.scala 29:58]
  wire [11:0] _T_278 = {io_dmi_reg_wdata[31:24],1'h0,io_dmi_reg_wdata[22:20]}; // @[Cat.scala 29:58]
  wire  rvclkhdr_5_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_5_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_5_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_5_io_scan_mode; // @[lib.scala 368:23]
  reg [31:0] command_reg; // @[lib.scala 374:16]
  wire  _T_281 = _T_83 & _T_199; // @[dbg.scala 248:58]
  wire  data0_reg_wren0 = _T_281 & _T_272; // @[dbg.scala 248:89]
  wire  _T_283 = dbg_state == 3'h4; // @[dbg.scala 249:59]
  wire  _T_284 = io_core_dbg_cmd_done & _T_283; // @[dbg.scala 249:46]
  wire  _T_286 = ~command_reg[16]; // @[dbg.scala 249:83]
  wire  data0_reg_wren1 = _T_284 & _T_286; // @[dbg.scala 249:81]
  wire [31:0] _T_288 = data0_reg_wren0 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_289 = _T_288 & io_dmi_reg_wdata; // @[dbg.scala 252:45]
  wire [31:0] _T_291 = data0_reg_wren1 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_292 = _T_291 & io_core_dbg_rddata; // @[dbg.scala 252:92]
  wire  rvclkhdr_6_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_6_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_6_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_6_io_scan_mode; // @[lib.scala 368:23]
  reg [31:0] data0_reg; // @[lib.scala 374:16]
  wire  _T_294 = io_dmi_reg_addr == 7'h5; // @[dbg.scala 257:77]
  wire  _T_295 = _T_83 & _T_294; // @[dbg.scala 257:58]
  wire  data1_reg_wren = _T_295 & _T_272; // @[dbg.scala 257:89]
  wire [31:0] _T_298 = data1_reg_wren ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire  rvclkhdr_7_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_7_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_7_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_7_io_scan_mode; // @[lib.scala 368:23]
  reg [31:0] _T_299; // @[lib.scala 374:16]
  wire [2:0] dbg_nxtstate;
  wire  _T_300 = 3'h0 == dbg_state; // @[Conditional.scala 37:30]
  wire  _T_302 = dmstatus_reg[9] | io_dec_tlu_mpc_halted_only; // @[dbg.scala 272:43]
  wire [2:0] _T_303 = _T_302 ? 3'h2 : 3'h1; // @[dbg.scala 272:26]
  wire  _T_305 = ~io_dec_tlu_debug_mode; // @[dbg.scala 273:45]
  wire  _T_306 = dmcontrol_reg[31] & _T_305; // @[dbg.scala 273:43]
  wire  _T_308 = _T_306 | dmstatus_reg[9]; // @[dbg.scala 273:69]
  wire  _T_309 = _T_308 | io_dec_tlu_mpc_halted_only; // @[dbg.scala 273:87]
  wire  _T_312 = _T_309 & _T_17; // @[dbg.scala 273:117]
  wire  _T_316 = dmcontrol_reg[31] & _T_17; // @[dbg.scala 274:45]
  wire  _T_318 = 3'h1 == dbg_state; // @[Conditional.scala 37:30]
  wire [2:0] _T_320 = dmcontrol_reg[1] ? 3'h0 : 3'h2; // @[dbg.scala 277:26]
  wire  _T_323 = dmstatus_reg[9] | dmcontrol_reg[1]; // @[dbg.scala 278:39]
  wire  _T_325 = dmcontrol_wren_Q & dmcontrol_reg[31]; // @[dbg.scala 279:44]
  wire  _T_328 = _T_325 & _T_17; // @[dbg.scala 279:64]
  wire  _T_330 = 3'h2 == dbg_state; // @[Conditional.scala 37:30]
  wire  _T_334 = dmstatus_reg[9] & _T_17; // @[dbg.scala 282:43]
  wire  _T_337 = ~dmcontrol_reg[31]; // @[dbg.scala 283:33]
  wire  _T_338 = dmcontrol_reg[30] & _T_337; // @[dbg.scala 283:31]
  wire [2:0] _T_339 = _T_338 ? 3'h6 : 3'h3; // @[dbg.scala 283:12]
  wire [2:0] _T_341 = dmcontrol_reg[31] ? 3'h1 : 3'h0; // @[dbg.scala 284:12]
  wire [2:0] _T_342 = _T_334 ? _T_339 : _T_341; // @[dbg.scala 282:26]
  wire  _T_345 = dmstatus_reg[9] & dmcontrol_reg[30]; // @[dbg.scala 285:39]
  wire  _T_348 = _T_345 & _T_337; // @[dbg.scala 285:59]
  wire  _T_349 = _T_348 & dmcontrol_wren_Q; // @[dbg.scala 285:80]
  wire  _T_350 = _T_349 | command_wren; // @[dbg.scala 285:99]
  wire  _T_352 = _T_350 | dmcontrol_reg[1]; // @[dbg.scala 285:114]
  wire  _T_355 = ~_T_302; // @[dbg.scala 286:28]
  wire  _T_356 = _T_352 | _T_355; // @[dbg.scala 286:26]
  wire  _T_357 = dbg_nxtstate == 3'h3; // @[dbg.scala 287:60]
  wire  _T_358 = dbg_state_en & _T_357; // @[dbg.scala 287:44]
  wire  _T_359 = dbg_nxtstate == 3'h6; // @[dbg.scala 289:58]
  wire  _T_360 = dbg_state_en & _T_359; // @[dbg.scala 289:42]
  wire  _T_368 = 3'h3 == dbg_state; // @[Conditional.scala 37:30]
  wire  _T_371 = |abstractcs_reg[10:8]; // @[dbg.scala 293:85]
  wire [2:0] _T_372 = _T_371 ? 3'h5 : 3'h4; // @[dbg.scala 293:62]
  wire [2:0] _T_373 = dmcontrol_reg[1] ? 3'h0 : _T_372; // @[dbg.scala 293:26]
  wire  _T_376 = io_dbg_dec_dbg_ib_dbg_cmd_valid | _T_371; // @[dbg.scala 294:55]
  wire  _T_378 = _T_376 | dmcontrol_reg[1]; // @[dbg.scala 294:83]
  wire  _T_385 = 3'h4 == dbg_state; // @[Conditional.scala 37:30]
  wire [2:0] _T_387 = dmcontrol_reg[1] ? 3'h0 : 3'h5; // @[dbg.scala 298:26]
  wire  _T_389 = io_core_dbg_cmd_done | dmcontrol_reg[1]; // @[dbg.scala 299:44]
  wire  _T_396 = 3'h5 == dbg_state; // @[Conditional.scala 37:30]
  wire  _T_405 = 3'h6 == dbg_state; // @[Conditional.scala 37:30]
  wire  _T_408 = dmstatus_reg[17] | dmcontrol_reg[1]; // @[dbg.scala 311:40]
  wire  _GEN_10 = _T_405 & _T_408; // @[Conditional.scala 39:67]
  wire  _GEN_11 = _T_405 & _T_328; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_12 = _T_396 ? _T_320 : 3'h0; // @[Conditional.scala 39:67]
  wire  _GEN_13 = _T_396 | _GEN_10; // @[Conditional.scala 39:67]
  wire  _GEN_14 = _T_396 & dbg_state_en; // @[Conditional.scala 39:67]
  wire  _GEN_16 = _T_396 ? _T_328 : _GEN_11; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_17 = _T_385 ? _T_387 : _GEN_12; // @[Conditional.scala 39:67]
  wire  _GEN_18 = _T_385 ? _T_389 : _GEN_13; // @[Conditional.scala 39:67]
  wire  _GEN_19 = _T_385 ? _T_328 : _GEN_16; // @[Conditional.scala 39:67]
  wire  _GEN_20 = _T_385 ? 1'h0 : _GEN_14; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_22 = _T_368 ? _T_373 : _GEN_17; // @[Conditional.scala 39:67]
  wire  _GEN_23 = _T_368 ? _T_378 : _GEN_18; // @[Conditional.scala 39:67]
  wire  _GEN_24 = _T_368 ? _T_328 : _GEN_19; // @[Conditional.scala 39:67]
  wire  _GEN_25 = _T_368 ? 1'h0 : _GEN_20; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_27 = _T_330 ? _T_342 : _GEN_22; // @[Conditional.scala 39:67]
  wire  _GEN_28 = _T_330 ? _T_356 : _GEN_23; // @[Conditional.scala 39:67]
  wire  _GEN_29 = _T_330 ? _T_358 : _GEN_25; // @[Conditional.scala 39:67]
  wire  _GEN_31 = _T_330 & _T_360; // @[Conditional.scala 39:67]
  wire  _GEN_32 = _T_330 ? _T_328 : _GEN_24; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_33 = _T_318 ? _T_320 : _GEN_27; // @[Conditional.scala 39:67]
  wire  _GEN_34 = _T_318 ? _T_323 : _GEN_28; // @[Conditional.scala 39:67]
  wire  _GEN_35 = _T_318 ? _T_328 : _GEN_32; // @[Conditional.scala 39:67]
  wire  _GEN_36 = _T_318 ? 1'h0 : _GEN_29; // @[Conditional.scala 39:67]
  wire  _GEN_38 = _T_318 ? 1'h0 : _GEN_31; // @[Conditional.scala 39:67]
  reg [2:0] _T_468; // @[Reg.scala 27:20]
  wire  _T_471 = command_reg[31:24] == 8'h2; // @[dbg.scala 331:62]
  wire [31:0] _T_473 = {data1_reg[31:2],2'h0}; // @[Cat.scala 29:58]
  wire [31:0] _T_475 = {20'h0,command_reg[11:0]}; // @[Cat.scala 29:58]
  wire  _T_478 = dbg_state == 3'h3; // @[dbg.scala 333:50]
  wire  _T_481 = ~_T_371; // @[dbg.scala 333:75]
  wire  _T_482 = _T_478 & _T_481; // @[dbg.scala 333:73]
  wire  _T_490 = command_reg[15:12] == 4'h0; // @[dbg.scala 335:122]
  wire [1:0] _T_491 = {1'h0,_T_490}; // @[Cat.scala 29:58]
  wire  _T_502 = 4'h0 == sb_state; // @[Conditional.scala 37:30]
  wire  _T_504 = sbdata0_reg_wren0 | sbreadondata_access; // @[dbg.scala 350:39]
  wire  _T_505 = _T_504 | sbreadonaddr_access; // @[dbg.scala 350:61]
  wire  _T_507 = |io_dmi_reg_wdata[14:12]; // @[dbg.scala 353:65]
  wire  _T_508 = sbcs_wren & _T_507; // @[dbg.scala 353:38]
  wire [2:0] _T_510 = ~io_dmi_reg_wdata[14:12]; // @[dbg.scala 354:27]
  wire [2:0] _T_512 = _T_510 & sbcs_reg[14:12]; // @[dbg.scala 354:53]
  wire  _T_513 = 4'h1 == sb_state; // @[Conditional.scala 37:30]
  wire  _T_514 = sbcs_unaligned | sbcs_illegal_size; // @[dbg.scala 357:41]
  wire  _T_516 = io_dbg_bus_clk_en | sbcs_unaligned; // @[dbg.scala 358:40]
  wire  _T_517 = _T_516 | sbcs_illegal_size; // @[dbg.scala 358:57]
  wire  _T_520 = 4'h2 == sb_state; // @[Conditional.scala 37:30]
  wire  _T_527 = 4'h3 == sb_state; // @[Conditional.scala 37:30]
  wire  _T_529 = 4'h4 == sb_state; // @[Conditional.scala 37:30]
  wire  _T_535 = 4'h5 == sb_state; // @[Conditional.scala 37:30]
  wire  _T_537 = 4'h6 == sb_state; // @[Conditional.scala 37:30]
  wire  _T_539 = 4'h7 == sb_state; // @[Conditional.scala 37:30]
  wire  _T_542 = 4'h8 == sb_state; // @[Conditional.scala 37:30]
  wire  _T_545 = 4'h9 == sb_state; // @[Conditional.scala 37:30]
  wire  _GEN_50 = _T_545 & sbcs_reg[16]; // @[Conditional.scala 39:67]
  wire  _GEN_52 = _T_542 ? 1'h0 : _T_545; // @[Conditional.scala 39:67]
  wire  _GEN_57 = _T_542 ? 1'h0 : _GEN_50; // @[Conditional.scala 39:67]
  wire  _GEN_59 = _T_539 ? 1'h0 : _GEN_52; // @[Conditional.scala 39:67]
  wire  _GEN_64 = _T_539 ? 1'h0 : _GEN_57; // @[Conditional.scala 39:67]
  wire  _GEN_66 = _T_537 ? 1'h0 : _GEN_59; // @[Conditional.scala 39:67]
  wire  _GEN_71 = _T_537 ? 1'h0 : _GEN_64; // @[Conditional.scala 39:67]
  wire  _GEN_73 = _T_535 ? 1'h0 : _GEN_66; // @[Conditional.scala 39:67]
  wire  _GEN_78 = _T_535 ? 1'h0 : _GEN_71; // @[Conditional.scala 39:67]
  wire  _GEN_80 = _T_529 ? 1'h0 : _GEN_73; // @[Conditional.scala 39:67]
  wire  _GEN_85 = _T_529 ? 1'h0 : _GEN_78; // @[Conditional.scala 39:67]
  wire  _GEN_87 = _T_527 ? 1'h0 : _GEN_80; // @[Conditional.scala 39:67]
  wire  _GEN_92 = _T_527 ? 1'h0 : _GEN_85; // @[Conditional.scala 39:67]
  wire  _GEN_94 = _T_520 ? _T_517 : _GEN_87; // @[Conditional.scala 39:67]
  wire  _GEN_95 = _T_520 & _T_514; // @[Conditional.scala 39:67]
  wire  _GEN_97 = _T_520 ? 1'h0 : _GEN_87; // @[Conditional.scala 39:67]
  wire  _GEN_99 = _T_520 ? 1'h0 : _GEN_92; // @[Conditional.scala 39:67]
  wire  _GEN_101 = _T_513 ? _T_517 : _GEN_94; // @[Conditional.scala 39:67]
  wire  _GEN_102 = _T_513 ? _T_514 : _GEN_95; // @[Conditional.scala 39:67]
  wire  _GEN_104 = _T_513 ? 1'h0 : _GEN_97; // @[Conditional.scala 39:67]
  wire  _GEN_106 = _T_513 ? 1'h0 : _GEN_99; // @[Conditional.scala 39:67]
  reg [3:0] _T_547; // @[Reg.scala 27:20]
  wire  _T_560 = sb_state == 4'h4; // @[dbg.scala 414:36]
  wire  _T_561 = sb_state == 4'h5; // @[dbg.scala 414:71]
  wire  _T_567 = sb_state == 4'h6; // @[dbg.scala 425:70]
  wire [7:0] _T_608 = _T_62 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [14:0] _T_610 = 15'h1 << sbaddress0_reg[2:0]; // @[dbg.scala 429:82]
  wire [14:0] _GEN_115 = {{7'd0}, _T_608}; // @[dbg.scala 429:67]
  wire [14:0] _T_611 = _GEN_115 & _T_610; // @[dbg.scala 429:67]
  wire [7:0] _T_615 = _T_47 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [2:0] _T_617 = {sbaddress0_reg[2:1],1'h0}; // @[Cat.scala 29:58]
  wire [14:0] _T_618 = 15'h3 << _T_617; // @[dbg.scala 430:59]
  wire [14:0] _GEN_116 = {{7'd0}, _T_615}; // @[dbg.scala 430:44]
  wire [14:0] _T_619 = _GEN_116 & _T_618; // @[dbg.scala 430:44]
  wire [14:0] _T_620 = _T_611 | _T_619; // @[dbg.scala 429:107]
  wire [7:0] _T_624 = _T_51 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [2:0] _T_626 = {sbaddress0_reg[2],2'h0}; // @[Cat.scala 29:58]
  wire [14:0] _T_627 = 15'hf << _T_626; // @[dbg.scala 431:59]
  wire [14:0] _GEN_117 = {{7'd0}, _T_624}; // @[dbg.scala 431:44]
  wire [14:0] _T_628 = _GEN_117 & _T_627; // @[dbg.scala 431:44]
  wire [14:0] _T_629 = _T_620 | _T_628; // @[dbg.scala 430:97]
  wire [7:0] _T_633 = _T_57 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [14:0] _GEN_118 = {{7'd0}, _T_633}; // @[dbg.scala 431:100]
  wire [14:0] _T_635 = _T_629 | _GEN_118; // @[dbg.scala 431:100]
  rvclkhdr rvclkhdr ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_io_l1clk),
    .io_clk(rvclkhdr_io_clk),
    .io_en(rvclkhdr_io_en),
    .io_scan_mode(rvclkhdr_io_scan_mode)
  );
  rvclkhdr rvclkhdr_1 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_1_io_l1clk),
    .io_clk(rvclkhdr_1_io_clk),
    .io_en(rvclkhdr_1_io_en),
    .io_scan_mode(rvclkhdr_1_io_scan_mode)
  );
  rvclkhdr rvclkhdr_2 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_2_io_l1clk),
    .io_clk(rvclkhdr_2_io_clk),
    .io_en(rvclkhdr_2_io_en),
    .io_scan_mode(rvclkhdr_2_io_scan_mode)
  );
  rvclkhdr rvclkhdr_3 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_3_io_l1clk),
    .io_clk(rvclkhdr_3_io_clk),
    .io_en(rvclkhdr_3_io_en),
    .io_scan_mode(rvclkhdr_3_io_scan_mode)
  );
  rvclkhdr rvclkhdr_4 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_4_io_l1clk),
    .io_clk(rvclkhdr_4_io_clk),
    .io_en(rvclkhdr_4_io_en),
    .io_scan_mode(rvclkhdr_4_io_scan_mode)
  );
  rvclkhdr rvclkhdr_5 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_5_io_l1clk),
    .io_clk(rvclkhdr_5_io_clk),
    .io_en(rvclkhdr_5_io_en),
    .io_scan_mode(rvclkhdr_5_io_scan_mode)
  );
  rvclkhdr rvclkhdr_6 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_6_io_l1clk),
    .io_clk(rvclkhdr_6_io_clk),
    .io_en(rvclkhdr_6_io_en),
    .io_scan_mode(rvclkhdr_6_io_scan_mode)
  );
  rvclkhdr rvclkhdr_7 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_7_io_l1clk),
    .io_clk(rvclkhdr_7_io_clk),
    .io_en(rvclkhdr_7_io_en),
    .io_scan_mode(rvclkhdr_7_io_scan_mode)
  );
  assign io_dbg_cmd_size = command_reg[21:20]; // @[dbg.scala 336:19]
  assign io_dbg_core_rst_l = ~dmcontrol_reg[1]; // @[dbg.scala 107:21]
  assign io_dbg_halt_req = _T_300 ? _T_316 : _GEN_35; // @[dbg.scala 268:19 dbg.scala 274:23 dbg.scala 279:23 dbg.scala 290:23 dbg.scala 295:23 dbg.scala 300:23 dbg.scala 307:23 dbg.scala 312:23]
  assign io_dbg_resume_req = _T_300 ? 1'h0 : _GEN_38; // @[dbg.scala 269:21 dbg.scala 289:25]
  assign io_sb_axi_aw_valid = _T_560 | _T_561; // @[dbg.scala 414:22]
  assign io_sb_axi_aw_bits_addr = sbaddress0_reg; // @[dbg.scala 415:26]
  assign io_sb_axi_aw_bits_size = sbcs_reg[19:17]; // @[dbg.scala 417:26]
  assign io_sb_axi_w_valid = _T_560 | _T_567; // @[dbg.scala 425:21]
  assign io_sb_axi_w_bits_strb = _T_635[7:0]; // @[dbg.scala 429:25]
  assign io_sb_axi_ar_valid = sb_state == 4'h3; // @[dbg.scala 435:22]
  assign io_sb_axi_ar_bits_addr = sbaddress0_reg; // @[dbg.scala 436:26]
  assign io_sb_axi_ar_bits_size = sbcs_reg[19:17]; // @[dbg.scala 438:26]
  assign io_dbg_dec_dbg_ib_dbg_cmd_valid = _T_482 & io_dbg_dma_io_dma_dbg_ready; // @[dbg.scala 333:35]
  assign io_dbg_dec_dbg_ib_dbg_cmd_write = command_reg[16]; // @[dbg.scala 334:35]
  assign io_dbg_dec_dbg_ib_dbg_cmd_type = _T_471 ? 2'h2 : _T_491; // @[dbg.scala 335:34]
  assign io_dbg_dec_dbg_ib_dbg_cmd_addr = _T_471 ? _T_473 : _T_475; // @[dbg.scala 331:34]
  assign io_dbg_dec_dbg_dctl_dbg_cmd_wrdata = data0_reg; // @[dbg.scala 332:38]
  assign io_dbg_dma_dbg_ib_dbg_cmd_valid = io_dbg_dec_dbg_ib_dbg_cmd_valid; // @[dbg.scala 456:39]
  assign io_dbg_dma_dbg_ib_dbg_cmd_write = io_dbg_dec_dbg_ib_dbg_cmd_write; // @[dbg.scala 457:39]
  assign io_dbg_dma_dbg_ib_dbg_cmd_type = io_dbg_dec_dbg_ib_dbg_cmd_type; // @[dbg.scala 458:39]
  assign io_dbg_dma_dbg_ib_dbg_cmd_addr = io_dbg_dec_dbg_ib_dbg_cmd_addr; // @[dbg.scala 454:39]
  assign io_dbg_dma_dbg_dctl_dbg_cmd_wrdata = io_dbg_dec_dbg_dctl_dbg_cmd_wrdata; // @[dbg.scala 455:39]
  assign io_dbg_dma_io_dbg_dma_bubble = _T_482 | _T_283; // @[dbg.scala 337:32]
  assign dbg_state = _T_468; // @[dbg.scala 322:13]
  assign dbg_state_en = _T_300 ? _T_312 : _GEN_34; // @[dbg.scala 265:16 dbg.scala 273:20 dbg.scala 278:20 dbg.scala 285:20 dbg.scala 294:20 dbg.scala 299:20 dbg.scala 304:20 dbg.scala 311:20]
  assign sb_state = _T_547; // @[dbg.scala 404:12]
  assign sb_state_en = _T_502 ? _T_505 : _GEN_101; // @[dbg.scala 350:19 dbg.scala 358:19 dbg.scala 364:19 dbg.scala 370:19 dbg.scala 374:19 dbg.scala 378:19 dbg.scala 382:19 dbg.scala 386:19 dbg.scala 392:19 dbg.scala 398:19]
  assign dmcontrol_reg = {_T_145,_T_143}; // @[dbg.scala 185:17]
  assign sbaddress0_reg = _T_118; // @[dbg.scala 166:18]
  assign sbcs_sbbusy_wren = _T_502 ? sb_state_en : _GEN_104; // @[dbg.scala 342:20 dbg.scala 351:24 dbg.scala 399:24]
  assign sbcs_sberror_wren = _T_502 ? _T_508 : _GEN_102; // @[dbg.scala 344:21 dbg.scala 353:25 dbg.scala 359:25 dbg.scala 365:25 dbg.scala 387:25 dbg.scala 393:25]
  assign sbaddress0_reg_wren1 = _T_502 ? 1'h0 : _GEN_106; // @[dbg.scala 346:24 dbg.scala 401:28]
  assign dmstatus_reg = {_T_163,_T_159}; // @[dbg.scala 191:16]
  assign dmstatus_havereset = _T_192; // @[dbg.scala 208:22]
  assign dmstatus_resumeack = _T_185; // @[dbg.scala 200:22]
  assign dmstatus_unavail = dmcontrol_reg[1] | _T_180; // @[dbg.scala 198:20]
  assign dmstatus_running = ~_T_183; // @[dbg.scala 199:20]
  assign dmstatus_halted = _T_188; // @[dbg.scala 204:19]
  assign abstractcs_busy_wren = _T_300 ? 1'h0 : _GEN_36; // @[dbg.scala 266:24 dbg.scala 287:28 dbg.scala 305:28]
  assign sbcs_sbbusy_din = 4'h0 == sb_state; // @[dbg.scala 343:19 dbg.scala 352:23 dbg.scala 400:23]
  assign data1_reg = _T_299; // @[dbg.scala 259:13]
  assign sbcs_reg = {_T_44,_T_40}; // @[dbg.scala 132:12]
  assign rvclkhdr_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_io_en = _T_3 | io_clk_override; // @[lib.scala 345:16]
  assign rvclkhdr_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_1_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_1_io_en = _T_6 | io_clk_override; // @[lib.scala 345:16]
  assign rvclkhdr_1_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_2_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_2_io_en = sbdata0_reg_wren0 | sbdata0_reg_wren1; // @[lib.scala 371:17]
  assign rvclkhdr_2_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_3_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_3_io_en = sbdata1_reg_wren0 | sbdata0_reg_wren1; // @[lib.scala 371:17]
  assign rvclkhdr_3_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_4_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_4_io_en = sbaddress0_reg_wren0 | sbaddress0_reg_wren1; // @[lib.scala 371:17]
  assign rvclkhdr_4_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign abstractcs_reg = {_T_267,_T_265}; // @[dbg.scala 240:18]
  assign rvclkhdr_5_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_5_io_en = _T_217 & _T_272; // @[lib.scala 371:17]
  assign rvclkhdr_5_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_6_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_6_io_en = data0_reg_wren0 | data0_reg_wren1; // @[lib.scala 371:17]
  assign rvclkhdr_6_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_7_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_7_io_en = _T_295 & _T_272; // @[lib.scala 371:17]
  assign rvclkhdr_7_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign dbg_nxtstate = _T_300 ? _T_303 : _GEN_33; // @[dbg.scala 264:16 dbg.scala 272:20 dbg.scala 277:20 dbg.scala 282:20 dbg.scala 293:20 dbg.scala 298:20 dbg.scala 303:20 dbg.scala 310:20]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  temp_sbcs_22 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  temp_sbcs_21 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  temp_sbcs_20 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  temp_sbcs_19_15 = _RAND_3[4:0];
  _RAND_4 = {1{`RANDOM}};
  temp_sbcs_14_12 = _RAND_4[2:0];
  _RAND_5 = {1{`RANDOM}};
  _T_118 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  dm_temp = _RAND_6[3:0];
  _RAND_7 = {1{`RANDOM}};
  dm_temp_0 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  dmcontrol_wren_Q = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  _T_185 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  _T_188 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  _T_192 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  abs_temp_12 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  abs_temp_10_8 = _RAND_13[2:0];
  _RAND_14 = {1{`RANDOM}};
  command_reg = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  data0_reg = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  _T_299 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  _T_468 = _RAND_17[2:0];
  _RAND_18 = {1{`RANDOM}};
  _T_547 = _RAND_18[3:0];
`endif // RANDOMIZE_REG_INIT
  if (dbg_dm_rst_l) begin
    temp_sbcs_22 = 1'h0;
  end
  if (dbg_dm_rst_l) begin
    temp_sbcs_21 = 1'h0;
  end
  if (dbg_dm_rst_l) begin
    temp_sbcs_20 = 1'h0;
  end
  if (dbg_dm_rst_l) begin
    temp_sbcs_19_15 = 5'h0;
  end
  if (rst_not) begin
    temp_sbcs_14_12 = 3'h0;
  end
  if (dbg_dm_rst_l) begin
    _T_118 = 32'h0;
  end
  if (dbg_dm_rst_l) begin
    dm_temp = 4'h0;
  end
  if (io_dbg_rst_l) begin
    dm_temp_0 = 1'h0;
  end
  if (dbg_dm_rst_l) begin
    dmcontrol_wren_Q = 1'h0;
  end
  if (dbg_dm_rst_l) begin
    _T_185 = 1'h0;
  end
  if (dbg_dm_rst_l) begin
    _T_188 = 1'h0;
  end
  if (dbg_dm_rst_l) begin
    _T_192 = 1'h0;
  end
  if (dbg_dm_rst_l) begin
    abs_temp_12 = 1'h0;
  end
  if (dbg_dm_rst_l) begin
    abs_temp_10_8 = 3'h0;
  end
  if (dbg_dm_rst_l) begin
    command_reg = 32'h0;
  end
  if (dbg_dm_rst_l) begin
    data0_reg = 32'h0;
  end
  if (dbg_dm_rst_l) begin
    _T_299 = 32'h0;
  end
  if (rst_temp) begin
    _T_468 = 3'h0;
  end
  if (dbg_dm_rst_l) begin
    _T_547 = 4'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge rvclkhdr_1_io_l1clk or posedge dbg_dm_rst_l) begin
    if (dbg_dm_rst_l) begin
      temp_sbcs_22 <= 1'h0;
    end else if (sbcs_sbbusyerror_wren) begin
      temp_sbcs_22 <= sbcs_sbbusyerror_din;
    end
  end
  always @(posedge rvclkhdr_1_io_l1clk or posedge dbg_dm_rst_l) begin
    if (dbg_dm_rst_l) begin
      temp_sbcs_21 <= 1'h0;
    end else if (sbcs_sbbusy_wren) begin
      temp_sbcs_21 <= sbcs_sbbusy_din;
    end
  end
  always @(posedge rvclkhdr_1_io_l1clk or posedge dbg_dm_rst_l) begin
    if (dbg_dm_rst_l) begin
      temp_sbcs_20 <= 1'h0;
    end else if (sbcs_wren) begin
      temp_sbcs_20 <= io_dmi_reg_wdata[20];
    end
  end
  always @(posedge rvclkhdr_1_io_l1clk or posedge dbg_dm_rst_l) begin
    if (dbg_dm_rst_l) begin
      temp_sbcs_19_15 <= 5'h0;
    end else if (sbcs_wren) begin
      temp_sbcs_19_15 <= io_dmi_reg_wdata[19:15];
    end
  end
  always @(posedge rvclkhdr_1_io_l1clk or posedge rst_not) begin
    if (rst_not) begin
      temp_sbcs_14_12 <= 3'h0;
    end else if (sbcs_sberror_wren) begin
      if (_T_502) begin
        temp_sbcs_14_12 <= _T_512;
      end else if (_T_513) begin
        if (sbcs_unaligned) begin
          temp_sbcs_14_12 <= 3'h3;
        end else begin
          temp_sbcs_14_12 <= 3'h4;
        end
      end else if (_T_520) begin
        if (sbcs_unaligned) begin
          temp_sbcs_14_12 <= 3'h3;
        end else begin
          temp_sbcs_14_12 <= 3'h4;
        end
      end else if (_T_527) begin
        temp_sbcs_14_12 <= 3'h0;
      end else if (_T_529) begin
        temp_sbcs_14_12 <= 3'h0;
      end else if (_T_535) begin
        temp_sbcs_14_12 <= 3'h0;
      end else if (_T_537) begin
        temp_sbcs_14_12 <= 3'h0;
      end else if (_T_539) begin
        temp_sbcs_14_12 <= 3'h2;
      end else if (_T_542) begin
        temp_sbcs_14_12 <= 3'h2;
      end else begin
        temp_sbcs_14_12 <= 3'h0;
      end
    end
  end
  always @(posedge rvclkhdr_4_io_l1clk or posedge dbg_dm_rst_l) begin
    if (dbg_dm_rst_l) begin
      _T_118 <= 32'h0;
    end else begin
      _T_118 <= _T_111 | _T_117;
    end
  end
  always @(posedge rvclkhdr_io_l1clk or posedge dbg_dm_rst_l) begin
    if (dbg_dm_rst_l) begin
      dm_temp <= 4'h0;
    end else if (dmcontrol_wren) begin
      dm_temp <= _T_136;
    end
  end
  always @(posedge rvclkhdr_io_l1clk or posedge io_dbg_rst_l) begin
    if (io_dbg_rst_l) begin
      dm_temp_0 <= 1'h0;
    end else if (dmcontrol_wren) begin
      dm_temp_0 <= io_dmi_reg_wdata[0];
    end
  end
  always @(posedge rvclkhdr_io_l1clk or posedge dbg_dm_rst_l) begin
    if (dbg_dm_rst_l) begin
      dmcontrol_wren_Q <= 1'h0;
    end else begin
      dmcontrol_wren_Q <= _T_131 & io_dmi_reg_wr_en;
    end
  end
  always @(posedge rvclkhdr_io_l1clk or posedge dbg_dm_rst_l) begin
    if (dbg_dm_rst_l) begin
      _T_185 <= 1'h0;
    end else if (dmstatus_resumeack_wren) begin
      _T_185 <= _T_166;
    end
  end
  always @(posedge rvclkhdr_io_l1clk or posedge dbg_dm_rst_l) begin
    if (dbg_dm_rst_l) begin
      _T_188 <= 1'h0;
    end else begin
      _T_188 <= io_dec_tlu_dbg_halted & _T_186;
    end
  end
  always @(posedge rvclkhdr_io_l1clk or posedge dbg_dm_rst_l) begin
    if (dbg_dm_rst_l) begin
      _T_192 <= 1'h0;
    end else begin
      _T_192 <= _T_189 & _T_190;
    end
  end
  always @(posedge rvclkhdr_io_l1clk or posedge dbg_dm_rst_l) begin
    if (dbg_dm_rst_l) begin
      abs_temp_12 <= 1'h0;
    end else if (abstractcs_busy_wren) begin
      if (_T_300) begin
        abs_temp_12 <= 1'h0;
      end else if (_T_318) begin
        abs_temp_12 <= 1'h0;
      end else begin
        abs_temp_12 <= _T_330;
      end
    end
  end
  always @(posedge rvclkhdr_io_l1clk or posedge dbg_dm_rst_l) begin
    if (dbg_dm_rst_l) begin
      abs_temp_10_8 <= 3'h0;
    end else begin
      abs_temp_10_8 <= _T_258 | _T_263;
    end
  end
  always @(posedge rvclkhdr_5_io_l1clk or posedge dbg_dm_rst_l) begin
    if (dbg_dm_rst_l) begin
      command_reg <= 32'h0;
    end else begin
      command_reg <= {_T_278,_T_276};
    end
  end
  always @(posedge rvclkhdr_6_io_l1clk or posedge dbg_dm_rst_l) begin
    if (dbg_dm_rst_l) begin
      data0_reg <= 32'h0;
    end else begin
      data0_reg <= _T_289 | _T_292;
    end
  end
  always @(posedge rvclkhdr_7_io_l1clk or posedge dbg_dm_rst_l) begin
    if (dbg_dm_rst_l) begin
      _T_299 <= 32'h0;
    end else begin
      _T_299 <= _T_298 & io_dmi_reg_wdata;
    end
  end
  always @(posedge rvclkhdr_io_l1clk or posedge rst_temp) begin
    if (rst_temp) begin
      _T_468 <= 3'h0;
    end else if (dbg_state_en) begin
      if (_T_300) begin
        if (_T_302) begin
          _T_468 <= 3'h2;
        end else begin
          _T_468 <= 3'h1;
        end
      end else if (_T_318) begin
        if (dmcontrol_reg[1]) begin
          _T_468 <= 3'h0;
        end else begin
          _T_468 <= 3'h2;
        end
      end else if (_T_330) begin
        if (_T_334) begin
          if (_T_338) begin
            _T_468 <= 3'h6;
          end else begin
            _T_468 <= 3'h3;
          end
        end else if (dmcontrol_reg[31]) begin
          _T_468 <= 3'h1;
        end else begin
          _T_468 <= 3'h0;
        end
      end else if (_T_368) begin
        if (dmcontrol_reg[1]) begin
          _T_468 <= 3'h0;
        end else if (_T_371) begin
          _T_468 <= 3'h5;
        end else begin
          _T_468 <= 3'h4;
        end
      end else if (_T_385) begin
        if (dmcontrol_reg[1]) begin
          _T_468 <= 3'h0;
        end else begin
          _T_468 <= 3'h5;
        end
      end else if (_T_396) begin
        if (dmcontrol_reg[1]) begin
          _T_468 <= 3'h0;
        end else begin
          _T_468 <= 3'h2;
        end
      end else begin
        _T_468 <= 3'h0;
      end
    end
  end
  always @(posedge rvclkhdr_1_io_l1clk or posedge dbg_dm_rst_l) begin
    if (dbg_dm_rst_l) begin
      _T_547 <= 4'h0;
    end else if (sb_state_en) begin
      if (_T_502) begin
        if (sbdata0_reg_wren0) begin
          _T_547 <= 4'h2;
        end else begin
          _T_547 <= 4'h1;
        end
      end else if (_T_513) begin
        if (_T_514) begin
          _T_547 <= 4'h9;
        end else begin
          _T_547 <= 4'h3;
        end
      end else if (_T_520) begin
        if (_T_514) begin
          _T_547 <= 4'h9;
        end else begin
          _T_547 <= 4'h4;
        end
      end else if (_T_527) begin
        _T_547 <= 4'h7;
      end else if (_T_529) begin
        _T_547 <= 4'h6;
      end else if (_T_535) begin
        _T_547 <= 4'h8;
      end else if (_T_537) begin
        _T_547 <= 4'h8;
      end else if (_T_539) begin
        _T_547 <= 4'h9;
      end else if (_T_542) begin
        _T_547 <= 4'h9;
      end else begin
        _T_547 <= 4'h0;
      end
    end
  end
endmodule
module exu_alu_ctl(
  input         clock,
  input         reset,
  input         io_dec_alu_dec_i0_alu_decode_d,
  input         io_dec_alu_dec_csr_ren_d,
  input  [11:0] io_dec_alu_dec_i0_br_immed_d,
  output [30:0] io_dec_alu_exu_i0_pc_x,
  input  [30:0] io_dec_i0_pc_d,
  input         io_scan_mode,
  input         io_flush_upper_x,
  input         io_dec_tlu_flush_lower_r,
  input         io_enable,
  input         io_i0_ap_land,
  input         io_i0_ap_lor,
  input         io_i0_ap_lxor,
  input         io_i0_ap_sll,
  input         io_i0_ap_srl,
  input         io_i0_ap_sra,
  input         io_i0_ap_beq,
  input         io_i0_ap_bne,
  input         io_i0_ap_blt,
  input         io_i0_ap_bge,
  input         io_i0_ap_add,
  input         io_i0_ap_sub,
  input         io_i0_ap_slt,
  input         io_i0_ap_unsign,
  input         io_i0_ap_jal,
  input         io_i0_ap_predict_t,
  input         io_i0_ap_predict_nt,
  input         io_i0_ap_csr_write,
  input         io_i0_ap_csr_imm,
  input  [31:0] io_a_in,
  input  [31:0] io_b_in,
  input         io_pp_in_valid,
  input         io_pp_in_bits_boffset,
  input         io_pp_in_bits_pc4,
  input  [1:0]  io_pp_in_bits_hist,
  input  [11:0] io_pp_in_bits_toffset,
  input         io_pp_in_bits_br_error,
  input         io_pp_in_bits_br_start_error,
  input  [30:0] io_pp_in_bits_prett,
  input         io_pp_in_bits_pcall,
  input         io_pp_in_bits_pret,
  input         io_pp_in_bits_pja,
  input         io_pp_in_bits_way,
  output [31:0] io_result_ff,
  output        io_flush_upper_out,
  output        io_flush_final_out,
  output [30:0] io_flush_path_out,
  output        io_pred_correct_out,
  output        io_predict_p_out_valid,
  output        io_predict_p_out_bits_misp,
  output        io_predict_p_out_bits_ataken,
  output        io_predict_p_out_bits_boffset,
  output        io_predict_p_out_bits_pc4,
  output [1:0]  io_predict_p_out_bits_hist,
  output [11:0] io_predict_p_out_bits_toffset,
  output        io_predict_p_out_bits_br_error,
  output        io_predict_p_out_bits_br_start_error,
  output        io_predict_p_out_bits_pcall,
  output        io_predict_p_out_bits_pret,
  output        io_predict_p_out_bits_pja,
  output        io_predict_p_out_bits_way
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  rvclkhdr_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_1_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_1_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_1_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_1_io_scan_mode; // @[lib.scala 368:23]
  reg [30:0] _T_1; // @[lib.scala 374:16]
  reg [31:0] _T_3; // @[lib.scala 374:16]
  wire [31:0] _T_5 = ~io_b_in; // @[exu_alu_ctl.scala 34:40]
  wire [31:0] bm = io_i0_ap_sub ? _T_5 : io_b_in; // @[exu_alu_ctl.scala 34:17]
  wire [32:0] _T_8 = {1'h0,io_a_in}; // @[Cat.scala 29:58]
  wire [32:0] _T_10 = {1'h0,_T_5}; // @[Cat.scala 29:58]
  wire [32:0] _T_12 = _T_8 + _T_10; // @[exu_alu_ctl.scala 37:58]
  wire [32:0] _T_13 = {32'h0,io_i0_ap_sub}; // @[Cat.scala 29:58]
  wire [32:0] _T_15 = _T_12 + _T_13; // @[exu_alu_ctl.scala 37:83]
  wire [32:0] _T_18 = {1'h0,io_b_in}; // @[Cat.scala 29:58]
  wire [32:0] _T_20 = _T_8 + _T_18; // @[exu_alu_ctl.scala 37:138]
  wire [32:0] _T_23 = _T_20 + _T_13; // @[exu_alu_ctl.scala 37:163]
  wire [32:0] aout = io_i0_ap_sub ? _T_15 : _T_23; // @[exu_alu_ctl.scala 37:14]
  wire  cout = aout[32]; // @[exu_alu_ctl.scala 38:18]
  wire  _T_26 = ~io_a_in[31]; // @[exu_alu_ctl.scala 40:14]
  wire  _T_28 = ~bm[31]; // @[exu_alu_ctl.scala 40:29]
  wire  _T_29 = _T_26 & _T_28; // @[exu_alu_ctl.scala 40:27]
  wire  _T_31 = _T_29 & aout[31]; // @[exu_alu_ctl.scala 40:37]
  wire  _T_34 = io_a_in[31] & bm[31]; // @[exu_alu_ctl.scala 40:66]
  wire  _T_36 = ~aout[31]; // @[exu_alu_ctl.scala 40:78]
  wire  _T_37 = _T_34 & _T_36; // @[exu_alu_ctl.scala 40:76]
  wire  ov = _T_31 | _T_37; // @[exu_alu_ctl.scala 40:50]
  wire  eq = $signed(io_a_in) == $signed(io_b_in); // @[exu_alu_ctl.scala 42:38]
  wire  ne = ~eq; // @[exu_alu_ctl.scala 43:29]
  wire  _T_39 = ~io_i0_ap_unsign; // @[exu_alu_ctl.scala 45:30]
  wire  _T_40 = aout[31] ^ ov; // @[exu_alu_ctl.scala 45:54]
  wire  _T_41 = _T_39 & _T_40; // @[exu_alu_ctl.scala 45:47]
  wire  _T_42 = ~cout; // @[exu_alu_ctl.scala 45:84]
  wire  _T_43 = io_i0_ap_unsign & _T_42; // @[exu_alu_ctl.scala 45:82]
  wire  lt = _T_41 | _T_43; // @[exu_alu_ctl.scala 45:61]
  wire  ge = ~lt; // @[exu_alu_ctl.scala 46:29]
  wire [31:0] _T_63 = $signed(io_a_in) & $signed(io_b_in); // @[Mux.scala 27:72]
  wire [31:0] _T_66 = $signed(io_a_in) | $signed(io_b_in); // @[Mux.scala 27:72]
  wire [31:0] _T_69 = $signed(io_a_in) ^ $signed(io_b_in); // @[Mux.scala 27:72]
  wire [31:0] _T_70 = io_dec_alu_dec_csr_ren_d ? $signed(io_b_in) : $signed(32'sh0); // @[Mux.scala 27:72]
  wire [31:0] _T_71 = io_i0_ap_land ? $signed(_T_63) : $signed(32'sh0); // @[Mux.scala 27:72]
  wire [31:0] _T_72 = io_i0_ap_lor ? $signed(_T_66) : $signed(32'sh0); // @[Mux.scala 27:72]
  wire [31:0] _T_73 = io_i0_ap_lxor ? $signed(_T_69) : $signed(32'sh0); // @[Mux.scala 27:72]
  wire [31:0] _T_75 = $signed(_T_70) | $signed(_T_71); // @[Mux.scala 27:72]
  wire [31:0] _T_77 = $signed(_T_75) | $signed(_T_72); // @[Mux.scala 27:72]
  wire [5:0] _T_84 = {1'h0,io_b_in[4:0]}; // @[Cat.scala 29:58]
  wire [5:0] _T_86 = 6'h20 - _T_84; // @[exu_alu_ctl.scala 56:41]
  wire [5:0] _T_93 = io_i0_ap_sll ? _T_86 : 6'h0; // @[Mux.scala 27:72]
  wire [5:0] _T_94 = io_i0_ap_srl ? _T_84 : 6'h0; // @[Mux.scala 27:72]
  wire [5:0] _T_95 = io_i0_ap_sra ? _T_84 : 6'h0; // @[Mux.scala 27:72]
  wire [5:0] _T_96 = _T_93 | _T_94; // @[Mux.scala 27:72]
  wire [5:0] shift_amount = _T_96 | _T_95; // @[Mux.scala 27:72]
  wire [4:0] _T_102 = {io_i0_ap_sll,io_i0_ap_sll,io_i0_ap_sll,io_i0_ap_sll,io_i0_ap_sll}; // @[Cat.scala 29:58]
  wire [4:0] _T_104 = _T_102 & io_b_in[4:0]; // @[exu_alu_ctl.scala 61:64]
  wire [62:0] _T_105 = 63'hffffffff << _T_104; // @[exu_alu_ctl.scala 61:39]
  wire [9:0] _T_115 = {io_i0_ap_sra,io_i0_ap_sra,io_i0_ap_sra,io_i0_ap_sra,io_i0_ap_sra,io_i0_ap_sra,io_i0_ap_sra,io_i0_ap_sra,io_i0_ap_sra,io_i0_ap_sra}; // @[Cat.scala 29:58]
  wire [18:0] _T_124 = {_T_115,io_i0_ap_sra,io_i0_ap_sra,io_i0_ap_sra,io_i0_ap_sra,io_i0_ap_sra,io_i0_ap_sra,io_i0_ap_sra,io_i0_ap_sra,io_i0_ap_sra}; // @[Cat.scala 29:58]
  wire [27:0] _T_133 = {_T_124,io_i0_ap_sra,io_i0_ap_sra,io_i0_ap_sra,io_i0_ap_sra,io_i0_ap_sra,io_i0_ap_sra,io_i0_ap_sra,io_i0_ap_sra,io_i0_ap_sra}; // @[Cat.scala 29:58]
  wire [30:0] _T_136 = {_T_133,io_i0_ap_sra,io_i0_ap_sra,io_i0_ap_sra}; // @[Cat.scala 29:58]
  wire [9:0] _T_147 = {io_a_in[31],io_a_in[31],io_a_in[31],io_a_in[31],io_a_in[31],io_a_in[31],io_a_in[31],io_a_in[31],io_a_in[31],io_a_in[31]}; // @[Cat.scala 29:58]
  wire [18:0] _T_156 = {_T_147,io_a_in[31],io_a_in[31],io_a_in[31],io_a_in[31],io_a_in[31],io_a_in[31],io_a_in[31],io_a_in[31],io_a_in[31]}; // @[Cat.scala 29:58]
  wire [27:0] _T_165 = {_T_156,io_a_in[31],io_a_in[31],io_a_in[31],io_a_in[31],io_a_in[31],io_a_in[31],io_a_in[31],io_a_in[31],io_a_in[31]}; // @[Cat.scala 29:58]
  wire [30:0] _T_168 = {_T_165,io_a_in[31],io_a_in[31],io_a_in[31]}; // @[Cat.scala 29:58]
  wire [30:0] _T_169 = _T_136 & _T_168; // @[exu_alu_ctl.scala 64:47]
  wire [9:0] _T_179 = {io_i0_ap_sll,io_i0_ap_sll,io_i0_ap_sll,io_i0_ap_sll,io_i0_ap_sll,io_i0_ap_sll,io_i0_ap_sll,io_i0_ap_sll,io_i0_ap_sll,io_i0_ap_sll}; // @[Cat.scala 29:58]
  wire [18:0] _T_188 = {_T_179,io_i0_ap_sll,io_i0_ap_sll,io_i0_ap_sll,io_i0_ap_sll,io_i0_ap_sll,io_i0_ap_sll,io_i0_ap_sll,io_i0_ap_sll,io_i0_ap_sll}; // @[Cat.scala 29:58]
  wire [27:0] _T_197 = {_T_188,io_i0_ap_sll,io_i0_ap_sll,io_i0_ap_sll,io_i0_ap_sll,io_i0_ap_sll,io_i0_ap_sll,io_i0_ap_sll,io_i0_ap_sll,io_i0_ap_sll}; // @[Cat.scala 29:58]
  wire [30:0] _T_200 = {_T_197,io_i0_ap_sll,io_i0_ap_sll,io_i0_ap_sll}; // @[Cat.scala 29:58]
  wire [30:0] _T_202 = _T_200 & io_a_in[30:0]; // @[exu_alu_ctl.scala 64:96]
  wire [30:0] _T_203 = _T_169 | _T_202; // @[exu_alu_ctl.scala 64:71]
  wire [62:0] shift_extend = {_T_203,io_a_in}; // @[Cat.scala 29:58]
  wire [62:0] shift_long = shift_extend >> shift_amount[4:0]; // @[exu_alu_ctl.scala 67:32]
  wire [31:0] shift_mask = _T_105[31:0]; // @[exu_alu_ctl.scala 61:14]
  wire [31:0] sout = shift_long[31:0] & shift_mask; // @[exu_alu_ctl.scala 69:34]
  wire  _T_210 = io_i0_ap_sll | io_i0_ap_srl; // @[exu_alu_ctl.scala 72:44]
  wire  sel_shift = _T_210 | io_i0_ap_sra; // @[exu_alu_ctl.scala 72:59]
  wire  _T_211 = io_i0_ap_add | io_i0_ap_sub; // @[exu_alu_ctl.scala 73:44]
  wire  _T_212 = ~io_i0_ap_slt; // @[exu_alu_ctl.scala 73:62]
  wire  sel_adder = _T_211 & _T_212; // @[exu_alu_ctl.scala 73:60]
  wire  _T_213 = io_i0_ap_jal | io_pp_in_bits_pcall; // @[exu_alu_ctl.scala 74:44]
  wire  _T_214 = _T_213 | io_pp_in_bits_pja; // @[exu_alu_ctl.scala 74:66]
  wire  sel_pc = _T_214 | io_pp_in_bits_pret; // @[exu_alu_ctl.scala 74:86]
  wire  slt_one = io_i0_ap_slt & lt; // @[exu_alu_ctl.scala 77:43]
  wire [31:0] _T_217 = {io_dec_i0_pc_d,1'h0}; // @[Cat.scala 29:58]
  wire [12:0] _T_218 = {io_dec_alu_dec_i0_br_immed_d,1'h0}; // @[Cat.scala 29:58]
  wire [12:0] _T_221 = _T_217[12:1] + _T_218[12:1]; // @[lib.scala 68:31]
  wire [18:0] _T_224 = _T_217[31:13] + 19'h1; // @[lib.scala 69:27]
  wire [18:0] _T_227 = _T_217[31:13] - 19'h1; // @[lib.scala 70:27]
  wire  _T_230 = ~_T_221[12]; // @[lib.scala 72:28]
  wire  _T_231 = _T_218[12] ^ _T_230; // @[lib.scala 72:26]
  wire  _T_234 = ~_T_218[12]; // @[lib.scala 73:20]
  wire  _T_236 = _T_234 & _T_221[12]; // @[lib.scala 73:26]
  wire  _T_240 = _T_218[12] & _T_230; // @[lib.scala 74:26]
  wire [18:0] _T_242 = _T_231 ? _T_217[31:13] : 19'h0; // @[Mux.scala 27:72]
  wire [18:0] _T_243 = _T_236 ? _T_224 : 19'h0; // @[Mux.scala 27:72]
  wire [18:0] _T_244 = _T_240 ? _T_227 : 19'h0; // @[Mux.scala 27:72]
  wire [18:0] _T_245 = _T_242 | _T_243; // @[Mux.scala 27:72]
  wire [18:0] _T_246 = _T_245 | _T_244; // @[Mux.scala 27:72]
  wire [31:0] pcout = {_T_246,_T_221[11:0],1'h0}; // @[Cat.scala 29:58]
  wire [31:0] _T_250 = $signed(_T_77) | $signed(_T_73); // @[exu_alu_ctl.scala 83:24]
  wire [31:0] _T_251 = {31'h0,slt_one}; // @[Cat.scala 29:58]
  wire [31:0] _T_252 = _T_250 | _T_251; // @[exu_alu_ctl.scala 83:31]
  wire [31:0] _T_259 = io_i0_ap_csr_imm ? $signed(io_b_in) : $signed(io_a_in); // @[exu_alu_ctl.scala 87:54]
  wire [31:0] _T_260 = sel_shift ? sout : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_261 = sel_adder ? aout[31:0] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_262 = sel_pc ? pcout : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_263 = io_i0_ap_csr_write ? _T_259 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_264 = _T_260 | _T_261; // @[Mux.scala 27:72]
  wire [31:0] _T_265 = _T_264 | _T_262; // @[Mux.scala 27:72]
  wire [31:0] _T_266 = _T_265 | _T_263; // @[Mux.scala 27:72]
  wire  _T_271 = io_i0_ap_beq & eq; // @[exu_alu_ctl.scala 96:43]
  wire  _T_272 = io_i0_ap_bne & ne; // @[exu_alu_ctl.scala 96:65]
  wire  _T_273 = _T_271 | _T_272; // @[exu_alu_ctl.scala 96:49]
  wire  _T_274 = io_i0_ap_blt & lt; // @[exu_alu_ctl.scala 96:94]
  wire  _T_275 = _T_273 | _T_274; // @[exu_alu_ctl.scala 96:78]
  wire  _T_276 = io_i0_ap_bge & ge; // @[exu_alu_ctl.scala 96:116]
  wire  _T_277 = _T_275 | _T_276; // @[exu_alu_ctl.scala 96:100]
  wire  actual_taken = _T_277 | sel_pc; // @[exu_alu_ctl.scala 96:122]
  wire  _T_278 = io_dec_alu_dec_i0_alu_decode_d & io_i0_ap_predict_nt; // @[exu_alu_ctl.scala 101:61]
  wire  _T_279 = ~actual_taken; // @[exu_alu_ctl.scala 101:85]
  wire  _T_280 = _T_278 & _T_279; // @[exu_alu_ctl.scala 101:83]
  wire  _T_281 = ~sel_pc; // @[exu_alu_ctl.scala 101:101]
  wire  _T_282 = _T_280 & _T_281; // @[exu_alu_ctl.scala 101:99]
  wire  _T_283 = io_dec_alu_dec_i0_alu_decode_d & io_i0_ap_predict_t; // @[exu_alu_ctl.scala 101:145]
  wire  _T_284 = _T_283 & actual_taken; // @[exu_alu_ctl.scala 101:167]
  wire  _T_286 = _T_284 & _T_281; // @[exu_alu_ctl.scala 101:183]
  wire  _T_293 = io_i0_ap_predict_t & _T_279; // @[exu_alu_ctl.scala 106:48]
  wire  _T_294 = io_i0_ap_predict_nt & actual_taken; // @[exu_alu_ctl.scala 106:88]
  wire  cond_mispredict = _T_293 | _T_294; // @[exu_alu_ctl.scala 106:65]
  wire  _T_296 = io_pp_in_bits_prett != aout[31:1]; // @[exu_alu_ctl.scala 109:72]
  wire  target_mispredict = io_pp_in_bits_pret & _T_296; // @[exu_alu_ctl.scala 109:49]
  wire  _T_297 = io_i0_ap_jal | cond_mispredict; // @[exu_alu_ctl.scala 111:45]
  wire  _T_298 = _T_297 | target_mispredict; // @[exu_alu_ctl.scala 111:63]
  wire  _T_299 = _T_298 & io_dec_alu_dec_i0_alu_decode_d; // @[exu_alu_ctl.scala 111:84]
  wire  _T_300 = ~io_flush_upper_x; // @[exu_alu_ctl.scala 111:119]
  wire  _T_301 = _T_299 & _T_300; // @[exu_alu_ctl.scala 111:117]
  wire  _T_302 = ~io_dec_tlu_flush_lower_r; // @[exu_alu_ctl.scala 111:141]
  wire  _T_312 = io_pp_in_bits_hist[1] & io_pp_in_bits_hist[0]; // @[exu_alu_ctl.scala 116:44]
  wire  _T_314 = ~io_pp_in_bits_hist[0]; // @[exu_alu_ctl.scala 116:73]
  wire  _T_315 = _T_314 & actual_taken; // @[exu_alu_ctl.scala 116:96]
  wire  _T_316 = _T_312 | _T_315; // @[exu_alu_ctl.scala 116:70]
  wire  _T_318 = ~io_pp_in_bits_hist[1]; // @[exu_alu_ctl.scala 117:6]
  wire  _T_320 = _T_318 & _T_279; // @[exu_alu_ctl.scala 117:29]
  wire  _T_322 = io_pp_in_bits_hist[1] & actual_taken; // @[exu_alu_ctl.scala 117:72]
  wire  _T_323 = _T_320 | _T_322; // @[exu_alu_ctl.scala 117:47]
  wire  _T_327 = _T_300 & _T_302; // @[exu_alu_ctl.scala 120:56]
  wire  _T_328 = cond_mispredict | target_mispredict; // @[exu_alu_ctl.scala 120:103]
  rvclkhdr rvclkhdr ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_io_l1clk),
    .io_clk(rvclkhdr_io_clk),
    .io_en(rvclkhdr_io_en),
    .io_scan_mode(rvclkhdr_io_scan_mode)
  );
  rvclkhdr rvclkhdr_1 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_1_io_l1clk),
    .io_clk(rvclkhdr_1_io_clk),
    .io_en(rvclkhdr_1_io_en),
    .io_scan_mode(rvclkhdr_1_io_scan_mode)
  );
  assign io_dec_alu_exu_i0_pc_x = _T_1; // @[exu_alu_ctl.scala 30:26]
  assign io_result_ff = _T_3; // @[exu_alu_ctl.scala 32:16]
  assign io_flush_upper_out = _T_301 & _T_302; // @[exu_alu_ctl.scala 111:26]
  assign io_flush_final_out = _T_301 | io_dec_tlu_flush_lower_r; // @[exu_alu_ctl.scala 112:26]
  assign io_flush_path_out = sel_pc ? aout[31:1] : pcout[31:1]; // @[exu_alu_ctl.scala 103:22]
  assign io_pred_correct_out = _T_282 | _T_286; // @[exu_alu_ctl.scala 101:26]
  assign io_predict_p_out_valid = io_pp_in_valid; // @[exu_alu_ctl.scala 119:30]
  assign io_predict_p_out_bits_misp = _T_327 & _T_328; // @[exu_alu_ctl.scala 119:30 exu_alu_ctl.scala 120:35]
  assign io_predict_p_out_bits_ataken = _T_277 | sel_pc; // @[exu_alu_ctl.scala 119:30 exu_alu_ctl.scala 121:35]
  assign io_predict_p_out_bits_boffset = io_pp_in_bits_boffset; // @[exu_alu_ctl.scala 119:30]
  assign io_predict_p_out_bits_pc4 = io_pp_in_bits_pc4; // @[exu_alu_ctl.scala 119:30]
  assign io_predict_p_out_bits_hist = {_T_316,_T_323}; // @[exu_alu_ctl.scala 119:30 exu_alu_ctl.scala 122:35]
  assign io_predict_p_out_bits_toffset = io_pp_in_bits_toffset; // @[exu_alu_ctl.scala 119:30]
  assign io_predict_p_out_bits_br_error = io_pp_in_bits_br_error; // @[exu_alu_ctl.scala 119:30]
  assign io_predict_p_out_bits_br_start_error = io_pp_in_bits_br_start_error; // @[exu_alu_ctl.scala 119:30]
  assign io_predict_p_out_bits_pcall = io_pp_in_bits_pcall; // @[exu_alu_ctl.scala 119:30]
  assign io_predict_p_out_bits_pret = io_pp_in_bits_pret; // @[exu_alu_ctl.scala 119:30]
  assign io_predict_p_out_bits_pja = io_pp_in_bits_pja; // @[exu_alu_ctl.scala 119:30]
  assign io_predict_p_out_bits_way = io_pp_in_bits_way; // @[exu_alu_ctl.scala 119:30]
  assign rvclkhdr_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_io_en = io_enable; // @[lib.scala 371:17]
  assign rvclkhdr_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_1_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_1_io_en = io_enable; // @[lib.scala 371:17]
  assign rvclkhdr_1_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_1 = _RAND_0[30:0];
  _RAND_1 = {1{`RANDOM}};
  _T_3 = _RAND_1[31:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    _T_1 = 31'h0;
  end
  if (reset) begin
    _T_3 = 32'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge rvclkhdr_io_l1clk or posedge reset) begin
    if (reset) begin
      _T_1 <= 31'h0;
    end else begin
      _T_1 <= io_dec_i0_pc_d;
    end
  end
  always @(posedge rvclkhdr_1_io_l1clk or posedge reset) begin
    if (reset) begin
      _T_3 <= 32'h0;
    end else begin
      _T_3 <= _T_252 | _T_266;
    end
  end
endmodule
module exu_mul_ctl(
  input         clock,
  input         reset,
  input         io_scan_mode,
  input         io_mul_p_valid,
  input         io_mul_p_bits_rs1_sign,
  input         io_mul_p_bits_rs2_sign,
  input         io_mul_p_bits_low,
  input  [31:0] io_rs1_in,
  input  [31:0] io_rs2_in,
  output [31:0] io_result_x
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire  rvclkhdr_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_1_io_l1clk; // @[lib.scala 388:23]
  wire  rvclkhdr_1_io_clk; // @[lib.scala 388:23]
  wire  rvclkhdr_1_io_en; // @[lib.scala 388:23]
  wire  rvclkhdr_1_io_scan_mode; // @[lib.scala 388:23]
  wire  rvclkhdr_2_io_l1clk; // @[lib.scala 388:23]
  wire  rvclkhdr_2_io_clk; // @[lib.scala 388:23]
  wire  rvclkhdr_2_io_en; // @[lib.scala 388:23]
  wire  rvclkhdr_2_io_scan_mode; // @[lib.scala 388:23]
  wire  _T_1 = io_mul_p_bits_rs1_sign & io_rs1_in[31]; // @[exu_mul_ctl.scala 26:44]
  wire  _T_5 = io_mul_p_bits_rs2_sign & io_rs2_in[31]; // @[exu_mul_ctl.scala 27:44]
  reg  low_x; // @[lib.scala 374:16]
  reg [32:0] rs1_x; // @[lib.scala 394:16]
  reg [32:0] rs2_x; // @[lib.scala 394:16]
  wire [65:0] prod_x = $signed(rs1_x) * $signed(rs2_x); // @[exu_mul_ctl.scala 33:20]
  wire  _T_16 = ~low_x; // @[exu_mul_ctl.scala 34:29]
  wire [31:0] _T_20 = _T_16 ? prod_x[63:32] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_21 = low_x ? prod_x[31:0] : 32'h0; // @[Mux.scala 27:72]
  rvclkhdr rvclkhdr ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_io_l1clk),
    .io_clk(rvclkhdr_io_clk),
    .io_en(rvclkhdr_io_en),
    .io_scan_mode(rvclkhdr_io_scan_mode)
  );
  rvclkhdr rvclkhdr_1 ( // @[lib.scala 388:23]
    .io_l1clk(rvclkhdr_1_io_l1clk),
    .io_clk(rvclkhdr_1_io_clk),
    .io_en(rvclkhdr_1_io_en),
    .io_scan_mode(rvclkhdr_1_io_scan_mode)
  );
  rvclkhdr rvclkhdr_2 ( // @[lib.scala 388:23]
    .io_l1clk(rvclkhdr_2_io_l1clk),
    .io_clk(rvclkhdr_2_io_clk),
    .io_en(rvclkhdr_2_io_en),
    .io_scan_mode(rvclkhdr_2_io_scan_mode)
  );
  assign io_result_x = _T_20 | _T_21; // @[exu_mul_ctl.scala 34:15]
  assign rvclkhdr_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_io_en = io_mul_p_valid; // @[lib.scala 371:17]
  assign rvclkhdr_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_1_io_clk = clock; // @[lib.scala 390:18]
  assign rvclkhdr_1_io_en = io_mul_p_valid; // @[lib.scala 391:17]
  assign rvclkhdr_1_io_scan_mode = io_scan_mode; // @[lib.scala 392:24]
  assign rvclkhdr_2_io_clk = clock; // @[lib.scala 390:18]
  assign rvclkhdr_2_io_en = io_mul_p_valid; // @[lib.scala 391:17]
  assign rvclkhdr_2_io_scan_mode = io_scan_mode; // @[lib.scala 392:24]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  low_x = _RAND_0[0:0];
  _RAND_1 = {2{`RANDOM}};
  rs1_x = _RAND_1[32:0];
  _RAND_2 = {2{`RANDOM}};
  rs2_x = _RAND_2[32:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    low_x = 1'h0;
  end
  if (reset) begin
    rs1_x = 33'sh0;
  end
  if (reset) begin
    rs2_x = 33'sh0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge rvclkhdr_io_l1clk or posedge reset) begin
    if (reset) begin
      low_x <= 1'h0;
    end else begin
      low_x <= io_mul_p_bits_low;
    end
  end
  always @(posedge rvclkhdr_1_io_l1clk or posedge reset) begin
    if (reset) begin
      rs1_x <= 33'sh0;
    end else begin
      rs1_x <= {_T_1,io_rs1_in};
    end
  end
  always @(posedge rvclkhdr_2_io_l1clk or posedge reset) begin
    if (reset) begin
      rs2_x <= 33'sh0;
    end else begin
      rs2_x <= {_T_5,io_rs2_in};
    end
  end
endmodule
module exu_div_ctl(
  input         clock,
  input         reset,
  input         io_scan_mode,
  input  [31:0] io_dividend,
  input  [31:0] io_divisor,
  output [31:0] io_exu_div_result,
  output        io_exu_div_wren,
  input         io_dec_div_div_p_valid,
  input         io_dec_div_div_p_bits_unsign,
  input         io_dec_div_div_p_bits_rem,
  input         io_dec_div_dec_div_cancel
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
`endif // RANDOMIZE_REG_INIT
  wire  rvclkhdr_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_1_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_1_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_1_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_1_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_2_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_2_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_2_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_2_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_3_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_3_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_3_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_3_io_scan_mode; // @[lib.scala 368:23]
  wire  _T = ~io_dec_div_dec_div_cancel; // @[exu_div_ctl.scala 46:30]
  reg  valid_ff_x; // @[exu_div_ctl.scala 195:26]
  wire  valid_x = valid_ff_x & _T; // @[exu_div_ctl.scala 46:28]
  reg [32:0] q_ff; // @[lib.scala 374:16]
  wire  _T_2 = q_ff[31:4] == 28'h0; // @[exu_div_ctl.scala 52:34]
  reg [32:0] m_ff; // @[lib.scala 374:16]
  wire  _T_4 = m_ff[31:4] == 28'h0; // @[exu_div_ctl.scala 52:57]
  wire  _T_5 = _T_2 & _T_4; // @[exu_div_ctl.scala 52:43]
  wire  _T_7 = m_ff[31:0] != 32'h0; // @[exu_div_ctl.scala 52:80]
  wire  _T_8 = _T_5 & _T_7; // @[exu_div_ctl.scala 52:66]
  reg  rem_ff; // @[Reg.scala 27:20]
  wire  _T_9 = ~rem_ff; // @[exu_div_ctl.scala 52:91]
  wire  _T_10 = _T_8 & _T_9; // @[exu_div_ctl.scala 52:89]
  wire  _T_11 = _T_10 & valid_x; // @[exu_div_ctl.scala 52:99]
  wire  _T_13 = q_ff[31:0] == 32'h0; // @[exu_div_ctl.scala 53:18]
  wire  _T_16 = _T_13 & _T_7; // @[exu_div_ctl.scala 53:27]
  wire  _T_18 = _T_16 & _T_9; // @[exu_div_ctl.scala 53:50]
  wire  _T_19 = _T_18 & valid_x; // @[exu_div_ctl.scala 53:60]
  wire  smallnum_case = _T_11 | _T_19; // @[exu_div_ctl.scala 52:110]
  wire  _T_23 = ~m_ff[3]; // @[exu_div_ctl.scala 57:69]
  wire  _T_25 = ~m_ff[2]; // @[exu_div_ctl.scala 57:69]
  wire  _T_27 = ~m_ff[1]; // @[exu_div_ctl.scala 57:69]
  wire  _T_28 = _T_23 & _T_25; // @[exu_div_ctl.scala 57:94]
  wire  _T_29 = _T_28 & _T_27; // @[exu_div_ctl.scala 57:94]
  wire  _T_30 = q_ff[3] & _T_29; // @[exu_div_ctl.scala 58:10]
  wire  _T_37 = q_ff[3] & _T_28; // @[exu_div_ctl.scala 58:10]
  wire  _T_39 = ~m_ff[0]; // @[exu_div_ctl.scala 64:32]
  wire  _T_40 = _T_37 & _T_39; // @[exu_div_ctl.scala 64:30]
  wire  _T_50 = q_ff[2] & _T_29; // @[exu_div_ctl.scala 58:10]
  wire  _T_51 = _T_40 | _T_50; // @[exu_div_ctl.scala 64:41]
  wire  _T_54 = q_ff[3] & q_ff[2]; // @[exu_div_ctl.scala 56:94]
  wire  _T_60 = _T_54 & _T_28; // @[exu_div_ctl.scala 58:10]
  wire  _T_61 = _T_51 | _T_60; // @[exu_div_ctl.scala 64:73]
  wire  _T_68 = q_ff[2] & _T_28; // @[exu_div_ctl.scala 58:10]
  wire  _T_71 = _T_68 & _T_39; // @[exu_div_ctl.scala 66:30]
  wire  _T_81 = q_ff[1] & _T_29; // @[exu_div_ctl.scala 58:10]
  wire  _T_82 = _T_71 | _T_81; // @[exu_div_ctl.scala 66:41]
  wire  _T_88 = _T_23 & _T_27; // @[exu_div_ctl.scala 57:94]
  wire  _T_89 = q_ff[3] & _T_88; // @[exu_div_ctl.scala 58:10]
  wire  _T_92 = _T_89 & _T_39; // @[exu_div_ctl.scala 66:103]
  wire  _T_93 = _T_82 | _T_92; // @[exu_div_ctl.scala 66:76]
  wire  _T_96 = ~q_ff[2]; // @[exu_div_ctl.scala 56:69]
  wire  _T_97 = q_ff[3] & _T_96; // @[exu_div_ctl.scala 56:94]
  wire  _T_105 = _T_28 & m_ff[1]; // @[exu_div_ctl.scala 57:94]
  wire  _T_106 = _T_105 & m_ff[0]; // @[exu_div_ctl.scala 57:94]
  wire  _T_107 = _T_97 & _T_106; // @[exu_div_ctl.scala 58:10]
  wire  _T_108 = _T_93 | _T_107; // @[exu_div_ctl.scala 66:114]
  wire  _T_110 = ~q_ff[3]; // @[exu_div_ctl.scala 56:69]
  wire  _T_113 = _T_110 & q_ff[2]; // @[exu_div_ctl.scala 56:94]
  wire  _T_114 = _T_113 & q_ff[1]; // @[exu_div_ctl.scala 56:94]
  wire  _T_120 = _T_114 & _T_28; // @[exu_div_ctl.scala 58:10]
  wire  _T_121 = _T_108 | _T_120; // @[exu_div_ctl.scala 67:43]
  wire  _T_127 = _T_54 & _T_23; // @[exu_div_ctl.scala 58:10]
  wire  _T_130 = _T_127 & _T_39; // @[exu_div_ctl.scala 67:104]
  wire  _T_131 = _T_121 | _T_130; // @[exu_div_ctl.scala 67:78]
  wire  _T_140 = _T_23 & m_ff[2]; // @[exu_div_ctl.scala 57:94]
  wire  _T_141 = _T_140 & _T_27; // @[exu_div_ctl.scala 57:94]
  wire  _T_142 = _T_54 & _T_141; // @[exu_div_ctl.scala 58:10]
  wire  _T_143 = _T_131 | _T_142; // @[exu_div_ctl.scala 67:116]
  wire  _T_146 = q_ff[3] & q_ff[1]; // @[exu_div_ctl.scala 56:94]
  wire  _T_152 = _T_146 & _T_88; // @[exu_div_ctl.scala 58:10]
  wire  _T_153 = _T_143 | _T_152; // @[exu_div_ctl.scala 68:43]
  wire  _T_158 = _T_54 & q_ff[1]; // @[exu_div_ctl.scala 56:94]
  wire  _T_163 = _T_158 & _T_140; // @[exu_div_ctl.scala 58:10]
  wire  _T_164 = _T_153 | _T_163; // @[exu_div_ctl.scala 68:77]
  wire  _T_168 = q_ff[2] & q_ff[1]; // @[exu_div_ctl.scala 56:94]
  wire  _T_169 = _T_168 & q_ff[0]; // @[exu_div_ctl.scala 56:94]
  wire  _T_175 = _T_169 & _T_88; // @[exu_div_ctl.scala 58:10]
  wire  _T_181 = _T_97 & q_ff[0]; // @[exu_div_ctl.scala 56:94]
  wire  _T_186 = _T_23 & m_ff[1]; // @[exu_div_ctl.scala 57:94]
  wire  _T_187 = _T_186 & m_ff[0]; // @[exu_div_ctl.scala 57:94]
  wire  _T_188 = _T_181 & _T_187; // @[exu_div_ctl.scala 58:10]
  wire  _T_189 = _T_175 | _T_188; // @[exu_div_ctl.scala 70:44]
  wire  _T_196 = q_ff[2] & _T_88; // @[exu_div_ctl.scala 58:10]
  wire  _T_199 = _T_196 & _T_39; // @[exu_div_ctl.scala 70:111]
  wire  _T_200 = _T_189 | _T_199; // @[exu_div_ctl.scala 70:84]
  wire  _T_207 = q_ff[1] & _T_28; // @[exu_div_ctl.scala 58:10]
  wire  _T_210 = _T_207 & _T_39; // @[exu_div_ctl.scala 71:32]
  wire  _T_211 = _T_200 | _T_210; // @[exu_div_ctl.scala 70:126]
  wire  _T_221 = q_ff[0] & _T_29; // @[exu_div_ctl.scala 58:10]
  wire  _T_222 = _T_211 | _T_221; // @[exu_div_ctl.scala 71:46]
  wire  _T_227 = ~q_ff[1]; // @[exu_div_ctl.scala 56:69]
  wire  _T_229 = _T_113 & _T_227; // @[exu_div_ctl.scala 56:94]
  wire  _T_239 = _T_229 & _T_106; // @[exu_div_ctl.scala 58:10]
  wire  _T_240 = _T_222 | _T_239; // @[exu_div_ctl.scala 71:86]
  wire  _T_249 = _T_114 & _T_23; // @[exu_div_ctl.scala 58:10]
  wire  _T_252 = _T_249 & _T_39; // @[exu_div_ctl.scala 72:35]
  wire  _T_253 = _T_240 | _T_252; // @[exu_div_ctl.scala 71:128]
  wire  _T_259 = _T_25 & _T_27; // @[exu_div_ctl.scala 57:94]
  wire  _T_260 = q_ff[3] & _T_259; // @[exu_div_ctl.scala 58:10]
  wire  _T_263 = _T_260 & _T_39; // @[exu_div_ctl.scala 72:74]
  wire  _T_264 = _T_253 | _T_263; // @[exu_div_ctl.scala 72:46]
  wire  _T_274 = _T_140 & m_ff[1]; // @[exu_div_ctl.scala 57:94]
  wire  _T_275 = _T_97 & _T_274; // @[exu_div_ctl.scala 58:10]
  wire  _T_276 = _T_264 | _T_275; // @[exu_div_ctl.scala 72:86]
  wire  _T_290 = _T_114 & _T_141; // @[exu_div_ctl.scala 58:10]
  wire  _T_291 = _T_276 | _T_290; // @[exu_div_ctl.scala 72:128]
  wire  _T_297 = _T_113 & q_ff[0]; // @[exu_div_ctl.scala 56:94]
  wire  _T_303 = _T_297 & _T_88; // @[exu_div_ctl.scala 58:10]
  wire  _T_304 = _T_291 | _T_303; // @[exu_div_ctl.scala 73:46]
  wire  _T_311 = _T_97 & _T_227; // @[exu_div_ctl.scala 56:94]
  wire  _T_317 = _T_140 & m_ff[0]; // @[exu_div_ctl.scala 57:94]
  wire  _T_318 = _T_311 & _T_317; // @[exu_div_ctl.scala 58:10]
  wire  _T_319 = _T_304 | _T_318; // @[exu_div_ctl.scala 73:86]
  wire  _T_324 = _T_96 & q_ff[1]; // @[exu_div_ctl.scala 56:94]
  wire  _T_325 = _T_324 & q_ff[0]; // @[exu_div_ctl.scala 56:94]
  wire  _T_331 = _T_325 & _T_28; // @[exu_div_ctl.scala 58:10]
  wire  _T_332 = _T_319 | _T_331; // @[exu_div_ctl.scala 73:128]
  wire  _T_338 = _T_54 & _T_27; // @[exu_div_ctl.scala 58:10]
  wire  _T_341 = _T_338 & _T_39; // @[exu_div_ctl.scala 74:73]
  wire  _T_342 = _T_332 | _T_341; // @[exu_div_ctl.scala 74:46]
  wire  _T_350 = _T_114 & q_ff[0]; // @[exu_div_ctl.scala 56:94]
  wire  _T_355 = _T_350 & _T_140; // @[exu_div_ctl.scala 58:10]
  wire  _T_356 = _T_342 | _T_355; // @[exu_div_ctl.scala 74:86]
  wire  _T_363 = m_ff[3] & _T_25; // @[exu_div_ctl.scala 57:94]
  wire  _T_364 = _T_54 & _T_363; // @[exu_div_ctl.scala 58:10]
  wire  _T_365 = _T_356 | _T_364; // @[exu_div_ctl.scala 74:128]
  wire  _T_375 = _T_363 & _T_27; // @[exu_div_ctl.scala 57:94]
  wire  _T_376 = _T_146 & _T_375; // @[exu_div_ctl.scala 58:10]
  wire  _T_377 = _T_365 | _T_376; // @[exu_div_ctl.scala 75:46]
  wire  _T_380 = q_ff[3] & q_ff[0]; // @[exu_div_ctl.scala 56:94]
  wire  _T_386 = _T_380 & _T_259; // @[exu_div_ctl.scala 58:10]
  wire  _T_387 = _T_377 | _T_386; // @[exu_div_ctl.scala 75:86]
  wire  _T_391 = q_ff[3] & _T_227; // @[exu_div_ctl.scala 56:94]
  wire  _T_399 = _T_274 & m_ff[0]; // @[exu_div_ctl.scala 57:94]
  wire  _T_400 = _T_391 & _T_399; // @[exu_div_ctl.scala 58:10]
  wire  _T_401 = _T_387 | _T_400; // @[exu_div_ctl.scala 75:128]
  wire  _T_408 = _T_158 & m_ff[3]; // @[exu_div_ctl.scala 58:10]
  wire  _T_411 = _T_408 & _T_39; // @[exu_div_ctl.scala 76:75]
  wire  _T_412 = _T_401 | _T_411; // @[exu_div_ctl.scala 76:46]
  wire  _T_421 = m_ff[3] & _T_27; // @[exu_div_ctl.scala 57:94]
  wire  _T_422 = _T_158 & _T_421; // @[exu_div_ctl.scala 58:10]
  wire  _T_423 = _T_412 | _T_422; // @[exu_div_ctl.scala 76:86]
  wire  _T_428 = _T_54 & q_ff[0]; // @[exu_div_ctl.scala 56:94]
  wire  _T_433 = _T_428 & _T_421; // @[exu_div_ctl.scala 58:10]
  wire  _T_434 = _T_423 | _T_433; // @[exu_div_ctl.scala 76:128]
  wire  _T_440 = _T_97 & q_ff[1]; // @[exu_div_ctl.scala 56:94]
  wire  _T_445 = _T_440 & _T_186; // @[exu_div_ctl.scala 58:10]
  wire  _T_446 = _T_434 | _T_445; // @[exu_div_ctl.scala 77:46]
  wire  _T_451 = _T_146 & q_ff[0]; // @[exu_div_ctl.scala 56:94]
  wire  _T_454 = _T_451 & _T_25; // @[exu_div_ctl.scala 58:10]
  wire  _T_455 = _T_446 | _T_454; // @[exu_div_ctl.scala 77:86]
  wire  _T_462 = _T_158 & q_ff[0]; // @[exu_div_ctl.scala 56:94]
  wire  _T_464 = _T_462 & m_ff[3]; // @[exu_div_ctl.scala 58:10]
  wire  _T_465 = _T_455 | _T_464; // @[exu_div_ctl.scala 77:128]
  wire  _T_471 = _T_146 & _T_25; // @[exu_div_ctl.scala 58:10]
  wire  _T_474 = _T_471 & _T_39; // @[exu_div_ctl.scala 78:72]
  wire  _T_475 = _T_465 | _T_474; // @[exu_div_ctl.scala 78:46]
  wire [1:0] _T_476 = {_T_164,_T_475}; // @[Cat.scala 29:58]
  wire [1:0] _T_477 = {_T_30,_T_61}; // @[Cat.scala 29:58]
  reg  sign_ff; // @[Reg.scala 27:20]
  wire  _T_479 = sign_ff & q_ff[31]; // @[exu_div_ctl.scala 87:34]
  wire [32:0] short_dividend = {_T_479,q_ff[31:0]}; // @[Cat.scala 29:58]
  wire  _T_484 = ~short_dividend[32]; // @[exu_div_ctl.scala 92:7]
  wire  _T_487 = short_dividend[31:24] != 8'h0; // @[exu_div_ctl.scala 92:60]
  wire  _T_492 = short_dividend[31:23] != 9'h1ff; // @[exu_div_ctl.scala 93:59]
  wire  _T_493 = _T_484 & _T_487; // @[Mux.scala 27:72]
  wire  _T_494 = short_dividend[32] & _T_492; // @[Mux.scala 27:72]
  wire  _T_495 = _T_493 | _T_494; // @[Mux.scala 27:72]
  wire  _T_502 = short_dividend[23:16] != 8'h0; // @[exu_div_ctl.scala 96:60]
  wire  _T_507 = short_dividend[22:15] != 8'hff; // @[exu_div_ctl.scala 97:59]
  wire  _T_508 = _T_484 & _T_502; // @[Mux.scala 27:72]
  wire  _T_509 = short_dividend[32] & _T_507; // @[Mux.scala 27:72]
  wire  _T_510 = _T_508 | _T_509; // @[Mux.scala 27:72]
  wire  _T_517 = short_dividend[15:8] != 8'h0; // @[exu_div_ctl.scala 100:59]
  wire  _T_522 = short_dividend[14:7] != 8'hff; // @[exu_div_ctl.scala 101:58]
  wire  _T_523 = _T_484 & _T_517; // @[Mux.scala 27:72]
  wire  _T_524 = short_dividend[32] & _T_522; // @[Mux.scala 27:72]
  wire  _T_525 = _T_523 | _T_524; // @[Mux.scala 27:72]
  wire [2:0] a_cls = {_T_495,_T_510,_T_525}; // @[Cat.scala 29:58]
  wire  _T_530 = ~m_ff[32]; // @[exu_div_ctl.scala 106:7]
  wire  _T_533 = m_ff[31:24] != 8'h0; // @[exu_div_ctl.scala 106:40]
  wire  _T_538 = m_ff[31:24] != 8'hff; // @[exu_div_ctl.scala 107:39]
  wire  _T_539 = _T_530 & _T_533; // @[Mux.scala 27:72]
  wire  _T_540 = m_ff[32] & _T_538; // @[Mux.scala 27:72]
  wire  _T_541 = _T_539 | _T_540; // @[Mux.scala 27:72]
  wire  _T_548 = m_ff[23:16] != 8'h0; // @[exu_div_ctl.scala 110:40]
  wire  _T_553 = m_ff[23:16] != 8'hff; // @[exu_div_ctl.scala 111:39]
  wire  _T_554 = _T_530 & _T_548; // @[Mux.scala 27:72]
  wire  _T_555 = m_ff[32] & _T_553; // @[Mux.scala 27:72]
  wire  _T_556 = _T_554 | _T_555; // @[Mux.scala 27:72]
  wire  _T_563 = m_ff[15:8] != 8'h0; // @[exu_div_ctl.scala 114:39]
  wire  _T_568 = m_ff[15:8] != 8'hff; // @[exu_div_ctl.scala 115:38]
  wire  _T_569 = _T_530 & _T_563; // @[Mux.scala 27:72]
  wire  _T_570 = m_ff[32] & _T_568; // @[Mux.scala 27:72]
  wire  _T_571 = _T_569 | _T_570; // @[Mux.scala 27:72]
  wire [2:0] b_cls = {_T_541,_T_556,_T_571}; // @[Cat.scala 29:58]
  wire  _T_575 = a_cls[2:1] == 2'h1; // @[exu_div_ctl.scala 119:19]
  wire  _T_578 = _T_575 & b_cls[2]; // @[exu_div_ctl.scala 119:34]
  wire  _T_580 = a_cls == 3'h1; // @[exu_div_ctl.scala 120:21]
  wire  _T_583 = _T_580 & b_cls[2]; // @[exu_div_ctl.scala 120:36]
  wire  _T_584 = _T_578 | _T_583; // @[exu_div_ctl.scala 119:65]
  wire  _T_586 = a_cls == 3'h0; // @[exu_div_ctl.scala 121:21]
  wire  _T_589 = _T_586 & b_cls[2]; // @[exu_div_ctl.scala 121:36]
  wire  _T_590 = _T_584 | _T_589; // @[exu_div_ctl.scala 120:67]
  wire  _T_594 = b_cls[2:1] == 2'h1; // @[exu_div_ctl.scala 122:50]
  wire  _T_595 = _T_580 & _T_594; // @[exu_div_ctl.scala 122:36]
  wire  _T_596 = _T_590 | _T_595; // @[exu_div_ctl.scala 121:67]
  wire  _T_601 = _T_586 & _T_594; // @[exu_div_ctl.scala 123:36]
  wire  _T_602 = _T_596 | _T_601; // @[exu_div_ctl.scala 122:67]
  wire  _T_606 = b_cls == 3'h1; // @[exu_div_ctl.scala 124:50]
  wire  _T_607 = _T_586 & _T_606; // @[exu_div_ctl.scala 124:36]
  wire  _T_608 = _T_602 | _T_607; // @[exu_div_ctl.scala 123:67]
  wire  _T_613 = a_cls[2] & b_cls[2]; // @[exu_div_ctl.scala 126:34]
  wire  _T_618 = _T_575 & _T_594; // @[exu_div_ctl.scala 127:36]
  wire  _T_619 = _T_613 | _T_618; // @[exu_div_ctl.scala 126:65]
  wire  _T_624 = _T_580 & _T_606; // @[exu_div_ctl.scala 128:36]
  wire  _T_625 = _T_619 | _T_624; // @[exu_div_ctl.scala 127:67]
  wire  _T_629 = b_cls == 3'h0; // @[exu_div_ctl.scala 129:50]
  wire  _T_630 = _T_586 & _T_629; // @[exu_div_ctl.scala 129:36]
  wire  _T_631 = _T_625 | _T_630; // @[exu_div_ctl.scala 128:67]
  wire  _T_636 = a_cls[2] & _T_594; // @[exu_div_ctl.scala 131:34]
  wire  _T_641 = _T_575 & _T_606; // @[exu_div_ctl.scala 132:36]
  wire  _T_642 = _T_636 | _T_641; // @[exu_div_ctl.scala 131:65]
  wire  _T_647 = _T_580 & _T_629; // @[exu_div_ctl.scala 133:36]
  wire  _T_648 = _T_642 | _T_647; // @[exu_div_ctl.scala 132:67]
  wire  _T_653 = a_cls[2] & _T_606; // @[exu_div_ctl.scala 135:34]
  wire  _T_658 = _T_575 & _T_629; // @[exu_div_ctl.scala 136:36]
  wire  _T_659 = _T_653 | _T_658; // @[exu_div_ctl.scala 135:65]
  wire [3:0] shortq_raw = {_T_608,_T_631,_T_648,_T_659}; // @[Cat.scala 29:58]
  wire  _T_664 = valid_ff_x & _T_7; // @[exu_div_ctl.scala 139:35]
  wire  _T_665 = shortq_raw != 4'h0; // @[exu_div_ctl.scala 139:78]
  wire  shortq_enable = _T_664 & _T_665; // @[exu_div_ctl.scala 139:64]
  wire [3:0] _T_667 = shortq_enable ? 4'hf : 4'h0; // @[Bitwise.scala 72:12]
  reg [3:0] shortq_shift_xx; // @[exu_div_ctl.scala 206:31]
  wire [4:0] _T_676 = shortq_shift_xx[3] ? 5'h1f : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_677 = shortq_shift_xx[2] ? 5'h18 : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_678 = shortq_shift_xx[1] ? 5'h10 : 5'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_679 = shortq_shift_xx[0] ? 4'h8 : 4'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_680 = _T_676 | _T_677; // @[Mux.scala 27:72]
  wire [4:0] _T_681 = _T_680 | _T_678; // @[Mux.scala 27:72]
  wire [4:0] _GEN_4 = {{1'd0}, _T_679}; // @[Mux.scala 27:72]
  wire [4:0] shortq_shift_ff = _T_681 | _GEN_4; // @[Mux.scala 27:72]
  reg [5:0] count; // @[exu_div_ctl.scala 198:21]
  wire  _T_684 = count == 6'h20; // @[exu_div_ctl.scala 150:55]
  wire  _T_685 = count == 6'h21; // @[exu_div_ctl.scala 150:76]
  wire  _T_686 = _T_9 ? _T_684 : _T_685; // @[exu_div_ctl.scala 150:39]
  wire  finish = smallnum_case | _T_686; // @[exu_div_ctl.scala 150:34]
  reg  run_state; // @[exu_div_ctl.scala 197:25]
  wire  _T_687 = io_dec_div_div_p_valid | run_state; // @[exu_div_ctl.scala 151:43]
  wire  _T_688 = _T_687 | finish; // @[exu_div_ctl.scala 151:55]
  reg  finish_ff; // @[exu_div_ctl.scala 196:25]
  wire  _T_690 = ~finish; // @[exu_div_ctl.scala 152:59]
  wire  _T_691 = _T_687 & _T_690; // @[exu_div_ctl.scala 152:57]
  wire  _T_694 = run_state & _T_690; // @[exu_div_ctl.scala 153:35]
  wire  _T_696 = _T_694 & _T; // @[exu_div_ctl.scala 153:45]
  wire  _T_697 = ~shortq_enable; // @[exu_div_ctl.scala 153:76]
  wire  _T_698 = _T_696 & _T_697; // @[exu_div_ctl.scala 153:74]
  wire [5:0] _T_700 = _T_698 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  wire [5:0] _T_701 = {1'h0,shortq_shift_ff}; // @[Cat.scala 29:58]
  wire [5:0] _T_703 = count + _T_701; // @[exu_div_ctl.scala 153:102]
  wire [5:0] _T_705 = _T_703 + 6'h1; // @[exu_div_ctl.scala 153:129]
  wire  _T_709 = ~io_dec_div_div_p_bits_unsign; // @[exu_div_ctl.scala 157:20]
  wire  _T_710 = io_divisor != 32'h0; // @[exu_div_ctl.scala 157:64]
  wire  sign_eff = _T_709 & _T_710; // @[exu_div_ctl.scala 157:50]
  wire  _T_711 = ~run_state; // @[exu_div_ctl.scala 161:6]
  wire [32:0] _T_713 = {1'h0,io_dividend}; // @[Cat.scala 29:58]
  reg  shortq_enable_ff; // @[exu_div_ctl.scala 205:32]
  wire  _T_714 = valid_ff_x | shortq_enable_ff; // @[exu_div_ctl.scala 162:30]
  wire  _T_715 = run_state & _T_714; // @[exu_div_ctl.scala 162:16]
  reg  dividend_neg_ff; // @[Reg.scala 27:20]
  wire  _T_738 = sign_ff & dividend_neg_ff; // @[exu_div_ctl.scala 166:32]
  wire  _T_923 = |q_ff[30:0]; // @[lib.scala 403:35]
  wire  _T_925 = ~q_ff[31]; // @[lib.scala 403:40]
  wire  _T_927 = _T_923 ? _T_925 : q_ff[31]; // @[lib.scala 403:23]
  wire  _T_917 = |q_ff[29:0]; // @[lib.scala 403:35]
  wire  _T_919 = ~q_ff[30]; // @[lib.scala 403:40]
  wire  _T_921 = _T_917 ? _T_919 : q_ff[30]; // @[lib.scala 403:23]
  wire  _T_911 = |q_ff[28:0]; // @[lib.scala 403:35]
  wire  _T_913 = ~q_ff[29]; // @[lib.scala 403:40]
  wire  _T_915 = _T_911 ? _T_913 : q_ff[29]; // @[lib.scala 403:23]
  wire  _T_905 = |q_ff[27:0]; // @[lib.scala 403:35]
  wire  _T_907 = ~q_ff[28]; // @[lib.scala 403:40]
  wire  _T_909 = _T_905 ? _T_907 : q_ff[28]; // @[lib.scala 403:23]
  wire  _T_899 = |q_ff[26:0]; // @[lib.scala 403:35]
  wire  _T_901 = ~q_ff[27]; // @[lib.scala 403:40]
  wire  _T_903 = _T_899 ? _T_901 : q_ff[27]; // @[lib.scala 403:23]
  wire  _T_893 = |q_ff[25:0]; // @[lib.scala 403:35]
  wire  _T_895 = ~q_ff[26]; // @[lib.scala 403:40]
  wire  _T_897 = _T_893 ? _T_895 : q_ff[26]; // @[lib.scala 403:23]
  wire  _T_887 = |q_ff[24:0]; // @[lib.scala 403:35]
  wire  _T_889 = ~q_ff[25]; // @[lib.scala 403:40]
  wire  _T_891 = _T_887 ? _T_889 : q_ff[25]; // @[lib.scala 403:23]
  wire  _T_881 = |q_ff[23:0]; // @[lib.scala 403:35]
  wire  _T_883 = ~q_ff[24]; // @[lib.scala 403:40]
  wire  _T_885 = _T_881 ? _T_883 : q_ff[24]; // @[lib.scala 403:23]
  wire  _T_875 = |q_ff[22:0]; // @[lib.scala 403:35]
  wire  _T_877 = ~q_ff[23]; // @[lib.scala 403:40]
  wire  _T_879 = _T_875 ? _T_877 : q_ff[23]; // @[lib.scala 403:23]
  wire  _T_869 = |q_ff[21:0]; // @[lib.scala 403:35]
  wire  _T_871 = ~q_ff[22]; // @[lib.scala 403:40]
  wire  _T_873 = _T_869 ? _T_871 : q_ff[22]; // @[lib.scala 403:23]
  wire  _T_863 = |q_ff[20:0]; // @[lib.scala 403:35]
  wire  _T_865 = ~q_ff[21]; // @[lib.scala 403:40]
  wire  _T_867 = _T_863 ? _T_865 : q_ff[21]; // @[lib.scala 403:23]
  wire  _T_857 = |q_ff[19:0]; // @[lib.scala 403:35]
  wire  _T_859 = ~q_ff[20]; // @[lib.scala 403:40]
  wire  _T_861 = _T_857 ? _T_859 : q_ff[20]; // @[lib.scala 403:23]
  wire  _T_851 = |q_ff[18:0]; // @[lib.scala 403:35]
  wire  _T_853 = ~q_ff[19]; // @[lib.scala 403:40]
  wire  _T_855 = _T_851 ? _T_853 : q_ff[19]; // @[lib.scala 403:23]
  wire  _T_845 = |q_ff[17:0]; // @[lib.scala 403:35]
  wire  _T_847 = ~q_ff[18]; // @[lib.scala 403:40]
  wire  _T_849 = _T_845 ? _T_847 : q_ff[18]; // @[lib.scala 403:23]
  wire  _T_839 = |q_ff[16:0]; // @[lib.scala 403:35]
  wire  _T_841 = ~q_ff[17]; // @[lib.scala 403:40]
  wire  _T_843 = _T_839 ? _T_841 : q_ff[17]; // @[lib.scala 403:23]
  wire  _T_833 = |q_ff[15:0]; // @[lib.scala 403:35]
  wire  _T_835 = ~q_ff[16]; // @[lib.scala 403:40]
  wire  _T_837 = _T_833 ? _T_835 : q_ff[16]; // @[lib.scala 403:23]
  wire [7:0] _T_948 = {_T_879,_T_873,_T_867,_T_861,_T_855,_T_849,_T_843,_T_837}; // @[lib.scala 405:14]
  wire  _T_827 = |q_ff[14:0]; // @[lib.scala 403:35]
  wire  _T_829 = ~q_ff[15]; // @[lib.scala 403:40]
  wire  _T_831 = _T_827 ? _T_829 : q_ff[15]; // @[lib.scala 403:23]
  wire  _T_821 = |q_ff[13:0]; // @[lib.scala 403:35]
  wire  _T_823 = ~q_ff[14]; // @[lib.scala 403:40]
  wire  _T_825 = _T_821 ? _T_823 : q_ff[14]; // @[lib.scala 403:23]
  wire  _T_815 = |q_ff[12:0]; // @[lib.scala 403:35]
  wire  _T_817 = ~q_ff[13]; // @[lib.scala 403:40]
  wire  _T_819 = _T_815 ? _T_817 : q_ff[13]; // @[lib.scala 403:23]
  wire  _T_809 = |q_ff[11:0]; // @[lib.scala 403:35]
  wire  _T_811 = ~q_ff[12]; // @[lib.scala 403:40]
  wire  _T_813 = _T_809 ? _T_811 : q_ff[12]; // @[lib.scala 403:23]
  wire  _T_803 = |q_ff[10:0]; // @[lib.scala 403:35]
  wire  _T_805 = ~q_ff[11]; // @[lib.scala 403:40]
  wire  _T_807 = _T_803 ? _T_805 : q_ff[11]; // @[lib.scala 403:23]
  wire  _T_797 = |q_ff[9:0]; // @[lib.scala 403:35]
  wire  _T_799 = ~q_ff[10]; // @[lib.scala 403:40]
  wire  _T_801 = _T_797 ? _T_799 : q_ff[10]; // @[lib.scala 403:23]
  wire  _T_791 = |q_ff[8:0]; // @[lib.scala 403:35]
  wire  _T_793 = ~q_ff[9]; // @[lib.scala 403:40]
  wire  _T_795 = _T_791 ? _T_793 : q_ff[9]; // @[lib.scala 403:23]
  wire  _T_785 = |q_ff[7:0]; // @[lib.scala 403:35]
  wire  _T_787 = ~q_ff[8]; // @[lib.scala 403:40]
  wire  _T_789 = _T_785 ? _T_787 : q_ff[8]; // @[lib.scala 403:23]
  wire  _T_779 = |q_ff[6:0]; // @[lib.scala 403:35]
  wire  _T_781 = ~q_ff[7]; // @[lib.scala 403:40]
  wire  _T_783 = _T_779 ? _T_781 : q_ff[7]; // @[lib.scala 403:23]
  wire  _T_773 = |q_ff[5:0]; // @[lib.scala 403:35]
  wire  _T_775 = ~q_ff[6]; // @[lib.scala 403:40]
  wire  _T_777 = _T_773 ? _T_775 : q_ff[6]; // @[lib.scala 403:23]
  wire  _T_767 = |q_ff[4:0]; // @[lib.scala 403:35]
  wire  _T_769 = ~q_ff[5]; // @[lib.scala 403:40]
  wire  _T_771 = _T_767 ? _T_769 : q_ff[5]; // @[lib.scala 403:23]
  wire  _T_761 = |q_ff[3:0]; // @[lib.scala 403:35]
  wire  _T_763 = ~q_ff[4]; // @[lib.scala 403:40]
  wire  _T_765 = _T_761 ? _T_763 : q_ff[4]; // @[lib.scala 403:23]
  wire  _T_755 = |q_ff[2:0]; // @[lib.scala 403:35]
  wire  _T_757 = ~q_ff[3]; // @[lib.scala 403:40]
  wire  _T_759 = _T_755 ? _T_757 : q_ff[3]; // @[lib.scala 403:23]
  wire  _T_749 = |q_ff[1:0]; // @[lib.scala 403:35]
  wire  _T_751 = ~q_ff[2]; // @[lib.scala 403:40]
  wire  _T_753 = _T_749 ? _T_751 : q_ff[2]; // @[lib.scala 403:23]
  wire  _T_743 = |q_ff[0]; // @[lib.scala 403:35]
  wire  _T_745 = ~q_ff[1]; // @[lib.scala 403:40]
  wire  _T_747 = _T_743 ? _T_745 : q_ff[1]; // @[lib.scala 403:23]
  wire [6:0] _T_933 = {_T_783,_T_777,_T_771,_T_765,_T_759,_T_753,_T_747}; // @[lib.scala 405:14]
  wire [14:0] _T_941 = {_T_831,_T_825,_T_819,_T_813,_T_807,_T_801,_T_795,_T_789,_T_933}; // @[lib.scala 405:14]
  wire [30:0] _T_957 = {_T_927,_T_921,_T_915,_T_909,_T_903,_T_897,_T_891,_T_885,_T_948,_T_941}; // @[lib.scala 405:14]
  wire [31:0] _T_959 = {_T_957,q_ff[0]}; // @[Cat.scala 29:58]
  wire [31:0] dividend_eff = _T_738 ? _T_959 : q_ff[31:0]; // @[exu_div_ctl.scala 166:22]
  wire [32:0] _T_995 = run_state ? 33'h1ffffffff : 33'h0; // @[Bitwise.scala 72:12]
  wire  _T_1007 = _T_685 & rem_ff; // @[exu_div_ctl.scala 182:41]
  reg [32:0] a_ff; // @[lib.scala 374:16]
  wire  rem_correct = _T_1007 & a_ff[32]; // @[exu_div_ctl.scala 182:50]
  wire [32:0] _T_980 = rem_correct ? a_ff : 33'h0; // @[Mux.scala 27:72]
  wire  _T_968 = ~rem_correct; // @[exu_div_ctl.scala 173:6]
  wire  _T_969 = ~shortq_enable_ff; // @[exu_div_ctl.scala 173:21]
  wire  _T_970 = _T_968 & _T_969; // @[exu_div_ctl.scala 173:19]
  wire [32:0] _T_974 = {a_ff[31:0],q_ff[32]}; // @[Cat.scala 29:58]
  wire [32:0] _T_981 = _T_970 ? _T_974 : 33'h0; // @[Mux.scala 27:72]
  wire [32:0] _T_983 = _T_980 | _T_981; // @[Mux.scala 27:72]
  wire  _T_976 = _T_968 & shortq_enable_ff; // @[exu_div_ctl.scala 174:19]
  wire [55:0] _T_965 = {24'h0,dividend_eff}; // @[Cat.scala 29:58]
  wire [86:0] _GEN_5 = {{31'd0}, _T_965}; // @[exu_div_ctl.scala 170:47]
  wire [86:0] _T_966 = _GEN_5 << shortq_shift_ff; // @[exu_div_ctl.scala 170:47]
  wire [55:0] a_eff_shift = _T_966[55:0]; // @[exu_div_ctl.scala 170:15]
  wire [32:0] _T_979 = {9'h0,a_eff_shift[55:32]}; // @[Cat.scala 29:58]
  wire [32:0] _T_982 = _T_976 ? _T_979 : 33'h0; // @[Mux.scala 27:72]
  wire [32:0] a_eff = _T_983 | _T_982; // @[Mux.scala 27:72]
  wire [32:0] a_shift = _T_995 & a_eff; // @[exu_div_ctl.scala 177:33]
  wire  _T_1004 = a_ff[32] | rem_correct; // @[exu_div_ctl.scala 181:21]
  reg  divisor_neg_ff; // @[Reg.scala 27:20]
  wire  m_already_comp = divisor_neg_ff & sign_ff; // @[exu_div_ctl.scala 179:48]
  wire  add = _T_1004 ^ m_already_comp; // @[exu_div_ctl.scala 181:36]
  wire [32:0] _T_963 = ~m_ff; // @[exu_div_ctl.scala 169:35]
  wire [32:0] m_eff = add ? m_ff : _T_963; // @[exu_div_ctl.scala 169:15]
  wire [32:0] _T_997 = a_shift + m_eff; // @[exu_div_ctl.scala 178:41]
  wire  _T_998 = ~add; // @[exu_div_ctl.scala 178:65]
  wire [32:0] _T_999 = {32'h0,_T_998}; // @[Cat.scala 29:58]
  wire [32:0] _T_1001 = _T_997 + _T_999; // @[exu_div_ctl.scala 178:49]
  wire [32:0] a_in = _T_995 & _T_1001; // @[exu_div_ctl.scala 178:30]
  wire  _T_719 = ~a_in[32]; // @[exu_div_ctl.scala 162:85]
  wire [32:0] _T_720 = {dividend_eff,_T_719}; // @[Cat.scala 29:58]
  wire [63:0] _GEN_6 = {{31'd0}, _T_720}; // @[exu_div_ctl.scala 162:96]
  wire [63:0] _T_721 = _GEN_6 << shortq_shift_ff; // @[exu_div_ctl.scala 162:96]
  wire  _T_723 = ~_T_714; // @[exu_div_ctl.scala 163:18]
  wire  _T_724 = run_state & _T_723; // @[exu_div_ctl.scala 163:16]
  wire [32:0] _T_729 = {q_ff[31:0],_T_719}; // @[Cat.scala 29:58]
  wire [32:0] _T_730 = _T_711 ? _T_713 : 33'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_731 = _T_715 ? _T_721 : 64'h0; // @[Mux.scala 27:72]
  wire [32:0] _T_732 = _T_724 ? _T_729 : 33'h0; // @[Mux.scala 27:72]
  wire [63:0] _GEN_7 = {{31'd0}, _T_730}; // @[Mux.scala 27:72]
  wire [63:0] _T_733 = _GEN_7 | _T_731; // @[Mux.scala 27:72]
  wire [63:0] _GEN_8 = {{31'd0}, _T_732}; // @[Mux.scala 27:72]
  wire [63:0] _T_734 = _T_733 | _GEN_8; // @[Mux.scala 27:72]
  wire  _T_737 = run_state & _T_697; // @[exu_div_ctl.scala 165:59]
  wire  _T_988 = count != 6'h21; // @[exu_div_ctl.scala 176:84]
  wire  _T_989 = _T_737 & _T_988; // @[exu_div_ctl.scala 176:75]
  wire  _T_990 = io_dec_div_div_p_valid | _T_989; // @[exu_div_ctl.scala 176:45]
  wire  _T_1010 = dividend_neg_ff ^ divisor_neg_ff; // @[exu_div_ctl.scala 183:50]
  wire  _T_1011 = sign_ff & _T_1010; // @[exu_div_ctl.scala 183:31]
  wire [31:0] q_ff_eff = _T_1011 ? _T_959 : q_ff[31:0]; // @[exu_div_ctl.scala 183:21]
  wire  _T_1239 = |a_ff[0]; // @[lib.scala 403:35]
  wire  _T_1241 = ~a_ff[1]; // @[lib.scala 403:40]
  wire  _T_1243 = _T_1239 ? _T_1241 : a_ff[1]; // @[lib.scala 403:23]
  wire  _T_1245 = |a_ff[1:0]; // @[lib.scala 403:35]
  wire  _T_1247 = ~a_ff[2]; // @[lib.scala 403:40]
  wire  _T_1249 = _T_1245 ? _T_1247 : a_ff[2]; // @[lib.scala 403:23]
  wire  _T_1251 = |a_ff[2:0]; // @[lib.scala 403:35]
  wire  _T_1253 = ~a_ff[3]; // @[lib.scala 403:40]
  wire  _T_1255 = _T_1251 ? _T_1253 : a_ff[3]; // @[lib.scala 403:23]
  wire  _T_1257 = |a_ff[3:0]; // @[lib.scala 403:35]
  wire  _T_1259 = ~a_ff[4]; // @[lib.scala 403:40]
  wire  _T_1261 = _T_1257 ? _T_1259 : a_ff[4]; // @[lib.scala 403:23]
  wire  _T_1263 = |a_ff[4:0]; // @[lib.scala 403:35]
  wire  _T_1265 = ~a_ff[5]; // @[lib.scala 403:40]
  wire  _T_1267 = _T_1263 ? _T_1265 : a_ff[5]; // @[lib.scala 403:23]
  wire  _T_1269 = |a_ff[5:0]; // @[lib.scala 403:35]
  wire  _T_1271 = ~a_ff[6]; // @[lib.scala 403:40]
  wire  _T_1273 = _T_1269 ? _T_1271 : a_ff[6]; // @[lib.scala 403:23]
  wire  _T_1275 = |a_ff[6:0]; // @[lib.scala 403:35]
  wire  _T_1277 = ~a_ff[7]; // @[lib.scala 403:40]
  wire  _T_1279 = _T_1275 ? _T_1277 : a_ff[7]; // @[lib.scala 403:23]
  wire  _T_1281 = |a_ff[7:0]; // @[lib.scala 403:35]
  wire  _T_1283 = ~a_ff[8]; // @[lib.scala 403:40]
  wire  _T_1285 = _T_1281 ? _T_1283 : a_ff[8]; // @[lib.scala 403:23]
  wire  _T_1287 = |a_ff[8:0]; // @[lib.scala 403:35]
  wire  _T_1289 = ~a_ff[9]; // @[lib.scala 403:40]
  wire  _T_1291 = _T_1287 ? _T_1289 : a_ff[9]; // @[lib.scala 403:23]
  wire  _T_1293 = |a_ff[9:0]; // @[lib.scala 403:35]
  wire  _T_1295 = ~a_ff[10]; // @[lib.scala 403:40]
  wire  _T_1297 = _T_1293 ? _T_1295 : a_ff[10]; // @[lib.scala 403:23]
  wire  _T_1299 = |a_ff[10:0]; // @[lib.scala 403:35]
  wire  _T_1301 = ~a_ff[11]; // @[lib.scala 403:40]
  wire  _T_1303 = _T_1299 ? _T_1301 : a_ff[11]; // @[lib.scala 403:23]
  wire  _T_1305 = |a_ff[11:0]; // @[lib.scala 403:35]
  wire  _T_1307 = ~a_ff[12]; // @[lib.scala 403:40]
  wire  _T_1309 = _T_1305 ? _T_1307 : a_ff[12]; // @[lib.scala 403:23]
  wire  _T_1311 = |a_ff[12:0]; // @[lib.scala 403:35]
  wire  _T_1313 = ~a_ff[13]; // @[lib.scala 403:40]
  wire  _T_1315 = _T_1311 ? _T_1313 : a_ff[13]; // @[lib.scala 403:23]
  wire  _T_1317 = |a_ff[13:0]; // @[lib.scala 403:35]
  wire  _T_1319 = ~a_ff[14]; // @[lib.scala 403:40]
  wire  _T_1321 = _T_1317 ? _T_1319 : a_ff[14]; // @[lib.scala 403:23]
  wire  _T_1323 = |a_ff[14:0]; // @[lib.scala 403:35]
  wire  _T_1325 = ~a_ff[15]; // @[lib.scala 403:40]
  wire  _T_1327 = _T_1323 ? _T_1325 : a_ff[15]; // @[lib.scala 403:23]
  wire  _T_1329 = |a_ff[15:0]; // @[lib.scala 403:35]
  wire  _T_1331 = ~a_ff[16]; // @[lib.scala 403:40]
  wire  _T_1333 = _T_1329 ? _T_1331 : a_ff[16]; // @[lib.scala 403:23]
  wire  _T_1335 = |a_ff[16:0]; // @[lib.scala 403:35]
  wire  _T_1337 = ~a_ff[17]; // @[lib.scala 403:40]
  wire  _T_1339 = _T_1335 ? _T_1337 : a_ff[17]; // @[lib.scala 403:23]
  wire  _T_1341 = |a_ff[17:0]; // @[lib.scala 403:35]
  wire  _T_1343 = ~a_ff[18]; // @[lib.scala 403:40]
  wire  _T_1345 = _T_1341 ? _T_1343 : a_ff[18]; // @[lib.scala 403:23]
  wire  _T_1347 = |a_ff[18:0]; // @[lib.scala 403:35]
  wire  _T_1349 = ~a_ff[19]; // @[lib.scala 403:40]
  wire  _T_1351 = _T_1347 ? _T_1349 : a_ff[19]; // @[lib.scala 403:23]
  wire  _T_1353 = |a_ff[19:0]; // @[lib.scala 403:35]
  wire  _T_1355 = ~a_ff[20]; // @[lib.scala 403:40]
  wire  _T_1357 = _T_1353 ? _T_1355 : a_ff[20]; // @[lib.scala 403:23]
  wire  _T_1359 = |a_ff[20:0]; // @[lib.scala 403:35]
  wire  _T_1361 = ~a_ff[21]; // @[lib.scala 403:40]
  wire  _T_1363 = _T_1359 ? _T_1361 : a_ff[21]; // @[lib.scala 403:23]
  wire  _T_1365 = |a_ff[21:0]; // @[lib.scala 403:35]
  wire  _T_1367 = ~a_ff[22]; // @[lib.scala 403:40]
  wire  _T_1369 = _T_1365 ? _T_1367 : a_ff[22]; // @[lib.scala 403:23]
  wire  _T_1371 = |a_ff[22:0]; // @[lib.scala 403:35]
  wire  _T_1373 = ~a_ff[23]; // @[lib.scala 403:40]
  wire  _T_1375 = _T_1371 ? _T_1373 : a_ff[23]; // @[lib.scala 403:23]
  wire  _T_1377 = |a_ff[23:0]; // @[lib.scala 403:35]
  wire  _T_1379 = ~a_ff[24]; // @[lib.scala 403:40]
  wire  _T_1381 = _T_1377 ? _T_1379 : a_ff[24]; // @[lib.scala 403:23]
  wire  _T_1383 = |a_ff[24:0]; // @[lib.scala 403:35]
  wire  _T_1385 = ~a_ff[25]; // @[lib.scala 403:40]
  wire  _T_1387 = _T_1383 ? _T_1385 : a_ff[25]; // @[lib.scala 403:23]
  wire  _T_1389 = |a_ff[25:0]; // @[lib.scala 403:35]
  wire  _T_1391 = ~a_ff[26]; // @[lib.scala 403:40]
  wire  _T_1393 = _T_1389 ? _T_1391 : a_ff[26]; // @[lib.scala 403:23]
  wire  _T_1395 = |a_ff[26:0]; // @[lib.scala 403:35]
  wire  _T_1397 = ~a_ff[27]; // @[lib.scala 403:40]
  wire  _T_1399 = _T_1395 ? _T_1397 : a_ff[27]; // @[lib.scala 403:23]
  wire  _T_1401 = |a_ff[27:0]; // @[lib.scala 403:35]
  wire  _T_1403 = ~a_ff[28]; // @[lib.scala 403:40]
  wire  _T_1405 = _T_1401 ? _T_1403 : a_ff[28]; // @[lib.scala 403:23]
  wire  _T_1407 = |a_ff[28:0]; // @[lib.scala 403:35]
  wire  _T_1409 = ~a_ff[29]; // @[lib.scala 403:40]
  wire  _T_1411 = _T_1407 ? _T_1409 : a_ff[29]; // @[lib.scala 403:23]
  wire  _T_1413 = |a_ff[29:0]; // @[lib.scala 403:35]
  wire  _T_1415 = ~a_ff[30]; // @[lib.scala 403:40]
  wire  _T_1417 = _T_1413 ? _T_1415 : a_ff[30]; // @[lib.scala 403:23]
  wire  _T_1419 = |a_ff[30:0]; // @[lib.scala 403:35]
  wire  _T_1421 = ~a_ff[31]; // @[lib.scala 403:40]
  wire  _T_1423 = _T_1419 ? _T_1421 : a_ff[31]; // @[lib.scala 403:23]
  wire [6:0] _T_1429 = {_T_1279,_T_1273,_T_1267,_T_1261,_T_1255,_T_1249,_T_1243}; // @[lib.scala 405:14]
  wire [14:0] _T_1437 = {_T_1327,_T_1321,_T_1315,_T_1309,_T_1303,_T_1297,_T_1291,_T_1285,_T_1429}; // @[lib.scala 405:14]
  wire [7:0] _T_1444 = {_T_1375,_T_1369,_T_1363,_T_1357,_T_1351,_T_1345,_T_1339,_T_1333}; // @[lib.scala 405:14]
  wire [30:0] _T_1453 = {_T_1423,_T_1417,_T_1411,_T_1405,_T_1399,_T_1393,_T_1387,_T_1381,_T_1444,_T_1437}; // @[lib.scala 405:14]
  wire [31:0] _T_1455 = {_T_1453,a_ff[0]}; // @[Cat.scala 29:58]
  wire [31:0] a_ff_eff = _T_738 ? _T_1455 : a_ff[31:0]; // @[exu_div_ctl.scala 184:21]
  reg  smallnum_case_ff; // @[exu_div_ctl.scala 203:32]
  reg [3:0] smallnum_ff; // @[exu_div_ctl.scala 204:27]
  wire [31:0] _T_1458 = {28'h0,smallnum_ff}; // @[Cat.scala 29:58]
  wire  _T_1460 = ~smallnum_case_ff; // @[exu_div_ctl.scala 189:6]
  wire  _T_1462 = _T_1460 & _T_9; // @[exu_div_ctl.scala 189:24]
  wire [31:0] _T_1464 = smallnum_case_ff ? _T_1458 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1465 = rem_ff ? a_ff_eff : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1466 = _T_1462 ? q_ff_eff : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1467 = _T_1464 | _T_1465; // @[Mux.scala 27:72]
  wire  _T_1499 = _T_709 & io_divisor[31]; // @[exu_div_ctl.scala 210:52]
  rvclkhdr rvclkhdr ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_io_l1clk),
    .io_clk(rvclkhdr_io_clk),
    .io_en(rvclkhdr_io_en),
    .io_scan_mode(rvclkhdr_io_scan_mode)
  );
  rvclkhdr rvclkhdr_1 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_1_io_l1clk),
    .io_clk(rvclkhdr_1_io_clk),
    .io_en(rvclkhdr_1_io_en),
    .io_scan_mode(rvclkhdr_1_io_scan_mode)
  );
  rvclkhdr rvclkhdr_2 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_2_io_l1clk),
    .io_clk(rvclkhdr_2_io_clk),
    .io_en(rvclkhdr_2_io_en),
    .io_scan_mode(rvclkhdr_2_io_scan_mode)
  );
  rvclkhdr rvclkhdr_3 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_3_io_l1clk),
    .io_clk(rvclkhdr_3_io_clk),
    .io_en(rvclkhdr_3_io_en),
    .io_scan_mode(rvclkhdr_3_io_scan_mode)
  );
  assign io_exu_div_result = _T_1467 | _T_1466; // @[exu_div_ctl.scala 186:21]
  assign io_exu_div_wren = finish_ff & _T; // @[exu_div_ctl.scala 156:20]
  assign rvclkhdr_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_io_en = _T_688 | finish_ff; // @[lib.scala 345:16]
  assign rvclkhdr_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_1_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_1_io_en = io_dec_div_div_p_valid | _T_737; // @[lib.scala 371:17]
  assign rvclkhdr_1_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_2_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_2_io_en = _T_990 | rem_correct; // @[lib.scala 371:17]
  assign rvclkhdr_2_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_3_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_3_io_en = io_dec_div_div_p_valid; // @[lib.scala 371:17]
  assign rvclkhdr_3_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  valid_ff_x = _RAND_0[0:0];
  _RAND_1 = {2{`RANDOM}};
  q_ff = _RAND_1[32:0];
  _RAND_2 = {2{`RANDOM}};
  m_ff = _RAND_2[32:0];
  _RAND_3 = {1{`RANDOM}};
  rem_ff = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  sign_ff = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  shortq_shift_xx = _RAND_5[3:0];
  _RAND_6 = {1{`RANDOM}};
  count = _RAND_6[5:0];
  _RAND_7 = {1{`RANDOM}};
  run_state = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  finish_ff = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  shortq_enable_ff = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  dividend_neg_ff = _RAND_10[0:0];
  _RAND_11 = {2{`RANDOM}};
  a_ff = _RAND_11[32:0];
  _RAND_12 = {1{`RANDOM}};
  divisor_neg_ff = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  smallnum_case_ff = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  smallnum_ff = _RAND_14[3:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    valid_ff_x = 1'h0;
  end
  if (reset) begin
    q_ff = 33'h0;
  end
  if (reset) begin
    m_ff = 33'h0;
  end
  if (reset) begin
    rem_ff = 1'h0;
  end
  if (reset) begin
    sign_ff = 1'h0;
  end
  if (reset) begin
    shortq_shift_xx = 4'h0;
  end
  if (reset) begin
    count = 6'h0;
  end
  if (reset) begin
    run_state = 1'h0;
  end
  if (reset) begin
    finish_ff = 1'h0;
  end
  if (reset) begin
    shortq_enable_ff = 1'h0;
  end
  if (reset) begin
    dividend_neg_ff = 1'h0;
  end
  if (reset) begin
    a_ff = 33'h0;
  end
  if (reset) begin
    divisor_neg_ff = 1'h0;
  end
  if (reset) begin
    smallnum_case_ff = 1'h0;
  end
  if (reset) begin
    smallnum_ff = 4'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge rvclkhdr_io_l1clk or posedge reset) begin
    if (reset) begin
      valid_ff_x <= 1'h0;
    end else begin
      valid_ff_x <= io_dec_div_div_p_valid & _T;
    end
  end
  always @(posedge rvclkhdr_1_io_l1clk or posedge reset) begin
    if (reset) begin
      q_ff <= 33'h0;
    end else begin
      q_ff <= _T_734[32:0];
    end
  end
  always @(posedge rvclkhdr_3_io_l1clk or posedge reset) begin
    if (reset) begin
      m_ff <= 33'h0;
    end else begin
      m_ff <= {_T_1499,io_divisor};
    end
  end
  always @(posedge rvclkhdr_io_l1clk or posedge reset) begin
    if (reset) begin
      rem_ff <= 1'h0;
    end else if (io_dec_div_div_p_valid) begin
      rem_ff <= io_dec_div_div_p_bits_rem;
    end
  end
  always @(posedge rvclkhdr_io_l1clk or posedge reset) begin
    if (reset) begin
      sign_ff <= 1'h0;
    end else if (io_dec_div_div_p_valid) begin
      sign_ff <= sign_eff;
    end
  end
  always @(posedge rvclkhdr_io_l1clk or posedge reset) begin
    if (reset) begin
      shortq_shift_xx <= 4'h0;
    end else begin
      shortq_shift_xx <= _T_667 & shortq_raw;
    end
  end
  always @(posedge rvclkhdr_io_l1clk or posedge reset) begin
    if (reset) begin
      count <= 6'h0;
    end else begin
      count <= _T_700 & _T_705;
    end
  end
  always @(posedge rvclkhdr_io_l1clk or posedge reset) begin
    if (reset) begin
      run_state <= 1'h0;
    end else begin
      run_state <= _T_691 & _T;
    end
  end
  always @(posedge rvclkhdr_io_l1clk or posedge reset) begin
    if (reset) begin
      finish_ff <= 1'h0;
    end else begin
      finish_ff <= finish & _T;
    end
  end
  always @(posedge rvclkhdr_io_l1clk or posedge reset) begin
    if (reset) begin
      shortq_enable_ff <= 1'h0;
    end else begin
      shortq_enable_ff <= _T_664 & _T_665;
    end
  end
  always @(posedge rvclkhdr_io_l1clk or posedge reset) begin
    if (reset) begin
      dividend_neg_ff <= 1'h0;
    end else if (io_dec_div_div_p_valid) begin
      dividend_neg_ff <= io_dividend[31];
    end
  end
  always @(posedge rvclkhdr_2_io_l1clk or posedge reset) begin
    if (reset) begin
      a_ff <= 33'h0;
    end else begin
      a_ff <= _T_995 & _T_1001;
    end
  end
  always @(posedge rvclkhdr_io_l1clk or posedge reset) begin
    if (reset) begin
      divisor_neg_ff <= 1'h0;
    end else if (io_dec_div_div_p_valid) begin
      divisor_neg_ff <= io_divisor[31];
    end
  end
  always @(posedge rvclkhdr_io_l1clk or posedge reset) begin
    if (reset) begin
      smallnum_case_ff <= 1'h0;
    end else begin
      smallnum_case_ff <= _T_11 | _T_19;
    end
  end
  always @(posedge rvclkhdr_io_l1clk or posedge reset) begin
    if (reset) begin
      smallnum_ff <= 4'h0;
    end else begin
      smallnum_ff <= {_T_477,_T_476};
    end
  end
endmodule
module exu(
  input         clock,
  input         reset,
  input         io_scan_mode,
  input         io_dec_exu_dec_alu_dec_i0_alu_decode_d,
  input         io_dec_exu_dec_alu_dec_csr_ren_d,
  input  [11:0] io_dec_exu_dec_alu_dec_i0_br_immed_d,
  output [30:0] io_dec_exu_dec_alu_exu_i0_pc_x,
  input         io_dec_exu_dec_div_div_p_valid,
  input         io_dec_exu_dec_div_div_p_bits_unsign,
  input         io_dec_exu_dec_div_div_p_bits_rem,
  input         io_dec_exu_dec_div_dec_div_cancel,
  input  [1:0]  io_dec_exu_decode_exu_dec_data_en,
  input  [1:0]  io_dec_exu_decode_exu_dec_ctl_en,
  input         io_dec_exu_decode_exu_i0_ap_land,
  input         io_dec_exu_decode_exu_i0_ap_lor,
  input         io_dec_exu_decode_exu_i0_ap_lxor,
  input         io_dec_exu_decode_exu_i0_ap_sll,
  input         io_dec_exu_decode_exu_i0_ap_srl,
  input         io_dec_exu_decode_exu_i0_ap_sra,
  input         io_dec_exu_decode_exu_i0_ap_beq,
  input         io_dec_exu_decode_exu_i0_ap_bne,
  input         io_dec_exu_decode_exu_i0_ap_blt,
  input         io_dec_exu_decode_exu_i0_ap_bge,
  input         io_dec_exu_decode_exu_i0_ap_add,
  input         io_dec_exu_decode_exu_i0_ap_sub,
  input         io_dec_exu_decode_exu_i0_ap_slt,
  input         io_dec_exu_decode_exu_i0_ap_unsign,
  input         io_dec_exu_decode_exu_i0_ap_jal,
  input         io_dec_exu_decode_exu_i0_ap_predict_t,
  input         io_dec_exu_decode_exu_i0_ap_predict_nt,
  input         io_dec_exu_decode_exu_i0_ap_csr_write,
  input         io_dec_exu_decode_exu_i0_ap_csr_imm,
  input         io_dec_exu_decode_exu_dec_i0_predict_p_d_valid,
  input         io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_pc4,
  input  [1:0]  io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_hist,
  input  [11:0] io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_toffset,
  input         io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_br_error,
  input         io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_br_start_error,
  input  [30:0] io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_prett,
  input         io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_pcall,
  input         io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_pret,
  input         io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_pja,
  input         io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_way,
  input  [7:0]  io_dec_exu_decode_exu_i0_predict_fghr_d,
  input  [7:0]  io_dec_exu_decode_exu_i0_predict_index_d,
  input  [4:0]  io_dec_exu_decode_exu_i0_predict_btag_d,
  input         io_dec_exu_decode_exu_dec_i0_rs1_en_d,
  input         io_dec_exu_decode_exu_dec_i0_rs2_en_d,
  input  [31:0] io_dec_exu_decode_exu_dec_i0_immed_d,
  input  [31:0] io_dec_exu_decode_exu_dec_i0_rs1_bypass_data_d,
  input  [31:0] io_dec_exu_decode_exu_dec_i0_rs2_bypass_data_d,
  input         io_dec_exu_decode_exu_dec_i0_select_pc_d,
  input  [1:0]  io_dec_exu_decode_exu_dec_i0_rs1_bypass_en_d,
  input  [1:0]  io_dec_exu_decode_exu_dec_i0_rs2_bypass_en_d,
  input         io_dec_exu_decode_exu_mul_p_valid,
  input         io_dec_exu_decode_exu_mul_p_bits_rs1_sign,
  input         io_dec_exu_decode_exu_mul_p_bits_rs2_sign,
  input         io_dec_exu_decode_exu_mul_p_bits_low,
  input  [30:0] io_dec_exu_decode_exu_pred_correct_npc_x,
  input         io_dec_exu_decode_exu_dec_extint_stall,
  output [31:0] io_dec_exu_decode_exu_exu_i0_result_x,
  output [31:0] io_dec_exu_decode_exu_exu_csr_rs1_x,
  input  [29:0] io_dec_exu_tlu_exu_dec_tlu_meihap,
  input         io_dec_exu_tlu_exu_dec_tlu_flush_lower_r,
  input  [30:0] io_dec_exu_tlu_exu_dec_tlu_flush_path_r,
  output [1:0]  io_dec_exu_tlu_exu_exu_i0_br_hist_r,
  output        io_dec_exu_tlu_exu_exu_i0_br_error_r,
  output        io_dec_exu_tlu_exu_exu_i0_br_start_error_r,
  output [7:0]  io_dec_exu_tlu_exu_exu_i0_br_index_r,
  output        io_dec_exu_tlu_exu_exu_i0_br_valid_r,
  output        io_dec_exu_tlu_exu_exu_i0_br_mp_r,
  output        io_dec_exu_tlu_exu_exu_i0_br_middle_r,
  output        io_dec_exu_tlu_exu_exu_pmu_i0_br_misp,
  output        io_dec_exu_tlu_exu_exu_pmu_i0_br_ataken,
  output        io_dec_exu_tlu_exu_exu_pmu_i0_pc4,
  output [30:0] io_dec_exu_tlu_exu_exu_npc_r,
  input  [30:0] io_dec_exu_ib_exu_dec_i0_pc_d,
  input         io_dec_exu_ib_exu_dec_debug_wdata_rs1_d,
  input  [31:0] io_dec_exu_gpr_exu_gpr_i0_rs1_d,
  input  [31:0] io_dec_exu_gpr_exu_gpr_i0_rs2_d,
  output [7:0]  io_exu_bp_exu_i0_br_fghr_r,
  output        io_exu_bp_exu_i0_br_way_r,
  output        io_exu_bp_exu_mp_pkt_bits_misp,
  output        io_exu_bp_exu_mp_pkt_bits_ataken,
  output        io_exu_bp_exu_mp_pkt_bits_boffset,
  output        io_exu_bp_exu_mp_pkt_bits_pc4,
  output [1:0]  io_exu_bp_exu_mp_pkt_bits_hist,
  output [11:0] io_exu_bp_exu_mp_pkt_bits_toffset,
  output        io_exu_bp_exu_mp_pkt_bits_pcall,
  output        io_exu_bp_exu_mp_pkt_bits_pret,
  output        io_exu_bp_exu_mp_pkt_bits_pja,
  output        io_exu_bp_exu_mp_pkt_bits_way,
  output [7:0]  io_exu_bp_exu_mp_eghr,
  output [7:0]  io_exu_bp_exu_mp_fghr,
  output [7:0]  io_exu_bp_exu_mp_index,
  output [4:0]  io_exu_bp_exu_mp_btag,
  output        io_exu_flush_final,
  output [31:0] io_exu_div_result,
  output        io_exu_div_wren,
  input  [31:0] io_dbg_cmd_wrdata,
  output [31:0] io_lsu_exu_exu_lsu_rs1_d,
  output [31:0] io_lsu_exu_exu_lsu_rs2_d,
  output [30:0] io_exu_flush_path_final
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
`endif // RANDOMIZE_REG_INIT
  wire  rvclkhdr_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_1_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_1_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_1_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_1_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_2_io_l1clk; // @[lib.scala 378:23]
  wire  rvclkhdr_2_io_clk; // @[lib.scala 378:23]
  wire  rvclkhdr_2_io_en; // @[lib.scala 378:23]
  wire  rvclkhdr_2_io_scan_mode; // @[lib.scala 378:23]
  wire  rvclkhdr_3_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_3_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_3_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_3_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_4_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_4_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_4_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_4_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_5_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_5_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_5_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_5_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_6_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_6_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_6_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_6_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_7_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_7_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_7_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_7_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_8_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_8_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_8_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_8_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_9_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_9_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_9_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_9_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_10_io_l1clk; // @[lib.scala 378:23]
  wire  rvclkhdr_10_io_clk; // @[lib.scala 378:23]
  wire  rvclkhdr_10_io_en; // @[lib.scala 378:23]
  wire  rvclkhdr_10_io_scan_mode; // @[lib.scala 378:23]
  wire  rvclkhdr_11_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_11_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_11_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_11_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_12_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_12_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_12_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_12_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_13_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_13_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_13_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_13_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_14_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_14_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_14_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_14_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_15_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_15_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_15_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_15_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_16_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_16_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_16_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_16_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_17_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_17_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_17_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_17_io_scan_mode; // @[lib.scala 368:23]
  wire  i_alu_clock; // @[exu.scala 144:19]
  wire  i_alu_reset; // @[exu.scala 144:19]
  wire  i_alu_io_dec_alu_dec_i0_alu_decode_d; // @[exu.scala 144:19]
  wire  i_alu_io_dec_alu_dec_csr_ren_d; // @[exu.scala 144:19]
  wire [11:0] i_alu_io_dec_alu_dec_i0_br_immed_d; // @[exu.scala 144:19]
  wire [30:0] i_alu_io_dec_alu_exu_i0_pc_x; // @[exu.scala 144:19]
  wire [30:0] i_alu_io_dec_i0_pc_d; // @[exu.scala 144:19]
  wire  i_alu_io_scan_mode; // @[exu.scala 144:19]
  wire  i_alu_io_flush_upper_x; // @[exu.scala 144:19]
  wire  i_alu_io_dec_tlu_flush_lower_r; // @[exu.scala 144:19]
  wire  i_alu_io_enable; // @[exu.scala 144:19]
  wire  i_alu_io_i0_ap_land; // @[exu.scala 144:19]
  wire  i_alu_io_i0_ap_lor; // @[exu.scala 144:19]
  wire  i_alu_io_i0_ap_lxor; // @[exu.scala 144:19]
  wire  i_alu_io_i0_ap_sll; // @[exu.scala 144:19]
  wire  i_alu_io_i0_ap_srl; // @[exu.scala 144:19]
  wire  i_alu_io_i0_ap_sra; // @[exu.scala 144:19]
  wire  i_alu_io_i0_ap_beq; // @[exu.scala 144:19]
  wire  i_alu_io_i0_ap_bne; // @[exu.scala 144:19]
  wire  i_alu_io_i0_ap_blt; // @[exu.scala 144:19]
  wire  i_alu_io_i0_ap_bge; // @[exu.scala 144:19]
  wire  i_alu_io_i0_ap_add; // @[exu.scala 144:19]
  wire  i_alu_io_i0_ap_sub; // @[exu.scala 144:19]
  wire  i_alu_io_i0_ap_slt; // @[exu.scala 144:19]
  wire  i_alu_io_i0_ap_unsign; // @[exu.scala 144:19]
  wire  i_alu_io_i0_ap_jal; // @[exu.scala 144:19]
  wire  i_alu_io_i0_ap_predict_t; // @[exu.scala 144:19]
  wire  i_alu_io_i0_ap_predict_nt; // @[exu.scala 144:19]
  wire  i_alu_io_i0_ap_csr_write; // @[exu.scala 144:19]
  wire  i_alu_io_i0_ap_csr_imm; // @[exu.scala 144:19]
  wire [31:0] i_alu_io_a_in; // @[exu.scala 144:19]
  wire [31:0] i_alu_io_b_in; // @[exu.scala 144:19]
  wire  i_alu_io_pp_in_valid; // @[exu.scala 144:19]
  wire  i_alu_io_pp_in_bits_boffset; // @[exu.scala 144:19]
  wire  i_alu_io_pp_in_bits_pc4; // @[exu.scala 144:19]
  wire [1:0] i_alu_io_pp_in_bits_hist; // @[exu.scala 144:19]
  wire [11:0] i_alu_io_pp_in_bits_toffset; // @[exu.scala 144:19]
  wire  i_alu_io_pp_in_bits_br_error; // @[exu.scala 144:19]
  wire  i_alu_io_pp_in_bits_br_start_error; // @[exu.scala 144:19]
  wire [30:0] i_alu_io_pp_in_bits_prett; // @[exu.scala 144:19]
  wire  i_alu_io_pp_in_bits_pcall; // @[exu.scala 144:19]
  wire  i_alu_io_pp_in_bits_pret; // @[exu.scala 144:19]
  wire  i_alu_io_pp_in_bits_pja; // @[exu.scala 144:19]
  wire  i_alu_io_pp_in_bits_way; // @[exu.scala 144:19]
  wire [31:0] i_alu_io_result_ff; // @[exu.scala 144:19]
  wire  i_alu_io_flush_upper_out; // @[exu.scala 144:19]
  wire  i_alu_io_flush_final_out; // @[exu.scala 144:19]
  wire [30:0] i_alu_io_flush_path_out; // @[exu.scala 144:19]
  wire  i_alu_io_pred_correct_out; // @[exu.scala 144:19]
  wire  i_alu_io_predict_p_out_valid; // @[exu.scala 144:19]
  wire  i_alu_io_predict_p_out_bits_misp; // @[exu.scala 144:19]
  wire  i_alu_io_predict_p_out_bits_ataken; // @[exu.scala 144:19]
  wire  i_alu_io_predict_p_out_bits_boffset; // @[exu.scala 144:19]
  wire  i_alu_io_predict_p_out_bits_pc4; // @[exu.scala 144:19]
  wire [1:0] i_alu_io_predict_p_out_bits_hist; // @[exu.scala 144:19]
  wire [11:0] i_alu_io_predict_p_out_bits_toffset; // @[exu.scala 144:19]
  wire  i_alu_io_predict_p_out_bits_br_error; // @[exu.scala 144:19]
  wire  i_alu_io_predict_p_out_bits_br_start_error; // @[exu.scala 144:19]
  wire  i_alu_io_predict_p_out_bits_pcall; // @[exu.scala 144:19]
  wire  i_alu_io_predict_p_out_bits_pret; // @[exu.scala 144:19]
  wire  i_alu_io_predict_p_out_bits_pja; // @[exu.scala 144:19]
  wire  i_alu_io_predict_p_out_bits_way; // @[exu.scala 144:19]
  wire  i_mul_clock; // @[exu.scala 162:19]
  wire  i_mul_reset; // @[exu.scala 162:19]
  wire  i_mul_io_scan_mode; // @[exu.scala 162:19]
  wire  i_mul_io_mul_p_valid; // @[exu.scala 162:19]
  wire  i_mul_io_mul_p_bits_rs1_sign; // @[exu.scala 162:19]
  wire  i_mul_io_mul_p_bits_rs2_sign; // @[exu.scala 162:19]
  wire  i_mul_io_mul_p_bits_low; // @[exu.scala 162:19]
  wire [31:0] i_mul_io_rs1_in; // @[exu.scala 162:19]
  wire [31:0] i_mul_io_rs2_in; // @[exu.scala 162:19]
  wire [31:0] i_mul_io_result_x; // @[exu.scala 162:19]
  wire  i_div_clock; // @[exu.scala 169:19]
  wire  i_div_reset; // @[exu.scala 169:19]
  wire  i_div_io_scan_mode; // @[exu.scala 169:19]
  wire [31:0] i_div_io_dividend; // @[exu.scala 169:19]
  wire [31:0] i_div_io_divisor; // @[exu.scala 169:19]
  wire [31:0] i_div_io_exu_div_result; // @[exu.scala 169:19]
  wire  i_div_io_exu_div_wren; // @[exu.scala 169:19]
  wire  i_div_io_dec_div_div_p_valid; // @[exu.scala 169:19]
  wire  i_div_io_dec_div_div_p_bits_unsign; // @[exu.scala 169:19]
  wire  i_div_io_dec_div_div_p_bits_rem; // @[exu.scala 169:19]
  wire  i_div_io_dec_div_dec_div_cancel; // @[exu.scala 169:19]
  wire [15:0] _T = {io_dec_exu_decode_exu_i0_predict_fghr_d,io_dec_exu_decode_exu_i0_predict_index_d}; // @[Cat.scala 29:58]
  reg [30:0] i0_flush_path_x; // @[lib.scala 374:16]
  reg [31:0] _T_3; // @[lib.scala 374:16]
  reg  i0_predict_p_x_valid; // @[lib.scala 384:16]
  reg  i0_predict_p_x_bits_misp; // @[lib.scala 384:16]
  reg  i0_predict_p_x_bits_ataken; // @[lib.scala 384:16]
  reg  i0_predict_p_x_bits_boffset; // @[lib.scala 384:16]
  reg  i0_predict_p_x_bits_pc4; // @[lib.scala 384:16]
  reg [1:0] i0_predict_p_x_bits_hist; // @[lib.scala 384:16]
  reg [11:0] i0_predict_p_x_bits_toffset; // @[lib.scala 384:16]
  reg  i0_predict_p_x_bits_br_error; // @[lib.scala 384:16]
  reg  i0_predict_p_x_bits_br_start_error; // @[lib.scala 384:16]
  reg  i0_predict_p_x_bits_pcall; // @[lib.scala 384:16]
  reg  i0_predict_p_x_bits_pret; // @[lib.scala 384:16]
  reg  i0_predict_p_x_bits_pja; // @[lib.scala 384:16]
  reg  i0_predict_p_x_bits_way; // @[lib.scala 384:16]
  reg [20:0] predpipe_x; // @[lib.scala 374:16]
  reg [20:0] predpipe_r; // @[lib.scala 374:16]
  reg [7:0] ghr_x; // @[lib.scala 374:16]
  reg  i0_pred_correct_upper_x; // @[lib.scala 374:16]
  reg  i0_flush_upper_x; // @[lib.scala 374:16]
  reg  i0_taken_x; // @[lib.scala 374:16]
  reg  i0_valid_x; // @[lib.scala 374:16]
  reg  i0_pp_r_valid; // @[lib.scala 384:16]
  reg  i0_pp_r_bits_misp; // @[lib.scala 384:16]
  reg  i0_pp_r_bits_ataken; // @[lib.scala 384:16]
  reg  i0_pp_r_bits_boffset; // @[lib.scala 384:16]
  reg  i0_pp_r_bits_pc4; // @[lib.scala 384:16]
  reg [1:0] i0_pp_r_bits_hist; // @[lib.scala 384:16]
  reg  i0_pp_r_bits_br_error; // @[lib.scala 384:16]
  reg  i0_pp_r_bits_br_start_error; // @[lib.scala 384:16]
  reg  i0_pp_r_bits_way; // @[lib.scala 384:16]
  reg [5:0] pred_temp1; // @[lib.scala 374:16]
  reg  i0_pred_correct_upper_r; // @[lib.scala 374:16]
  reg [30:0] i0_flush_path_upper_r; // @[lib.scala 374:16]
  reg [24:0] pred_temp2; // @[lib.scala 374:16]
  wire [30:0] _T_23 = {pred_temp2,pred_temp1}; // @[Cat.scala 29:58]
  wire  _T_149 = ~io_dec_exu_tlu_exu_dec_tlu_flush_lower_r; // @[exu.scala 194:6]
  wire  i0_predict_p_d_valid = i_alu_io_predict_p_out_valid; // @[exu.scala 43:53 exu.scala 159:41]
  wire  _T_145 = i0_predict_p_d_valid & io_dec_exu_dec_alu_dec_i0_alu_decode_d; // @[exu.scala 187:54]
  wire  i0_valid_d = _T_145 & _T_149; // @[exu.scala 187:95]
  wire  _T_150 = _T_149 & i0_valid_d; // @[exu.scala 194:48]
  reg [7:0] ghr_d; // @[lib.scala 374:16]
  wire  i0_predict_p_d_bits_ataken = i_alu_io_predict_p_out_bits_ataken; // @[exu.scala 43:53 exu.scala 159:41]
  wire  i0_taken_d = i0_predict_p_d_bits_ataken & io_dec_exu_dec_alu_dec_i0_alu_decode_d; // @[exu.scala 188:59]
  wire [7:0] _T_153 = {ghr_d[6:0],i0_taken_d}; // @[Cat.scala 29:58]
  wire [7:0] _T_159 = _T_150 ? _T_153 : 8'h0; // @[Mux.scala 27:72]
  wire  _T_155 = ~i0_valid_d; // @[exu.scala 195:50]
  wire  _T_156 = _T_149 & _T_155; // @[exu.scala 195:48]
  wire [7:0] _T_160 = _T_156 ? ghr_d : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_162 = _T_159 | _T_160; // @[Mux.scala 27:72]
  wire [7:0] _T_161 = io_dec_exu_tlu_exu_dec_tlu_flush_lower_r ? ghr_x : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] ghr_d_ns = _T_162 | _T_161; // @[Mux.scala 27:72]
  wire  _T_39 = ghr_d_ns != ghr_d; // @[exu.scala 91:39]
  reg  mul_valid_x; // @[lib.scala 374:16]
  wire  _T_40 = io_dec_exu_decode_exu_mul_p_valid != mul_valid_x; // @[exu.scala 91:89]
  wire  _T_41 = _T_39 | _T_40; // @[exu.scala 91:50]
  reg  flush_lower_ff; // @[lib.scala 374:16]
  wire  _T_42 = io_dec_exu_tlu_exu_dec_tlu_flush_lower_r != flush_lower_ff; // @[exu.scala 91:151]
  wire  i0_rs1_bypass_en_d = io_dec_exu_decode_exu_dec_i0_rs1_bypass_en_d[0] | io_dec_exu_decode_exu_dec_i0_rs1_bypass_en_d[1]; // @[exu.scala 92:84]
  wire  i0_rs2_bypass_en_d = io_dec_exu_decode_exu_dec_i0_rs2_bypass_en_d[0] | io_dec_exu_decode_exu_dec_i0_rs2_bypass_en_d[1]; // @[exu.scala 93:84]
  wire [31:0] _T_52 = io_dec_exu_decode_exu_dec_i0_rs1_bypass_en_d[0] ? io_dec_exu_decode_exu_dec_i0_rs1_bypass_data_d : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_53 = io_dec_exu_decode_exu_dec_i0_rs1_bypass_en_d[1] ? io_dec_exu_decode_exu_exu_i0_result_x : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] i0_rs1_bypass_data_d = _T_52 | _T_53; // @[Mux.scala 27:72]
  wire [31:0] _T_59 = io_dec_exu_decode_exu_dec_i0_rs2_bypass_en_d[0] ? io_dec_exu_decode_exu_dec_i0_rs2_bypass_data_d : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_60 = io_dec_exu_decode_exu_dec_i0_rs2_bypass_en_d[1] ? io_dec_exu_decode_exu_exu_i0_result_x : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] i0_rs2_bypass_data_d = _T_59 | _T_60; // @[Mux.scala 27:72]
  wire  _T_63 = ~i0_rs1_bypass_en_d; // @[exu.scala 107:6]
  wire  _T_64 = _T_63 & io_dec_exu_decode_exu_dec_i0_select_pc_d; // @[exu.scala 107:26]
  wire [31:0] _T_66 = {io_dec_exu_ib_exu_dec_i0_pc_d,1'h0}; // @[Cat.scala 29:58]
  wire  _T_68 = _T_63 & io_dec_exu_ib_exu_dec_debug_wdata_rs1_d; // @[exu.scala 108:26]
  wire  _T_71 = ~io_dec_exu_ib_exu_dec_debug_wdata_rs1_d; // @[exu.scala 109:28]
  wire  _T_72 = _T_63 & _T_71; // @[exu.scala 109:26]
  wire  _T_73 = _T_72 & io_dec_exu_decode_exu_dec_i0_rs1_en_d; // @[exu.scala 109:69]
  wire [31:0] _T_75 = i0_rs1_bypass_en_d ? i0_rs1_bypass_data_d : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_76 = _T_64 ? _T_66 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_77 = _T_68 ? io_dbg_cmd_wrdata : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_78 = _T_73 ? io_dec_exu_gpr_exu_gpr_i0_rs1_d : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_79 = _T_75 | _T_76; // @[Mux.scala 27:72]
  wire [31:0] _T_80 = _T_79 | _T_77; // @[Mux.scala 27:72]
  wire [31:0] i0_rs1_d = _T_80 | _T_78; // @[Mux.scala 27:72]
  wire  _T_82 = ~i0_rs2_bypass_en_d; // @[exu.scala 113:6]
  wire  _T_83 = _T_82 & io_dec_exu_decode_exu_dec_i0_rs2_en_d; // @[exu.scala 113:26]
  wire [31:0] _T_88 = _T_83 ? io_dec_exu_gpr_exu_gpr_i0_rs2_d : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_89 = _T_82 ? io_dec_exu_decode_exu_dec_i0_immed_d : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_90 = i0_rs2_bypass_en_d ? i0_rs2_bypass_data_d : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_91 = _T_88 | _T_89; // @[Mux.scala 27:72]
  wire [31:0] _T_92 = _T_91 | _T_90; // @[Mux.scala 27:72]
  wire  _T_94 = ~io_dec_exu_decode_exu_dec_extint_stall; // @[exu.scala 120:28]
  wire  _T_95 = _T_63 & _T_94; // @[exu.scala 120:26]
  wire  _T_96 = _T_95 & io_dec_exu_decode_exu_dec_i0_rs1_en_d; // @[exu.scala 120:68]
  wire  _T_99 = i0_rs1_bypass_en_d & _T_94; // @[exu.scala 121:25]
  wire [31:0] _T_102 = {io_dec_exu_tlu_exu_dec_tlu_meihap,2'h0}; // @[Cat.scala 29:58]
  wire [31:0] _T_103 = _T_96 ? io_dec_exu_gpr_exu_gpr_i0_rs1_d : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_104 = _T_99 ? i0_rs1_bypass_data_d : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_105 = io_dec_exu_decode_exu_dec_extint_stall ? _T_102 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_106 = _T_103 | _T_104; // @[Mux.scala 27:72]
  wire  _T_111 = _T_82 & _T_94; // @[exu.scala 126:26]
  wire  _T_112 = _T_111 & io_dec_exu_decode_exu_dec_i0_rs2_en_d; // @[exu.scala 126:68]
  wire  _T_115 = i0_rs2_bypass_en_d & _T_94; // @[exu.scala 127:25]
  wire [31:0] _T_117 = _T_112 ? io_dec_exu_gpr_exu_gpr_i0_rs2_d : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_118 = _T_115 ? i0_rs2_bypass_data_d : 32'h0; // @[Mux.scala 27:72]
  wire  _T_122 = _T_63 & io_dec_exu_decode_exu_dec_i0_rs1_en_d; // @[exu.scala 131:26]
  wire [31:0] _T_125 = _T_122 ? io_dec_exu_gpr_exu_gpr_i0_rs1_d : 32'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_167 = {ghr_x[6:0],i0_taken_x}; // @[Cat.scala 29:58]
  wire [20:0] final_predpipe_mp = i0_flush_upper_x ? predpipe_x : 21'h0; // @[exu.scala 213:49]
  wire  _T_179 = i0_flush_upper_x & _T_149; // @[exu.scala 215:67]
  wire [30:0] i0_flush_path_d = i_alu_io_flush_path_out; // @[exu.scala 42:53 exu.scala 157:41]
  wire [31:0] pred_correct_npc_r = {{1'd0}, _T_23}; // @[exu.scala 47:51 exu.scala 78:41]
  wire [31:0] _T_188 = i0_pred_correct_upper_r ? pred_correct_npc_r : {{1'd0}, i0_flush_path_upper_r}; // @[exu.scala 233:72]
  wire [31:0] i0_rs2_d = _T_92; // @[Mux.scala 27:72 Mux.scala 27:72]
  rvclkhdr rvclkhdr ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_io_l1clk),
    .io_clk(rvclkhdr_io_clk),
    .io_en(rvclkhdr_io_en),
    .io_scan_mode(rvclkhdr_io_scan_mode)
  );
  rvclkhdr rvclkhdr_1 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_1_io_l1clk),
    .io_clk(rvclkhdr_1_io_clk),
    .io_en(rvclkhdr_1_io_en),
    .io_scan_mode(rvclkhdr_1_io_scan_mode)
  );
  rvclkhdr rvclkhdr_2 ( // @[lib.scala 378:23]
    .io_l1clk(rvclkhdr_2_io_l1clk),
    .io_clk(rvclkhdr_2_io_clk),
    .io_en(rvclkhdr_2_io_en),
    .io_scan_mode(rvclkhdr_2_io_scan_mode)
  );
  rvclkhdr rvclkhdr_3 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_3_io_l1clk),
    .io_clk(rvclkhdr_3_io_clk),
    .io_en(rvclkhdr_3_io_en),
    .io_scan_mode(rvclkhdr_3_io_scan_mode)
  );
  rvclkhdr rvclkhdr_4 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_4_io_l1clk),
    .io_clk(rvclkhdr_4_io_clk),
    .io_en(rvclkhdr_4_io_en),
    .io_scan_mode(rvclkhdr_4_io_scan_mode)
  );
  rvclkhdr rvclkhdr_5 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_5_io_l1clk),
    .io_clk(rvclkhdr_5_io_clk),
    .io_en(rvclkhdr_5_io_en),
    .io_scan_mode(rvclkhdr_5_io_scan_mode)
  );
  rvclkhdr rvclkhdr_6 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_6_io_l1clk),
    .io_clk(rvclkhdr_6_io_clk),
    .io_en(rvclkhdr_6_io_en),
    .io_scan_mode(rvclkhdr_6_io_scan_mode)
  );
  rvclkhdr rvclkhdr_7 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_7_io_l1clk),
    .io_clk(rvclkhdr_7_io_clk),
    .io_en(rvclkhdr_7_io_en),
    .io_scan_mode(rvclkhdr_7_io_scan_mode)
  );
  rvclkhdr rvclkhdr_8 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_8_io_l1clk),
    .io_clk(rvclkhdr_8_io_clk),
    .io_en(rvclkhdr_8_io_en),
    .io_scan_mode(rvclkhdr_8_io_scan_mode)
  );
  rvclkhdr rvclkhdr_9 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_9_io_l1clk),
    .io_clk(rvclkhdr_9_io_clk),
    .io_en(rvclkhdr_9_io_en),
    .io_scan_mode(rvclkhdr_9_io_scan_mode)
  );
  rvclkhdr rvclkhdr_10 ( // @[lib.scala 378:23]
    .io_l1clk(rvclkhdr_10_io_l1clk),
    .io_clk(rvclkhdr_10_io_clk),
    .io_en(rvclkhdr_10_io_en),
    .io_scan_mode(rvclkhdr_10_io_scan_mode)
  );
  rvclkhdr rvclkhdr_11 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_11_io_l1clk),
    .io_clk(rvclkhdr_11_io_clk),
    .io_en(rvclkhdr_11_io_en),
    .io_scan_mode(rvclkhdr_11_io_scan_mode)
  );
  rvclkhdr rvclkhdr_12 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_12_io_l1clk),
    .io_clk(rvclkhdr_12_io_clk),
    .io_en(rvclkhdr_12_io_en),
    .io_scan_mode(rvclkhdr_12_io_scan_mode)
  );
  rvclkhdr rvclkhdr_13 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_13_io_l1clk),
    .io_clk(rvclkhdr_13_io_clk),
    .io_en(rvclkhdr_13_io_en),
    .io_scan_mode(rvclkhdr_13_io_scan_mode)
  );
  rvclkhdr rvclkhdr_14 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_14_io_l1clk),
    .io_clk(rvclkhdr_14_io_clk),
    .io_en(rvclkhdr_14_io_en),
    .io_scan_mode(rvclkhdr_14_io_scan_mode)
  );
  rvclkhdr rvclkhdr_15 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_15_io_l1clk),
    .io_clk(rvclkhdr_15_io_clk),
    .io_en(rvclkhdr_15_io_en),
    .io_scan_mode(rvclkhdr_15_io_scan_mode)
  );
  rvclkhdr rvclkhdr_16 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_16_io_l1clk),
    .io_clk(rvclkhdr_16_io_clk),
    .io_en(rvclkhdr_16_io_en),
    .io_scan_mode(rvclkhdr_16_io_scan_mode)
  );
  rvclkhdr rvclkhdr_17 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_17_io_l1clk),
    .io_clk(rvclkhdr_17_io_clk),
    .io_en(rvclkhdr_17_io_en),
    .io_scan_mode(rvclkhdr_17_io_scan_mode)
  );
  exu_alu_ctl i_alu ( // @[exu.scala 144:19]
    .clock(i_alu_clock),
    .reset(i_alu_reset),
    .io_dec_alu_dec_i0_alu_decode_d(i_alu_io_dec_alu_dec_i0_alu_decode_d),
    .io_dec_alu_dec_csr_ren_d(i_alu_io_dec_alu_dec_csr_ren_d),
    .io_dec_alu_dec_i0_br_immed_d(i_alu_io_dec_alu_dec_i0_br_immed_d),
    .io_dec_alu_exu_i0_pc_x(i_alu_io_dec_alu_exu_i0_pc_x),
    .io_dec_i0_pc_d(i_alu_io_dec_i0_pc_d),
    .io_scan_mode(i_alu_io_scan_mode),
    .io_flush_upper_x(i_alu_io_flush_upper_x),
    .io_dec_tlu_flush_lower_r(i_alu_io_dec_tlu_flush_lower_r),
    .io_enable(i_alu_io_enable),
    .io_i0_ap_land(i_alu_io_i0_ap_land),
    .io_i0_ap_lor(i_alu_io_i0_ap_lor),
    .io_i0_ap_lxor(i_alu_io_i0_ap_lxor),
    .io_i0_ap_sll(i_alu_io_i0_ap_sll),
    .io_i0_ap_srl(i_alu_io_i0_ap_srl),
    .io_i0_ap_sra(i_alu_io_i0_ap_sra),
    .io_i0_ap_beq(i_alu_io_i0_ap_beq),
    .io_i0_ap_bne(i_alu_io_i0_ap_bne),
    .io_i0_ap_blt(i_alu_io_i0_ap_blt),
    .io_i0_ap_bge(i_alu_io_i0_ap_bge),
    .io_i0_ap_add(i_alu_io_i0_ap_add),
    .io_i0_ap_sub(i_alu_io_i0_ap_sub),
    .io_i0_ap_slt(i_alu_io_i0_ap_slt),
    .io_i0_ap_unsign(i_alu_io_i0_ap_unsign),
    .io_i0_ap_jal(i_alu_io_i0_ap_jal),
    .io_i0_ap_predict_t(i_alu_io_i0_ap_predict_t),
    .io_i0_ap_predict_nt(i_alu_io_i0_ap_predict_nt),
    .io_i0_ap_csr_write(i_alu_io_i0_ap_csr_write),
    .io_i0_ap_csr_imm(i_alu_io_i0_ap_csr_imm),
    .io_a_in(i_alu_io_a_in),
    .io_b_in(i_alu_io_b_in),
    .io_pp_in_valid(i_alu_io_pp_in_valid),
    .io_pp_in_bits_boffset(i_alu_io_pp_in_bits_boffset),
    .io_pp_in_bits_pc4(i_alu_io_pp_in_bits_pc4),
    .io_pp_in_bits_hist(i_alu_io_pp_in_bits_hist),
    .io_pp_in_bits_toffset(i_alu_io_pp_in_bits_toffset),
    .io_pp_in_bits_br_error(i_alu_io_pp_in_bits_br_error),
    .io_pp_in_bits_br_start_error(i_alu_io_pp_in_bits_br_start_error),
    .io_pp_in_bits_prett(i_alu_io_pp_in_bits_prett),
    .io_pp_in_bits_pcall(i_alu_io_pp_in_bits_pcall),
    .io_pp_in_bits_pret(i_alu_io_pp_in_bits_pret),
    .io_pp_in_bits_pja(i_alu_io_pp_in_bits_pja),
    .io_pp_in_bits_way(i_alu_io_pp_in_bits_way),
    .io_result_ff(i_alu_io_result_ff),
    .io_flush_upper_out(i_alu_io_flush_upper_out),
    .io_flush_final_out(i_alu_io_flush_final_out),
    .io_flush_path_out(i_alu_io_flush_path_out),
    .io_pred_correct_out(i_alu_io_pred_correct_out),
    .io_predict_p_out_valid(i_alu_io_predict_p_out_valid),
    .io_predict_p_out_bits_misp(i_alu_io_predict_p_out_bits_misp),
    .io_predict_p_out_bits_ataken(i_alu_io_predict_p_out_bits_ataken),
    .io_predict_p_out_bits_boffset(i_alu_io_predict_p_out_bits_boffset),
    .io_predict_p_out_bits_pc4(i_alu_io_predict_p_out_bits_pc4),
    .io_predict_p_out_bits_hist(i_alu_io_predict_p_out_bits_hist),
    .io_predict_p_out_bits_toffset(i_alu_io_predict_p_out_bits_toffset),
    .io_predict_p_out_bits_br_error(i_alu_io_predict_p_out_bits_br_error),
    .io_predict_p_out_bits_br_start_error(i_alu_io_predict_p_out_bits_br_start_error),
    .io_predict_p_out_bits_pcall(i_alu_io_predict_p_out_bits_pcall),
    .io_predict_p_out_bits_pret(i_alu_io_predict_p_out_bits_pret),
    .io_predict_p_out_bits_pja(i_alu_io_predict_p_out_bits_pja),
    .io_predict_p_out_bits_way(i_alu_io_predict_p_out_bits_way)
  );
  exu_mul_ctl i_mul ( // @[exu.scala 162:19]
    .clock(i_mul_clock),
    .reset(i_mul_reset),
    .io_scan_mode(i_mul_io_scan_mode),
    .io_mul_p_valid(i_mul_io_mul_p_valid),
    .io_mul_p_bits_rs1_sign(i_mul_io_mul_p_bits_rs1_sign),
    .io_mul_p_bits_rs2_sign(i_mul_io_mul_p_bits_rs2_sign),
    .io_mul_p_bits_low(i_mul_io_mul_p_bits_low),
    .io_rs1_in(i_mul_io_rs1_in),
    .io_rs2_in(i_mul_io_rs2_in),
    .io_result_x(i_mul_io_result_x)
  );
  exu_div_ctl i_div ( // @[exu.scala 169:19]
    .clock(i_div_clock),
    .reset(i_div_reset),
    .io_scan_mode(i_div_io_scan_mode),
    .io_dividend(i_div_io_dividend),
    .io_divisor(i_div_io_divisor),
    .io_exu_div_result(i_div_io_exu_div_result),
    .io_exu_div_wren(i_div_io_exu_div_wren),
    .io_dec_div_div_p_valid(i_div_io_dec_div_div_p_valid),
    .io_dec_div_div_p_bits_unsign(i_div_io_dec_div_div_p_bits_unsign),
    .io_dec_div_div_p_bits_rem(i_div_io_dec_div_div_p_bits_rem),
    .io_dec_div_dec_div_cancel(i_div_io_dec_div_dec_div_cancel)
  );
  assign io_dec_exu_dec_alu_exu_i0_pc_x = i_alu_io_dec_alu_exu_i0_pc_x; // @[exu.scala 145:20]
  assign io_dec_exu_decode_exu_exu_i0_result_x = mul_valid_x ? i_mul_io_result_x : i_alu_io_result_ff; // @[exu.scala 178:58]
  assign io_dec_exu_decode_exu_exu_csr_rs1_x = _T_3; // @[exu.scala 64:57]
  assign io_dec_exu_tlu_exu_exu_i0_br_hist_r = i0_pp_r_bits_hist; // @[exu.scala 205:66]
  assign io_dec_exu_tlu_exu_exu_i0_br_error_r = i0_pp_r_bits_br_error; // @[exu.scala 206:58]
  assign io_dec_exu_tlu_exu_exu_i0_br_start_error_r = i0_pp_r_bits_br_start_error; // @[exu.scala 208:52]
  assign io_dec_exu_tlu_exu_exu_i0_br_index_r = predpipe_r[12:5]; // @[exu.scala 210:58]
  assign io_dec_exu_tlu_exu_exu_i0_br_valid_r = i0_pp_r_valid; // @[exu.scala 202:52]
  assign io_dec_exu_tlu_exu_exu_i0_br_mp_r = i0_pp_r_bits_misp; // @[exu.scala 203:52]
  assign io_dec_exu_tlu_exu_exu_i0_br_middle_r = i0_pp_r_bits_pc4 ^ i0_pp_r_bits_boffset; // @[exu.scala 207:52]
  assign io_dec_exu_tlu_exu_exu_pmu_i0_br_misp = i0_pp_r_bits_misp; // @[exu.scala 182:47]
  assign io_dec_exu_tlu_exu_exu_pmu_i0_br_ataken = i0_pp_r_bits_ataken; // @[exu.scala 183:47]
  assign io_dec_exu_tlu_exu_exu_pmu_i0_pc4 = i0_pp_r_bits_pc4; // @[exu.scala 184:47]
  assign io_dec_exu_tlu_exu_exu_npc_r = _T_188[30:0]; // @[exu.scala 233:66]
  assign io_exu_bp_exu_i0_br_fghr_r = predpipe_r[20:13]; // @[exu.scala 209:58]
  assign io_exu_bp_exu_i0_br_way_r = i0_pp_r_bits_way; // @[exu.scala 204:43]
  assign io_exu_bp_exu_mp_pkt_bits_misp = i0_flush_upper_x & i0_predict_p_x_bits_misp; // @[exu.scala 219:48]
  assign io_exu_bp_exu_mp_pkt_bits_ataken = i0_flush_upper_x & i0_predict_p_x_bits_ataken; // @[exu.scala 223:48]
  assign io_exu_bp_exu_mp_pkt_bits_boffset = i0_flush_upper_x & i0_predict_p_x_bits_boffset; // @[exu.scala 224:48]
  assign io_exu_bp_exu_mp_pkt_bits_pc4 = i0_flush_upper_x & i0_predict_p_x_bits_pc4; // @[exu.scala 225:48]
  assign io_exu_bp_exu_mp_pkt_bits_hist = i0_flush_upper_x ? i0_predict_p_x_bits_hist : 2'h0; // @[exu.scala 226:66]
  assign io_exu_bp_exu_mp_pkt_bits_toffset = i0_flush_upper_x ? i0_predict_p_x_bits_toffset : 12'h0; // @[exu.scala 227:58]
  assign io_exu_bp_exu_mp_pkt_bits_pcall = i0_flush_upper_x & i0_predict_p_x_bits_pcall; // @[exu.scala 220:48]
  assign io_exu_bp_exu_mp_pkt_bits_pret = i0_flush_upper_x & i0_predict_p_x_bits_pret; // @[exu.scala 222:48]
  assign io_exu_bp_exu_mp_pkt_bits_pja = i0_flush_upper_x & i0_predict_p_x_bits_pja; // @[exu.scala 221:48]
  assign io_exu_bp_exu_mp_pkt_bits_way = i0_flush_upper_x & i0_predict_p_x_bits_way; // @[exu.scala 218:48]
  assign io_exu_bp_exu_mp_eghr = final_predpipe_mp[20:13]; // @[exu.scala 231:43]
  assign io_exu_bp_exu_mp_fghr = _T_179 ? ghr_d : ghr_x; // @[exu.scala 228:43]
  assign io_exu_bp_exu_mp_index = final_predpipe_mp[12:5]; // @[exu.scala 229:66]
  assign io_exu_bp_exu_mp_btag = final_predpipe_mp[4:0]; // @[exu.scala 230:58]
  assign io_exu_flush_final = i_alu_io_flush_final_out; // @[exu.scala 158:22]
  assign io_exu_div_result = i_div_io_exu_div_result; // @[exu.scala 176:33]
  assign io_exu_div_wren = i_div_io_exu_div_wren; // @[exu.scala 175:41]
  assign io_lsu_exu_exu_lsu_rs1_d = _T_106 | _T_105; // @[exu.scala 119:27]
  assign io_lsu_exu_exu_lsu_rs2_d = _T_117 | _T_118; // @[exu.scala 125:27]
  assign io_exu_flush_path_final = io_dec_exu_tlu_exu_dec_tlu_flush_lower_r ? io_dec_exu_tlu_exu_dec_tlu_flush_path_r : i0_flush_path_d; // @[exu.scala 232:50]
  assign rvclkhdr_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_io_en = io_dec_exu_decode_exu_dec_data_en[1]; // @[lib.scala 371:17]
  assign rvclkhdr_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_1_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_1_io_en = io_dec_exu_decode_exu_dec_data_en[1]; // @[lib.scala 371:17]
  assign rvclkhdr_1_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_2_io_clk = clock; // @[lib.scala 380:18]
  assign rvclkhdr_2_io_en = io_dec_exu_decode_exu_dec_data_en[1]; // @[lib.scala 381:17]
  assign rvclkhdr_2_io_scan_mode = io_scan_mode; // @[lib.scala 382:24]
  assign rvclkhdr_3_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_3_io_en = io_dec_exu_decode_exu_dec_data_en[1]; // @[lib.scala 371:17]
  assign rvclkhdr_3_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_4_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_4_io_en = io_dec_exu_decode_exu_dec_data_en[0]; // @[lib.scala 371:17]
  assign rvclkhdr_4_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_5_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_5_io_en = io_dec_exu_decode_exu_dec_ctl_en[1]; // @[lib.scala 371:17]
  assign rvclkhdr_5_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_6_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_6_io_en = io_dec_exu_decode_exu_dec_ctl_en[1]; // @[lib.scala 371:17]
  assign rvclkhdr_6_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_7_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_7_io_en = io_dec_exu_decode_exu_dec_ctl_en[1]; // @[lib.scala 371:17]
  assign rvclkhdr_7_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_8_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_8_io_en = io_dec_exu_decode_exu_dec_ctl_en[1]; // @[lib.scala 371:17]
  assign rvclkhdr_8_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_9_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_9_io_en = io_dec_exu_decode_exu_dec_ctl_en[1]; // @[lib.scala 371:17]
  assign rvclkhdr_9_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_10_io_clk = clock; // @[lib.scala 380:18]
  assign rvclkhdr_10_io_en = io_dec_exu_decode_exu_dec_ctl_en[0]; // @[lib.scala 381:17]
  assign rvclkhdr_10_io_scan_mode = io_scan_mode; // @[lib.scala 382:24]
  assign rvclkhdr_11_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_11_io_en = io_dec_exu_decode_exu_dec_ctl_en[0]; // @[lib.scala 371:17]
  assign rvclkhdr_11_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_12_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_12_io_en = io_dec_exu_decode_exu_dec_ctl_en[0]; // @[lib.scala 371:17]
  assign rvclkhdr_12_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_13_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_13_io_en = io_dec_exu_decode_exu_dec_data_en[0]; // @[lib.scala 371:17]
  assign rvclkhdr_13_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_14_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_14_io_en = io_dec_exu_decode_exu_dec_data_en[0]; // @[lib.scala 371:17]
  assign rvclkhdr_14_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_15_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_15_io_en = _T_41 | _T_42; // @[lib.scala 371:17]
  assign rvclkhdr_15_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_16_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_16_io_en = _T_41 | _T_42; // @[lib.scala 371:17]
  assign rvclkhdr_16_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_17_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_17_io_en = _T_41 | _T_42; // @[lib.scala 371:17]
  assign rvclkhdr_17_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign i_alu_clock = clock;
  assign i_alu_reset = reset;
  assign i_alu_io_dec_alu_dec_i0_alu_decode_d = io_dec_exu_dec_alu_dec_i0_alu_decode_d; // @[exu.scala 145:20]
  assign i_alu_io_dec_alu_dec_csr_ren_d = io_dec_exu_dec_alu_dec_csr_ren_d; // @[exu.scala 145:20]
  assign i_alu_io_dec_alu_dec_i0_br_immed_d = io_dec_exu_dec_alu_dec_i0_br_immed_d; // @[exu.scala 145:20]
  assign i_alu_io_dec_i0_pc_d = io_dec_exu_ib_exu_dec_i0_pc_d; // @[exu.scala 153:41]
  assign i_alu_io_scan_mode = io_scan_mode; // @[exu.scala 146:33]
  assign i_alu_io_flush_upper_x = i0_flush_upper_x; // @[exu.scala 149:33]
  assign i_alu_io_dec_tlu_flush_lower_r = io_dec_exu_tlu_exu_dec_tlu_flush_lower_r; // @[exu.scala 150:41]
  assign i_alu_io_enable = io_dec_exu_decode_exu_dec_ctl_en[1]; // @[exu.scala 147:41]
  assign i_alu_io_i0_ap_land = io_dec_exu_decode_exu_i0_ap_land; // @[exu.scala 154:49]
  assign i_alu_io_i0_ap_lor = io_dec_exu_decode_exu_i0_ap_lor; // @[exu.scala 154:49]
  assign i_alu_io_i0_ap_lxor = io_dec_exu_decode_exu_i0_ap_lxor; // @[exu.scala 154:49]
  assign i_alu_io_i0_ap_sll = io_dec_exu_decode_exu_i0_ap_sll; // @[exu.scala 154:49]
  assign i_alu_io_i0_ap_srl = io_dec_exu_decode_exu_i0_ap_srl; // @[exu.scala 154:49]
  assign i_alu_io_i0_ap_sra = io_dec_exu_decode_exu_i0_ap_sra; // @[exu.scala 154:49]
  assign i_alu_io_i0_ap_beq = io_dec_exu_decode_exu_i0_ap_beq; // @[exu.scala 154:49]
  assign i_alu_io_i0_ap_bne = io_dec_exu_decode_exu_i0_ap_bne; // @[exu.scala 154:49]
  assign i_alu_io_i0_ap_blt = io_dec_exu_decode_exu_i0_ap_blt; // @[exu.scala 154:49]
  assign i_alu_io_i0_ap_bge = io_dec_exu_decode_exu_i0_ap_bge; // @[exu.scala 154:49]
  assign i_alu_io_i0_ap_add = io_dec_exu_decode_exu_i0_ap_add; // @[exu.scala 154:49]
  assign i_alu_io_i0_ap_sub = io_dec_exu_decode_exu_i0_ap_sub; // @[exu.scala 154:49]
  assign i_alu_io_i0_ap_slt = io_dec_exu_decode_exu_i0_ap_slt; // @[exu.scala 154:49]
  assign i_alu_io_i0_ap_unsign = io_dec_exu_decode_exu_i0_ap_unsign; // @[exu.scala 154:49]
  assign i_alu_io_i0_ap_jal = io_dec_exu_decode_exu_i0_ap_jal; // @[exu.scala 154:49]
  assign i_alu_io_i0_ap_predict_t = io_dec_exu_decode_exu_i0_ap_predict_t; // @[exu.scala 154:49]
  assign i_alu_io_i0_ap_predict_nt = io_dec_exu_decode_exu_i0_ap_predict_nt; // @[exu.scala 154:49]
  assign i_alu_io_i0_ap_csr_write = io_dec_exu_decode_exu_i0_ap_csr_write; // @[exu.scala 154:49]
  assign i_alu_io_i0_ap_csr_imm = io_dec_exu_decode_exu_i0_ap_csr_imm; // @[exu.scala 154:49]
  assign i_alu_io_a_in = _T_80 | _T_78; // @[exu.scala 151:33]
  assign i_alu_io_b_in = i0_rs2_d; // @[exu.scala 152:33]
  assign i_alu_io_pp_in_valid = io_dec_exu_decode_exu_dec_i0_predict_p_d_valid; // @[exu.scala 148:41]
  assign i_alu_io_pp_in_bits_boffset = io_dec_exu_ib_exu_dec_i0_pc_d[0]; // @[exu.scala 148:41]
  assign i_alu_io_pp_in_bits_pc4 = io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_pc4; // @[exu.scala 148:41]
  assign i_alu_io_pp_in_bits_hist = io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_hist; // @[exu.scala 148:41]
  assign i_alu_io_pp_in_bits_toffset = io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_toffset; // @[exu.scala 148:41]
  assign i_alu_io_pp_in_bits_br_error = io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_br_error; // @[exu.scala 148:41]
  assign i_alu_io_pp_in_bits_br_start_error = io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_br_start_error; // @[exu.scala 148:41]
  assign i_alu_io_pp_in_bits_prett = io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_prett; // @[exu.scala 148:41]
  assign i_alu_io_pp_in_bits_pcall = io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_pcall; // @[exu.scala 148:41]
  assign i_alu_io_pp_in_bits_pret = io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_pret; // @[exu.scala 148:41]
  assign i_alu_io_pp_in_bits_pja = io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_pja; // @[exu.scala 148:41]
  assign i_alu_io_pp_in_bits_way = io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_way; // @[exu.scala 148:41]
  assign i_mul_clock = clock;
  assign i_mul_reset = reset;
  assign i_mul_io_scan_mode = io_scan_mode; // @[exu.scala 163:33]
  assign i_mul_io_mul_p_valid = io_dec_exu_decode_exu_mul_p_valid; // @[exu.scala 164:41]
  assign i_mul_io_mul_p_bits_rs1_sign = io_dec_exu_decode_exu_mul_p_bits_rs1_sign; // @[exu.scala 164:41]
  assign i_mul_io_mul_p_bits_rs2_sign = io_dec_exu_decode_exu_mul_p_bits_rs2_sign; // @[exu.scala 164:41]
  assign i_mul_io_mul_p_bits_low = io_dec_exu_decode_exu_mul_p_bits_low; // @[exu.scala 164:41]
  assign i_mul_io_rs1_in = _T_125 | _T_75; // @[exu.scala 165:41]
  assign i_mul_io_rs2_in = _T_91 | _T_90; // @[exu.scala 166:41]
  assign i_div_clock = clock;
  assign i_div_reset = reset;
  assign i_div_io_scan_mode = io_scan_mode; // @[exu.scala 171:33]
  assign i_div_io_dividend = _T_125 | _T_75; // @[exu.scala 173:33]
  assign i_div_io_divisor = _T_91 | _T_90; // @[exu.scala 174:33]
  assign i_div_io_dec_div_div_p_valid = io_dec_exu_dec_div_div_p_valid; // @[exu.scala 170:20]
  assign i_div_io_dec_div_div_p_bits_unsign = io_dec_exu_dec_div_div_p_bits_unsign; // @[exu.scala 170:20]
  assign i_div_io_dec_div_div_p_bits_rem = io_dec_exu_dec_div_div_p_bits_rem; // @[exu.scala 170:20]
  assign i_div_io_dec_div_dec_div_cancel = io_dec_exu_dec_div_dec_div_cancel; // @[exu.scala 170:20]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  i0_flush_path_x = _RAND_0[30:0];
  _RAND_1 = {1{`RANDOM}};
  _T_3 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  i0_predict_p_x_valid = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  i0_predict_p_x_bits_misp = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  i0_predict_p_x_bits_ataken = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  i0_predict_p_x_bits_boffset = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  i0_predict_p_x_bits_pc4 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  i0_predict_p_x_bits_hist = _RAND_7[1:0];
  _RAND_8 = {1{`RANDOM}};
  i0_predict_p_x_bits_toffset = _RAND_8[11:0];
  _RAND_9 = {1{`RANDOM}};
  i0_predict_p_x_bits_br_error = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  i0_predict_p_x_bits_br_start_error = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  i0_predict_p_x_bits_pcall = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  i0_predict_p_x_bits_pret = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  i0_predict_p_x_bits_pja = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  i0_predict_p_x_bits_way = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  predpipe_x = _RAND_15[20:0];
  _RAND_16 = {1{`RANDOM}};
  predpipe_r = _RAND_16[20:0];
  _RAND_17 = {1{`RANDOM}};
  ghr_x = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  i0_pred_correct_upper_x = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  i0_flush_upper_x = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  i0_taken_x = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  i0_valid_x = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  i0_pp_r_valid = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  i0_pp_r_bits_misp = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  i0_pp_r_bits_ataken = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  i0_pp_r_bits_boffset = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  i0_pp_r_bits_pc4 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  i0_pp_r_bits_hist = _RAND_27[1:0];
  _RAND_28 = {1{`RANDOM}};
  i0_pp_r_bits_br_error = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  i0_pp_r_bits_br_start_error = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  i0_pp_r_bits_way = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  pred_temp1 = _RAND_31[5:0];
  _RAND_32 = {1{`RANDOM}};
  i0_pred_correct_upper_r = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  i0_flush_path_upper_r = _RAND_33[30:0];
  _RAND_34 = {1{`RANDOM}};
  pred_temp2 = _RAND_34[24:0];
  _RAND_35 = {1{`RANDOM}};
  ghr_d = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  mul_valid_x = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  flush_lower_ff = _RAND_37[0:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    i0_flush_path_x = 31'h0;
  end
  if (reset) begin
    _T_3 = 32'h0;
  end
  if (reset) begin
    i0_predict_p_x_valid = 1'h0;
  end
  if (reset) begin
    i0_predict_p_x_bits_misp = 1'h0;
  end
  if (reset) begin
    i0_predict_p_x_bits_ataken = 1'h0;
  end
  if (reset) begin
    i0_predict_p_x_bits_boffset = 1'h0;
  end
  if (reset) begin
    i0_predict_p_x_bits_pc4 = 1'h0;
  end
  if (reset) begin
    i0_predict_p_x_bits_hist = 2'h0;
  end
  if (reset) begin
    i0_predict_p_x_bits_toffset = 12'h0;
  end
  if (reset) begin
    i0_predict_p_x_bits_br_error = 1'h0;
  end
  if (reset) begin
    i0_predict_p_x_bits_br_start_error = 1'h0;
  end
  if (reset) begin
    i0_predict_p_x_bits_pcall = 1'h0;
  end
  if (reset) begin
    i0_predict_p_x_bits_pret = 1'h0;
  end
  if (reset) begin
    i0_predict_p_x_bits_pja = 1'h0;
  end
  if (reset) begin
    i0_predict_p_x_bits_way = 1'h0;
  end
  if (reset) begin
    predpipe_x = 21'h0;
  end
  if (reset) begin
    predpipe_r = 21'h0;
  end
  if (reset) begin
    ghr_x = 8'h0;
  end
  if (reset) begin
    i0_pred_correct_upper_x = 1'h0;
  end
  if (reset) begin
    i0_flush_upper_x = 1'h0;
  end
  if (reset) begin
    i0_taken_x = 1'h0;
  end
  if (reset) begin
    i0_valid_x = 1'h0;
  end
  if (reset) begin
    i0_pp_r_valid = 1'h0;
  end
  if (reset) begin
    i0_pp_r_bits_misp = 1'h0;
  end
  if (reset) begin
    i0_pp_r_bits_ataken = 1'h0;
  end
  if (reset) begin
    i0_pp_r_bits_boffset = 1'h0;
  end
  if (reset) begin
    i0_pp_r_bits_pc4 = 1'h0;
  end
  if (reset) begin
    i0_pp_r_bits_hist = 2'h0;
  end
  if (reset) begin
    i0_pp_r_bits_br_error = 1'h0;
  end
  if (reset) begin
    i0_pp_r_bits_br_start_error = 1'h0;
  end
  if (reset) begin
    i0_pp_r_bits_way = 1'h0;
  end
  if (reset) begin
    pred_temp1 = 6'h0;
  end
  if (reset) begin
    i0_pred_correct_upper_r = 1'h0;
  end
  if (reset) begin
    i0_flush_path_upper_r = 31'h0;
  end
  if (reset) begin
    pred_temp2 = 25'h0;
  end
  if (reset) begin
    ghr_d = 8'h0;
  end
  if (reset) begin
    mul_valid_x = 1'h0;
  end
  if (reset) begin
    flush_lower_ff = 1'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge rvclkhdr_io_l1clk or posedge reset) begin
    if (reset) begin
      i0_flush_path_x <= 31'h0;
    end else begin
      i0_flush_path_x <= i_alu_io_flush_path_out;
    end
  end
  always @(posedge rvclkhdr_1_io_l1clk or posedge reset) begin
    if (reset) begin
      _T_3 <= 32'h0;
    end else if (io_dec_exu_dec_alu_dec_csr_ren_d) begin
      _T_3 <= i0_rs1_d;
    end else begin
      _T_3 <= io_dec_exu_decode_exu_exu_csr_rs1_x;
    end
  end
  always @(posedge rvclkhdr_2_io_l1clk or posedge reset) begin
    if (reset) begin
      i0_predict_p_x_valid <= 1'h0;
    end else begin
      i0_predict_p_x_valid <= i_alu_io_predict_p_out_valid;
    end
  end
  always @(posedge rvclkhdr_2_io_l1clk or posedge reset) begin
    if (reset) begin
      i0_predict_p_x_bits_misp <= 1'h0;
    end else begin
      i0_predict_p_x_bits_misp <= i_alu_io_predict_p_out_bits_misp;
    end
  end
  always @(posedge rvclkhdr_2_io_l1clk or posedge reset) begin
    if (reset) begin
      i0_predict_p_x_bits_ataken <= 1'h0;
    end else begin
      i0_predict_p_x_bits_ataken <= i_alu_io_predict_p_out_bits_ataken;
    end
  end
  always @(posedge rvclkhdr_2_io_l1clk or posedge reset) begin
    if (reset) begin
      i0_predict_p_x_bits_boffset <= 1'h0;
    end else begin
      i0_predict_p_x_bits_boffset <= i_alu_io_predict_p_out_bits_boffset;
    end
  end
  always @(posedge rvclkhdr_2_io_l1clk or posedge reset) begin
    if (reset) begin
      i0_predict_p_x_bits_pc4 <= 1'h0;
    end else begin
      i0_predict_p_x_bits_pc4 <= i_alu_io_predict_p_out_bits_pc4;
    end
  end
  always @(posedge rvclkhdr_2_io_l1clk or posedge reset) begin
    if (reset) begin
      i0_predict_p_x_bits_hist <= 2'h0;
    end else begin
      i0_predict_p_x_bits_hist <= i_alu_io_predict_p_out_bits_hist;
    end
  end
  always @(posedge rvclkhdr_2_io_l1clk or posedge reset) begin
    if (reset) begin
      i0_predict_p_x_bits_toffset <= 12'h0;
    end else begin
      i0_predict_p_x_bits_toffset <= i_alu_io_predict_p_out_bits_toffset;
    end
  end
  always @(posedge rvclkhdr_2_io_l1clk or posedge reset) begin
    if (reset) begin
      i0_predict_p_x_bits_br_error <= 1'h0;
    end else begin
      i0_predict_p_x_bits_br_error <= i_alu_io_predict_p_out_bits_br_error;
    end
  end
  always @(posedge rvclkhdr_2_io_l1clk or posedge reset) begin
    if (reset) begin
      i0_predict_p_x_bits_br_start_error <= 1'h0;
    end else begin
      i0_predict_p_x_bits_br_start_error <= i_alu_io_predict_p_out_bits_br_start_error;
    end
  end
  always @(posedge rvclkhdr_2_io_l1clk or posedge reset) begin
    if (reset) begin
      i0_predict_p_x_bits_pcall <= 1'h0;
    end else begin
      i0_predict_p_x_bits_pcall <= i_alu_io_predict_p_out_bits_pcall;
    end
  end
  always @(posedge rvclkhdr_2_io_l1clk or posedge reset) begin
    if (reset) begin
      i0_predict_p_x_bits_pret <= 1'h0;
    end else begin
      i0_predict_p_x_bits_pret <= i_alu_io_predict_p_out_bits_pret;
    end
  end
  always @(posedge rvclkhdr_2_io_l1clk or posedge reset) begin
    if (reset) begin
      i0_predict_p_x_bits_pja <= 1'h0;
    end else begin
      i0_predict_p_x_bits_pja <= i_alu_io_predict_p_out_bits_pja;
    end
  end
  always @(posedge rvclkhdr_2_io_l1clk or posedge reset) begin
    if (reset) begin
      i0_predict_p_x_bits_way <= 1'h0;
    end else begin
      i0_predict_p_x_bits_way <= i_alu_io_predict_p_out_bits_way;
    end
  end
  always @(posedge rvclkhdr_3_io_l1clk or posedge reset) begin
    if (reset) begin
      predpipe_x <= 21'h0;
    end else begin
      predpipe_x <= {_T,io_dec_exu_decode_exu_i0_predict_btag_d};
    end
  end
  always @(posedge rvclkhdr_4_io_l1clk or posedge reset) begin
    if (reset) begin
      predpipe_r <= 21'h0;
    end else begin
      predpipe_r <= predpipe_x;
    end
  end
  always @(posedge rvclkhdr_5_io_l1clk or posedge reset) begin
    if (reset) begin
      ghr_x <= 8'h0;
    end else if (i0_valid_x) begin
      ghr_x <= _T_167;
    end
  end
  always @(posedge rvclkhdr_6_io_l1clk or posedge reset) begin
    if (reset) begin
      i0_pred_correct_upper_x <= 1'h0;
    end else begin
      i0_pred_correct_upper_x <= i_alu_io_pred_correct_out;
    end
  end
  always @(posedge rvclkhdr_7_io_l1clk or posedge reset) begin
    if (reset) begin
      i0_flush_upper_x <= 1'h0;
    end else begin
      i0_flush_upper_x <= i_alu_io_flush_upper_out;
    end
  end
  always @(posedge rvclkhdr_8_io_l1clk or posedge reset) begin
    if (reset) begin
      i0_taken_x <= 1'h0;
    end else begin
      i0_taken_x <= i0_predict_p_d_bits_ataken & io_dec_exu_dec_alu_dec_i0_alu_decode_d;
    end
  end
  always @(posedge rvclkhdr_9_io_l1clk or posedge reset) begin
    if (reset) begin
      i0_valid_x <= 1'h0;
    end else begin
      i0_valid_x <= _T_145 & _T_149;
    end
  end
  always @(posedge rvclkhdr_10_io_l1clk or posedge reset) begin
    if (reset) begin
      i0_pp_r_valid <= 1'h0;
    end else begin
      i0_pp_r_valid <= i0_predict_p_x_valid;
    end
  end
  always @(posedge rvclkhdr_10_io_l1clk or posedge reset) begin
    if (reset) begin
      i0_pp_r_bits_misp <= 1'h0;
    end else begin
      i0_pp_r_bits_misp <= i0_predict_p_x_bits_misp;
    end
  end
  always @(posedge rvclkhdr_10_io_l1clk or posedge reset) begin
    if (reset) begin
      i0_pp_r_bits_ataken <= 1'h0;
    end else begin
      i0_pp_r_bits_ataken <= i0_predict_p_x_bits_ataken;
    end
  end
  always @(posedge rvclkhdr_10_io_l1clk or posedge reset) begin
    if (reset) begin
      i0_pp_r_bits_boffset <= 1'h0;
    end else begin
      i0_pp_r_bits_boffset <= i0_predict_p_x_bits_boffset;
    end
  end
  always @(posedge rvclkhdr_10_io_l1clk or posedge reset) begin
    if (reset) begin
      i0_pp_r_bits_pc4 <= 1'h0;
    end else begin
      i0_pp_r_bits_pc4 <= i0_predict_p_x_bits_pc4;
    end
  end
  always @(posedge rvclkhdr_10_io_l1clk or posedge reset) begin
    if (reset) begin
      i0_pp_r_bits_hist <= 2'h0;
    end else begin
      i0_pp_r_bits_hist <= i0_predict_p_x_bits_hist;
    end
  end
  always @(posedge rvclkhdr_10_io_l1clk or posedge reset) begin
    if (reset) begin
      i0_pp_r_bits_br_error <= 1'h0;
    end else begin
      i0_pp_r_bits_br_error <= i0_predict_p_x_bits_br_error;
    end
  end
  always @(posedge rvclkhdr_10_io_l1clk or posedge reset) begin
    if (reset) begin
      i0_pp_r_bits_br_start_error <= 1'h0;
    end else begin
      i0_pp_r_bits_br_start_error <= i0_predict_p_x_bits_br_start_error;
    end
  end
  always @(posedge rvclkhdr_10_io_l1clk or posedge reset) begin
    if (reset) begin
      i0_pp_r_bits_way <= 1'h0;
    end else begin
      i0_pp_r_bits_way <= i0_predict_p_x_bits_way;
    end
  end
  always @(posedge rvclkhdr_11_io_l1clk or posedge reset) begin
    if (reset) begin
      pred_temp1 <= 6'h0;
    end else begin
      pred_temp1 <= io_dec_exu_decode_exu_pred_correct_npc_x[5:0];
    end
  end
  always @(posedge rvclkhdr_12_io_l1clk or posedge reset) begin
    if (reset) begin
      i0_pred_correct_upper_r <= 1'h0;
    end else begin
      i0_pred_correct_upper_r <= i0_pred_correct_upper_x;
    end
  end
  always @(posedge rvclkhdr_13_io_l1clk or posedge reset) begin
    if (reset) begin
      i0_flush_path_upper_r <= 31'h0;
    end else begin
      i0_flush_path_upper_r <= i0_flush_path_x;
    end
  end
  always @(posedge rvclkhdr_14_io_l1clk or posedge reset) begin
    if (reset) begin
      pred_temp2 <= 25'h0;
    end else begin
      pred_temp2 <= io_dec_exu_decode_exu_pred_correct_npc_x[30:6];
    end
  end
  always @(posedge rvclkhdr_15_io_l1clk or posedge reset) begin
    if (reset) begin
      ghr_d <= 8'h0;
    end else begin
      ghr_d <= _T_162 | _T_161;
    end
  end
  always @(posedge rvclkhdr_16_io_l1clk or posedge reset) begin
    if (reset) begin
      mul_valid_x <= 1'h0;
    end else begin
      mul_valid_x <= io_dec_exu_decode_exu_mul_p_valid;
    end
  end
  always @(posedge rvclkhdr_17_io_l1clk or posedge reset) begin
    if (reset) begin
      flush_lower_ff <= 1'h0;
    end else begin
      flush_lower_ff <= io_dec_exu_tlu_exu_dec_tlu_flush_lower_r;
    end
  end
endmodule
module lsu_addrcheck(
  input         reset,
  input         io_lsu_c2_m_clk,
  input  [31:0] io_start_addr_d,
  input  [31:0] io_end_addr_d,
  input         io_lsu_pkt_d_valid,
  input         io_lsu_pkt_d_bits_fast_int,
  input         io_lsu_pkt_d_bits_by,
  input         io_lsu_pkt_d_bits_half,
  input         io_lsu_pkt_d_bits_word,
  input         io_lsu_pkt_d_bits_load,
  input         io_lsu_pkt_d_bits_store,
  input         io_lsu_pkt_d_bits_dma,
  input  [31:0] io_dec_tlu_mrac_ff,
  input  [3:0]  io_rs1_region_d,
  output        io_is_sideeffects_m,
  output        io_addr_in_dccm_d,
  output        io_addr_in_pic_d,
  output        io_addr_external_d,
  output        io_access_fault_d,
  output        io_misaligned_fault_d,
  output [3:0]  io_exc_mscause_d,
  output        io_fir_dccm_access_error_d,
  output        io_fir_nondccm_access_error_d
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  start_addr_in_dccm_region_d = io_start_addr_d[31:28] == 4'hf; // @[lib.scala 356:49]
  wire  start_addr_in_dccm_d = io_start_addr_d[31:16] == 16'hf004; // @[lib.scala 361:39]
  wire  end_addr_in_dccm_region_d = io_end_addr_d[31:28] == 4'hf; // @[lib.scala 356:49]
  wire  end_addr_in_dccm_d = io_end_addr_d[31:16] == 16'hf004; // @[lib.scala 361:39]
  wire  addr_in_iccm = io_start_addr_d[31:28] == 4'he; // @[lsu_addrcheck.scala 42:45]
  wire  start_addr_in_pic_d = io_start_addr_d[31:15] == 17'h1e018; // @[lib.scala 361:39]
  wire  end_addr_in_pic_d = io_end_addr_d[31:15] == 17'h1e018; // @[lib.scala 361:39]
  wire  start_addr_dccm_or_pic = start_addr_in_dccm_region_d | start_addr_in_dccm_region_d; // @[lsu_addrcheck.scala 54:60]
  wire  _T_17 = io_rs1_region_d == 4'hf; // @[lsu_addrcheck.scala 55:54]
  wire  base_reg_dccm_or_pic = _T_17 | _T_17; // @[lsu_addrcheck.scala 55:73]
  wire [4:0] csr_idx = {io_start_addr_d[31:28],1'h1}; // @[Cat.scala 29:58]
  wire [31:0] _T_25 = io_dec_tlu_mrac_ff >> csr_idx; // @[lsu_addrcheck.scala 61:50]
  wire  _T_28 = start_addr_dccm_or_pic | addr_in_iccm; // @[lsu_addrcheck.scala 61:121]
  wire  _T_29 = ~_T_28; // @[lsu_addrcheck.scala 61:62]
  wire  _T_30 = _T_25[0] & _T_29; // @[lsu_addrcheck.scala 61:60]
  wire  _T_31 = _T_30 & io_lsu_pkt_d_valid; // @[lsu_addrcheck.scala 61:137]
  wire  _T_32 = io_lsu_pkt_d_bits_store | io_lsu_pkt_d_bits_load; // @[lsu_addrcheck.scala 61:185]
  wire  is_sideeffects_d = _T_31 & _T_32; // @[lsu_addrcheck.scala 61:158]
  wire  _T_34 = io_start_addr_d[1:0] == 2'h0; // @[lsu_addrcheck.scala 62:80]
  wire  _T_35 = io_lsu_pkt_d_bits_word & _T_34; // @[lsu_addrcheck.scala 62:56]
  wire  _T_37 = ~io_start_addr_d[0]; // @[lsu_addrcheck.scala 62:138]
  wire  _T_38 = io_lsu_pkt_d_bits_half & _T_37; // @[lsu_addrcheck.scala 62:116]
  wire  _T_39 = _T_35 | _T_38; // @[lsu_addrcheck.scala 62:90]
  wire  is_aligned_d = _T_39 | io_lsu_pkt_d_bits_by; // @[lsu_addrcheck.scala 62:148]
  wire [31:0] _T_50 = io_start_addr_d | 32'h7fffffff; // @[lsu_addrcheck.scala 67:56]
  wire  _T_52 = _T_50 == 32'h7fffffff; // @[lsu_addrcheck.scala 67:88]
  wire [31:0] _T_55 = io_start_addr_d | 32'h3fffffff; // @[lsu_addrcheck.scala 68:56]
  wire  _T_57 = _T_55 == 32'hffffffff; // @[lsu_addrcheck.scala 68:88]
  wire  _T_59 = _T_52 | _T_57; // @[lsu_addrcheck.scala 67:153]
  wire [31:0] _T_61 = io_start_addr_d | 32'h1fffffff; // @[lsu_addrcheck.scala 69:56]
  wire  _T_63 = _T_61 == 32'hbfffffff; // @[lsu_addrcheck.scala 69:88]
  wire  _T_65 = _T_59 | _T_63; // @[lsu_addrcheck.scala 68:153]
  wire [31:0] _T_67 = io_start_addr_d | 32'hfffffff; // @[lsu_addrcheck.scala 70:56]
  wire  _T_69 = _T_67 == 32'h8fffffff; // @[lsu_addrcheck.scala 70:88]
  wire  _T_71 = _T_65 | _T_69; // @[lsu_addrcheck.scala 69:153]
  wire [31:0] _T_97 = io_end_addr_d | 32'h7fffffff; // @[lsu_addrcheck.scala 76:57]
  wire  _T_99 = _T_97 == 32'h7fffffff; // @[lsu_addrcheck.scala 76:89]
  wire [31:0] _T_102 = io_end_addr_d | 32'h3fffffff; // @[lsu_addrcheck.scala 77:58]
  wire  _T_104 = _T_102 == 32'hffffffff; // @[lsu_addrcheck.scala 77:90]
  wire  _T_106 = _T_99 | _T_104; // @[lsu_addrcheck.scala 76:154]
  wire [31:0] _T_108 = io_end_addr_d | 32'h1fffffff; // @[lsu_addrcheck.scala 78:58]
  wire  _T_110 = _T_108 == 32'hbfffffff; // @[lsu_addrcheck.scala 78:90]
  wire  _T_112 = _T_106 | _T_110; // @[lsu_addrcheck.scala 77:155]
  wire [31:0] _T_114 = io_end_addr_d | 32'hfffffff; // @[lsu_addrcheck.scala 79:58]
  wire  _T_116 = _T_114 == 32'h8fffffff; // @[lsu_addrcheck.scala 79:90]
  wire  _T_118 = _T_112 | _T_116; // @[lsu_addrcheck.scala 78:155]
  wire  non_dccm_access_ok = _T_71 & _T_118; // @[lsu_addrcheck.scala 75:7]
  wire  regpred_access_fault_d = start_addr_dccm_or_pic ^ base_reg_dccm_or_pic; // @[lsu_addrcheck.scala 85:57]
  wire  _T_145 = io_start_addr_d[1:0] != 2'h0; // @[lsu_addrcheck.scala 86:76]
  wire  _T_146 = ~io_lsu_pkt_d_bits_word; // @[lsu_addrcheck.scala 86:92]
  wire  _T_147 = _T_145 | _T_146; // @[lsu_addrcheck.scala 86:90]
  wire  picm_access_fault_d = io_addr_in_pic_d & _T_147; // @[lsu_addrcheck.scala 86:51]
  wire  _T_148 = start_addr_in_dccm_d | start_addr_in_pic_d; // @[lsu_addrcheck.scala 91:87]
  wire  _T_149 = ~_T_148; // @[lsu_addrcheck.scala 91:64]
  wire  _T_150 = start_addr_in_dccm_region_d & _T_149; // @[lsu_addrcheck.scala 91:62]
  wire  _T_151 = end_addr_in_dccm_d | end_addr_in_pic_d; // @[lsu_addrcheck.scala 93:57]
  wire  _T_152 = ~_T_151; // @[lsu_addrcheck.scala 93:36]
  wire  _T_153 = end_addr_in_dccm_region_d & _T_152; // @[lsu_addrcheck.scala 93:34]
  wire  _T_154 = _T_150 | _T_153; // @[lsu_addrcheck.scala 91:112]
  wire  _T_155 = start_addr_in_dccm_d & end_addr_in_pic_d; // @[lsu_addrcheck.scala 95:29]
  wire  _T_156 = _T_154 | _T_155; // @[lsu_addrcheck.scala 93:85]
  wire  _T_157 = start_addr_in_pic_d & end_addr_in_dccm_d; // @[lsu_addrcheck.scala 97:29]
  wire  unmapped_access_fault_d = _T_156 | _T_157; // @[lsu_addrcheck.scala 95:85]
  wire  _T_159 = ~start_addr_in_dccm_region_d; // @[lsu_addrcheck.scala 99:33]
  wire  _T_160 = ~non_dccm_access_ok; // @[lsu_addrcheck.scala 99:64]
  wire  mpu_access_fault_d = _T_159 & _T_160; // @[lsu_addrcheck.scala 99:62]
  wire  _T_162 = unmapped_access_fault_d | mpu_access_fault_d; // @[lsu_addrcheck.scala 111:49]
  wire  _T_163 = _T_162 | picm_access_fault_d; // @[lsu_addrcheck.scala 111:70]
  wire  _T_164 = _T_163 | regpred_access_fault_d; // @[lsu_addrcheck.scala 111:92]
  wire  _T_165 = _T_164 & io_lsu_pkt_d_valid; // @[lsu_addrcheck.scala 111:118]
  wire  _T_166 = ~io_lsu_pkt_d_bits_dma; // @[lsu_addrcheck.scala 111:141]
  wire [3:0] _T_172 = picm_access_fault_d ? 4'h6 : 4'h0; // @[lsu_addrcheck.scala 112:164]
  wire [3:0] _T_173 = regpred_access_fault_d ? 4'h5 : _T_172; // @[lsu_addrcheck.scala 112:120]
  wire [3:0] _T_174 = mpu_access_fault_d ? 4'h3 : _T_173; // @[lsu_addrcheck.scala 112:80]
  wire [3:0] access_fault_mscause_d = unmapped_access_fault_d ? 4'h2 : _T_174; // @[lsu_addrcheck.scala 112:35]
  wire  regcross_misaligned_fault_d = io_start_addr_d[31:28] != io_end_addr_d[31:28]; // @[lsu_addrcheck.scala 113:61]
  wire  _T_177 = ~is_aligned_d; // @[lsu_addrcheck.scala 114:59]
  wire  sideeffect_misaligned_fault_d = is_sideeffects_d & _T_177; // @[lsu_addrcheck.scala 114:57]
  wire  _T_178 = sideeffect_misaligned_fault_d & io_addr_external_d; // @[lsu_addrcheck.scala 115:90]
  wire  _T_179 = regcross_misaligned_fault_d | _T_178; // @[lsu_addrcheck.scala 115:57]
  wire  _T_180 = _T_179 & io_lsu_pkt_d_valid; // @[lsu_addrcheck.scala 115:113]
  wire [3:0] _T_184 = sideeffect_misaligned_fault_d ? 4'h1 : 4'h0; // @[lsu_addrcheck.scala 116:80]
  wire [3:0] misaligned_fault_mscause_d = regcross_misaligned_fault_d ? 4'h2 : _T_184; // @[lsu_addrcheck.scala 116:39]
  wire  _T_189 = ~start_addr_in_dccm_d; // @[lsu_addrcheck.scala 118:66]
  wire  _T_190 = start_addr_in_dccm_region_d & _T_189; // @[lsu_addrcheck.scala 118:64]
  wire  _T_191 = ~end_addr_in_dccm_d; // @[lsu_addrcheck.scala 118:120]
  wire  _T_192 = end_addr_in_dccm_region_d & _T_191; // @[lsu_addrcheck.scala 118:118]
  wire  _T_193 = _T_190 | _T_192; // @[lsu_addrcheck.scala 118:88]
  wire  _T_194 = _T_193 & io_lsu_pkt_d_valid; // @[lsu_addrcheck.scala 118:142]
  wire  _T_196 = start_addr_in_dccm_region_d & end_addr_in_dccm_region_d; // @[lsu_addrcheck.scala 119:66]
  wire  _T_197 = ~_T_196; // @[lsu_addrcheck.scala 119:36]
  wire  _T_198 = _T_197 & io_lsu_pkt_d_valid; // @[lsu_addrcheck.scala 119:95]
  reg  _T_200; // @[lsu_addrcheck.scala 121:60]
  assign io_is_sideeffects_m = _T_200; // @[lsu_addrcheck.scala 121:50]
  assign io_addr_in_dccm_d = start_addr_in_dccm_d & end_addr_in_dccm_d; // @[lsu_addrcheck.scala 56:32]
  assign io_addr_in_pic_d = start_addr_in_pic_d & end_addr_in_pic_d; // @[lsu_addrcheck.scala 57:32]
  assign io_addr_external_d = ~start_addr_dccm_or_pic; // @[lsu_addrcheck.scala 59:30]
  assign io_access_fault_d = _T_165 & _T_166; // @[lsu_addrcheck.scala 111:21]
  assign io_misaligned_fault_d = _T_180 & _T_166; // @[lsu_addrcheck.scala 115:25]
  assign io_exc_mscause_d = io_misaligned_fault_d ? misaligned_fault_mscause_d : access_fault_mscause_d; // @[lsu_addrcheck.scala 117:21]
  assign io_fir_dccm_access_error_d = _T_194 & io_lsu_pkt_d_bits_fast_int; // @[lsu_addrcheck.scala 118:31]
  assign io_fir_nondccm_access_error_d = _T_198 & io_lsu_pkt_d_bits_fast_int; // @[lsu_addrcheck.scala 119:33]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_200 = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    _T_200 = 1'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge io_lsu_c2_m_clk or posedge reset) begin
    if (reset) begin
      _T_200 <= 1'h0;
    end else begin
      _T_200 <= _T_31 & _T_32;
    end
  end
endmodule
module lsu_lsc_ctl(
  input         reset,
  input         io_lsu_c1_m_clk,
  input         io_lsu_c1_r_clk,
  input         io_lsu_c2_m_clk,
  input         io_lsu_c2_r_clk,
  input         io_lsu_store_c1_m_clk,
  input  [31:0] io_lsu_ld_data_corr_r,
  input         io_lsu_single_ecc_error_r,
  input         io_lsu_double_ecc_error_r,
  input  [31:0] io_lsu_ld_data_m,
  input         io_lsu_single_ecc_error_m,
  input         io_lsu_double_ecc_error_m,
  input         io_flush_m_up,
  input         io_flush_r,
  input  [31:0] io_lsu_exu_exu_lsu_rs1_d,
  input  [31:0] io_lsu_exu_exu_lsu_rs2_d,
  input         io_lsu_p_valid,
  input         io_lsu_p_bits_fast_int,
  input         io_lsu_p_bits_by,
  input         io_lsu_p_bits_half,
  input         io_lsu_p_bits_word,
  input         io_lsu_p_bits_load,
  input         io_lsu_p_bits_store,
  input         io_lsu_p_bits_unsign,
  input         io_lsu_p_bits_store_data_bypass_d,
  input         io_lsu_p_bits_load_ldst_bypass_d,
  input         io_dec_lsu_valid_raw_d,
  input  [11:0] io_dec_lsu_offset_d,
  input  [31:0] io_picm_mask_data_m,
  input  [31:0] io_bus_read_data_m,
  output [31:0] io_lsu_result_m,
  output [31:0] io_lsu_result_corr_r,
  output [31:0] io_lsu_addr_d,
  output [31:0] io_lsu_addr_m,
  output [31:0] io_lsu_addr_r,
  output [31:0] io_end_addr_d,
  output [31:0] io_end_addr_m,
  output [31:0] io_end_addr_r,
  output [31:0] io_store_data_m,
  input  [31:0] io_dec_tlu_mrac_ff,
  output        io_lsu_exc_m,
  output        io_is_sideeffects_m,
  output        io_lsu_commit_r,
  output        io_lsu_single_ecc_error_incr,
  output        io_lsu_error_pkt_r_valid,
  output        io_lsu_error_pkt_r_bits_single_ecc_error,
  output        io_lsu_error_pkt_r_bits_inst_type,
  output        io_lsu_error_pkt_r_bits_exc_type,
  output [3:0]  io_lsu_error_pkt_r_bits_mscause,
  output [31:0] io_lsu_error_pkt_r_bits_addr,
  output [30:0] io_lsu_fir_addr,
  output [1:0]  io_lsu_fir_error,
  output        io_addr_in_dccm_d,
  output        io_addr_in_dccm_m,
  output        io_addr_in_dccm_r,
  output        io_addr_in_pic_d,
  output        io_addr_in_pic_m,
  output        io_addr_in_pic_r,
  output        io_addr_external_m,
  input         io_dma_lsc_ctl_dma_dccm_req,
  input  [31:0] io_dma_lsc_ctl_dma_mem_addr,
  input  [2:0]  io_dma_lsc_ctl_dma_mem_sz,
  input         io_dma_lsc_ctl_dma_mem_write,
  input  [63:0] io_dma_lsc_ctl_dma_mem_wdata,
  output        io_lsu_pkt_d_valid,
  output        io_lsu_pkt_d_bits_fast_int,
  output        io_lsu_pkt_d_bits_by,
  output        io_lsu_pkt_d_bits_half,
  output        io_lsu_pkt_d_bits_word,
  output        io_lsu_pkt_d_bits_dword,
  output        io_lsu_pkt_d_bits_load,
  output        io_lsu_pkt_d_bits_store,
  output        io_lsu_pkt_d_bits_unsign,
  output        io_lsu_pkt_d_bits_dma,
  output        io_lsu_pkt_d_bits_store_data_bypass_d,
  output        io_lsu_pkt_d_bits_load_ldst_bypass_d,
  output        io_lsu_pkt_d_bits_store_data_bypass_m,
  output        io_lsu_pkt_m_valid,
  output        io_lsu_pkt_m_bits_fast_int,
  output        io_lsu_pkt_m_bits_by,
  output        io_lsu_pkt_m_bits_half,
  output        io_lsu_pkt_m_bits_word,
  output        io_lsu_pkt_m_bits_dword,
  output        io_lsu_pkt_m_bits_load,
  output        io_lsu_pkt_m_bits_store,
  output        io_lsu_pkt_m_bits_unsign,
  output        io_lsu_pkt_m_bits_dma,
  output        io_lsu_pkt_m_bits_store_data_bypass_m,
  output        io_lsu_pkt_r_valid,
  output        io_lsu_pkt_r_bits_by,
  output        io_lsu_pkt_r_bits_half,
  output        io_lsu_pkt_r_bits_word,
  output        io_lsu_pkt_r_bits_dword,
  output        io_lsu_pkt_r_bits_load,
  output        io_lsu_pkt_r_bits_store,
  output        io_lsu_pkt_r_bits_unsign,
  output        io_lsu_pkt_r_bits_dma
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
`endif // RANDOMIZE_REG_INIT
  wire  addrcheck_reset; // @[lsu_lsc_ctl.scala 113:25]
  wire  addrcheck_io_lsu_c2_m_clk; // @[lsu_lsc_ctl.scala 113:25]
  wire [31:0] addrcheck_io_start_addr_d; // @[lsu_lsc_ctl.scala 113:25]
  wire [31:0] addrcheck_io_end_addr_d; // @[lsu_lsc_ctl.scala 113:25]
  wire  addrcheck_io_lsu_pkt_d_valid; // @[lsu_lsc_ctl.scala 113:25]
  wire  addrcheck_io_lsu_pkt_d_bits_fast_int; // @[lsu_lsc_ctl.scala 113:25]
  wire  addrcheck_io_lsu_pkt_d_bits_by; // @[lsu_lsc_ctl.scala 113:25]
  wire  addrcheck_io_lsu_pkt_d_bits_half; // @[lsu_lsc_ctl.scala 113:25]
  wire  addrcheck_io_lsu_pkt_d_bits_word; // @[lsu_lsc_ctl.scala 113:25]
  wire  addrcheck_io_lsu_pkt_d_bits_load; // @[lsu_lsc_ctl.scala 113:25]
  wire  addrcheck_io_lsu_pkt_d_bits_store; // @[lsu_lsc_ctl.scala 113:25]
  wire  addrcheck_io_lsu_pkt_d_bits_dma; // @[lsu_lsc_ctl.scala 113:25]
  wire [31:0] addrcheck_io_dec_tlu_mrac_ff; // @[lsu_lsc_ctl.scala 113:25]
  wire [3:0] addrcheck_io_rs1_region_d; // @[lsu_lsc_ctl.scala 113:25]
  wire  addrcheck_io_is_sideeffects_m; // @[lsu_lsc_ctl.scala 113:25]
  wire  addrcheck_io_addr_in_dccm_d; // @[lsu_lsc_ctl.scala 113:25]
  wire  addrcheck_io_addr_in_pic_d; // @[lsu_lsc_ctl.scala 113:25]
  wire  addrcheck_io_addr_external_d; // @[lsu_lsc_ctl.scala 113:25]
  wire  addrcheck_io_access_fault_d; // @[lsu_lsc_ctl.scala 113:25]
  wire  addrcheck_io_misaligned_fault_d; // @[lsu_lsc_ctl.scala 113:25]
  wire [3:0] addrcheck_io_exc_mscause_d; // @[lsu_lsc_ctl.scala 113:25]
  wire  addrcheck_io_fir_dccm_access_error_d; // @[lsu_lsc_ctl.scala 113:25]
  wire  addrcheck_io_fir_nondccm_access_error_d; // @[lsu_lsc_ctl.scala 113:25]
  wire [31:0] lsu_rs1_d = io_dec_lsu_valid_raw_d ? io_lsu_exu_exu_lsu_rs1_d : io_dma_lsc_ctl_dma_mem_addr; // @[lsu_lsc_ctl.scala 95:28]
  wire [11:0] _T_3 = io_dec_lsu_valid_raw_d ? 12'hfff : 12'h0; // @[Bitwise.scala 72:12]
  wire [11:0] lsu_offset_d = io_dec_lsu_offset_d & _T_3; // @[lsu_lsc_ctl.scala 96:51]
  wire [31:0] rs1_d = io_lsu_pkt_d_bits_load_ldst_bypass_d ? io_lsu_result_m : lsu_rs1_d; // @[lsu_lsc_ctl.scala 99:28]
  wire [12:0] _T_6 = {1'h0,rs1_d[11:0]}; // @[Cat.scala 29:58]
  wire [12:0] _T_8 = {1'h0,lsu_offset_d}; // @[Cat.scala 29:58]
  wire [12:0] _T_10 = _T_6 + _T_8; // @[lib.scala 92:39]
  wire  _T_13 = lsu_offset_d[11] ^ _T_10[12]; // @[lib.scala 93:46]
  wire  _T_14 = ~_T_13; // @[lib.scala 93:33]
  wire [19:0] _T_16 = _T_14 ? 20'hfffff : 20'h0; // @[Bitwise.scala 72:12]
  wire [19:0] _T_18 = _T_16 & rs1_d[31:12]; // @[lib.scala 93:58]
  wire  _T_20 = ~lsu_offset_d[11]; // @[lib.scala 94:18]
  wire  _T_22 = _T_20 & _T_10[12]; // @[lib.scala 94:30]
  wire [19:0] _T_24 = _T_22 ? 20'hfffff : 20'h0; // @[Bitwise.scala 72:12]
  wire [19:0] _T_27 = rs1_d[31:12] + 20'h1; // @[lib.scala 94:54]
  wire [19:0] _T_28 = _T_24 & _T_27; // @[lib.scala 94:41]
  wire [19:0] _T_29 = _T_18 | _T_28; // @[lib.scala 93:72]
  wire  _T_32 = ~_T_10[12]; // @[lib.scala 95:31]
  wire  _T_33 = lsu_offset_d[11] & _T_32; // @[lib.scala 95:29]
  wire [19:0] _T_35 = _T_33 ? 20'hfffff : 20'h0; // @[Bitwise.scala 72:12]
  wire [19:0] _T_38 = rs1_d[31:12] - 20'h1; // @[lib.scala 95:54]
  wire [19:0] _T_39 = _T_35 & _T_38; // @[lib.scala 95:41]
  wire [19:0] _T_40 = _T_29 | _T_39; // @[lib.scala 94:61]
  wire [2:0] _T_43 = io_lsu_pkt_d_bits_half ? 3'h7 : 3'h0; // @[Bitwise.scala 72:12]
  wire [2:0] _T_44 = _T_43 & 3'h1; // @[lsu_lsc_ctl.scala 104:58]
  wire [2:0] _T_46 = io_lsu_pkt_d_bits_word ? 3'h7 : 3'h0; // @[Bitwise.scala 72:12]
  wire [2:0] _T_47 = _T_46 & 3'h3; // @[lsu_lsc_ctl.scala 105:40]
  wire [2:0] _T_48 = _T_44 | _T_47; // @[lsu_lsc_ctl.scala 104:70]
  wire [2:0] _T_50 = io_lsu_pkt_d_bits_dword ? 3'h7 : 3'h0; // @[Bitwise.scala 72:12]
  wire [2:0] addr_offset_d = _T_48 | _T_50; // @[lsu_lsc_ctl.scala 105:52]
  wire [12:0] _T_54 = {lsu_offset_d[11],lsu_offset_d}; // @[Cat.scala 29:58]
  wire [11:0] _T_57 = {9'h0,addr_offset_d}; // @[Cat.scala 29:58]
  wire [12:0] _GEN_0 = {{1'd0}, _T_57}; // @[lsu_lsc_ctl.scala 108:60]
  wire [12:0] end_addr_offset_d = _T_54 + _GEN_0; // @[lsu_lsc_ctl.scala 108:60]
  wire [18:0] _T_62 = end_addr_offset_d[12] ? 19'h7ffff : 19'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_64 = {_T_62,end_addr_offset_d}; // @[Cat.scala 29:58]
  reg  access_fault_m; // @[lsu_lsc_ctl.scala 144:75]
  reg  misaligned_fault_m; // @[lsu_lsc_ctl.scala 145:75]
  reg [3:0] exc_mscause_m; // @[lsu_lsc_ctl.scala 146:75]
  reg  fir_dccm_access_error_m; // @[lsu_lsc_ctl.scala 147:75]
  reg  fir_nondccm_access_error_m; // @[lsu_lsc_ctl.scala 148:75]
  wire  _T_69 = access_fault_m | misaligned_fault_m; // @[lsu_lsc_ctl.scala 150:34]
  wire  _T_70 = ~io_lsu_double_ecc_error_r; // @[lsu_lsc_ctl.scala 151:64]
  wire  _T_71 = io_lsu_single_ecc_error_r & _T_70; // @[lsu_lsc_ctl.scala 151:62]
  wire  _T_72 = io_lsu_commit_r | io_lsu_pkt_r_bits_dma; // @[lsu_lsc_ctl.scala 151:111]
  wire  _T_73 = _T_71 & _T_72; // @[lsu_lsc_ctl.scala 151:92]
  wire  _T_76 = _T_69 | io_lsu_double_ecc_error_m; // @[lsu_lsc_ctl.scala 173:67]
  wire  _T_77 = _T_76 & io_lsu_pkt_m_valid; // @[lsu_lsc_ctl.scala 173:96]
  wire  _T_78 = ~io_lsu_pkt_m_bits_dma; // @[lsu_lsc_ctl.scala 173:119]
  wire  _T_79 = _T_77 & _T_78; // @[lsu_lsc_ctl.scala 173:117]
  wire  _T_80 = ~io_lsu_pkt_m_bits_fast_int; // @[lsu_lsc_ctl.scala 173:144]
  wire  _T_81 = _T_79 & _T_80; // @[lsu_lsc_ctl.scala 173:142]
  wire  _T_82 = ~io_flush_m_up; // @[lsu_lsc_ctl.scala 173:174]
  wire  lsu_error_pkt_m_valid = _T_81 & _T_82; // @[lsu_lsc_ctl.scala 173:172]
  wire  _T_84 = ~lsu_error_pkt_m_valid; // @[lsu_lsc_ctl.scala 174:75]
  wire  _T_85 = io_lsu_single_ecc_error_m & _T_84; // @[lsu_lsc_ctl.scala 174:73]
  wire  lsu_error_pkt_m_bits_exc_type = ~misaligned_fault_m; // @[lsu_lsc_ctl.scala 176:46]
  wire  _T_90 = io_lsu_double_ecc_error_m & lsu_error_pkt_m_bits_exc_type; // @[lsu_lsc_ctl.scala 177:78]
  wire  _T_91 = ~access_fault_m; // @[lsu_lsc_ctl.scala 177:102]
  wire  _T_92 = _T_90 & _T_91; // @[lsu_lsc_ctl.scala 177:100]
  wire  _T_99 = io_lsu_pkt_m_bits_fast_int & io_lsu_double_ecc_error_m; // @[lsu_lsc_ctl.scala 179:166]
  reg  _T_105_valid; // @[lsu_lsc_ctl.scala 180:75]
  reg  _T_105_bits_single_ecc_error; // @[lsu_lsc_ctl.scala 180:75]
  reg  _T_105_bits_inst_type; // @[lsu_lsc_ctl.scala 180:75]
  reg  _T_105_bits_exc_type; // @[lsu_lsc_ctl.scala 180:75]
  reg [3:0] _T_105_bits_mscause; // @[lsu_lsc_ctl.scala 180:75]
  reg [31:0] _T_105_bits_addr; // @[lsu_lsc_ctl.scala 180:75]
  reg [1:0] _T_106; // @[lsu_lsc_ctl.scala 181:75]
  wire  dma_pkt_d_bits_load = ~io_dma_lsc_ctl_dma_mem_write; // @[lsu_lsc_ctl.scala 188:30]
  wire  dma_pkt_d_bits_by = io_dma_lsc_ctl_dma_mem_sz == 3'h0; // @[lsu_lsc_ctl.scala 189:62]
  wire  dma_pkt_d_bits_half = io_dma_lsc_ctl_dma_mem_sz == 3'h1; // @[lsu_lsc_ctl.scala 190:62]
  wire  dma_pkt_d_bits_word = io_dma_lsc_ctl_dma_mem_sz == 3'h2; // @[lsu_lsc_ctl.scala 191:62]
  wire  dma_pkt_d_bits_dword = io_dma_lsc_ctl_dma_mem_sz == 3'h3; // @[lsu_lsc_ctl.scala 192:62]
  wire  _T_118 = ~io_lsu_p_bits_fast_int; // @[lsu_lsc_ctl.scala 205:64]
  wire  _T_119 = io_flush_m_up & _T_118; // @[lsu_lsc_ctl.scala 205:61]
  wire  _T_120 = ~_T_119; // @[lsu_lsc_ctl.scala 205:45]
  wire  _T_121 = io_lsu_p_valid & _T_120; // @[lsu_lsc_ctl.scala 205:43]
  wire  _T_123 = ~io_lsu_pkt_d_bits_dma; // @[lsu_lsc_ctl.scala 206:68]
  wire  _T_124 = io_flush_m_up & _T_123; // @[lsu_lsc_ctl.scala 206:65]
  wire  _T_125 = ~_T_124; // @[lsu_lsc_ctl.scala 206:49]
  wire  _T_128 = io_flush_m_up & _T_78; // @[lsu_lsc_ctl.scala 207:65]
  wire  _T_129 = ~_T_128; // @[lsu_lsc_ctl.scala 207:49]
  reg  _T_132_bits_fast_int; // @[lsu_lsc_ctl.scala 209:65]
  reg  _T_132_bits_by; // @[lsu_lsc_ctl.scala 209:65]
  reg  _T_132_bits_half; // @[lsu_lsc_ctl.scala 209:65]
  reg  _T_132_bits_word; // @[lsu_lsc_ctl.scala 209:65]
  reg  _T_132_bits_dword; // @[lsu_lsc_ctl.scala 209:65]
  reg  _T_132_bits_load; // @[lsu_lsc_ctl.scala 209:65]
  reg  _T_132_bits_store; // @[lsu_lsc_ctl.scala 209:65]
  reg  _T_132_bits_unsign; // @[lsu_lsc_ctl.scala 209:65]
  reg  _T_132_bits_dma; // @[lsu_lsc_ctl.scala 209:65]
  reg  _T_132_bits_store_data_bypass_m; // @[lsu_lsc_ctl.scala 209:65]
  reg  _T_134_bits_by; // @[lsu_lsc_ctl.scala 210:65]
  reg  _T_134_bits_half; // @[lsu_lsc_ctl.scala 210:65]
  reg  _T_134_bits_word; // @[lsu_lsc_ctl.scala 210:65]
  reg  _T_134_bits_dword; // @[lsu_lsc_ctl.scala 210:65]
  reg  _T_134_bits_load; // @[lsu_lsc_ctl.scala 210:65]
  reg  _T_134_bits_store; // @[lsu_lsc_ctl.scala 210:65]
  reg  _T_134_bits_unsign; // @[lsu_lsc_ctl.scala 210:65]
  reg  _T_134_bits_dma; // @[lsu_lsc_ctl.scala 210:65]
  reg  _T_135; // @[lsu_lsc_ctl.scala 211:65]
  reg  _T_136; // @[lsu_lsc_ctl.scala 212:65]
  wire [5:0] _T_139 = {io_dma_lsc_ctl_dma_mem_addr[2:0],3'h0}; // @[Cat.scala 29:58]
  wire [63:0] dma_mem_wdata_shifted = io_dma_lsc_ctl_dma_mem_wdata >> _T_139; // @[lsu_lsc_ctl.scala 214:66]
  reg [31:0] store_data_pre_m; // @[lsu_lsc_ctl.scala 218:72]
  reg [31:0] _T_146; // @[lsu_lsc_ctl.scala 219:62]
  reg [31:0] _T_147; // @[lsu_lsc_ctl.scala 220:62]
  reg [31:0] _T_148; // @[lsu_lsc_ctl.scala 221:62]
  reg [31:0] _T_149; // @[lsu_lsc_ctl.scala 222:62]
  reg  _T_150; // @[lsu_lsc_ctl.scala 223:62]
  reg  _T_151; // @[lsu_lsc_ctl.scala 224:62]
  reg  _T_152; // @[lsu_lsc_ctl.scala 225:62]
  reg  _T_153; // @[lsu_lsc_ctl.scala 226:62]
  reg  _T_154; // @[lsu_lsc_ctl.scala 227:62]
  reg  addr_external_r; // @[lsu_lsc_ctl.scala 228:66]
  reg [31:0] bus_read_data_r; // @[lsu_lsc_ctl.scala 229:66]
  wire  _T_156 = io_lsu_pkt_r_bits_store | io_lsu_pkt_r_bits_load; // @[lsu_lsc_ctl.scala 235:68]
  wire  _T_157 = io_lsu_pkt_r_valid & _T_156; // @[lsu_lsc_ctl.scala 235:41]
  wire  _T_158 = ~io_flush_r; // @[lsu_lsc_ctl.scala 235:96]
  wire  _T_159 = _T_157 & _T_158; // @[lsu_lsc_ctl.scala 235:94]
  wire  _T_160 = ~io_lsu_pkt_r_bits_dma; // @[lsu_lsc_ctl.scala 235:110]
  wire  _T_163 = ~io_addr_in_pic_m; // @[lsu_lsc_ctl.scala 236:69]
  wire [31:0] _T_165 = _T_163 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_166 = io_picm_mask_data_m | _T_165; // @[lsu_lsc_ctl.scala 236:59]
  wire [31:0] _T_168 = io_lsu_pkt_m_bits_store_data_bypass_m ? io_lsu_result_m : store_data_pre_m; // @[lsu_lsc_ctl.scala 236:94]
  wire [31:0] lsu_ld_datafn_m = io_addr_external_m ? io_bus_read_data_m : io_lsu_ld_data_m; // @[lsu_lsc_ctl.scala 257:33]
  wire [31:0] lsu_ld_datafn_corr_r = addr_external_r ? bus_read_data_r : io_lsu_ld_data_corr_r; // @[lsu_lsc_ctl.scala 258:33]
  wire  _T_174 = io_lsu_pkt_m_bits_unsign & io_lsu_pkt_m_bits_by; // @[lsu_lsc_ctl.scala 259:66]
  wire [31:0] _T_176 = _T_174 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_178 = {24'h0,lsu_ld_datafn_m[7:0]}; // @[Cat.scala 29:58]
  wire [31:0] _T_179 = _T_176 & _T_178; // @[lsu_lsc_ctl.scala 259:94]
  wire  _T_180 = io_lsu_pkt_m_bits_unsign & io_lsu_pkt_m_bits_half; // @[lsu_lsc_ctl.scala 260:43]
  wire [31:0] _T_182 = _T_180 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_184 = {16'h0,lsu_ld_datafn_m[15:0]}; // @[Cat.scala 29:58]
  wire [31:0] _T_185 = _T_182 & _T_184; // @[lsu_lsc_ctl.scala 260:71]
  wire [31:0] _T_186 = _T_179 | _T_185; // @[lsu_lsc_ctl.scala 259:133]
  wire  _T_187 = ~io_lsu_pkt_m_bits_unsign; // @[lsu_lsc_ctl.scala 261:17]
  wire  _T_188 = _T_187 & io_lsu_pkt_m_bits_by; // @[lsu_lsc_ctl.scala 261:43]
  wire [31:0] _T_190 = _T_188 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [23:0] _T_193 = lsu_ld_datafn_m[7] ? 24'hffffff : 24'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_195 = {_T_193,lsu_ld_datafn_m[7:0]}; // @[Cat.scala 29:58]
  wire [31:0] _T_196 = _T_190 & _T_195; // @[lsu_lsc_ctl.scala 261:71]
  wire [31:0] _T_197 = _T_186 | _T_196; // @[lsu_lsc_ctl.scala 260:114]
  wire  _T_199 = _T_187 & io_lsu_pkt_m_bits_half; // @[lsu_lsc_ctl.scala 262:43]
  wire [31:0] _T_201 = _T_199 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _T_204 = lsu_ld_datafn_m[15] ? 16'hffff : 16'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_206 = {_T_204,lsu_ld_datafn_m[15:0]}; // @[Cat.scala 29:58]
  wire [31:0] _T_207 = _T_201 & _T_206; // @[lsu_lsc_ctl.scala 262:71]
  wire [31:0] _T_208 = _T_197 | _T_207; // @[lsu_lsc_ctl.scala 261:134]
  wire [31:0] _T_210 = io_lsu_pkt_m_bits_word ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_212 = _T_210 & lsu_ld_datafn_m; // @[lsu_lsc_ctl.scala 263:43]
  wire  _T_214 = io_lsu_pkt_r_bits_unsign & io_lsu_pkt_r_bits_by; // @[lsu_lsc_ctl.scala 264:66]
  wire [31:0] _T_216 = _T_214 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_218 = {24'h0,lsu_ld_datafn_corr_r[7:0]}; // @[Cat.scala 29:58]
  wire [31:0] _T_219 = _T_216 & _T_218; // @[lsu_lsc_ctl.scala 264:94]
  wire  _T_220 = io_lsu_pkt_r_bits_unsign & io_lsu_pkt_r_bits_half; // @[lsu_lsc_ctl.scala 265:43]
  wire [31:0] _T_222 = _T_220 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_224 = {16'h0,lsu_ld_datafn_corr_r[15:0]}; // @[Cat.scala 29:58]
  wire [31:0] _T_225 = _T_222 & _T_224; // @[lsu_lsc_ctl.scala 265:71]
  wire [31:0] _T_226 = _T_219 | _T_225; // @[lsu_lsc_ctl.scala 264:138]
  wire  _T_227 = ~io_lsu_pkt_r_bits_unsign; // @[lsu_lsc_ctl.scala 266:17]
  wire  _T_228 = _T_227 & io_lsu_pkt_r_bits_by; // @[lsu_lsc_ctl.scala 266:43]
  wire [31:0] _T_230 = _T_228 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [23:0] _T_233 = lsu_ld_datafn_corr_r[7] ? 24'hffffff : 24'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_235 = {_T_233,lsu_ld_datafn_corr_r[7:0]}; // @[Cat.scala 29:58]
  wire [31:0] _T_236 = _T_230 & _T_235; // @[lsu_lsc_ctl.scala 266:71]
  wire [31:0] _T_237 = _T_226 | _T_236; // @[lsu_lsc_ctl.scala 265:119]
  wire  _T_239 = _T_227 & io_lsu_pkt_r_bits_half; // @[lsu_lsc_ctl.scala 267:43]
  wire [31:0] _T_241 = _T_239 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _T_244 = lsu_ld_datafn_corr_r[15] ? 16'hffff : 16'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_246 = {_T_244,lsu_ld_datafn_corr_r[15:0]}; // @[Cat.scala 29:58]
  wire [31:0] _T_247 = _T_241 & _T_246; // @[lsu_lsc_ctl.scala 267:71]
  wire [31:0] _T_248 = _T_237 | _T_247; // @[lsu_lsc_ctl.scala 266:144]
  wire [31:0] _T_250 = io_lsu_pkt_r_bits_word ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_252 = _T_250 & lsu_ld_datafn_corr_r; // @[lsu_lsc_ctl.scala 268:43]
  lsu_addrcheck addrcheck ( // @[lsu_lsc_ctl.scala 113:25]
    .reset(addrcheck_reset),
    .io_lsu_c2_m_clk(addrcheck_io_lsu_c2_m_clk),
    .io_start_addr_d(addrcheck_io_start_addr_d),
    .io_end_addr_d(addrcheck_io_end_addr_d),
    .io_lsu_pkt_d_valid(addrcheck_io_lsu_pkt_d_valid),
    .io_lsu_pkt_d_bits_fast_int(addrcheck_io_lsu_pkt_d_bits_fast_int),
    .io_lsu_pkt_d_bits_by(addrcheck_io_lsu_pkt_d_bits_by),
    .io_lsu_pkt_d_bits_half(addrcheck_io_lsu_pkt_d_bits_half),
    .io_lsu_pkt_d_bits_word(addrcheck_io_lsu_pkt_d_bits_word),
    .io_lsu_pkt_d_bits_load(addrcheck_io_lsu_pkt_d_bits_load),
    .io_lsu_pkt_d_bits_store(addrcheck_io_lsu_pkt_d_bits_store),
    .io_lsu_pkt_d_bits_dma(addrcheck_io_lsu_pkt_d_bits_dma),
    .io_dec_tlu_mrac_ff(addrcheck_io_dec_tlu_mrac_ff),
    .io_rs1_region_d(addrcheck_io_rs1_region_d),
    .io_is_sideeffects_m(addrcheck_io_is_sideeffects_m),
    .io_addr_in_dccm_d(addrcheck_io_addr_in_dccm_d),
    .io_addr_in_pic_d(addrcheck_io_addr_in_pic_d),
    .io_addr_external_d(addrcheck_io_addr_external_d),
    .io_access_fault_d(addrcheck_io_access_fault_d),
    .io_misaligned_fault_d(addrcheck_io_misaligned_fault_d),
    .io_exc_mscause_d(addrcheck_io_exc_mscause_d),
    .io_fir_dccm_access_error_d(addrcheck_io_fir_dccm_access_error_d),
    .io_fir_nondccm_access_error_d(addrcheck_io_fir_nondccm_access_error_d)
  );
  assign io_lsu_result_m = _T_208 | _T_212; // @[lsu_lsc_ctl.scala 259:27]
  assign io_lsu_result_corr_r = _T_248 | _T_252; // @[lsu_lsc_ctl.scala 264:27]
  assign io_lsu_addr_d = {_T_40,_T_10[11:0]}; // @[lsu_lsc_ctl.scala 233:28]
  assign io_lsu_addr_m = _T_146; // @[lsu_lsc_ctl.scala 219:24]
  assign io_lsu_addr_r = _T_147; // @[lsu_lsc_ctl.scala 220:24]
  assign io_end_addr_d = rs1_d + _T_64; // @[lsu_lsc_ctl.scala 110:24]
  assign io_end_addr_m = _T_148; // @[lsu_lsc_ctl.scala 221:24]
  assign io_end_addr_r = _T_149; // @[lsu_lsc_ctl.scala 222:24]
  assign io_store_data_m = _T_166 & _T_168; // @[lsu_lsc_ctl.scala 236:29]
  assign io_lsu_exc_m = access_fault_m | misaligned_fault_m; // @[lsu_lsc_ctl.scala 150:16]
  assign io_is_sideeffects_m = addrcheck_io_is_sideeffects_m; // @[lsu_lsc_ctl.scala 123:42]
  assign io_lsu_commit_r = _T_159 & _T_160; // @[lsu_lsc_ctl.scala 235:19]
  assign io_lsu_single_ecc_error_incr = _T_73 & io_lsu_pkt_r_valid; // @[lsu_lsc_ctl.scala 151:32]
  assign io_lsu_error_pkt_r_valid = _T_105_valid; // @[lsu_lsc_ctl.scala 180:38]
  assign io_lsu_error_pkt_r_bits_single_ecc_error = _T_105_bits_single_ecc_error; // @[lsu_lsc_ctl.scala 180:38]
  assign io_lsu_error_pkt_r_bits_inst_type = _T_105_bits_inst_type; // @[lsu_lsc_ctl.scala 180:38]
  assign io_lsu_error_pkt_r_bits_exc_type = _T_105_bits_exc_type; // @[lsu_lsc_ctl.scala 180:38]
  assign io_lsu_error_pkt_r_bits_mscause = _T_105_bits_mscause; // @[lsu_lsc_ctl.scala 180:38]
  assign io_lsu_error_pkt_r_bits_addr = _T_105_bits_addr; // @[lsu_lsc_ctl.scala 180:38]
  assign io_lsu_fir_addr = io_lsu_ld_data_corr_r[31:1]; // @[lsu_lsc_ctl.scala 231:28]
  assign io_lsu_fir_error = _T_106; // @[lsu_lsc_ctl.scala 181:38]
  assign io_addr_in_dccm_d = addrcheck_io_addr_in_dccm_d; // @[lsu_lsc_ctl.scala 124:42]
  assign io_addr_in_dccm_m = _T_150; // @[lsu_lsc_ctl.scala 223:24]
  assign io_addr_in_dccm_r = _T_151; // @[lsu_lsc_ctl.scala 224:24]
  assign io_addr_in_pic_d = addrcheck_io_addr_in_pic_d; // @[lsu_lsc_ctl.scala 125:42]
  assign io_addr_in_pic_m = _T_152; // @[lsu_lsc_ctl.scala 225:24]
  assign io_addr_in_pic_r = _T_153; // @[lsu_lsc_ctl.scala 226:24]
  assign io_addr_external_m = _T_154; // @[lsu_lsc_ctl.scala 227:24]
  assign io_lsu_pkt_d_valid = _T_121 | io_dma_lsc_ctl_dma_dccm_req; // @[lsu_lsc_ctl.scala 201:20 lsu_lsc_ctl.scala 205:24]
  assign io_lsu_pkt_d_bits_fast_int = io_dec_lsu_valid_raw_d & io_lsu_p_bits_fast_int; // @[lsu_lsc_ctl.scala 201:20]
  assign io_lsu_pkt_d_bits_by = io_dec_lsu_valid_raw_d ? io_lsu_p_bits_by : dma_pkt_d_bits_by; // @[lsu_lsc_ctl.scala 201:20]
  assign io_lsu_pkt_d_bits_half = io_dec_lsu_valid_raw_d ? io_lsu_p_bits_half : dma_pkt_d_bits_half; // @[lsu_lsc_ctl.scala 201:20]
  assign io_lsu_pkt_d_bits_word = io_dec_lsu_valid_raw_d ? io_lsu_p_bits_word : dma_pkt_d_bits_word; // @[lsu_lsc_ctl.scala 201:20]
  assign io_lsu_pkt_d_bits_dword = io_dec_lsu_valid_raw_d ? 1'h0 : dma_pkt_d_bits_dword; // @[lsu_lsc_ctl.scala 201:20]
  assign io_lsu_pkt_d_bits_load = io_dec_lsu_valid_raw_d ? io_lsu_p_bits_load : dma_pkt_d_bits_load; // @[lsu_lsc_ctl.scala 201:20]
  assign io_lsu_pkt_d_bits_store = io_dec_lsu_valid_raw_d ? io_lsu_p_bits_store : io_dma_lsc_ctl_dma_mem_write; // @[lsu_lsc_ctl.scala 201:20]
  assign io_lsu_pkt_d_bits_unsign = io_dec_lsu_valid_raw_d & io_lsu_p_bits_unsign; // @[lsu_lsc_ctl.scala 201:20]
  assign io_lsu_pkt_d_bits_dma = io_dec_lsu_valid_raw_d ? 1'h0 : 1'h1; // @[lsu_lsc_ctl.scala 201:20]
  assign io_lsu_pkt_d_bits_store_data_bypass_d = io_dec_lsu_valid_raw_d & io_lsu_p_bits_store_data_bypass_d; // @[lsu_lsc_ctl.scala 201:20]
  assign io_lsu_pkt_d_bits_load_ldst_bypass_d = io_dec_lsu_valid_raw_d & io_lsu_p_bits_load_ldst_bypass_d; // @[lsu_lsc_ctl.scala 201:20]
  assign io_lsu_pkt_d_bits_store_data_bypass_m = 1'h0; // @[lsu_lsc_ctl.scala 201:20]
  assign io_lsu_pkt_m_valid = _T_135; // @[lsu_lsc_ctl.scala 209:28 lsu_lsc_ctl.scala 211:28]
  assign io_lsu_pkt_m_bits_fast_int = _T_132_bits_fast_int; // @[lsu_lsc_ctl.scala 209:28]
  assign io_lsu_pkt_m_bits_by = _T_132_bits_by; // @[lsu_lsc_ctl.scala 209:28]
  assign io_lsu_pkt_m_bits_half = _T_132_bits_half; // @[lsu_lsc_ctl.scala 209:28]
  assign io_lsu_pkt_m_bits_word = _T_132_bits_word; // @[lsu_lsc_ctl.scala 209:28]
  assign io_lsu_pkt_m_bits_dword = _T_132_bits_dword; // @[lsu_lsc_ctl.scala 209:28]
  assign io_lsu_pkt_m_bits_load = _T_132_bits_load; // @[lsu_lsc_ctl.scala 209:28]
  assign io_lsu_pkt_m_bits_store = _T_132_bits_store; // @[lsu_lsc_ctl.scala 209:28]
  assign io_lsu_pkt_m_bits_unsign = _T_132_bits_unsign; // @[lsu_lsc_ctl.scala 209:28]
  assign io_lsu_pkt_m_bits_dma = _T_132_bits_dma; // @[lsu_lsc_ctl.scala 209:28]
  assign io_lsu_pkt_m_bits_store_data_bypass_m = _T_132_bits_store_data_bypass_m; // @[lsu_lsc_ctl.scala 209:28]
  assign io_lsu_pkt_r_valid = _T_136; // @[lsu_lsc_ctl.scala 210:28 lsu_lsc_ctl.scala 212:28]
  assign io_lsu_pkt_r_bits_by = _T_134_bits_by; // @[lsu_lsc_ctl.scala 210:28]
  assign io_lsu_pkt_r_bits_half = _T_134_bits_half; // @[lsu_lsc_ctl.scala 210:28]
  assign io_lsu_pkt_r_bits_word = _T_134_bits_word; // @[lsu_lsc_ctl.scala 210:28]
  assign io_lsu_pkt_r_bits_dword = _T_134_bits_dword; // @[lsu_lsc_ctl.scala 210:28]
  assign io_lsu_pkt_r_bits_load = _T_134_bits_load; // @[lsu_lsc_ctl.scala 210:28]
  assign io_lsu_pkt_r_bits_store = _T_134_bits_store; // @[lsu_lsc_ctl.scala 210:28]
  assign io_lsu_pkt_r_bits_unsign = _T_134_bits_unsign; // @[lsu_lsc_ctl.scala 210:28]
  assign io_lsu_pkt_r_bits_dma = _T_134_bits_dma; // @[lsu_lsc_ctl.scala 210:28]
  assign addrcheck_reset = reset;
  assign addrcheck_io_lsu_c2_m_clk = io_lsu_c2_m_clk; // @[lsu_lsc_ctl.scala 115:42]
  assign addrcheck_io_start_addr_d = {_T_40,_T_10[11:0]}; // @[lsu_lsc_ctl.scala 117:42]
  assign addrcheck_io_end_addr_d = rs1_d + _T_64; // @[lsu_lsc_ctl.scala 118:42]
  assign addrcheck_io_lsu_pkt_d_valid = io_lsu_pkt_d_valid; // @[lsu_lsc_ctl.scala 119:42]
  assign addrcheck_io_lsu_pkt_d_bits_fast_int = io_lsu_pkt_d_bits_fast_int; // @[lsu_lsc_ctl.scala 119:42]
  assign addrcheck_io_lsu_pkt_d_bits_by = io_lsu_pkt_d_bits_by; // @[lsu_lsc_ctl.scala 119:42]
  assign addrcheck_io_lsu_pkt_d_bits_half = io_lsu_pkt_d_bits_half; // @[lsu_lsc_ctl.scala 119:42]
  assign addrcheck_io_lsu_pkt_d_bits_word = io_lsu_pkt_d_bits_word; // @[lsu_lsc_ctl.scala 119:42]
  assign addrcheck_io_lsu_pkt_d_bits_load = io_lsu_pkt_d_bits_load; // @[lsu_lsc_ctl.scala 119:42]
  assign addrcheck_io_lsu_pkt_d_bits_store = io_lsu_pkt_d_bits_store; // @[lsu_lsc_ctl.scala 119:42]
  assign addrcheck_io_lsu_pkt_d_bits_dma = io_lsu_pkt_d_bits_dma; // @[lsu_lsc_ctl.scala 119:42]
  assign addrcheck_io_dec_tlu_mrac_ff = io_dec_tlu_mrac_ff; // @[lsu_lsc_ctl.scala 120:42]
  assign addrcheck_io_rs1_region_d = rs1_d[31:28]; // @[lsu_lsc_ctl.scala 121:42]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  access_fault_m = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  misaligned_fault_m = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  exc_mscause_m = _RAND_2[3:0];
  _RAND_3 = {1{`RANDOM}};
  fir_dccm_access_error_m = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  fir_nondccm_access_error_m = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  _T_105_valid = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  _T_105_bits_single_ecc_error = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  _T_105_bits_inst_type = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  _T_105_bits_exc_type = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  _T_105_bits_mscause = _RAND_9[3:0];
  _RAND_10 = {1{`RANDOM}};
  _T_105_bits_addr = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  _T_106 = _RAND_11[1:0];
  _RAND_12 = {1{`RANDOM}};
  _T_132_bits_fast_int = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  _T_132_bits_by = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  _T_132_bits_half = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  _T_132_bits_word = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  _T_132_bits_dword = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  _T_132_bits_load = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  _T_132_bits_store = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  _T_132_bits_unsign = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  _T_132_bits_dma = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  _T_132_bits_store_data_bypass_m = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  _T_134_bits_by = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  _T_134_bits_half = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  _T_134_bits_word = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  _T_134_bits_dword = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  _T_134_bits_load = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  _T_134_bits_store = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  _T_134_bits_unsign = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  _T_134_bits_dma = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  _T_135 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  _T_136 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  store_data_pre_m = _RAND_32[31:0];
  _RAND_33 = {1{`RANDOM}};
  _T_146 = _RAND_33[31:0];
  _RAND_34 = {1{`RANDOM}};
  _T_147 = _RAND_34[31:0];
  _RAND_35 = {1{`RANDOM}};
  _T_148 = _RAND_35[31:0];
  _RAND_36 = {1{`RANDOM}};
  _T_149 = _RAND_36[31:0];
  _RAND_37 = {1{`RANDOM}};
  _T_150 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  _T_151 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  _T_152 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  _T_153 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  _T_154 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  addr_external_r = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  bus_read_data_r = _RAND_43[31:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    access_fault_m = 1'h0;
  end
  if (reset) begin
    misaligned_fault_m = 1'h0;
  end
  if (reset) begin
    exc_mscause_m = 4'h0;
  end
  if (reset) begin
    fir_dccm_access_error_m = 1'h0;
  end
  if (reset) begin
    fir_nondccm_access_error_m = 1'h0;
  end
  if (reset) begin
    _T_105_valid = 1'h0;
  end
  if (reset) begin
    _T_105_bits_single_ecc_error = 1'h0;
  end
  if (reset) begin
    _T_105_bits_inst_type = 1'h0;
  end
  if (reset) begin
    _T_105_bits_exc_type = 1'h0;
  end
  if (reset) begin
    _T_105_bits_mscause = 4'h0;
  end
  if (reset) begin
    _T_105_bits_addr = 32'h0;
  end
  if (reset) begin
    _T_106 = 2'h0;
  end
  if (reset) begin
    _T_132_bits_fast_int = 1'h0;
  end
  if (reset) begin
    _T_132_bits_by = 1'h0;
  end
  if (reset) begin
    _T_132_bits_half = 1'h0;
  end
  if (reset) begin
    _T_132_bits_word = 1'h0;
  end
  if (reset) begin
    _T_132_bits_dword = 1'h0;
  end
  if (reset) begin
    _T_132_bits_load = 1'h0;
  end
  if (reset) begin
    _T_132_bits_store = 1'h0;
  end
  if (reset) begin
    _T_132_bits_unsign = 1'h0;
  end
  if (reset) begin
    _T_132_bits_dma = 1'h0;
  end
  if (reset) begin
    _T_132_bits_store_data_bypass_m = 1'h0;
  end
  if (reset) begin
    _T_134_bits_by = 1'h0;
  end
  if (reset) begin
    _T_134_bits_half = 1'h0;
  end
  if (reset) begin
    _T_134_bits_word = 1'h0;
  end
  if (reset) begin
    _T_134_bits_dword = 1'h0;
  end
  if (reset) begin
    _T_134_bits_load = 1'h0;
  end
  if (reset) begin
    _T_134_bits_store = 1'h0;
  end
  if (reset) begin
    _T_134_bits_unsign = 1'h0;
  end
  if (reset) begin
    _T_134_bits_dma = 1'h0;
  end
  if (reset) begin
    _T_135 = 1'h0;
  end
  if (reset) begin
    _T_136 = 1'h0;
  end
  if (reset) begin
    store_data_pre_m = 32'h0;
  end
  if (reset) begin
    _T_146 = 32'h0;
  end
  if (reset) begin
    _T_147 = 32'h0;
  end
  if (reset) begin
    _T_148 = 32'h0;
  end
  if (reset) begin
    _T_149 = 32'h0;
  end
  if (reset) begin
    _T_150 = 1'h0;
  end
  if (reset) begin
    _T_151 = 1'h0;
  end
  if (reset) begin
    _T_152 = 1'h0;
  end
  if (reset) begin
    _T_153 = 1'h0;
  end
  if (reset) begin
    _T_154 = 1'h0;
  end
  if (reset) begin
    addr_external_r = 1'h0;
  end
  if (reset) begin
    bus_read_data_r = 32'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge io_lsu_c1_m_clk or posedge reset) begin
    if (reset) begin
      access_fault_m <= 1'h0;
    end else begin
      access_fault_m <= addrcheck_io_access_fault_d;
    end
  end
  always @(posedge io_lsu_c1_m_clk or posedge reset) begin
    if (reset) begin
      misaligned_fault_m <= 1'h0;
    end else begin
      misaligned_fault_m <= addrcheck_io_misaligned_fault_d;
    end
  end
  always @(posedge io_lsu_c1_m_clk or posedge reset) begin
    if (reset) begin
      exc_mscause_m <= 4'h0;
    end else begin
      exc_mscause_m <= addrcheck_io_exc_mscause_d;
    end
  end
  always @(posedge io_lsu_c1_m_clk or posedge reset) begin
    if (reset) begin
      fir_dccm_access_error_m <= 1'h0;
    end else begin
      fir_dccm_access_error_m <= addrcheck_io_fir_dccm_access_error_d;
    end
  end
  always @(posedge io_lsu_c1_m_clk or posedge reset) begin
    if (reset) begin
      fir_nondccm_access_error_m <= 1'h0;
    end else begin
      fir_nondccm_access_error_m <= addrcheck_io_fir_nondccm_access_error_d;
    end
  end
  always @(posedge io_lsu_c2_r_clk or posedge reset) begin
    if (reset) begin
      _T_105_valid <= 1'h0;
    end else begin
      _T_105_valid <= _T_81 & _T_82;
    end
  end
  always @(posedge io_lsu_c2_r_clk or posedge reset) begin
    if (reset) begin
      _T_105_bits_single_ecc_error <= 1'h0;
    end else begin
      _T_105_bits_single_ecc_error <= _T_85 & _T_78;
    end
  end
  always @(posedge io_lsu_c2_r_clk or posedge reset) begin
    if (reset) begin
      _T_105_bits_inst_type <= 1'h0;
    end else begin
      _T_105_bits_inst_type <= io_lsu_pkt_m_bits_store;
    end
  end
  always @(posedge io_lsu_c2_r_clk or posedge reset) begin
    if (reset) begin
      _T_105_bits_exc_type <= 1'h0;
    end else begin
      _T_105_bits_exc_type <= ~misaligned_fault_m;
    end
  end
  always @(posedge io_lsu_c2_r_clk or posedge reset) begin
    if (reset) begin
      _T_105_bits_mscause <= 4'h0;
    end else if (_T_92) begin
      _T_105_bits_mscause <= 4'h1;
    end else begin
      _T_105_bits_mscause <= exc_mscause_m;
    end
  end
  always @(posedge io_lsu_c2_r_clk or posedge reset) begin
    if (reset) begin
      _T_105_bits_addr <= 32'h0;
    end else begin
      _T_105_bits_addr <= io_lsu_addr_m;
    end
  end
  always @(posedge io_lsu_c2_r_clk or posedge reset) begin
    if (reset) begin
      _T_106 <= 2'h0;
    end else if (fir_nondccm_access_error_m) begin
      _T_106 <= 2'h3;
    end else if (fir_dccm_access_error_m) begin
      _T_106 <= 2'h2;
    end else if (_T_99) begin
      _T_106 <= 2'h1;
    end else begin
      _T_106 <= 2'h0;
    end
  end
  always @(posedge io_lsu_c1_m_clk or posedge reset) begin
    if (reset) begin
      _T_132_bits_fast_int <= 1'h0;
    end else begin
      _T_132_bits_fast_int <= io_lsu_pkt_d_bits_fast_int;
    end
  end
  always @(posedge io_lsu_c1_m_clk or posedge reset) begin
    if (reset) begin
      _T_132_bits_by <= 1'h0;
    end else begin
      _T_132_bits_by <= io_lsu_pkt_d_bits_by;
    end
  end
  always @(posedge io_lsu_c1_m_clk or posedge reset) begin
    if (reset) begin
      _T_132_bits_half <= 1'h0;
    end else begin
      _T_132_bits_half <= io_lsu_pkt_d_bits_half;
    end
  end
  always @(posedge io_lsu_c1_m_clk or posedge reset) begin
    if (reset) begin
      _T_132_bits_word <= 1'h0;
    end else begin
      _T_132_bits_word <= io_lsu_pkt_d_bits_word;
    end
  end
  always @(posedge io_lsu_c1_m_clk or posedge reset) begin
    if (reset) begin
      _T_132_bits_dword <= 1'h0;
    end else begin
      _T_132_bits_dword <= io_lsu_pkt_d_bits_dword;
    end
  end
  always @(posedge io_lsu_c1_m_clk or posedge reset) begin
    if (reset) begin
      _T_132_bits_load <= 1'h0;
    end else begin
      _T_132_bits_load <= io_lsu_pkt_d_bits_load;
    end
  end
  always @(posedge io_lsu_c1_m_clk or posedge reset) begin
    if (reset) begin
      _T_132_bits_store <= 1'h0;
    end else begin
      _T_132_bits_store <= io_lsu_pkt_d_bits_store;
    end
  end
  always @(posedge io_lsu_c1_m_clk or posedge reset) begin
    if (reset) begin
      _T_132_bits_unsign <= 1'h0;
    end else begin
      _T_132_bits_unsign <= io_lsu_pkt_d_bits_unsign;
    end
  end
  always @(posedge io_lsu_c1_m_clk or posedge reset) begin
    if (reset) begin
      _T_132_bits_dma <= 1'h0;
    end else begin
      _T_132_bits_dma <= io_lsu_pkt_d_bits_dma;
    end
  end
  always @(posedge io_lsu_c1_m_clk or posedge reset) begin
    if (reset) begin
      _T_132_bits_store_data_bypass_m <= 1'h0;
    end else begin
      _T_132_bits_store_data_bypass_m <= io_lsu_pkt_d_bits_store_data_bypass_m;
    end
  end
  always @(posedge io_lsu_c1_r_clk or posedge reset) begin
    if (reset) begin
      _T_134_bits_by <= 1'h0;
    end else begin
      _T_134_bits_by <= io_lsu_pkt_m_bits_by;
    end
  end
  always @(posedge io_lsu_c1_r_clk or posedge reset) begin
    if (reset) begin
      _T_134_bits_half <= 1'h0;
    end else begin
      _T_134_bits_half <= io_lsu_pkt_m_bits_half;
    end
  end
  always @(posedge io_lsu_c1_r_clk or posedge reset) begin
    if (reset) begin
      _T_134_bits_word <= 1'h0;
    end else begin
      _T_134_bits_word <= io_lsu_pkt_m_bits_word;
    end
  end
  always @(posedge io_lsu_c1_r_clk or posedge reset) begin
    if (reset) begin
      _T_134_bits_dword <= 1'h0;
    end else begin
      _T_134_bits_dword <= io_lsu_pkt_m_bits_dword;
    end
  end
  always @(posedge io_lsu_c1_r_clk or posedge reset) begin
    if (reset) begin
      _T_134_bits_load <= 1'h0;
    end else begin
      _T_134_bits_load <= io_lsu_pkt_m_bits_load;
    end
  end
  always @(posedge io_lsu_c1_r_clk or posedge reset) begin
    if (reset) begin
      _T_134_bits_store <= 1'h0;
    end else begin
      _T_134_bits_store <= io_lsu_pkt_m_bits_store;
    end
  end
  always @(posedge io_lsu_c1_r_clk or posedge reset) begin
    if (reset) begin
      _T_134_bits_unsign <= 1'h0;
    end else begin
      _T_134_bits_unsign <= io_lsu_pkt_m_bits_unsign;
    end
  end
  always @(posedge io_lsu_c1_r_clk or posedge reset) begin
    if (reset) begin
      _T_134_bits_dma <= 1'h0;
    end else begin
      _T_134_bits_dma <= io_lsu_pkt_m_bits_dma;
    end
  end
  always @(posedge io_lsu_c2_m_clk or posedge reset) begin
    if (reset) begin
      _T_135 <= 1'h0;
    end else begin
      _T_135 <= io_lsu_pkt_d_valid & _T_125;
    end
  end
  always @(posedge io_lsu_c2_r_clk or posedge reset) begin
    if (reset) begin
      _T_136 <= 1'h0;
    end else begin
      _T_136 <= io_lsu_pkt_m_valid & _T_129;
    end
  end
  always @(posedge io_lsu_store_c1_m_clk or posedge reset) begin
    if (reset) begin
      store_data_pre_m <= 32'h0;
    end else if (io_lsu_pkt_d_bits_store_data_bypass_d) begin
      store_data_pre_m <= io_lsu_result_m;
    end else if (io_dma_lsc_ctl_dma_dccm_req) begin
      store_data_pre_m <= dma_mem_wdata_shifted[31:0];
    end else begin
      store_data_pre_m <= io_lsu_exu_exu_lsu_rs2_d;
    end
  end
  always @(posedge io_lsu_c1_m_clk or posedge reset) begin
    if (reset) begin
      _T_146 <= 32'h0;
    end else begin
      _T_146 <= io_lsu_addr_d;
    end
  end
  always @(posedge io_lsu_c1_r_clk or posedge reset) begin
    if (reset) begin
      _T_147 <= 32'h0;
    end else begin
      _T_147 <= io_lsu_addr_m;
    end
  end
  always @(posedge io_lsu_c1_m_clk or posedge reset) begin
    if (reset) begin
      _T_148 <= 32'h0;
    end else begin
      _T_148 <= io_end_addr_d;
    end
  end
  always @(posedge io_lsu_c1_r_clk or posedge reset) begin
    if (reset) begin
      _T_149 <= 32'h0;
    end else begin
      _T_149 <= io_end_addr_m;
    end
  end
  always @(posedge io_lsu_c1_m_clk or posedge reset) begin
    if (reset) begin
      _T_150 <= 1'h0;
    end else begin
      _T_150 <= io_addr_in_dccm_d;
    end
  end
  always @(posedge io_lsu_c1_r_clk or posedge reset) begin
    if (reset) begin
      _T_151 <= 1'h0;
    end else begin
      _T_151 <= io_addr_in_dccm_m;
    end
  end
  always @(posedge io_lsu_c1_m_clk or posedge reset) begin
    if (reset) begin
      _T_152 <= 1'h0;
    end else begin
      _T_152 <= io_addr_in_pic_d;
    end
  end
  always @(posedge io_lsu_c1_r_clk or posedge reset) begin
    if (reset) begin
      _T_153 <= 1'h0;
    end else begin
      _T_153 <= io_addr_in_pic_m;
    end
  end
  always @(posedge io_lsu_c1_m_clk or posedge reset) begin
    if (reset) begin
      _T_154 <= 1'h0;
    end else begin
      _T_154 <= addrcheck_io_addr_external_d;
    end
  end
  always @(posedge io_lsu_c1_r_clk or posedge reset) begin
    if (reset) begin
      addr_external_r <= 1'h0;
    end else begin
      addr_external_r <= io_addr_external_m;
    end
  end
  always @(posedge io_lsu_c1_r_clk or posedge reset) begin
    if (reset) begin
      bus_read_data_r <= 32'h0;
    end else begin
      bus_read_data_r <= io_bus_read_data_m;
    end
  end
endmodule
module lsu_dccm_ctl(
  input         clock,
  input         reset,
  input         io_lsu_c2_m_clk,
  input         io_lsu_c2_r_clk,
  input         io_lsu_free_c2_clk,
  input         io_lsu_store_c1_r_clk,
  input         io_lsu_pkt_d_valid,
  input         io_lsu_pkt_d_bits_word,
  input         io_lsu_pkt_d_bits_dword,
  input         io_lsu_pkt_d_bits_load,
  input         io_lsu_pkt_d_bits_store,
  input         io_lsu_pkt_d_bits_dma,
  input         io_lsu_pkt_m_valid,
  input         io_lsu_pkt_m_bits_by,
  input         io_lsu_pkt_m_bits_half,
  input         io_lsu_pkt_m_bits_word,
  input         io_lsu_pkt_m_bits_load,
  input         io_lsu_pkt_m_bits_store,
  input         io_lsu_pkt_m_bits_dma,
  input         io_lsu_pkt_r_valid,
  input         io_lsu_pkt_r_bits_by,
  input         io_lsu_pkt_r_bits_half,
  input         io_lsu_pkt_r_bits_word,
  input         io_lsu_pkt_r_bits_load,
  input         io_lsu_pkt_r_bits_store,
  input         io_lsu_pkt_r_bits_dma,
  input         io_addr_in_dccm_d,
  input         io_addr_in_dccm_m,
  input         io_addr_in_dccm_r,
  input         io_addr_in_pic_d,
  input         io_addr_in_pic_m,
  input         io_addr_in_pic_r,
  input         io_lsu_raw_fwd_lo_r,
  input         io_lsu_raw_fwd_hi_r,
  input         io_lsu_commit_r,
  input  [31:0] io_lsu_addr_d,
  input  [15:0] io_lsu_addr_m,
  input  [31:0] io_lsu_addr_r,
  input  [15:0] io_end_addr_d,
  input  [15:0] io_end_addr_m,
  input  [15:0] io_end_addr_r,
  input         io_stbuf_reqvld_any,
  input  [15:0] io_stbuf_addr_any,
  input  [31:0] io_stbuf_data_any,
  input  [6:0]  io_stbuf_ecc_any,
  input  [31:0] io_stbuf_fwddata_hi_m,
  input  [31:0] io_stbuf_fwddata_lo_m,
  input  [3:0]  io_stbuf_fwdbyteen_lo_m,
  input  [3:0]  io_stbuf_fwdbyteen_hi_m,
  output [31:0] io_lsu_ld_data_corr_r,
  input         io_lsu_double_ecc_error_r,
  input         io_single_ecc_error_hi_r,
  input         io_single_ecc_error_lo_r,
  input  [31:0] io_sec_data_hi_r_ff,
  input  [31:0] io_sec_data_lo_r_ff,
  input  [6:0]  io_sec_data_ecc_hi_r_ff,
  input  [6:0]  io_sec_data_ecc_lo_r_ff,
  output [31:0] io_dccm_rdata_hi_m,
  output [31:0] io_dccm_rdata_lo_m,
  output [6:0]  io_dccm_data_ecc_hi_m,
  output [6:0]  io_dccm_data_ecc_lo_m,
  output [31:0] io_lsu_ld_data_m,
  input         io_lsu_double_ecc_error_m,
  input  [31:0] io_sec_data_hi_m,
  input  [31:0] io_sec_data_lo_m,
  input  [31:0] io_store_data_m,
  input         io_dma_dccm_wen,
  input         io_dma_pic_wen,
  input  [2:0]  io_dma_mem_tag_m,
  input  [31:0] io_dma_dccm_wdata_lo,
  input  [31:0] io_dma_dccm_wdata_hi,
  input  [6:0]  io_dma_dccm_wdata_ecc_hi,
  input  [6:0]  io_dma_dccm_wdata_ecc_lo,
  output [31:0] io_store_data_hi_r,
  output [31:0] io_store_data_lo_r,
  output [31:0] io_store_datafn_hi_r,
  output [31:0] io_store_datafn_lo_r,
  output [31:0] io_store_data_r,
  output        io_ld_single_ecc_error_r,
  output        io_ld_single_ecc_error_r_ff,
  output [31:0] io_picm_mask_data_m,
  output        io_lsu_stbuf_commit_any,
  output        io_lsu_dccm_rden_m,
  input  [31:0] io_dma_dccm_ctl_dma_mem_addr,
  input  [63:0] io_dma_dccm_ctl_dma_mem_wdata,
  output        io_dma_dccm_ctl_dccm_dma_rvalid,
  output        io_dma_dccm_ctl_dccm_dma_ecc_error,
  output [2:0]  io_dma_dccm_ctl_dccm_dma_rtag,
  output [63:0] io_dma_dccm_ctl_dccm_dma_rdata,
  output        io_dccm_wren,
  output        io_dccm_rden,
  output [15:0] io_dccm_wr_addr_lo,
  output [15:0] io_dccm_wr_addr_hi,
  output [15:0] io_dccm_rd_addr_lo,
  output [15:0] io_dccm_rd_addr_hi,
  output [38:0] io_dccm_wr_data_lo,
  output [38:0] io_dccm_wr_data_hi,
  input  [38:0] io_dccm_rd_data_lo,
  input  [38:0] io_dccm_rd_data_hi,
  output        io_lsu_pic_picm_wren,
  output        io_lsu_pic_picm_rden,
  output        io_lsu_pic_picm_mken,
  output [31:0] io_lsu_pic_picm_rdaddr,
  output [31:0] io_lsu_pic_picm_wraddr,
  output [31:0] io_lsu_pic_picm_wr_data,
  input  [31:0] io_lsu_pic_picm_rd_data,
  input         io_scan_mode
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
`endif // RANDOMIZE_REG_INIT
  wire  rvclkhdr_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_1_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_1_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_1_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_1_io_scan_mode; // @[lib.scala 368:23]
  wire [63:0] picm_rd_data_m = {io_lsu_pic_picm_rd_data,io_lsu_pic_picm_rd_data}; // @[Cat.scala 29:58]
  wire [63:0] dccm_rdata_corr_m = {io_sec_data_hi_m,io_sec_data_lo_m}; // @[Cat.scala 29:58]
  wire [63:0] dccm_rdata_m = {io_dccm_rdata_hi_m,io_dccm_rdata_lo_m}; // @[Cat.scala 29:58]
  wire  _T = io_lsu_pkt_m_valid & io_lsu_pkt_m_bits_load; // @[lsu_dccm_ctl.scala 137:63]
  reg [63:0] _T_2; // @[lsu_dccm_ctl.scala 147:65]
  wire [7:0] _T_3 = {io_stbuf_fwdbyteen_hi_m,io_stbuf_fwdbyteen_lo_m}; // @[Cat.scala 29:58]
  wire [63:0] _T_6 = {io_stbuf_fwddata_hi_m,io_stbuf_fwddata_lo_m}; // @[Cat.scala 29:58]
  wire [7:0] _T_11 = io_addr_in_pic_m ? picm_rd_data_m[7:0] : dccm_rdata_corr_m[7:0]; // @[lsu_dccm_ctl.scala 148:213]
  wire [7:0] _T_12 = _T_3[0] ? _T_6[7:0] : _T_11; // @[lsu_dccm_ctl.scala 148:78]
  wire [7:0] _T_16 = {{4'd0}, _T_12[7:4]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_18 = {_T_12[3:0], 4'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_20 = _T_18 & 8'hf0; // @[Bitwise.scala 103:75]
  wire [7:0] _T_21 = _T_16 | _T_20; // @[Bitwise.scala 103:39]
  wire [7:0] _GEN_0 = {{2'd0}, _T_21[7:2]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_26 = _GEN_0 & 8'h33; // @[Bitwise.scala 103:31]
  wire [7:0] _T_28 = {_T_21[5:0], 2'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_30 = _T_28 & 8'hcc; // @[Bitwise.scala 103:75]
  wire [7:0] _T_31 = _T_26 | _T_30; // @[Bitwise.scala 103:39]
  wire [7:0] _GEN_1 = {{1'd0}, _T_31[7:1]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_36 = _GEN_1 & 8'h55; // @[Bitwise.scala 103:31]
  wire [7:0] _T_38 = {_T_31[6:0], 1'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_40 = _T_38 & 8'haa; // @[Bitwise.scala 103:75]
  wire [7:0] _T_41 = _T_36 | _T_40; // @[Bitwise.scala 103:39]
  wire [7:0] _T_50 = io_addr_in_pic_m ? picm_rd_data_m[15:8] : dccm_rdata_corr_m[15:8]; // @[lsu_dccm_ctl.scala 148:213]
  wire [7:0] _T_51 = _T_3[1] ? _T_6[15:8] : _T_50; // @[lsu_dccm_ctl.scala 148:78]
  wire [7:0] _T_55 = {{4'd0}, _T_51[7:4]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_57 = {_T_51[3:0], 4'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_59 = _T_57 & 8'hf0; // @[Bitwise.scala 103:75]
  wire [7:0] _T_60 = _T_55 | _T_59; // @[Bitwise.scala 103:39]
  wire [7:0] _GEN_2 = {{2'd0}, _T_60[7:2]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_65 = _GEN_2 & 8'h33; // @[Bitwise.scala 103:31]
  wire [7:0] _T_67 = {_T_60[5:0], 2'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_69 = _T_67 & 8'hcc; // @[Bitwise.scala 103:75]
  wire [7:0] _T_70 = _T_65 | _T_69; // @[Bitwise.scala 103:39]
  wire [7:0] _GEN_3 = {{1'd0}, _T_70[7:1]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_75 = _GEN_3 & 8'h55; // @[Bitwise.scala 103:31]
  wire [7:0] _T_77 = {_T_70[6:0], 1'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_79 = _T_77 & 8'haa; // @[Bitwise.scala 103:75]
  wire [7:0] _T_80 = _T_75 | _T_79; // @[Bitwise.scala 103:39]
  wire [7:0] _T_89 = io_addr_in_pic_m ? picm_rd_data_m[23:16] : dccm_rdata_corr_m[23:16]; // @[lsu_dccm_ctl.scala 148:213]
  wire [7:0] _T_90 = _T_3[2] ? _T_6[23:16] : _T_89; // @[lsu_dccm_ctl.scala 148:78]
  wire [7:0] _T_94 = {{4'd0}, _T_90[7:4]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_96 = {_T_90[3:0], 4'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_98 = _T_96 & 8'hf0; // @[Bitwise.scala 103:75]
  wire [7:0] _T_99 = _T_94 | _T_98; // @[Bitwise.scala 103:39]
  wire [7:0] _GEN_4 = {{2'd0}, _T_99[7:2]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_104 = _GEN_4 & 8'h33; // @[Bitwise.scala 103:31]
  wire [7:0] _T_106 = {_T_99[5:0], 2'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_108 = _T_106 & 8'hcc; // @[Bitwise.scala 103:75]
  wire [7:0] _T_109 = _T_104 | _T_108; // @[Bitwise.scala 103:39]
  wire [7:0] _GEN_5 = {{1'd0}, _T_109[7:1]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_114 = _GEN_5 & 8'h55; // @[Bitwise.scala 103:31]
  wire [7:0] _T_116 = {_T_109[6:0], 1'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_118 = _T_116 & 8'haa; // @[Bitwise.scala 103:75]
  wire [7:0] _T_119 = _T_114 | _T_118; // @[Bitwise.scala 103:39]
  wire [7:0] _T_128 = io_addr_in_pic_m ? picm_rd_data_m[31:24] : dccm_rdata_corr_m[31:24]; // @[lsu_dccm_ctl.scala 148:213]
  wire [7:0] _T_129 = _T_3[3] ? _T_6[31:24] : _T_128; // @[lsu_dccm_ctl.scala 148:78]
  wire [7:0] _T_133 = {{4'd0}, _T_129[7:4]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_135 = {_T_129[3:0], 4'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_137 = _T_135 & 8'hf0; // @[Bitwise.scala 103:75]
  wire [7:0] _T_138 = _T_133 | _T_137; // @[Bitwise.scala 103:39]
  wire [7:0] _GEN_6 = {{2'd0}, _T_138[7:2]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_143 = _GEN_6 & 8'h33; // @[Bitwise.scala 103:31]
  wire [7:0] _T_145 = {_T_138[5:0], 2'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_147 = _T_145 & 8'hcc; // @[Bitwise.scala 103:75]
  wire [7:0] _T_148 = _T_143 | _T_147; // @[Bitwise.scala 103:39]
  wire [7:0] _GEN_7 = {{1'd0}, _T_148[7:1]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_153 = _GEN_7 & 8'h55; // @[Bitwise.scala 103:31]
  wire [7:0] _T_155 = {_T_148[6:0], 1'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_157 = _T_155 & 8'haa; // @[Bitwise.scala 103:75]
  wire [7:0] _T_158 = _T_153 | _T_157; // @[Bitwise.scala 103:39]
  wire [7:0] _T_167 = io_addr_in_pic_m ? picm_rd_data_m[39:32] : dccm_rdata_corr_m[39:32]; // @[lsu_dccm_ctl.scala 148:213]
  wire [7:0] _T_168 = _T_3[4] ? _T_6[39:32] : _T_167; // @[lsu_dccm_ctl.scala 148:78]
  wire [7:0] _T_172 = {{4'd0}, _T_168[7:4]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_174 = {_T_168[3:0], 4'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_176 = _T_174 & 8'hf0; // @[Bitwise.scala 103:75]
  wire [7:0] _T_177 = _T_172 | _T_176; // @[Bitwise.scala 103:39]
  wire [7:0] _GEN_8 = {{2'd0}, _T_177[7:2]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_182 = _GEN_8 & 8'h33; // @[Bitwise.scala 103:31]
  wire [7:0] _T_184 = {_T_177[5:0], 2'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_186 = _T_184 & 8'hcc; // @[Bitwise.scala 103:75]
  wire [7:0] _T_187 = _T_182 | _T_186; // @[Bitwise.scala 103:39]
  wire [7:0] _GEN_9 = {{1'd0}, _T_187[7:1]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_192 = _GEN_9 & 8'h55; // @[Bitwise.scala 103:31]
  wire [7:0] _T_194 = {_T_187[6:0], 1'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_196 = _T_194 & 8'haa; // @[Bitwise.scala 103:75]
  wire [7:0] _T_197 = _T_192 | _T_196; // @[Bitwise.scala 103:39]
  wire [7:0] _T_206 = io_addr_in_pic_m ? picm_rd_data_m[47:40] : dccm_rdata_corr_m[47:40]; // @[lsu_dccm_ctl.scala 148:213]
  wire [7:0] _T_207 = _T_3[5] ? _T_6[47:40] : _T_206; // @[lsu_dccm_ctl.scala 148:78]
  wire [7:0] _T_211 = {{4'd0}, _T_207[7:4]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_213 = {_T_207[3:0], 4'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_215 = _T_213 & 8'hf0; // @[Bitwise.scala 103:75]
  wire [7:0] _T_216 = _T_211 | _T_215; // @[Bitwise.scala 103:39]
  wire [7:0] _GEN_10 = {{2'd0}, _T_216[7:2]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_221 = _GEN_10 & 8'h33; // @[Bitwise.scala 103:31]
  wire [7:0] _T_223 = {_T_216[5:0], 2'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_225 = _T_223 & 8'hcc; // @[Bitwise.scala 103:75]
  wire [7:0] _T_226 = _T_221 | _T_225; // @[Bitwise.scala 103:39]
  wire [7:0] _GEN_11 = {{1'd0}, _T_226[7:1]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_231 = _GEN_11 & 8'h55; // @[Bitwise.scala 103:31]
  wire [7:0] _T_233 = {_T_226[6:0], 1'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_235 = _T_233 & 8'haa; // @[Bitwise.scala 103:75]
  wire [7:0] _T_236 = _T_231 | _T_235; // @[Bitwise.scala 103:39]
  wire [7:0] _T_245 = io_addr_in_pic_m ? picm_rd_data_m[55:48] : dccm_rdata_corr_m[55:48]; // @[lsu_dccm_ctl.scala 148:213]
  wire [7:0] _T_246 = _T_3[6] ? _T_6[55:48] : _T_245; // @[lsu_dccm_ctl.scala 148:78]
  wire [7:0] _T_250 = {{4'd0}, _T_246[7:4]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_252 = {_T_246[3:0], 4'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_254 = _T_252 & 8'hf0; // @[Bitwise.scala 103:75]
  wire [7:0] _T_255 = _T_250 | _T_254; // @[Bitwise.scala 103:39]
  wire [7:0] _GEN_12 = {{2'd0}, _T_255[7:2]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_260 = _GEN_12 & 8'h33; // @[Bitwise.scala 103:31]
  wire [7:0] _T_262 = {_T_255[5:0], 2'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_264 = _T_262 & 8'hcc; // @[Bitwise.scala 103:75]
  wire [7:0] _T_265 = _T_260 | _T_264; // @[Bitwise.scala 103:39]
  wire [7:0] _GEN_13 = {{1'd0}, _T_265[7:1]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_270 = _GEN_13 & 8'h55; // @[Bitwise.scala 103:31]
  wire [7:0] _T_272 = {_T_265[6:0], 1'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_274 = _T_272 & 8'haa; // @[Bitwise.scala 103:75]
  wire [7:0] _T_275 = _T_270 | _T_274; // @[Bitwise.scala 103:39]
  wire [7:0] _T_284 = io_addr_in_pic_m ? picm_rd_data_m[63:56] : dccm_rdata_corr_m[63:56]; // @[lsu_dccm_ctl.scala 148:213]
  wire [7:0] _T_285 = _T_3[7] ? _T_6[63:56] : _T_284; // @[lsu_dccm_ctl.scala 148:78]
  wire [7:0] _T_289 = {{4'd0}, _T_285[7:4]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_291 = {_T_285[3:0], 4'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_293 = _T_291 & 8'hf0; // @[Bitwise.scala 103:75]
  wire [7:0] _T_294 = _T_289 | _T_293; // @[Bitwise.scala 103:39]
  wire [7:0] _GEN_14 = {{2'd0}, _T_294[7:2]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_299 = _GEN_14 & 8'h33; // @[Bitwise.scala 103:31]
  wire [7:0] _T_301 = {_T_294[5:0], 2'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_303 = _T_301 & 8'hcc; // @[Bitwise.scala 103:75]
  wire [7:0] _T_304 = _T_299 | _T_303; // @[Bitwise.scala 103:39]
  wire [7:0] _GEN_15 = {{1'd0}, _T_304[7:1]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_309 = _GEN_15 & 8'h55; // @[Bitwise.scala 103:31]
  wire [7:0] _T_311 = {_T_304[6:0], 1'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_313 = _T_311 & 8'haa; // @[Bitwise.scala 103:75]
  wire [7:0] _T_314 = _T_309 | _T_313; // @[Bitwise.scala 103:39]
  wire [63:0] _T_322 = {_T_41,_T_80,_T_119,_T_158,_T_197,_T_236,_T_275,_T_314}; // @[Cat.scala 29:58]
  wire [63:0] _T_326 = {{32'd0}, _T_322[63:32]}; // @[Bitwise.scala 103:31]
  wire [63:0] _T_328 = {_T_322[31:0], 32'h0}; // @[Bitwise.scala 103:65]
  wire [63:0] _T_330 = _T_328 & 64'hffffffff00000000; // @[Bitwise.scala 103:75]
  wire [63:0] _T_331 = _T_326 | _T_330; // @[Bitwise.scala 103:39]
  wire [63:0] _GEN_16 = {{16'd0}, _T_331[63:16]}; // @[Bitwise.scala 103:31]
  wire [63:0] _T_336 = _GEN_16 & 64'hffff0000ffff; // @[Bitwise.scala 103:31]
  wire [63:0] _T_338 = {_T_331[47:0], 16'h0}; // @[Bitwise.scala 103:65]
  wire [63:0] _T_340 = _T_338 & 64'hffff0000ffff0000; // @[Bitwise.scala 103:75]
  wire [63:0] _T_341 = _T_336 | _T_340; // @[Bitwise.scala 103:39]
  wire [63:0] _GEN_17 = {{8'd0}, _T_341[63:8]}; // @[Bitwise.scala 103:31]
  wire [63:0] _T_346 = _GEN_17 & 64'hff00ff00ff00ff; // @[Bitwise.scala 103:31]
  wire [63:0] _T_348 = {_T_341[55:0], 8'h0}; // @[Bitwise.scala 103:65]
  wire [63:0] _T_350 = _T_348 & 64'hff00ff00ff00ff00; // @[Bitwise.scala 103:75]
  wire [63:0] _T_351 = _T_346 | _T_350; // @[Bitwise.scala 103:39]
  wire [63:0] _GEN_18 = {{4'd0}, _T_351[63:4]}; // @[Bitwise.scala 103:31]
  wire [63:0] _T_356 = _GEN_18 & 64'hf0f0f0f0f0f0f0f; // @[Bitwise.scala 103:31]
  wire [63:0] _T_358 = {_T_351[59:0], 4'h0}; // @[Bitwise.scala 103:65]
  wire [63:0] _T_360 = _T_358 & 64'hf0f0f0f0f0f0f0f0; // @[Bitwise.scala 103:75]
  wire [63:0] _T_361 = _T_356 | _T_360; // @[Bitwise.scala 103:39]
  wire [63:0] _GEN_19 = {{2'd0}, _T_361[63:2]}; // @[Bitwise.scala 103:31]
  wire [63:0] _T_366 = _GEN_19 & 64'h3333333333333333; // @[Bitwise.scala 103:31]
  wire [63:0] _T_368 = {_T_361[61:0], 2'h0}; // @[Bitwise.scala 103:65]
  wire [63:0] _T_370 = _T_368 & 64'hcccccccccccccccc; // @[Bitwise.scala 103:75]
  wire [63:0] _T_371 = _T_366 | _T_370; // @[Bitwise.scala 103:39]
  wire [63:0] _GEN_20 = {{1'd0}, _T_371[63:1]}; // @[Bitwise.scala 103:31]
  wire [63:0] _T_376 = _GEN_20 & 64'h5555555555555555; // @[Bitwise.scala 103:31]
  wire [63:0] _T_378 = {_T_371[62:0], 1'h0}; // @[Bitwise.scala 103:65]
  wire [63:0] _T_380 = _T_378 & 64'haaaaaaaaaaaaaaaa; // @[Bitwise.scala 103:75]
  wire [63:0] lsu_rdata_corr_m = _T_376 | _T_380; // @[Bitwise.scala 103:39]
  wire [7:0] _T_390 = io_addr_in_pic_m ? picm_rd_data_m[7:0] : dccm_rdata_m[7:0]; // @[lsu_dccm_ctl.scala 149:213]
  wire [7:0] _T_391 = _T_3[0] ? _T_6[7:0] : _T_390; // @[lsu_dccm_ctl.scala 149:78]
  wire [7:0] _T_395 = {{4'd0}, _T_391[7:4]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_397 = {_T_391[3:0], 4'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_399 = _T_397 & 8'hf0; // @[Bitwise.scala 103:75]
  wire [7:0] _T_400 = _T_395 | _T_399; // @[Bitwise.scala 103:39]
  wire [7:0] _GEN_21 = {{2'd0}, _T_400[7:2]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_405 = _GEN_21 & 8'h33; // @[Bitwise.scala 103:31]
  wire [7:0] _T_407 = {_T_400[5:0], 2'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_409 = _T_407 & 8'hcc; // @[Bitwise.scala 103:75]
  wire [7:0] _T_410 = _T_405 | _T_409; // @[Bitwise.scala 103:39]
  wire [7:0] _GEN_22 = {{1'd0}, _T_410[7:1]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_415 = _GEN_22 & 8'h55; // @[Bitwise.scala 103:31]
  wire [7:0] _T_417 = {_T_410[6:0], 1'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_419 = _T_417 & 8'haa; // @[Bitwise.scala 103:75]
  wire [7:0] _T_420 = _T_415 | _T_419; // @[Bitwise.scala 103:39]
  wire [7:0] _T_429 = io_addr_in_pic_m ? picm_rd_data_m[15:8] : dccm_rdata_m[15:8]; // @[lsu_dccm_ctl.scala 149:213]
  wire [7:0] _T_430 = _T_3[1] ? _T_6[15:8] : _T_429; // @[lsu_dccm_ctl.scala 149:78]
  wire [7:0] _T_434 = {{4'd0}, _T_430[7:4]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_436 = {_T_430[3:0], 4'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_438 = _T_436 & 8'hf0; // @[Bitwise.scala 103:75]
  wire [7:0] _T_439 = _T_434 | _T_438; // @[Bitwise.scala 103:39]
  wire [7:0] _GEN_23 = {{2'd0}, _T_439[7:2]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_444 = _GEN_23 & 8'h33; // @[Bitwise.scala 103:31]
  wire [7:0] _T_446 = {_T_439[5:0], 2'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_448 = _T_446 & 8'hcc; // @[Bitwise.scala 103:75]
  wire [7:0] _T_449 = _T_444 | _T_448; // @[Bitwise.scala 103:39]
  wire [7:0] _GEN_24 = {{1'd0}, _T_449[7:1]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_454 = _GEN_24 & 8'h55; // @[Bitwise.scala 103:31]
  wire [7:0] _T_456 = {_T_449[6:0], 1'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_458 = _T_456 & 8'haa; // @[Bitwise.scala 103:75]
  wire [7:0] _T_459 = _T_454 | _T_458; // @[Bitwise.scala 103:39]
  wire [7:0] _T_468 = io_addr_in_pic_m ? picm_rd_data_m[23:16] : dccm_rdata_m[23:16]; // @[lsu_dccm_ctl.scala 149:213]
  wire [7:0] _T_469 = _T_3[2] ? _T_6[23:16] : _T_468; // @[lsu_dccm_ctl.scala 149:78]
  wire [7:0] _T_473 = {{4'd0}, _T_469[7:4]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_475 = {_T_469[3:0], 4'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_477 = _T_475 & 8'hf0; // @[Bitwise.scala 103:75]
  wire [7:0] _T_478 = _T_473 | _T_477; // @[Bitwise.scala 103:39]
  wire [7:0] _GEN_25 = {{2'd0}, _T_478[7:2]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_483 = _GEN_25 & 8'h33; // @[Bitwise.scala 103:31]
  wire [7:0] _T_485 = {_T_478[5:0], 2'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_487 = _T_485 & 8'hcc; // @[Bitwise.scala 103:75]
  wire [7:0] _T_488 = _T_483 | _T_487; // @[Bitwise.scala 103:39]
  wire [7:0] _GEN_26 = {{1'd0}, _T_488[7:1]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_493 = _GEN_26 & 8'h55; // @[Bitwise.scala 103:31]
  wire [7:0] _T_495 = {_T_488[6:0], 1'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_497 = _T_495 & 8'haa; // @[Bitwise.scala 103:75]
  wire [7:0] _T_498 = _T_493 | _T_497; // @[Bitwise.scala 103:39]
  wire [7:0] _T_507 = io_addr_in_pic_m ? picm_rd_data_m[31:24] : dccm_rdata_m[31:24]; // @[lsu_dccm_ctl.scala 149:213]
  wire [7:0] _T_508 = _T_3[3] ? _T_6[31:24] : _T_507; // @[lsu_dccm_ctl.scala 149:78]
  wire [7:0] _T_512 = {{4'd0}, _T_508[7:4]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_514 = {_T_508[3:0], 4'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_516 = _T_514 & 8'hf0; // @[Bitwise.scala 103:75]
  wire [7:0] _T_517 = _T_512 | _T_516; // @[Bitwise.scala 103:39]
  wire [7:0] _GEN_27 = {{2'd0}, _T_517[7:2]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_522 = _GEN_27 & 8'h33; // @[Bitwise.scala 103:31]
  wire [7:0] _T_524 = {_T_517[5:0], 2'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_526 = _T_524 & 8'hcc; // @[Bitwise.scala 103:75]
  wire [7:0] _T_527 = _T_522 | _T_526; // @[Bitwise.scala 103:39]
  wire [7:0] _GEN_28 = {{1'd0}, _T_527[7:1]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_532 = _GEN_28 & 8'h55; // @[Bitwise.scala 103:31]
  wire [7:0] _T_534 = {_T_527[6:0], 1'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_536 = _T_534 & 8'haa; // @[Bitwise.scala 103:75]
  wire [7:0] _T_537 = _T_532 | _T_536; // @[Bitwise.scala 103:39]
  wire [7:0] _T_546 = io_addr_in_pic_m ? picm_rd_data_m[39:32] : dccm_rdata_m[39:32]; // @[lsu_dccm_ctl.scala 149:213]
  wire [7:0] _T_547 = _T_3[4] ? _T_6[39:32] : _T_546; // @[lsu_dccm_ctl.scala 149:78]
  wire [7:0] _T_551 = {{4'd0}, _T_547[7:4]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_553 = {_T_547[3:0], 4'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_555 = _T_553 & 8'hf0; // @[Bitwise.scala 103:75]
  wire [7:0] _T_556 = _T_551 | _T_555; // @[Bitwise.scala 103:39]
  wire [7:0] _GEN_29 = {{2'd0}, _T_556[7:2]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_561 = _GEN_29 & 8'h33; // @[Bitwise.scala 103:31]
  wire [7:0] _T_563 = {_T_556[5:0], 2'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_565 = _T_563 & 8'hcc; // @[Bitwise.scala 103:75]
  wire [7:0] _T_566 = _T_561 | _T_565; // @[Bitwise.scala 103:39]
  wire [7:0] _GEN_30 = {{1'd0}, _T_566[7:1]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_571 = _GEN_30 & 8'h55; // @[Bitwise.scala 103:31]
  wire [7:0] _T_573 = {_T_566[6:0], 1'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_575 = _T_573 & 8'haa; // @[Bitwise.scala 103:75]
  wire [7:0] _T_576 = _T_571 | _T_575; // @[Bitwise.scala 103:39]
  wire [7:0] _T_585 = io_addr_in_pic_m ? picm_rd_data_m[47:40] : dccm_rdata_m[47:40]; // @[lsu_dccm_ctl.scala 149:213]
  wire [7:0] _T_586 = _T_3[5] ? _T_6[47:40] : _T_585; // @[lsu_dccm_ctl.scala 149:78]
  wire [7:0] _T_590 = {{4'd0}, _T_586[7:4]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_592 = {_T_586[3:0], 4'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_594 = _T_592 & 8'hf0; // @[Bitwise.scala 103:75]
  wire [7:0] _T_595 = _T_590 | _T_594; // @[Bitwise.scala 103:39]
  wire [7:0] _GEN_31 = {{2'd0}, _T_595[7:2]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_600 = _GEN_31 & 8'h33; // @[Bitwise.scala 103:31]
  wire [7:0] _T_602 = {_T_595[5:0], 2'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_604 = _T_602 & 8'hcc; // @[Bitwise.scala 103:75]
  wire [7:0] _T_605 = _T_600 | _T_604; // @[Bitwise.scala 103:39]
  wire [7:0] _GEN_32 = {{1'd0}, _T_605[7:1]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_610 = _GEN_32 & 8'h55; // @[Bitwise.scala 103:31]
  wire [7:0] _T_612 = {_T_605[6:0], 1'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_614 = _T_612 & 8'haa; // @[Bitwise.scala 103:75]
  wire [7:0] _T_615 = _T_610 | _T_614; // @[Bitwise.scala 103:39]
  wire [7:0] _T_624 = io_addr_in_pic_m ? picm_rd_data_m[55:48] : dccm_rdata_m[55:48]; // @[lsu_dccm_ctl.scala 149:213]
  wire [7:0] _T_625 = _T_3[6] ? _T_6[55:48] : _T_624; // @[lsu_dccm_ctl.scala 149:78]
  wire [7:0] _T_629 = {{4'd0}, _T_625[7:4]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_631 = {_T_625[3:0], 4'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_633 = _T_631 & 8'hf0; // @[Bitwise.scala 103:75]
  wire [7:0] _T_634 = _T_629 | _T_633; // @[Bitwise.scala 103:39]
  wire [7:0] _GEN_33 = {{2'd0}, _T_634[7:2]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_639 = _GEN_33 & 8'h33; // @[Bitwise.scala 103:31]
  wire [7:0] _T_641 = {_T_634[5:0], 2'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_643 = _T_641 & 8'hcc; // @[Bitwise.scala 103:75]
  wire [7:0] _T_644 = _T_639 | _T_643; // @[Bitwise.scala 103:39]
  wire [7:0] _GEN_34 = {{1'd0}, _T_644[7:1]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_649 = _GEN_34 & 8'h55; // @[Bitwise.scala 103:31]
  wire [7:0] _T_651 = {_T_644[6:0], 1'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_653 = _T_651 & 8'haa; // @[Bitwise.scala 103:75]
  wire [7:0] _T_654 = _T_649 | _T_653; // @[Bitwise.scala 103:39]
  wire [7:0] _T_663 = io_addr_in_pic_m ? picm_rd_data_m[63:56] : dccm_rdata_m[63:56]; // @[lsu_dccm_ctl.scala 149:213]
  wire [7:0] _T_664 = _T_3[7] ? _T_6[63:56] : _T_663; // @[lsu_dccm_ctl.scala 149:78]
  wire [7:0] _T_668 = {{4'd0}, _T_664[7:4]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_670 = {_T_664[3:0], 4'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_672 = _T_670 & 8'hf0; // @[Bitwise.scala 103:75]
  wire [7:0] _T_673 = _T_668 | _T_672; // @[Bitwise.scala 103:39]
  wire [7:0] _GEN_35 = {{2'd0}, _T_673[7:2]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_678 = _GEN_35 & 8'h33; // @[Bitwise.scala 103:31]
  wire [7:0] _T_680 = {_T_673[5:0], 2'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_682 = _T_680 & 8'hcc; // @[Bitwise.scala 103:75]
  wire [7:0] _T_683 = _T_678 | _T_682; // @[Bitwise.scala 103:39]
  wire [7:0] _GEN_36 = {{1'd0}, _T_683[7:1]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_688 = _GEN_36 & 8'h55; // @[Bitwise.scala 103:31]
  wire [7:0] _T_690 = {_T_683[6:0], 1'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_692 = _T_690 & 8'haa; // @[Bitwise.scala 103:75]
  wire [7:0] _T_693 = _T_688 | _T_692; // @[Bitwise.scala 103:39]
  wire [63:0] _T_701 = {_T_420,_T_459,_T_498,_T_537,_T_576,_T_615,_T_654,_T_693}; // @[Cat.scala 29:58]
  wire [63:0] _T_705 = {{32'd0}, _T_701[63:32]}; // @[Bitwise.scala 103:31]
  wire [63:0] _T_707 = {_T_701[31:0], 32'h0}; // @[Bitwise.scala 103:65]
  wire [63:0] _T_709 = _T_707 & 64'hffffffff00000000; // @[Bitwise.scala 103:75]
  wire [63:0] _T_710 = _T_705 | _T_709; // @[Bitwise.scala 103:39]
  wire [63:0] _GEN_37 = {{16'd0}, _T_710[63:16]}; // @[Bitwise.scala 103:31]
  wire [63:0] _T_715 = _GEN_37 & 64'hffff0000ffff; // @[Bitwise.scala 103:31]
  wire [63:0] _T_717 = {_T_710[47:0], 16'h0}; // @[Bitwise.scala 103:65]
  wire [63:0] _T_719 = _T_717 & 64'hffff0000ffff0000; // @[Bitwise.scala 103:75]
  wire [63:0] _T_720 = _T_715 | _T_719; // @[Bitwise.scala 103:39]
  wire [63:0] _GEN_38 = {{8'd0}, _T_720[63:8]}; // @[Bitwise.scala 103:31]
  wire [63:0] _T_725 = _GEN_38 & 64'hff00ff00ff00ff; // @[Bitwise.scala 103:31]
  wire [63:0] _T_727 = {_T_720[55:0], 8'h0}; // @[Bitwise.scala 103:65]
  wire [63:0] _T_729 = _T_727 & 64'hff00ff00ff00ff00; // @[Bitwise.scala 103:75]
  wire [63:0] _T_730 = _T_725 | _T_729; // @[Bitwise.scala 103:39]
  wire [63:0] _GEN_39 = {{4'd0}, _T_730[63:4]}; // @[Bitwise.scala 103:31]
  wire [63:0] _T_735 = _GEN_39 & 64'hf0f0f0f0f0f0f0f; // @[Bitwise.scala 103:31]
  wire [63:0] _T_737 = {_T_730[59:0], 4'h0}; // @[Bitwise.scala 103:65]
  wire [63:0] _T_739 = _T_737 & 64'hf0f0f0f0f0f0f0f0; // @[Bitwise.scala 103:75]
  wire [63:0] _T_740 = _T_735 | _T_739; // @[Bitwise.scala 103:39]
  wire [63:0] _GEN_40 = {{2'd0}, _T_740[63:2]}; // @[Bitwise.scala 103:31]
  wire [63:0] _T_745 = _GEN_40 & 64'h3333333333333333; // @[Bitwise.scala 103:31]
  wire [63:0] _T_747 = {_T_740[61:0], 2'h0}; // @[Bitwise.scala 103:65]
  wire [63:0] _T_749 = _T_747 & 64'hcccccccccccccccc; // @[Bitwise.scala 103:75]
  wire [63:0] _T_750 = _T_745 | _T_749; // @[Bitwise.scala 103:39]
  wire [63:0] _GEN_41 = {{1'd0}, _T_750[63:1]}; // @[Bitwise.scala 103:31]
  wire [63:0] _T_755 = _GEN_41 & 64'h5555555555555555; // @[Bitwise.scala 103:31]
  wire [63:0] _T_757 = {_T_750[62:0], 1'h0}; // @[Bitwise.scala 103:65]
  wire [63:0] _T_759 = _T_757 & 64'haaaaaaaaaaaaaaaa; // @[Bitwise.scala 103:75]
  wire [63:0] lsu_rdata_m = _T_755 | _T_759; // @[Bitwise.scala 103:39]
  wire [3:0] _GEN_42 = {{2'd0}, io_lsu_addr_m[1:0]}; // @[lsu_dccm_ctl.scala 150:49]
  wire [5:0] _T_762 = 4'h8 * _GEN_42; // @[lsu_dccm_ctl.scala 150:49]
  wire [63:0] _T_763 = lsu_rdata_m >> _T_762; // @[lsu_dccm_ctl.scala 150:43]
  wire  _T_769 = io_lsu_addr_d[15:2] == io_lsu_addr_r[15:2]; // @[lsu_dccm_ctl.scala 155:60]
  wire  _T_772 = io_end_addr_d[15:2] == io_lsu_addr_r[15:2]; // @[lsu_dccm_ctl.scala 155:133]
  wire  _T_773 = _T_769 | _T_772; // @[lsu_dccm_ctl.scala 155:101]
  wire  _T_774 = _T_773 & io_lsu_pkt_d_valid; // @[lsu_dccm_ctl.scala 155:175]
  wire  _T_775 = _T_774 & io_lsu_pkt_d_bits_store; // @[lsu_dccm_ctl.scala 155:196]
  wire  _T_776 = _T_775 & io_lsu_pkt_d_bits_dma; // @[lsu_dccm_ctl.scala 155:222]
  wire  _T_777 = _T_776 & io_addr_in_dccm_d; // @[lsu_dccm_ctl.scala 155:246]
  wire  _T_780 = io_lsu_addr_m[15:2] == io_lsu_addr_r[15:2]; // @[lsu_dccm_ctl.scala 156:37]
  wire  _T_783 = io_end_addr_m[15:2] == io_lsu_addr_r[15:2]; // @[lsu_dccm_ctl.scala 156:110]
  wire  _T_784 = _T_780 | _T_783; // @[lsu_dccm_ctl.scala 156:78]
  wire  _T_785 = _T_784 & io_lsu_pkt_m_valid; // @[lsu_dccm_ctl.scala 156:152]
  wire  _T_786 = _T_785 & io_lsu_pkt_m_bits_store; // @[lsu_dccm_ctl.scala 156:173]
  wire  _T_787 = _T_786 & io_lsu_pkt_m_bits_dma; // @[lsu_dccm_ctl.scala 156:199]
  wire  _T_788 = _T_787 & io_addr_in_dccm_m; // @[lsu_dccm_ctl.scala 156:223]
  wire  kill_ecc_corr_lo_r = _T_777 | _T_788; // @[lsu_dccm_ctl.scala 155:267]
  wire  _T_791 = io_lsu_addr_d[15:2] == io_end_addr_r[15:2]; // @[lsu_dccm_ctl.scala 158:60]
  wire  _T_794 = io_end_addr_d[15:2] == io_end_addr_r[15:2]; // @[lsu_dccm_ctl.scala 158:133]
  wire  _T_795 = _T_791 | _T_794; // @[lsu_dccm_ctl.scala 158:101]
  wire  _T_796 = _T_795 & io_lsu_pkt_d_valid; // @[lsu_dccm_ctl.scala 158:175]
  wire  _T_797 = _T_796 & io_lsu_pkt_d_bits_store; // @[lsu_dccm_ctl.scala 158:196]
  wire  _T_798 = _T_797 & io_lsu_pkt_d_bits_dma; // @[lsu_dccm_ctl.scala 158:222]
  wire  _T_799 = _T_798 & io_addr_in_dccm_d; // @[lsu_dccm_ctl.scala 158:246]
  wire  _T_802 = io_lsu_addr_m[15:2] == io_end_addr_r[15:2]; // @[lsu_dccm_ctl.scala 159:37]
  wire  _T_805 = io_end_addr_m[15:2] == io_end_addr_r[15:2]; // @[lsu_dccm_ctl.scala 159:110]
  wire  _T_806 = _T_802 | _T_805; // @[lsu_dccm_ctl.scala 159:78]
  wire  _T_807 = _T_806 & io_lsu_pkt_m_valid; // @[lsu_dccm_ctl.scala 159:152]
  wire  _T_808 = _T_807 & io_lsu_pkt_m_bits_store; // @[lsu_dccm_ctl.scala 159:173]
  wire  _T_809 = _T_808 & io_lsu_pkt_m_bits_dma; // @[lsu_dccm_ctl.scala 159:199]
  wire  _T_810 = _T_809 & io_addr_in_dccm_m; // @[lsu_dccm_ctl.scala 159:223]
  wire  kill_ecc_corr_hi_r = _T_799 | _T_810; // @[lsu_dccm_ctl.scala 158:267]
  wire  _T_811 = io_lsu_pkt_r_bits_load & io_single_ecc_error_lo_r; // @[lsu_dccm_ctl.scala 161:60]
  wire  _T_812 = ~io_lsu_raw_fwd_lo_r; // @[lsu_dccm_ctl.scala 161:89]
  wire  ld_single_ecc_error_lo_r = _T_811 & _T_812; // @[lsu_dccm_ctl.scala 161:87]
  wire  _T_813 = io_lsu_pkt_r_bits_load & io_single_ecc_error_hi_r; // @[lsu_dccm_ctl.scala 162:60]
  wire  _T_814 = ~io_lsu_raw_fwd_hi_r; // @[lsu_dccm_ctl.scala 162:89]
  wire  ld_single_ecc_error_hi_r = _T_813 & _T_814; // @[lsu_dccm_ctl.scala 162:87]
  wire  _T_815 = ld_single_ecc_error_lo_r | ld_single_ecc_error_hi_r; // @[lsu_dccm_ctl.scala 163:63]
  wire  _T_816 = ~io_lsu_double_ecc_error_r; // @[lsu_dccm_ctl.scala 163:93]
  wire  _T_818 = io_lsu_commit_r | io_lsu_pkt_r_bits_dma; // @[lsu_dccm_ctl.scala 164:81]
  wire  _T_819 = ld_single_ecc_error_lo_r & _T_818; // @[lsu_dccm_ctl.scala 164:62]
  wire  _T_820 = ~kill_ecc_corr_lo_r; // @[lsu_dccm_ctl.scala 164:108]
  wire  _T_822 = ld_single_ecc_error_hi_r & _T_818; // @[lsu_dccm_ctl.scala 165:62]
  wire  _T_823 = ~kill_ecc_corr_hi_r; // @[lsu_dccm_ctl.scala 165:108]
  reg  lsu_double_ecc_error_r_ff; // @[lsu_dccm_ctl.scala 167:74]
  reg  ld_single_ecc_error_hi_r_ff; // @[lsu_dccm_ctl.scala 168:74]
  reg  ld_single_ecc_error_lo_r_ff; // @[lsu_dccm_ctl.scala 169:74]
  reg [15:0] ld_sec_addr_hi_r_ff; // @[lib.scala 374:16]
  reg [15:0] ld_sec_addr_lo_r_ff; // @[lib.scala 374:16]
  wire  _T_830 = io_lsu_pkt_d_bits_word | io_lsu_pkt_d_bits_dword; // @[lsu_dccm_ctl.scala 173:125]
  wire  _T_831 = ~_T_830; // @[lsu_dccm_ctl.scala 173:100]
  wire  _T_833 = io_lsu_addr_d[1:0] != 2'h0; // @[lsu_dccm_ctl.scala 173:174]
  wire  _T_834 = _T_831 | _T_833; // @[lsu_dccm_ctl.scala 173:152]
  wire  _T_835 = io_lsu_pkt_d_bits_store & _T_834; // @[lsu_dccm_ctl.scala 173:97]
  wire  _T_836 = io_lsu_pkt_d_bits_load | _T_835; // @[lsu_dccm_ctl.scala 173:70]
  wire  _T_837 = io_lsu_pkt_d_valid & _T_836; // @[lsu_dccm_ctl.scala 173:44]
  wire  lsu_dccm_rden_d = _T_837 & io_addr_in_dccm_d; // @[lsu_dccm_ctl.scala 173:191]
  wire  _T_838 = ld_single_ecc_error_lo_r_ff | ld_single_ecc_error_hi_r_ff; // @[lsu_dccm_ctl.scala 176:63]
  wire  _T_839 = ~lsu_double_ecc_error_r_ff; // @[lsu_dccm_ctl.scala 176:96]
  wire  _T_841 = lsu_dccm_rden_d | io_dma_dccm_wen; // @[lsu_dccm_ctl.scala 177:75]
  wire  _T_842 = _T_841 | io_ld_single_ecc_error_r_ff; // @[lsu_dccm_ctl.scala 177:93]
  wire  _T_843 = ~_T_842; // @[lsu_dccm_ctl.scala 177:57]
  wire  _T_846 = io_stbuf_addr_any[3:2] == io_lsu_addr_d[3:2]; // @[lsu_dccm_ctl.scala 178:95]
  wire  _T_849 = io_stbuf_addr_any[3:2] == io_end_addr_d[3:2]; // @[lsu_dccm_ctl.scala 179:76]
  wire  _T_850 = _T_846 | _T_849; // @[lsu_dccm_ctl.scala 178:171]
  wire  _T_851 = ~_T_850; // @[lsu_dccm_ctl.scala 178:24]
  wire  _T_852 = lsu_dccm_rden_d & _T_851; // @[lsu_dccm_ctl.scala 178:22]
  wire  _T_853 = _T_843 | _T_852; // @[lsu_dccm_ctl.scala 177:124]
  wire  _T_855 = io_dma_dccm_wen | io_lsu_stbuf_commit_any; // @[lsu_dccm_ctl.scala 183:41]
  wire [15:0] _T_862 = ld_single_ecc_error_lo_r_ff ? ld_sec_addr_lo_r_ff : ld_sec_addr_hi_r_ff; // @[lsu_dccm_ctl.scala 187:8]
  wire [15:0] _T_866 = io_dma_dccm_wen ? io_lsu_addr_d[15:0] : io_stbuf_addr_any; // @[lsu_dccm_ctl.scala 188:8]
  wire [15:0] _T_872 = ld_single_ecc_error_hi_r_ff ? ld_sec_addr_hi_r_ff : ld_sec_addr_lo_r_ff; // @[lsu_dccm_ctl.scala 191:8]
  wire [15:0] _T_876 = io_dma_dccm_wen ? io_end_addr_d : io_stbuf_addr_any; // @[lsu_dccm_ctl.scala 192:8]
  wire [38:0] _T_884 = {io_sec_data_ecc_lo_r_ff,io_sec_data_lo_r_ff}; // @[Cat.scala 29:58]
  wire [38:0] _T_887 = {io_sec_data_ecc_hi_r_ff,io_sec_data_hi_r_ff}; // @[Cat.scala 29:58]
  wire [38:0] _T_888 = ld_single_ecc_error_lo_r_ff ? _T_884 : _T_887; // @[lsu_dccm_ctl.scala 198:8]
  wire [38:0] _T_892 = {io_dma_dccm_wdata_ecc_lo,io_dma_dccm_wdata_lo}; // @[Cat.scala 29:58]
  wire [38:0] _T_895 = {io_stbuf_ecc_any,io_stbuf_data_any}; // @[Cat.scala 29:58]
  wire [38:0] _T_896 = io_dma_dccm_wen ? _T_892 : _T_895; // @[lsu_dccm_ctl.scala 200:8]
  wire [38:0] _T_906 = ld_single_ecc_error_hi_r_ff ? _T_887 : _T_884; // @[lsu_dccm_ctl.scala 204:8]
  wire [38:0] _T_910 = {io_dma_dccm_wdata_ecc_hi,io_dma_dccm_wdata_hi}; // @[Cat.scala 29:58]
  wire [38:0] _T_914 = io_dma_dccm_wen ? _T_910 : _T_895; // @[lsu_dccm_ctl.scala 206:8]
  wire [3:0] _T_917 = io_lsu_pkt_m_bits_store ? 4'hf : 4'h0; // @[Bitwise.scala 72:12]
  wire [3:0] _T_919 = io_lsu_pkt_m_bits_by ? 4'hf : 4'h0; // @[Bitwise.scala 72:12]
  wire [3:0] _T_920 = _T_919 & 4'h1; // @[lsu_dccm_ctl.scala 210:94]
  wire [3:0] _T_922 = io_lsu_pkt_m_bits_half ? 4'hf : 4'h0; // @[Bitwise.scala 72:12]
  wire [3:0] _T_923 = _T_922 & 4'h3; // @[lsu_dccm_ctl.scala 211:38]
  wire [3:0] _T_924 = _T_920 | _T_923; // @[lsu_dccm_ctl.scala 210:107]
  wire [3:0] _T_926 = io_lsu_pkt_m_bits_word ? 4'hf : 4'h0; // @[Bitwise.scala 72:12]
  wire [3:0] _T_928 = _T_924 | _T_926; // @[lsu_dccm_ctl.scala 211:51]
  wire [3:0] store_byteen_m = _T_917 & _T_928; // @[lsu_dccm_ctl.scala 210:58]
  wire [3:0] _T_930 = io_lsu_pkt_r_bits_store ? 4'hf : 4'h0; // @[Bitwise.scala 72:12]
  wire [3:0] _T_932 = io_lsu_pkt_r_bits_by ? 4'hf : 4'h0; // @[Bitwise.scala 72:12]
  wire [3:0] _T_933 = _T_932 & 4'h1; // @[lsu_dccm_ctl.scala 214:94]
  wire [3:0] _T_935 = io_lsu_pkt_r_bits_half ? 4'hf : 4'h0; // @[Bitwise.scala 72:12]
  wire [3:0] _T_936 = _T_935 & 4'h3; // @[lsu_dccm_ctl.scala 215:38]
  wire [3:0] _T_937 = _T_933 | _T_936; // @[lsu_dccm_ctl.scala 214:107]
  wire [3:0] _T_939 = io_lsu_pkt_r_bits_word ? 4'hf : 4'h0; // @[Bitwise.scala 72:12]
  wire [3:0] _T_941 = _T_937 | _T_939; // @[lsu_dccm_ctl.scala 215:51]
  wire [3:0] store_byteen_r = _T_930 & _T_941; // @[lsu_dccm_ctl.scala 214:58]
  wire [6:0] _GEN_44 = {{3'd0}, store_byteen_m}; // @[lsu_dccm_ctl.scala 218:45]
  wire [6:0] _T_944 = _GEN_44 << io_lsu_addr_m[1:0]; // @[lsu_dccm_ctl.scala 218:45]
  wire [6:0] _GEN_45 = {{3'd0}, store_byteen_r}; // @[lsu_dccm_ctl.scala 220:45]
  wire [6:0] _T_947 = _GEN_45 << io_lsu_addr_r[1:0]; // @[lsu_dccm_ctl.scala 220:45]
  wire  _T_950 = io_stbuf_addr_any[15:2] == io_lsu_addr_m[15:2]; // @[lsu_dccm_ctl.scala 223:67]
  wire  dccm_wr_bypass_d_m_lo = _T_950 & io_addr_in_dccm_m; // @[lsu_dccm_ctl.scala 223:101]
  wire  _T_953 = io_stbuf_addr_any[15:2] == io_end_addr_m[15:2]; // @[lsu_dccm_ctl.scala 224:67]
  wire  dccm_wr_bypass_d_m_hi = _T_953 & io_addr_in_dccm_m; // @[lsu_dccm_ctl.scala 224:101]
  wire  _T_956 = io_stbuf_addr_any[15:2] == io_lsu_addr_r[15:2]; // @[lsu_dccm_ctl.scala 226:67]
  wire  dccm_wr_bypass_d_r_lo = _T_956 & io_addr_in_dccm_r; // @[lsu_dccm_ctl.scala 226:101]
  wire  _T_959 = io_stbuf_addr_any[15:2] == io_end_addr_r[15:2]; // @[lsu_dccm_ctl.scala 227:67]
  wire  dccm_wr_bypass_d_r_hi = _T_959 & io_addr_in_dccm_r; // @[lsu_dccm_ctl.scala 227:101]
  wire [63:0] _T_962 = {32'h0,io_store_data_m}; // @[Cat.scala 29:58]
  wire [126:0] _GEN_47 = {{63'd0}, _T_962}; // @[lsu_dccm_ctl.scala 256:72]
  wire [126:0] _T_965 = _GEN_47 << _T_762; // @[lsu_dccm_ctl.scala 256:72]
  wire [63:0] store_data_pre_m = _T_965[63:0]; // @[lsu_dccm_ctl.scala 256:29]
  wire [31:0] store_data_hi_m = store_data_pre_m[63:32]; // @[lsu_dccm_ctl.scala 257:48]
  wire [31:0] store_data_lo_m = store_data_pre_m[31:0]; // @[lsu_dccm_ctl.scala 258:48]
  wire [7:0] store_byteen_ext_m = {{1'd0}, _T_944}; // @[lsu_dccm_ctl.scala 218:22]
  wire  _T_971 = io_lsu_stbuf_commit_any & dccm_wr_bypass_d_m_lo; // @[lsu_dccm_ctl.scala 259:211]
  wire [7:0] _T_975 = _T_971 ? io_stbuf_data_any[7:0] : io_sec_data_lo_m[7:0]; // @[lsu_dccm_ctl.scala 259:185]
  wire [7:0] _T_976 = store_byteen_ext_m[0] ? store_data_lo_m[7:0] : _T_975; // @[lsu_dccm_ctl.scala 259:120]
  wire [7:0] _T_980 = {{4'd0}, _T_976[7:4]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_982 = {_T_976[3:0], 4'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_984 = _T_982 & 8'hf0; // @[Bitwise.scala 103:75]
  wire [7:0] _T_985 = _T_980 | _T_984; // @[Bitwise.scala 103:39]
  wire [7:0] _GEN_48 = {{2'd0}, _T_985[7:2]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_990 = _GEN_48 & 8'h33; // @[Bitwise.scala 103:31]
  wire [7:0] _T_992 = {_T_985[5:0], 2'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_994 = _T_992 & 8'hcc; // @[Bitwise.scala 103:75]
  wire [7:0] _T_995 = _T_990 | _T_994; // @[Bitwise.scala 103:39]
  wire [7:0] _GEN_49 = {{1'd0}, _T_995[7:1]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_1000 = _GEN_49 & 8'h55; // @[Bitwise.scala 103:31]
  wire [7:0] _T_1002 = {_T_995[6:0], 1'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_1004 = _T_1002 & 8'haa; // @[Bitwise.scala 103:75]
  wire [7:0] _T_1005 = _T_1000 | _T_1004; // @[Bitwise.scala 103:39]
  wire [7:0] _T_1013 = _T_971 ? io_stbuf_data_any[15:8] : io_sec_data_lo_m[15:8]; // @[lsu_dccm_ctl.scala 259:185]
  wire [7:0] _T_1014 = store_byteen_ext_m[1] ? store_data_lo_m[15:8] : _T_1013; // @[lsu_dccm_ctl.scala 259:120]
  wire [7:0] _T_1018 = {{4'd0}, _T_1014[7:4]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_1020 = {_T_1014[3:0], 4'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_1022 = _T_1020 & 8'hf0; // @[Bitwise.scala 103:75]
  wire [7:0] _T_1023 = _T_1018 | _T_1022; // @[Bitwise.scala 103:39]
  wire [7:0] _GEN_50 = {{2'd0}, _T_1023[7:2]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_1028 = _GEN_50 & 8'h33; // @[Bitwise.scala 103:31]
  wire [7:0] _T_1030 = {_T_1023[5:0], 2'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_1032 = _T_1030 & 8'hcc; // @[Bitwise.scala 103:75]
  wire [7:0] _T_1033 = _T_1028 | _T_1032; // @[Bitwise.scala 103:39]
  wire [7:0] _GEN_51 = {{1'd0}, _T_1033[7:1]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_1038 = _GEN_51 & 8'h55; // @[Bitwise.scala 103:31]
  wire [7:0] _T_1040 = {_T_1033[6:0], 1'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_1042 = _T_1040 & 8'haa; // @[Bitwise.scala 103:75]
  wire [7:0] _T_1043 = _T_1038 | _T_1042; // @[Bitwise.scala 103:39]
  wire [7:0] _T_1051 = _T_971 ? io_stbuf_data_any[23:16] : io_sec_data_lo_m[23:16]; // @[lsu_dccm_ctl.scala 259:185]
  wire [7:0] _T_1052 = store_byteen_ext_m[2] ? store_data_lo_m[23:16] : _T_1051; // @[lsu_dccm_ctl.scala 259:120]
  wire [7:0] _T_1056 = {{4'd0}, _T_1052[7:4]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_1058 = {_T_1052[3:0], 4'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_1060 = _T_1058 & 8'hf0; // @[Bitwise.scala 103:75]
  wire [7:0] _T_1061 = _T_1056 | _T_1060; // @[Bitwise.scala 103:39]
  wire [7:0] _GEN_52 = {{2'd0}, _T_1061[7:2]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_1066 = _GEN_52 & 8'h33; // @[Bitwise.scala 103:31]
  wire [7:0] _T_1068 = {_T_1061[5:0], 2'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_1070 = _T_1068 & 8'hcc; // @[Bitwise.scala 103:75]
  wire [7:0] _T_1071 = _T_1066 | _T_1070; // @[Bitwise.scala 103:39]
  wire [7:0] _GEN_53 = {{1'd0}, _T_1071[7:1]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_1076 = _GEN_53 & 8'h55; // @[Bitwise.scala 103:31]
  wire [7:0] _T_1078 = {_T_1071[6:0], 1'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_1080 = _T_1078 & 8'haa; // @[Bitwise.scala 103:75]
  wire [7:0] _T_1081 = _T_1076 | _T_1080; // @[Bitwise.scala 103:39]
  wire [7:0] _T_1089 = _T_971 ? io_stbuf_data_any[31:24] : io_sec_data_lo_m[31:24]; // @[lsu_dccm_ctl.scala 259:185]
  wire [7:0] _T_1090 = store_byteen_ext_m[3] ? store_data_lo_m[31:24] : _T_1089; // @[lsu_dccm_ctl.scala 259:120]
  wire [7:0] _T_1094 = {{4'd0}, _T_1090[7:4]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_1096 = {_T_1090[3:0], 4'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_1098 = _T_1096 & 8'hf0; // @[Bitwise.scala 103:75]
  wire [7:0] _T_1099 = _T_1094 | _T_1098; // @[Bitwise.scala 103:39]
  wire [7:0] _GEN_54 = {{2'd0}, _T_1099[7:2]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_1104 = _GEN_54 & 8'h33; // @[Bitwise.scala 103:31]
  wire [7:0] _T_1106 = {_T_1099[5:0], 2'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_1108 = _T_1106 & 8'hcc; // @[Bitwise.scala 103:75]
  wire [7:0] _T_1109 = _T_1104 | _T_1108; // @[Bitwise.scala 103:39]
  wire [7:0] _GEN_55 = {{1'd0}, _T_1109[7:1]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_1114 = _GEN_55 & 8'h55; // @[Bitwise.scala 103:31]
  wire [7:0] _T_1116 = {_T_1109[6:0], 1'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_1118 = _T_1116 & 8'haa; // @[Bitwise.scala 103:75]
  wire [7:0] _T_1119 = _T_1114 | _T_1118; // @[Bitwise.scala 103:39]
  wire [31:0] _T_1123 = {_T_1005,_T_1043,_T_1081,_T_1119}; // @[Cat.scala 29:58]
  wire [31:0] _T_1127 = {{16'd0}, _T_1123[31:16]}; // @[Bitwise.scala 103:31]
  wire [31:0] _T_1129 = {_T_1123[15:0], 16'h0}; // @[Bitwise.scala 103:65]
  wire [31:0] _T_1131 = _T_1129 & 32'hffff0000; // @[Bitwise.scala 103:75]
  wire [31:0] _T_1132 = _T_1127 | _T_1131; // @[Bitwise.scala 103:39]
  wire [31:0] _GEN_56 = {{8'd0}, _T_1132[31:8]}; // @[Bitwise.scala 103:31]
  wire [31:0] _T_1137 = _GEN_56 & 32'hff00ff; // @[Bitwise.scala 103:31]
  wire [31:0] _T_1139 = {_T_1132[23:0], 8'h0}; // @[Bitwise.scala 103:65]
  wire [31:0] _T_1141 = _T_1139 & 32'hff00ff00; // @[Bitwise.scala 103:75]
  wire [31:0] _T_1142 = _T_1137 | _T_1141; // @[Bitwise.scala 103:39]
  wire [31:0] _GEN_57 = {{4'd0}, _T_1142[31:4]}; // @[Bitwise.scala 103:31]
  wire [31:0] _T_1147 = _GEN_57 & 32'hf0f0f0f; // @[Bitwise.scala 103:31]
  wire [31:0] _T_1149 = {_T_1142[27:0], 4'h0}; // @[Bitwise.scala 103:65]
  wire [31:0] _T_1151 = _T_1149 & 32'hf0f0f0f0; // @[Bitwise.scala 103:75]
  wire [31:0] _T_1152 = _T_1147 | _T_1151; // @[Bitwise.scala 103:39]
  wire [31:0] _GEN_58 = {{2'd0}, _T_1152[31:2]}; // @[Bitwise.scala 103:31]
  wire [31:0] _T_1157 = _GEN_58 & 32'h33333333; // @[Bitwise.scala 103:31]
  wire [31:0] _T_1159 = {_T_1152[29:0], 2'h0}; // @[Bitwise.scala 103:65]
  wire [31:0] _T_1161 = _T_1159 & 32'hcccccccc; // @[Bitwise.scala 103:75]
  wire [31:0] _T_1162 = _T_1157 | _T_1161; // @[Bitwise.scala 103:39]
  wire [31:0] _GEN_59 = {{1'd0}, _T_1162[31:1]}; // @[Bitwise.scala 103:31]
  wire [31:0] _T_1167 = _GEN_59 & 32'h55555555; // @[Bitwise.scala 103:31]
  wire [31:0] _T_1169 = {_T_1162[30:0], 1'h0}; // @[Bitwise.scala 103:65]
  wire [31:0] _T_1171 = _T_1169 & 32'haaaaaaaa; // @[Bitwise.scala 103:75]
  reg [31:0] _T_1173; // @[lsu_dccm_ctl.scala 259:72]
  wire  _T_1177 = io_lsu_stbuf_commit_any & dccm_wr_bypass_d_m_hi; // @[lsu_dccm_ctl.scala 260:211]
  wire [7:0] _T_1181 = _T_1177 ? io_stbuf_data_any[7:0] : io_sec_data_hi_m[7:0]; // @[lsu_dccm_ctl.scala 260:185]
  wire [7:0] _T_1182 = store_byteen_ext_m[4] ? store_data_hi_m[7:0] : _T_1181; // @[lsu_dccm_ctl.scala 260:120]
  wire [7:0] _T_1186 = {{4'd0}, _T_1182[7:4]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_1188 = {_T_1182[3:0], 4'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_1190 = _T_1188 & 8'hf0; // @[Bitwise.scala 103:75]
  wire [7:0] _T_1191 = _T_1186 | _T_1190; // @[Bitwise.scala 103:39]
  wire [7:0] _GEN_60 = {{2'd0}, _T_1191[7:2]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_1196 = _GEN_60 & 8'h33; // @[Bitwise.scala 103:31]
  wire [7:0] _T_1198 = {_T_1191[5:0], 2'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_1200 = _T_1198 & 8'hcc; // @[Bitwise.scala 103:75]
  wire [7:0] _T_1201 = _T_1196 | _T_1200; // @[Bitwise.scala 103:39]
  wire [7:0] _GEN_61 = {{1'd0}, _T_1201[7:1]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_1206 = _GEN_61 & 8'h55; // @[Bitwise.scala 103:31]
  wire [7:0] _T_1208 = {_T_1201[6:0], 1'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_1210 = _T_1208 & 8'haa; // @[Bitwise.scala 103:75]
  wire [7:0] _T_1211 = _T_1206 | _T_1210; // @[Bitwise.scala 103:39]
  wire [7:0] _T_1219 = _T_1177 ? io_stbuf_data_any[15:8] : io_sec_data_hi_m[15:8]; // @[lsu_dccm_ctl.scala 260:185]
  wire [7:0] _T_1220 = store_byteen_ext_m[5] ? store_data_hi_m[15:8] : _T_1219; // @[lsu_dccm_ctl.scala 260:120]
  wire [7:0] _T_1224 = {{4'd0}, _T_1220[7:4]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_1226 = {_T_1220[3:0], 4'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_1228 = _T_1226 & 8'hf0; // @[Bitwise.scala 103:75]
  wire [7:0] _T_1229 = _T_1224 | _T_1228; // @[Bitwise.scala 103:39]
  wire [7:0] _GEN_62 = {{2'd0}, _T_1229[7:2]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_1234 = _GEN_62 & 8'h33; // @[Bitwise.scala 103:31]
  wire [7:0] _T_1236 = {_T_1229[5:0], 2'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_1238 = _T_1236 & 8'hcc; // @[Bitwise.scala 103:75]
  wire [7:0] _T_1239 = _T_1234 | _T_1238; // @[Bitwise.scala 103:39]
  wire [7:0] _GEN_63 = {{1'd0}, _T_1239[7:1]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_1244 = _GEN_63 & 8'h55; // @[Bitwise.scala 103:31]
  wire [7:0] _T_1246 = {_T_1239[6:0], 1'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_1248 = _T_1246 & 8'haa; // @[Bitwise.scala 103:75]
  wire [7:0] _T_1249 = _T_1244 | _T_1248; // @[Bitwise.scala 103:39]
  wire [7:0] _T_1257 = _T_1177 ? io_stbuf_data_any[23:16] : io_sec_data_hi_m[23:16]; // @[lsu_dccm_ctl.scala 260:185]
  wire [7:0] _T_1258 = store_byteen_ext_m[6] ? store_data_hi_m[23:16] : _T_1257; // @[lsu_dccm_ctl.scala 260:120]
  wire [7:0] _T_1262 = {{4'd0}, _T_1258[7:4]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_1264 = {_T_1258[3:0], 4'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_1266 = _T_1264 & 8'hf0; // @[Bitwise.scala 103:75]
  wire [7:0] _T_1267 = _T_1262 | _T_1266; // @[Bitwise.scala 103:39]
  wire [7:0] _GEN_64 = {{2'd0}, _T_1267[7:2]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_1272 = _GEN_64 & 8'h33; // @[Bitwise.scala 103:31]
  wire [7:0] _T_1274 = {_T_1267[5:0], 2'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_1276 = _T_1274 & 8'hcc; // @[Bitwise.scala 103:75]
  wire [7:0] _T_1277 = _T_1272 | _T_1276; // @[Bitwise.scala 103:39]
  wire [7:0] _GEN_65 = {{1'd0}, _T_1277[7:1]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_1282 = _GEN_65 & 8'h55; // @[Bitwise.scala 103:31]
  wire [7:0] _T_1284 = {_T_1277[6:0], 1'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_1286 = _T_1284 & 8'haa; // @[Bitwise.scala 103:75]
  wire [7:0] _T_1287 = _T_1282 | _T_1286; // @[Bitwise.scala 103:39]
  wire [7:0] _T_1295 = _T_1177 ? io_stbuf_data_any[31:24] : io_sec_data_hi_m[31:24]; // @[lsu_dccm_ctl.scala 260:185]
  wire [7:0] _T_1296 = store_byteen_ext_m[7] ? store_data_hi_m[31:24] : _T_1295; // @[lsu_dccm_ctl.scala 260:120]
  wire [7:0] _T_1300 = {{4'd0}, _T_1296[7:4]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_1302 = {_T_1296[3:0], 4'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_1304 = _T_1302 & 8'hf0; // @[Bitwise.scala 103:75]
  wire [7:0] _T_1305 = _T_1300 | _T_1304; // @[Bitwise.scala 103:39]
  wire [7:0] _GEN_66 = {{2'd0}, _T_1305[7:2]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_1310 = _GEN_66 & 8'h33; // @[Bitwise.scala 103:31]
  wire [7:0] _T_1312 = {_T_1305[5:0], 2'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_1314 = _T_1312 & 8'hcc; // @[Bitwise.scala 103:75]
  wire [7:0] _T_1315 = _T_1310 | _T_1314; // @[Bitwise.scala 103:39]
  wire [7:0] _GEN_67 = {{1'd0}, _T_1315[7:1]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_1320 = _GEN_67 & 8'h55; // @[Bitwise.scala 103:31]
  wire [7:0] _T_1322 = {_T_1315[6:0], 1'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_1324 = _T_1322 & 8'haa; // @[Bitwise.scala 103:75]
  wire [7:0] _T_1325 = _T_1320 | _T_1324; // @[Bitwise.scala 103:39]
  wire [31:0] _T_1329 = {_T_1211,_T_1249,_T_1287,_T_1325}; // @[Cat.scala 29:58]
  wire [31:0] _T_1333 = {{16'd0}, _T_1329[31:16]}; // @[Bitwise.scala 103:31]
  wire [31:0] _T_1335 = {_T_1329[15:0], 16'h0}; // @[Bitwise.scala 103:65]
  wire [31:0] _T_1337 = _T_1335 & 32'hffff0000; // @[Bitwise.scala 103:75]
  wire [31:0] _T_1338 = _T_1333 | _T_1337; // @[Bitwise.scala 103:39]
  wire [31:0] _GEN_68 = {{8'd0}, _T_1338[31:8]}; // @[Bitwise.scala 103:31]
  wire [31:0] _T_1343 = _GEN_68 & 32'hff00ff; // @[Bitwise.scala 103:31]
  wire [31:0] _T_1345 = {_T_1338[23:0], 8'h0}; // @[Bitwise.scala 103:65]
  wire [31:0] _T_1347 = _T_1345 & 32'hff00ff00; // @[Bitwise.scala 103:75]
  wire [31:0] _T_1348 = _T_1343 | _T_1347; // @[Bitwise.scala 103:39]
  wire [31:0] _GEN_69 = {{4'd0}, _T_1348[31:4]}; // @[Bitwise.scala 103:31]
  wire [31:0] _T_1353 = _GEN_69 & 32'hf0f0f0f; // @[Bitwise.scala 103:31]
  wire [31:0] _T_1355 = {_T_1348[27:0], 4'h0}; // @[Bitwise.scala 103:65]
  wire [31:0] _T_1357 = _T_1355 & 32'hf0f0f0f0; // @[Bitwise.scala 103:75]
  wire [31:0] _T_1358 = _T_1353 | _T_1357; // @[Bitwise.scala 103:39]
  wire [31:0] _GEN_70 = {{2'd0}, _T_1358[31:2]}; // @[Bitwise.scala 103:31]
  wire [31:0] _T_1363 = _GEN_70 & 32'h33333333; // @[Bitwise.scala 103:31]
  wire [31:0] _T_1365 = {_T_1358[29:0], 2'h0}; // @[Bitwise.scala 103:65]
  wire [31:0] _T_1367 = _T_1365 & 32'hcccccccc; // @[Bitwise.scala 103:75]
  wire [31:0] _T_1368 = _T_1363 | _T_1367; // @[Bitwise.scala 103:39]
  wire [31:0] _GEN_71 = {{1'd0}, _T_1368[31:1]}; // @[Bitwise.scala 103:31]
  wire [31:0] _T_1373 = _GEN_71 & 32'h55555555; // @[Bitwise.scala 103:31]
  wire [31:0] _T_1375 = {_T_1368[30:0], 1'h0}; // @[Bitwise.scala 103:65]
  wire [31:0] _T_1377 = _T_1375 & 32'haaaaaaaa; // @[Bitwise.scala 103:75]
  reg [31:0] _T_1379; // @[lsu_dccm_ctl.scala 260:72]
  wire  _T_1380 = io_lsu_stbuf_commit_any & dccm_wr_bypass_d_r_lo; // @[lsu_dccm_ctl.scala 261:105]
  wire [7:0] store_byteen_ext_r = {{1'd0}, _T_947}; // @[lsu_dccm_ctl.scala 220:22]
  wire  _T_1382 = ~store_byteen_ext_r[0]; // @[lsu_dccm_ctl.scala 261:131]
  wire  _T_1383 = _T_1380 & _T_1382; // @[lsu_dccm_ctl.scala 261:129]
  wire [7:0] _T_1387 = _T_1383 ? io_stbuf_data_any[7:0] : io_store_data_lo_r[7:0]; // @[lsu_dccm_ctl.scala 261:79]
  wire [7:0] _T_1391 = {{4'd0}, _T_1387[7:4]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_1393 = {_T_1387[3:0], 4'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_1395 = _T_1393 & 8'hf0; // @[Bitwise.scala 103:75]
  wire [7:0] _T_1396 = _T_1391 | _T_1395; // @[Bitwise.scala 103:39]
  wire [7:0] _GEN_72 = {{2'd0}, _T_1396[7:2]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_1401 = _GEN_72 & 8'h33; // @[Bitwise.scala 103:31]
  wire [7:0] _T_1403 = {_T_1396[5:0], 2'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_1405 = _T_1403 & 8'hcc; // @[Bitwise.scala 103:75]
  wire [7:0] _T_1406 = _T_1401 | _T_1405; // @[Bitwise.scala 103:39]
  wire [7:0] _GEN_73 = {{1'd0}, _T_1406[7:1]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_1411 = _GEN_73 & 8'h55; // @[Bitwise.scala 103:31]
  wire [7:0] _T_1413 = {_T_1406[6:0], 1'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_1415 = _T_1413 & 8'haa; // @[Bitwise.scala 103:75]
  wire [7:0] _T_1416 = _T_1411 | _T_1415; // @[Bitwise.scala 103:39]
  wire  _T_1419 = ~store_byteen_ext_r[1]; // @[lsu_dccm_ctl.scala 261:131]
  wire  _T_1420 = _T_1380 & _T_1419; // @[lsu_dccm_ctl.scala 261:129]
  wire [7:0] _T_1424 = _T_1420 ? io_stbuf_data_any[15:8] : io_store_data_lo_r[15:8]; // @[lsu_dccm_ctl.scala 261:79]
  wire [7:0] _T_1428 = {{4'd0}, _T_1424[7:4]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_1430 = {_T_1424[3:0], 4'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_1432 = _T_1430 & 8'hf0; // @[Bitwise.scala 103:75]
  wire [7:0] _T_1433 = _T_1428 | _T_1432; // @[Bitwise.scala 103:39]
  wire [7:0] _GEN_74 = {{2'd0}, _T_1433[7:2]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_1438 = _GEN_74 & 8'h33; // @[Bitwise.scala 103:31]
  wire [7:0] _T_1440 = {_T_1433[5:0], 2'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_1442 = _T_1440 & 8'hcc; // @[Bitwise.scala 103:75]
  wire [7:0] _T_1443 = _T_1438 | _T_1442; // @[Bitwise.scala 103:39]
  wire [7:0] _GEN_75 = {{1'd0}, _T_1443[7:1]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_1448 = _GEN_75 & 8'h55; // @[Bitwise.scala 103:31]
  wire [7:0] _T_1450 = {_T_1443[6:0], 1'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_1452 = _T_1450 & 8'haa; // @[Bitwise.scala 103:75]
  wire [7:0] _T_1453 = _T_1448 | _T_1452; // @[Bitwise.scala 103:39]
  wire  _T_1456 = ~store_byteen_ext_r[2]; // @[lsu_dccm_ctl.scala 261:131]
  wire  _T_1457 = _T_1380 & _T_1456; // @[lsu_dccm_ctl.scala 261:129]
  wire [7:0] _T_1461 = _T_1457 ? io_stbuf_data_any[23:16] : io_store_data_lo_r[23:16]; // @[lsu_dccm_ctl.scala 261:79]
  wire [7:0] _T_1465 = {{4'd0}, _T_1461[7:4]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_1467 = {_T_1461[3:0], 4'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_1469 = _T_1467 & 8'hf0; // @[Bitwise.scala 103:75]
  wire [7:0] _T_1470 = _T_1465 | _T_1469; // @[Bitwise.scala 103:39]
  wire [7:0] _GEN_76 = {{2'd0}, _T_1470[7:2]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_1475 = _GEN_76 & 8'h33; // @[Bitwise.scala 103:31]
  wire [7:0] _T_1477 = {_T_1470[5:0], 2'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_1479 = _T_1477 & 8'hcc; // @[Bitwise.scala 103:75]
  wire [7:0] _T_1480 = _T_1475 | _T_1479; // @[Bitwise.scala 103:39]
  wire [7:0] _GEN_77 = {{1'd0}, _T_1480[7:1]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_1485 = _GEN_77 & 8'h55; // @[Bitwise.scala 103:31]
  wire [7:0] _T_1487 = {_T_1480[6:0], 1'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_1489 = _T_1487 & 8'haa; // @[Bitwise.scala 103:75]
  wire [7:0] _T_1490 = _T_1485 | _T_1489; // @[Bitwise.scala 103:39]
  wire  _T_1493 = ~store_byteen_ext_r[3]; // @[lsu_dccm_ctl.scala 261:131]
  wire  _T_1494 = _T_1380 & _T_1493; // @[lsu_dccm_ctl.scala 261:129]
  wire [7:0] _T_1498 = _T_1494 ? io_stbuf_data_any[31:24] : io_store_data_lo_r[31:24]; // @[lsu_dccm_ctl.scala 261:79]
  wire [7:0] _T_1502 = {{4'd0}, _T_1498[7:4]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_1504 = {_T_1498[3:0], 4'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_1506 = _T_1504 & 8'hf0; // @[Bitwise.scala 103:75]
  wire [7:0] _T_1507 = _T_1502 | _T_1506; // @[Bitwise.scala 103:39]
  wire [7:0] _GEN_78 = {{2'd0}, _T_1507[7:2]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_1512 = _GEN_78 & 8'h33; // @[Bitwise.scala 103:31]
  wire [7:0] _T_1514 = {_T_1507[5:0], 2'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_1516 = _T_1514 & 8'hcc; // @[Bitwise.scala 103:75]
  wire [7:0] _T_1517 = _T_1512 | _T_1516; // @[Bitwise.scala 103:39]
  wire [7:0] _GEN_79 = {{1'd0}, _T_1517[7:1]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_1522 = _GEN_79 & 8'h55; // @[Bitwise.scala 103:31]
  wire [7:0] _T_1524 = {_T_1517[6:0], 1'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_1526 = _T_1524 & 8'haa; // @[Bitwise.scala 103:75]
  wire [7:0] _T_1527 = _T_1522 | _T_1526; // @[Bitwise.scala 103:39]
  wire [31:0] _T_1531 = {_T_1416,_T_1453,_T_1490,_T_1527}; // @[Cat.scala 29:58]
  wire [31:0] _T_1535 = {{16'd0}, _T_1531[31:16]}; // @[Bitwise.scala 103:31]
  wire [31:0] _T_1537 = {_T_1531[15:0], 16'h0}; // @[Bitwise.scala 103:65]
  wire [31:0] _T_1539 = _T_1537 & 32'hffff0000; // @[Bitwise.scala 103:75]
  wire [31:0] _T_1540 = _T_1535 | _T_1539; // @[Bitwise.scala 103:39]
  wire [31:0] _GEN_80 = {{8'd0}, _T_1540[31:8]}; // @[Bitwise.scala 103:31]
  wire [31:0] _T_1545 = _GEN_80 & 32'hff00ff; // @[Bitwise.scala 103:31]
  wire [31:0] _T_1547 = {_T_1540[23:0], 8'h0}; // @[Bitwise.scala 103:65]
  wire [31:0] _T_1549 = _T_1547 & 32'hff00ff00; // @[Bitwise.scala 103:75]
  wire [31:0] _T_1550 = _T_1545 | _T_1549; // @[Bitwise.scala 103:39]
  wire [31:0] _GEN_81 = {{4'd0}, _T_1550[31:4]}; // @[Bitwise.scala 103:31]
  wire [31:0] _T_1555 = _GEN_81 & 32'hf0f0f0f; // @[Bitwise.scala 103:31]
  wire [31:0] _T_1557 = {_T_1550[27:0], 4'h0}; // @[Bitwise.scala 103:65]
  wire [31:0] _T_1559 = _T_1557 & 32'hf0f0f0f0; // @[Bitwise.scala 103:75]
  wire [31:0] _T_1560 = _T_1555 | _T_1559; // @[Bitwise.scala 103:39]
  wire [31:0] _GEN_82 = {{2'd0}, _T_1560[31:2]}; // @[Bitwise.scala 103:31]
  wire [31:0] _T_1565 = _GEN_82 & 32'h33333333; // @[Bitwise.scala 103:31]
  wire [31:0] _T_1567 = {_T_1560[29:0], 2'h0}; // @[Bitwise.scala 103:65]
  wire [31:0] _T_1569 = _T_1567 & 32'hcccccccc; // @[Bitwise.scala 103:75]
  wire [31:0] _T_1570 = _T_1565 | _T_1569; // @[Bitwise.scala 103:39]
  wire [31:0] _GEN_83 = {{1'd0}, _T_1570[31:1]}; // @[Bitwise.scala 103:31]
  wire [31:0] _T_1575 = _GEN_83 & 32'h55555555; // @[Bitwise.scala 103:31]
  wire [31:0] _T_1577 = {_T_1570[30:0], 1'h0}; // @[Bitwise.scala 103:65]
  wire [31:0] _T_1579 = _T_1577 & 32'haaaaaaaa; // @[Bitwise.scala 103:75]
  wire  _T_1581 = io_lsu_stbuf_commit_any & dccm_wr_bypass_d_r_hi; // @[lsu_dccm_ctl.scala 262:105]
  wire  _T_1583 = ~store_byteen_ext_r[4]; // @[lsu_dccm_ctl.scala 262:131]
  wire  _T_1584 = _T_1581 & _T_1583; // @[lsu_dccm_ctl.scala 262:129]
  wire [7:0] _T_1588 = _T_1584 ? io_stbuf_data_any[7:0] : io_store_data_hi_r[7:0]; // @[lsu_dccm_ctl.scala 262:79]
  wire [7:0] _T_1592 = {{4'd0}, _T_1588[7:4]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_1594 = {_T_1588[3:0], 4'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_1596 = _T_1594 & 8'hf0; // @[Bitwise.scala 103:75]
  wire [7:0] _T_1597 = _T_1592 | _T_1596; // @[Bitwise.scala 103:39]
  wire [7:0] _GEN_84 = {{2'd0}, _T_1597[7:2]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_1602 = _GEN_84 & 8'h33; // @[Bitwise.scala 103:31]
  wire [7:0] _T_1604 = {_T_1597[5:0], 2'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_1606 = _T_1604 & 8'hcc; // @[Bitwise.scala 103:75]
  wire [7:0] _T_1607 = _T_1602 | _T_1606; // @[Bitwise.scala 103:39]
  wire [7:0] _GEN_85 = {{1'd0}, _T_1607[7:1]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_1612 = _GEN_85 & 8'h55; // @[Bitwise.scala 103:31]
  wire [7:0] _T_1614 = {_T_1607[6:0], 1'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_1616 = _T_1614 & 8'haa; // @[Bitwise.scala 103:75]
  wire [7:0] _T_1617 = _T_1612 | _T_1616; // @[Bitwise.scala 103:39]
  wire  _T_1620 = ~store_byteen_ext_r[5]; // @[lsu_dccm_ctl.scala 262:131]
  wire  _T_1621 = _T_1581 & _T_1620; // @[lsu_dccm_ctl.scala 262:129]
  wire [7:0] _T_1625 = _T_1621 ? io_stbuf_data_any[15:8] : io_store_data_hi_r[15:8]; // @[lsu_dccm_ctl.scala 262:79]
  wire [7:0] _T_1629 = {{4'd0}, _T_1625[7:4]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_1631 = {_T_1625[3:0], 4'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_1633 = _T_1631 & 8'hf0; // @[Bitwise.scala 103:75]
  wire [7:0] _T_1634 = _T_1629 | _T_1633; // @[Bitwise.scala 103:39]
  wire [7:0] _GEN_86 = {{2'd0}, _T_1634[7:2]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_1639 = _GEN_86 & 8'h33; // @[Bitwise.scala 103:31]
  wire [7:0] _T_1641 = {_T_1634[5:0], 2'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_1643 = _T_1641 & 8'hcc; // @[Bitwise.scala 103:75]
  wire [7:0] _T_1644 = _T_1639 | _T_1643; // @[Bitwise.scala 103:39]
  wire [7:0] _GEN_87 = {{1'd0}, _T_1644[7:1]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_1649 = _GEN_87 & 8'h55; // @[Bitwise.scala 103:31]
  wire [7:0] _T_1651 = {_T_1644[6:0], 1'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_1653 = _T_1651 & 8'haa; // @[Bitwise.scala 103:75]
  wire [7:0] _T_1654 = _T_1649 | _T_1653; // @[Bitwise.scala 103:39]
  wire  _T_1657 = ~store_byteen_ext_r[6]; // @[lsu_dccm_ctl.scala 262:131]
  wire  _T_1658 = _T_1581 & _T_1657; // @[lsu_dccm_ctl.scala 262:129]
  wire [7:0] _T_1662 = _T_1658 ? io_stbuf_data_any[23:16] : io_store_data_hi_r[23:16]; // @[lsu_dccm_ctl.scala 262:79]
  wire [7:0] _T_1666 = {{4'd0}, _T_1662[7:4]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_1668 = {_T_1662[3:0], 4'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_1670 = _T_1668 & 8'hf0; // @[Bitwise.scala 103:75]
  wire [7:0] _T_1671 = _T_1666 | _T_1670; // @[Bitwise.scala 103:39]
  wire [7:0] _GEN_88 = {{2'd0}, _T_1671[7:2]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_1676 = _GEN_88 & 8'h33; // @[Bitwise.scala 103:31]
  wire [7:0] _T_1678 = {_T_1671[5:0], 2'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_1680 = _T_1678 & 8'hcc; // @[Bitwise.scala 103:75]
  wire [7:0] _T_1681 = _T_1676 | _T_1680; // @[Bitwise.scala 103:39]
  wire [7:0] _GEN_89 = {{1'd0}, _T_1681[7:1]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_1686 = _GEN_89 & 8'h55; // @[Bitwise.scala 103:31]
  wire [7:0] _T_1688 = {_T_1681[6:0], 1'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_1690 = _T_1688 & 8'haa; // @[Bitwise.scala 103:75]
  wire [7:0] _T_1691 = _T_1686 | _T_1690; // @[Bitwise.scala 103:39]
  wire  _T_1694 = ~store_byteen_ext_r[7]; // @[lsu_dccm_ctl.scala 262:131]
  wire  _T_1695 = _T_1581 & _T_1694; // @[lsu_dccm_ctl.scala 262:129]
  wire [7:0] _T_1699 = _T_1695 ? io_stbuf_data_any[31:24] : io_store_data_hi_r[31:24]; // @[lsu_dccm_ctl.scala 262:79]
  wire [7:0] _T_1703 = {{4'd0}, _T_1699[7:4]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_1705 = {_T_1699[3:0], 4'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_1707 = _T_1705 & 8'hf0; // @[Bitwise.scala 103:75]
  wire [7:0] _T_1708 = _T_1703 | _T_1707; // @[Bitwise.scala 103:39]
  wire [7:0] _GEN_90 = {{2'd0}, _T_1708[7:2]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_1713 = _GEN_90 & 8'h33; // @[Bitwise.scala 103:31]
  wire [7:0] _T_1715 = {_T_1708[5:0], 2'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_1717 = _T_1715 & 8'hcc; // @[Bitwise.scala 103:75]
  wire [7:0] _T_1718 = _T_1713 | _T_1717; // @[Bitwise.scala 103:39]
  wire [7:0] _GEN_91 = {{1'd0}, _T_1718[7:1]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_1723 = _GEN_91 & 8'h55; // @[Bitwise.scala 103:31]
  wire [7:0] _T_1725 = {_T_1718[6:0], 1'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_1727 = _T_1725 & 8'haa; // @[Bitwise.scala 103:75]
  wire [7:0] _T_1728 = _T_1723 | _T_1727; // @[Bitwise.scala 103:39]
  wire [31:0] _T_1732 = {_T_1617,_T_1654,_T_1691,_T_1728}; // @[Cat.scala 29:58]
  wire [31:0] _T_1736 = {{16'd0}, _T_1732[31:16]}; // @[Bitwise.scala 103:31]
  wire [31:0] _T_1738 = {_T_1732[15:0], 16'h0}; // @[Bitwise.scala 103:65]
  wire [31:0] _T_1740 = _T_1738 & 32'hffff0000; // @[Bitwise.scala 103:75]
  wire [31:0] _T_1741 = _T_1736 | _T_1740; // @[Bitwise.scala 103:39]
  wire [31:0] _GEN_92 = {{8'd0}, _T_1741[31:8]}; // @[Bitwise.scala 103:31]
  wire [31:0] _T_1746 = _GEN_92 & 32'hff00ff; // @[Bitwise.scala 103:31]
  wire [31:0] _T_1748 = {_T_1741[23:0], 8'h0}; // @[Bitwise.scala 103:65]
  wire [31:0] _T_1750 = _T_1748 & 32'hff00ff00; // @[Bitwise.scala 103:75]
  wire [31:0] _T_1751 = _T_1746 | _T_1750; // @[Bitwise.scala 103:39]
  wire [31:0] _GEN_93 = {{4'd0}, _T_1751[31:4]}; // @[Bitwise.scala 103:31]
  wire [31:0] _T_1756 = _GEN_93 & 32'hf0f0f0f; // @[Bitwise.scala 103:31]
  wire [31:0] _T_1758 = {_T_1751[27:0], 4'h0}; // @[Bitwise.scala 103:65]
  wire [31:0] _T_1760 = _T_1758 & 32'hf0f0f0f0; // @[Bitwise.scala 103:75]
  wire [31:0] _T_1761 = _T_1756 | _T_1760; // @[Bitwise.scala 103:39]
  wire [31:0] _GEN_94 = {{2'd0}, _T_1761[31:2]}; // @[Bitwise.scala 103:31]
  wire [31:0] _T_1766 = _GEN_94 & 32'h33333333; // @[Bitwise.scala 103:31]
  wire [31:0] _T_1768 = {_T_1761[29:0], 2'h0}; // @[Bitwise.scala 103:65]
  wire [31:0] _T_1770 = _T_1768 & 32'hcccccccc; // @[Bitwise.scala 103:75]
  wire [31:0] _T_1771 = _T_1766 | _T_1770; // @[Bitwise.scala 103:39]
  wire [31:0] _GEN_95 = {{1'd0}, _T_1771[31:1]}; // @[Bitwise.scala 103:31]
  wire [31:0] _T_1776 = _GEN_95 & 32'h55555555; // @[Bitwise.scala 103:31]
  wire [31:0] _T_1778 = {_T_1771[30:0], 1'h0}; // @[Bitwise.scala 103:65]
  wire [31:0] _T_1780 = _T_1778 & 32'haaaaaaaa; // @[Bitwise.scala 103:75]
  wire [63:0] _T_1784 = {io_store_data_hi_r,io_store_data_lo_r}; // @[Cat.scala 29:58]
  wire [3:0] _GEN_96 = {{2'd0}, io_lsu_addr_r[1:0]}; // @[lsu_dccm_ctl.scala 263:94]
  wire [5:0] _T_1786 = 4'h8 * _GEN_96; // @[lsu_dccm_ctl.scala 263:94]
  wire [63:0] _T_1787 = _T_1784 >> _T_1786; // @[lsu_dccm_ctl.scala 263:88]
  wire [7:0] _T_1790 = store_byteen_r[0] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_1793 = store_byteen_r[1] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_1796 = store_byteen_r[2] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_1799 = store_byteen_r[3] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_1803 = {_T_1790,_T_1793,_T_1796,_T_1799}; // @[Cat.scala 29:58]
  wire [31:0] _T_1807 = {{16'd0}, _T_1803[31:16]}; // @[Bitwise.scala 103:31]
  wire [31:0] _T_1809 = {_T_1803[15:0], 16'h0}; // @[Bitwise.scala 103:65]
  wire [31:0] _T_1811 = _T_1809 & 32'hffff0000; // @[Bitwise.scala 103:75]
  wire [31:0] _T_1812 = _T_1807 | _T_1811; // @[Bitwise.scala 103:39]
  wire [31:0] _GEN_97 = {{8'd0}, _T_1812[31:8]}; // @[Bitwise.scala 103:31]
  wire [31:0] _T_1817 = _GEN_97 & 32'hff00ff; // @[Bitwise.scala 103:31]
  wire [31:0] _T_1819 = {_T_1812[23:0], 8'h0}; // @[Bitwise.scala 103:65]
  wire [31:0] _T_1821 = _T_1819 & 32'hff00ff00; // @[Bitwise.scala 103:75]
  wire [31:0] _T_1822 = _T_1817 | _T_1821; // @[Bitwise.scala 103:39]
  wire [31:0] _GEN_98 = {{4'd0}, _T_1822[31:4]}; // @[Bitwise.scala 103:31]
  wire [31:0] _T_1827 = _GEN_98 & 32'hf0f0f0f; // @[Bitwise.scala 103:31]
  wire [31:0] _T_1829 = {_T_1822[27:0], 4'h0}; // @[Bitwise.scala 103:65]
  wire [31:0] _T_1831 = _T_1829 & 32'hf0f0f0f0; // @[Bitwise.scala 103:75]
  wire [31:0] _T_1832 = _T_1827 | _T_1831; // @[Bitwise.scala 103:39]
  wire [31:0] _GEN_99 = {{2'd0}, _T_1832[31:2]}; // @[Bitwise.scala 103:31]
  wire [31:0] _T_1837 = _GEN_99 & 32'h33333333; // @[Bitwise.scala 103:31]
  wire [31:0] _T_1839 = {_T_1832[29:0], 2'h0}; // @[Bitwise.scala 103:65]
  wire [31:0] _T_1841 = _T_1839 & 32'hcccccccc; // @[Bitwise.scala 103:75]
  wire [31:0] _T_1842 = _T_1837 | _T_1841; // @[Bitwise.scala 103:39]
  wire [31:0] _GEN_100 = {{1'd0}, _T_1842[31:1]}; // @[Bitwise.scala 103:31]
  wire [31:0] _T_1847 = _GEN_100 & 32'h55555555; // @[Bitwise.scala 103:31]
  wire [31:0] _T_1849 = {_T_1842[30:0], 1'h0}; // @[Bitwise.scala 103:65]
  wire [31:0] _T_1851 = _T_1849 & 32'haaaaaaaa; // @[Bitwise.scala 103:75]
  wire [31:0] _T_1852 = _T_1847 | _T_1851; // @[Bitwise.scala 103:39]
  wire [63:0] _GEN_101 = {{32'd0}, _T_1852}; // @[lsu_dccm_ctl.scala 263:115]
  wire [63:0] _T_1853 = _T_1787 & _GEN_101; // @[lsu_dccm_ctl.scala 263:115]
  wire  _T_1858 = io_lsu_pkt_r_valid & io_lsu_pkt_r_bits_store; // @[lsu_dccm_ctl.scala 270:58]
  wire  _T_1859 = _T_1858 & io_addr_in_pic_r; // @[lsu_dccm_ctl.scala 270:84]
  wire  _T_1860 = _T_1859 & io_lsu_commit_r; // @[lsu_dccm_ctl.scala 270:103]
  wire  _T_1862 = io_lsu_pkt_d_valid & io_lsu_pkt_d_bits_load; // @[lsu_dccm_ctl.scala 271:58]
  wire  _T_1864 = io_lsu_pkt_d_valid & io_lsu_pkt_d_bits_store; // @[lsu_dccm_ctl.scala 272:58]
  wire [31:0] _T_1868 = {17'h0,io_lsu_addr_d[14:0]}; // @[Cat.scala 29:58]
  wire [14:0] _T_1874 = io_dma_pic_wen ? io_dma_dccm_ctl_dma_mem_addr[14:0] : io_lsu_addr_r[14:0]; // @[lsu_dccm_ctl.scala 274:93]
  wire [31:0] _T_1875 = {17'h0,_T_1874}; // @[Cat.scala 29:58]
  reg  _T_1882; // @[lsu_dccm_ctl.scala 279:61]
  rvclkhdr rvclkhdr ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_io_l1clk),
    .io_clk(rvclkhdr_io_clk),
    .io_en(rvclkhdr_io_en),
    .io_scan_mode(rvclkhdr_io_scan_mode)
  );
  rvclkhdr rvclkhdr_1 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_1_io_l1clk),
    .io_clk(rvclkhdr_1_io_clk),
    .io_en(rvclkhdr_1_io_en),
    .io_scan_mode(rvclkhdr_1_io_scan_mode)
  );
  assign io_lsu_ld_data_corr_r = _T_2[31:0]; // @[lsu_dccm_ctl.scala 147:28]
  assign io_dccm_rdata_hi_m = io_dccm_rd_data_hi[31:0]; // @[lsu_dccm_ctl.scala 266:27]
  assign io_dccm_rdata_lo_m = io_dccm_rd_data_lo[31:0]; // @[lsu_dccm_ctl.scala 265:27]
  assign io_dccm_data_ecc_hi_m = io_dccm_rd_data_hi[38:32]; // @[lsu_dccm_ctl.scala 268:27]
  assign io_dccm_data_ecc_lo_m = io_dccm_rd_data_lo[38:32]; // @[lsu_dccm_ctl.scala 267:27]
  assign io_lsu_ld_data_m = _T_763[31:0]; // @[lsu_dccm_ctl.scala 150:28]
  assign io_store_data_hi_r = _T_1379; // @[lsu_dccm_ctl.scala 260:29]
  assign io_store_data_lo_r = _T_1173; // @[lsu_dccm_ctl.scala 259:29]
  assign io_store_datafn_hi_r = _T_1776 | _T_1780; // @[lsu_dccm_ctl.scala 262:29]
  assign io_store_datafn_lo_r = _T_1575 | _T_1579; // @[lsu_dccm_ctl.scala 261:29]
  assign io_store_data_r = _T_1853[31:0]; // @[lsu_dccm_ctl.scala 263:29]
  assign io_ld_single_ecc_error_r = _T_815 & _T_816; // @[lsu_dccm_ctl.scala 163:34]
  assign io_ld_single_ecc_error_r_ff = _T_838 & _T_839; // @[lsu_dccm_ctl.scala 176:31]
  assign io_picm_mask_data_m = picm_rd_data_m[31:0]; // @[lsu_dccm_ctl.scala 275:27]
  assign io_lsu_stbuf_commit_any = io_stbuf_reqvld_any & _T_853; // @[lsu_dccm_ctl.scala 177:31]
  assign io_lsu_dccm_rden_m = _T_1882; // @[lsu_dccm_ctl.scala 279:24]
  assign io_dma_dccm_ctl_dccm_dma_rvalid = _T & io_lsu_pkt_m_bits_dma; // @[lsu_dccm_ctl.scala 137:41]
  assign io_dma_dccm_ctl_dccm_dma_ecc_error = io_lsu_double_ecc_error_m; // @[lsu_dccm_ctl.scala 138:41]
  assign io_dma_dccm_ctl_dccm_dma_rtag = io_dma_mem_tag_m; // @[lsu_dccm_ctl.scala 140:41]
  assign io_dma_dccm_ctl_dccm_dma_rdata = _T_376 | _T_380; // @[lsu_dccm_ctl.scala 139:41]
  assign io_dccm_wren = _T_855 | io_ld_single_ecc_error_r_ff; // @[lsu_dccm_ctl.scala 183:22]
  assign io_dccm_rden = lsu_dccm_rden_d & io_addr_in_dccm_d; // @[lsu_dccm_ctl.scala 184:22]
  assign io_dccm_wr_addr_lo = io_ld_single_ecc_error_r_ff ? _T_862 : _T_866; // @[lsu_dccm_ctl.scala 186:22]
  assign io_dccm_wr_addr_hi = io_ld_single_ecc_error_r_ff ? _T_872 : _T_876; // @[lsu_dccm_ctl.scala 190:22]
  assign io_dccm_rd_addr_lo = io_lsu_addr_d[15:0]; // @[lsu_dccm_ctl.scala 194:22]
  assign io_dccm_rd_addr_hi = io_end_addr_d; // @[lsu_dccm_ctl.scala 195:22]
  assign io_dccm_wr_data_lo = io_ld_single_ecc_error_r_ff ? _T_888 : _T_896; // @[lsu_dccm_ctl.scala 197:22]
  assign io_dccm_wr_data_hi = io_ld_single_ecc_error_r_ff ? _T_906 : _T_914; // @[lsu_dccm_ctl.scala 203:22]
  assign io_lsu_pic_picm_wren = _T_1860 | io_dma_pic_wen; // @[lsu_dccm_ctl.scala 270:35]
  assign io_lsu_pic_picm_rden = _T_1862 & io_addr_in_pic_d; // @[lsu_dccm_ctl.scala 271:35]
  assign io_lsu_pic_picm_mken = _T_1864 & io_addr_in_pic_d; // @[lsu_dccm_ctl.scala 272:35]
  assign io_lsu_pic_picm_rdaddr = 32'hf00c0000 | _T_1868; // @[lsu_dccm_ctl.scala 273:35]
  assign io_lsu_pic_picm_wraddr = 32'hf00c0000 | _T_1875; // @[lsu_dccm_ctl.scala 274:35]
  assign io_lsu_pic_picm_wr_data = io_dma_pic_wen ? io_dma_dccm_ctl_dma_mem_wdata[31:0] : io_store_datafn_lo_r; // @[lsu_dccm_ctl.scala 276:35]
  assign rvclkhdr_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_io_en = io_ld_single_ecc_error_r; // @[lib.scala 371:17]
  assign rvclkhdr_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_1_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_1_io_en = io_ld_single_ecc_error_r; // @[lib.scala 371:17]
  assign rvclkhdr_1_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  _T_2 = _RAND_0[63:0];
  _RAND_1 = {1{`RANDOM}};
  lsu_double_ecc_error_r_ff = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  ld_single_ecc_error_hi_r_ff = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  ld_single_ecc_error_lo_r_ff = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  ld_sec_addr_hi_r_ff = _RAND_4[15:0];
  _RAND_5 = {1{`RANDOM}};
  ld_sec_addr_lo_r_ff = _RAND_5[15:0];
  _RAND_6 = {1{`RANDOM}};
  _T_1173 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  _T_1379 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  _T_1882 = _RAND_8[0:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    _T_2 = 64'h0;
  end
  if (reset) begin
    lsu_double_ecc_error_r_ff = 1'h0;
  end
  if (reset) begin
    ld_single_ecc_error_hi_r_ff = 1'h0;
  end
  if (reset) begin
    ld_single_ecc_error_lo_r_ff = 1'h0;
  end
  if (reset) begin
    ld_sec_addr_hi_r_ff = 16'h0;
  end
  if (reset) begin
    ld_sec_addr_lo_r_ff = 16'h0;
  end
  if (reset) begin
    _T_1173 = 32'h0;
  end
  if (reset) begin
    _T_1379 = 32'h0;
  end
  if (reset) begin
    _T_1882 = 1'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge io_lsu_c2_r_clk or posedge reset) begin
    if (reset) begin
      _T_2 <= 64'h0;
    end else begin
      _T_2 <= lsu_rdata_corr_m >> _T_762;
    end
  end
  always @(posedge io_lsu_free_c2_clk or posedge reset) begin
    if (reset) begin
      lsu_double_ecc_error_r_ff <= 1'h0;
    end else begin
      lsu_double_ecc_error_r_ff <= io_lsu_double_ecc_error_r;
    end
  end
  always @(posedge io_lsu_free_c2_clk or posedge reset) begin
    if (reset) begin
      ld_single_ecc_error_hi_r_ff <= 1'h0;
    end else begin
      ld_single_ecc_error_hi_r_ff <= _T_822 & _T_823;
    end
  end
  always @(posedge io_lsu_free_c2_clk or posedge reset) begin
    if (reset) begin
      ld_single_ecc_error_lo_r_ff <= 1'h0;
    end else begin
      ld_single_ecc_error_lo_r_ff <= _T_819 & _T_820;
    end
  end
  always @(posedge rvclkhdr_io_l1clk or posedge reset) begin
    if (reset) begin
      ld_sec_addr_hi_r_ff <= 16'h0;
    end else begin
      ld_sec_addr_hi_r_ff <= io_end_addr_r;
    end
  end
  always @(posedge rvclkhdr_1_io_l1clk or posedge reset) begin
    if (reset) begin
      ld_sec_addr_lo_r_ff <= 16'h0;
    end else begin
      ld_sec_addr_lo_r_ff <= io_lsu_addr_r[15:0];
    end
  end
  always @(posedge io_lsu_store_c1_r_clk or posedge reset) begin
    if (reset) begin
      _T_1173 <= 32'h0;
    end else begin
      _T_1173 <= _T_1167 | _T_1171;
    end
  end
  always @(posedge io_lsu_store_c1_r_clk or posedge reset) begin
    if (reset) begin
      _T_1379 <= 32'h0;
    end else begin
      _T_1379 <= _T_1373 | _T_1377;
    end
  end
  always @(posedge io_lsu_c2_m_clk or posedge reset) begin
    if (reset) begin
      _T_1882 <= 1'h0;
    end else begin
      _T_1882 <= _T_837 & io_addr_in_dccm_d;
    end
  end
endmodule
module lsu_stbuf(
  input         clock,
  input         reset,
  input         io_lsu_c1_m_clk,
  input         io_lsu_c1_r_clk,
  input         io_lsu_stbuf_c1_clk,
  input         io_lsu_free_c2_clk,
  input         io_lsu_pkt_m_valid,
  input         io_lsu_pkt_m_bits_store,
  input         io_lsu_pkt_m_bits_dma,
  input         io_lsu_pkt_r_valid,
  input         io_lsu_pkt_r_bits_by,
  input         io_lsu_pkt_r_bits_half,
  input         io_lsu_pkt_r_bits_word,
  input         io_lsu_pkt_r_bits_dword,
  input         io_lsu_pkt_r_bits_store,
  input         io_lsu_pkt_r_bits_dma,
  input         io_store_stbuf_reqvld_r,
  input         io_lsu_commit_r,
  input         io_dec_lsu_valid_raw_d,
  input  [31:0] io_store_data_hi_r,
  input  [31:0] io_store_data_lo_r,
  input  [31:0] io_store_datafn_hi_r,
  input  [31:0] io_store_datafn_lo_r,
  input         io_lsu_stbuf_commit_any,
  input  [15:0] io_lsu_addr_d,
  input  [31:0] io_lsu_addr_m,
  input  [31:0] io_lsu_addr_r,
  input  [15:0] io_end_addr_d,
  input  [31:0] io_end_addr_m,
  input  [31:0] io_end_addr_r,
  input         io_addr_in_dccm_m,
  input         io_addr_in_dccm_r,
  input         io_scan_mode,
  output        io_stbuf_reqvld_any,
  output        io_stbuf_reqvld_flushed_any,
  output [15:0] io_stbuf_addr_any,
  output [31:0] io_stbuf_data_any,
  output        io_lsu_stbuf_full_any,
  output        io_lsu_stbuf_empty_any,
  output        io_ldst_stbuf_reqvld_r,
  output [31:0] io_stbuf_fwddata_hi_m,
  output [31:0] io_stbuf_fwddata_lo_m,
  output [3:0]  io_stbuf_fwdbyteen_hi_m,
  output [3:0]  io_stbuf_fwdbyteen_lo_m
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
`endif // RANDOMIZE_REG_INIT
  wire  rvclkhdr_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_1_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_1_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_1_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_1_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_2_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_2_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_2_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_2_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_3_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_3_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_3_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_3_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_4_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_4_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_4_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_4_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_5_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_5_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_5_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_5_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_6_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_6_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_6_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_6_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_7_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_7_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_7_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_7_io_scan_mode; // @[lib.scala 368:23]
  wire [1:0] _T_5 = io_lsu_pkt_r_bits_half ? 2'h3 : 2'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_6 = io_lsu_pkt_r_bits_word ? 4'hf : 4'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_7 = io_lsu_pkt_r_bits_dword ? 8'hff : 8'h0; // @[Mux.scala 27:72]
  wire [1:0] _GEN_10 = {{1'd0}, io_lsu_pkt_r_bits_by}; // @[Mux.scala 27:72]
  wire [1:0] _T_8 = _GEN_10 | _T_5; // @[Mux.scala 27:72]
  wire [3:0] _GEN_11 = {{2'd0}, _T_8}; // @[Mux.scala 27:72]
  wire [3:0] _T_9 = _GEN_11 | _T_6; // @[Mux.scala 27:72]
  wire [7:0] _GEN_12 = {{4'd0}, _T_9}; // @[Mux.scala 27:72]
  wire [7:0] ldst_byteen_r = _GEN_12 | _T_7; // @[Mux.scala 27:72]
  wire  ldst_dual_d = io_lsu_addr_d[2] != io_end_addr_d[2]; // @[lsu_stbuf.scala 117:39]
  reg  ldst_dual_r; // @[lsu_stbuf.scala 171:52]
  wire  dual_stbuf_write_r = ldst_dual_r & io_store_stbuf_reqvld_r; // @[lsu_stbuf.scala 118:40]
  wire [10:0] _GEN_13 = {{3'd0}, ldst_byteen_r}; // @[lsu_stbuf.scala 120:39]
  wire [10:0] _T_14 = _GEN_13 << io_lsu_addr_r[1:0]; // @[lsu_stbuf.scala 120:39]
  wire [7:0] store_byteen_ext_r = _T_14[7:0]; // @[lsu_stbuf.scala 120:22]
  wire [3:0] _T_17 = io_lsu_pkt_r_bits_store ? 4'hf : 4'h0; // @[Bitwise.scala 72:12]
  wire [3:0] store_byteen_hi_r = store_byteen_ext_r[7:4] & _T_17; // @[lsu_stbuf.scala 121:52]
  wire [3:0] store_byteen_lo_r = store_byteen_ext_r[3:0] & _T_17; // @[lsu_stbuf.scala 122:52]
  reg [1:0] RdPtr; // @[Reg.scala 27:20]
  wire [1:0] RdPtrPlus1 = RdPtr + 2'h1; // @[lsu_stbuf.scala 124:26]
  reg [1:0] WrPtr; // @[Reg.scala 27:20]
  wire [1:0] WrPtrPlus1 = WrPtr + 2'h1; // @[lsu_stbuf.scala 125:26]
  wire [1:0] WrPtrPlus2 = WrPtr + 2'h2; // @[lsu_stbuf.scala 126:26]
  reg [15:0] stbuf_addr_0; // @[lib.scala 374:16]
  wire  _T_27 = stbuf_addr_0[15:2] == io_lsu_addr_r[15:2]; // @[lsu_stbuf.scala 130:120]
  reg  _T_588; // @[lsu_stbuf.scala 163:88]
  reg  _T_580; // @[lsu_stbuf.scala 163:88]
  reg  _T_572; // @[lsu_stbuf.scala 163:88]
  reg  _T_564; // @[lsu_stbuf.scala 163:88]
  wire [3:0] stbuf_vld = {_T_588,_T_580,_T_572,_T_564}; // @[Cat.scala 29:58]
  wire  _T_29 = _T_27 & stbuf_vld[0]; // @[lsu_stbuf.scala 130:179]
  reg  _T_623; // @[lsu_stbuf.scala 164:92]
  reg  _T_615; // @[lsu_stbuf.scala 164:92]
  reg  _T_607; // @[lsu_stbuf.scala 164:92]
  reg  _T_599; // @[lsu_stbuf.scala 164:92]
  wire [3:0] stbuf_dma_kill = {_T_623,_T_615,_T_607,_T_599}; // @[Cat.scala 29:58]
  wire  _T_31 = ~stbuf_dma_kill[0]; // @[lsu_stbuf.scala 130:197]
  wire  _T_32 = _T_29 & _T_31; // @[lsu_stbuf.scala 130:195]
  wire  _T_212 = io_lsu_stbuf_commit_any | io_stbuf_reqvld_flushed_any; // @[lsu_stbuf.scala 141:78]
  wire  _T_213 = 2'h3 == RdPtr; // @[lsu_stbuf.scala 141:121]
  wire  _T_215 = _T_212 & _T_213; // @[lsu_stbuf.scala 141:109]
  wire  _T_209 = 2'h2 == RdPtr; // @[lsu_stbuf.scala 141:121]
  wire  _T_211 = _T_212 & _T_209; // @[lsu_stbuf.scala 141:109]
  wire  _T_205 = 2'h1 == RdPtr; // @[lsu_stbuf.scala 141:121]
  wire  _T_207 = _T_212 & _T_205; // @[lsu_stbuf.scala 141:109]
  wire  _T_201 = 2'h0 == RdPtr; // @[lsu_stbuf.scala 141:121]
  wire  _T_203 = _T_212 & _T_201; // @[lsu_stbuf.scala 141:109]
  wire [3:0] stbuf_reset = {_T_215,_T_211,_T_207,_T_203}; // @[Cat.scala 29:58]
  wire  _T_34 = ~stbuf_reset[0]; // @[lsu_stbuf.scala 130:218]
  wire  _T_35 = _T_32 & _T_34; // @[lsu_stbuf.scala 130:216]
  reg [15:0] stbuf_addr_1; // @[lib.scala 374:16]
  wire  _T_38 = stbuf_addr_1[15:2] == io_lsu_addr_r[15:2]; // @[lsu_stbuf.scala 130:120]
  wire  _T_40 = _T_38 & stbuf_vld[1]; // @[lsu_stbuf.scala 130:179]
  wire  _T_42 = ~stbuf_dma_kill[1]; // @[lsu_stbuf.scala 130:197]
  wire  _T_43 = _T_40 & _T_42; // @[lsu_stbuf.scala 130:195]
  wire  _T_45 = ~stbuf_reset[1]; // @[lsu_stbuf.scala 130:218]
  wire  _T_46 = _T_43 & _T_45; // @[lsu_stbuf.scala 130:216]
  reg [15:0] stbuf_addr_2; // @[lib.scala 374:16]
  wire  _T_49 = stbuf_addr_2[15:2] == io_lsu_addr_r[15:2]; // @[lsu_stbuf.scala 130:120]
  wire  _T_51 = _T_49 & stbuf_vld[2]; // @[lsu_stbuf.scala 130:179]
  wire  _T_53 = ~stbuf_dma_kill[2]; // @[lsu_stbuf.scala 130:197]
  wire  _T_54 = _T_51 & _T_53; // @[lsu_stbuf.scala 130:195]
  wire  _T_56 = ~stbuf_reset[2]; // @[lsu_stbuf.scala 130:218]
  wire  _T_57 = _T_54 & _T_56; // @[lsu_stbuf.scala 130:216]
  reg [15:0] stbuf_addr_3; // @[lib.scala 374:16]
  wire  _T_60 = stbuf_addr_3[15:2] == io_lsu_addr_r[15:2]; // @[lsu_stbuf.scala 130:120]
  wire  _T_62 = _T_60 & stbuf_vld[3]; // @[lsu_stbuf.scala 130:179]
  wire  _T_64 = ~stbuf_dma_kill[3]; // @[lsu_stbuf.scala 130:197]
  wire  _T_65 = _T_62 & _T_64; // @[lsu_stbuf.scala 130:195]
  wire  _T_67 = ~stbuf_reset[3]; // @[lsu_stbuf.scala 130:218]
  wire  _T_68 = _T_65 & _T_67; // @[lsu_stbuf.scala 130:216]
  wire [3:0] store_matchvec_lo_r = {_T_68,_T_57,_T_46,_T_35}; // @[Cat.scala 29:58]
  wire  _T_73 = stbuf_addr_0[15:2] == io_end_addr_r[15:2]; // @[lsu_stbuf.scala 131:120]
  wire  _T_75 = _T_73 & stbuf_vld[0]; // @[lsu_stbuf.scala 131:179]
  wire  _T_78 = _T_75 & _T_31; // @[lsu_stbuf.scala 131:194]
  wire  _T_79 = _T_78 & dual_stbuf_write_r; // @[lsu_stbuf.scala 131:215]
  wire  _T_82 = _T_79 & _T_34; // @[lsu_stbuf.scala 131:236]
  wire  _T_85 = stbuf_addr_1[15:2] == io_end_addr_r[15:2]; // @[lsu_stbuf.scala 131:120]
  wire  _T_87 = _T_85 & stbuf_vld[1]; // @[lsu_stbuf.scala 131:179]
  wire  _T_90 = _T_87 & _T_42; // @[lsu_stbuf.scala 131:194]
  wire  _T_91 = _T_90 & dual_stbuf_write_r; // @[lsu_stbuf.scala 131:215]
  wire  _T_94 = _T_91 & _T_45; // @[lsu_stbuf.scala 131:236]
  wire  _T_97 = stbuf_addr_2[15:2] == io_end_addr_r[15:2]; // @[lsu_stbuf.scala 131:120]
  wire  _T_99 = _T_97 & stbuf_vld[2]; // @[lsu_stbuf.scala 131:179]
  wire  _T_102 = _T_99 & _T_53; // @[lsu_stbuf.scala 131:194]
  wire  _T_103 = _T_102 & dual_stbuf_write_r; // @[lsu_stbuf.scala 131:215]
  wire  _T_106 = _T_103 & _T_56; // @[lsu_stbuf.scala 131:236]
  wire  _T_109 = stbuf_addr_3[15:2] == io_end_addr_r[15:2]; // @[lsu_stbuf.scala 131:120]
  wire  _T_111 = _T_109 & stbuf_vld[3]; // @[lsu_stbuf.scala 131:179]
  wire  _T_114 = _T_111 & _T_64; // @[lsu_stbuf.scala 131:194]
  wire  _T_115 = _T_114 & dual_stbuf_write_r; // @[lsu_stbuf.scala 131:215]
  wire  _T_118 = _T_115 & _T_67; // @[lsu_stbuf.scala 131:236]
  wire [3:0] store_matchvec_hi_r = {_T_118,_T_106,_T_94,_T_82}; // @[Cat.scala 29:58]
  wire  store_coalesce_lo_r = |store_matchvec_lo_r; // @[lsu_stbuf.scala 133:49]
  wire  store_coalesce_hi_r = |store_matchvec_hi_r; // @[lsu_stbuf.scala 134:49]
  wire  _T_121 = 2'h0 == WrPtr; // @[lsu_stbuf.scala 137:16]
  wire  _T_122 = ~store_coalesce_lo_r; // @[lsu_stbuf.scala 137:29]
  wire  _T_123 = _T_121 & _T_122; // @[lsu_stbuf.scala 137:27]
  wire  _T_125 = _T_121 & dual_stbuf_write_r; // @[lsu_stbuf.scala 138:29]
  wire  _T_126 = ~store_coalesce_hi_r; // @[lsu_stbuf.scala 138:52]
  wire  _T_127 = _T_125 & _T_126; // @[lsu_stbuf.scala 138:50]
  wire  _T_128 = _T_123 | _T_127; // @[lsu_stbuf.scala 137:51]
  wire  _T_129 = 2'h0 == WrPtrPlus1; // @[lsu_stbuf.scala 139:18]
  wire  _T_130 = _T_129 & dual_stbuf_write_r; // @[lsu_stbuf.scala 139:34]
  wire  _T_131 = store_coalesce_lo_r | store_coalesce_hi_r; // @[lsu_stbuf.scala 139:79]
  wire  _T_132 = ~_T_131; // @[lsu_stbuf.scala 139:57]
  wire  _T_133 = _T_130 & _T_132; // @[lsu_stbuf.scala 139:55]
  wire  _T_134 = _T_128 | _T_133; // @[lsu_stbuf.scala 138:74]
  wire  _T_136 = _T_134 | store_matchvec_lo_r[0]; // @[lsu_stbuf.scala 139:103]
  wire  _T_138 = _T_136 | store_matchvec_hi_r[0]; // @[lsu_stbuf.scala 140:30]
  wire  _T_139 = io_ldst_stbuf_reqvld_r & _T_138; // @[lsu_stbuf.scala 136:76]
  wire  _T_140 = 2'h1 == WrPtr; // @[lsu_stbuf.scala 137:16]
  wire  _T_142 = _T_140 & _T_122; // @[lsu_stbuf.scala 137:27]
  wire  _T_144 = _T_140 & dual_stbuf_write_r; // @[lsu_stbuf.scala 138:29]
  wire  _T_146 = _T_144 & _T_126; // @[lsu_stbuf.scala 138:50]
  wire  _T_147 = _T_142 | _T_146; // @[lsu_stbuf.scala 137:51]
  wire  _T_148 = 2'h1 == WrPtrPlus1; // @[lsu_stbuf.scala 139:18]
  wire  _T_149 = _T_148 & dual_stbuf_write_r; // @[lsu_stbuf.scala 139:34]
  wire  _T_152 = _T_149 & _T_132; // @[lsu_stbuf.scala 139:55]
  wire  _T_153 = _T_147 | _T_152; // @[lsu_stbuf.scala 138:74]
  wire  _T_155 = _T_153 | store_matchvec_lo_r[1]; // @[lsu_stbuf.scala 139:103]
  wire  _T_157 = _T_155 | store_matchvec_hi_r[1]; // @[lsu_stbuf.scala 140:30]
  wire  _T_158 = io_ldst_stbuf_reqvld_r & _T_157; // @[lsu_stbuf.scala 136:76]
  wire  _T_159 = 2'h2 == WrPtr; // @[lsu_stbuf.scala 137:16]
  wire  _T_161 = _T_159 & _T_122; // @[lsu_stbuf.scala 137:27]
  wire  _T_163 = _T_159 & dual_stbuf_write_r; // @[lsu_stbuf.scala 138:29]
  wire  _T_165 = _T_163 & _T_126; // @[lsu_stbuf.scala 138:50]
  wire  _T_166 = _T_161 | _T_165; // @[lsu_stbuf.scala 137:51]
  wire  _T_167 = 2'h2 == WrPtrPlus1; // @[lsu_stbuf.scala 139:18]
  wire  _T_168 = _T_167 & dual_stbuf_write_r; // @[lsu_stbuf.scala 139:34]
  wire  _T_171 = _T_168 & _T_132; // @[lsu_stbuf.scala 139:55]
  wire  _T_172 = _T_166 | _T_171; // @[lsu_stbuf.scala 138:74]
  wire  _T_174 = _T_172 | store_matchvec_lo_r[2]; // @[lsu_stbuf.scala 139:103]
  wire  _T_176 = _T_174 | store_matchvec_hi_r[2]; // @[lsu_stbuf.scala 140:30]
  wire  _T_177 = io_ldst_stbuf_reqvld_r & _T_176; // @[lsu_stbuf.scala 136:76]
  wire  _T_178 = 2'h3 == WrPtr; // @[lsu_stbuf.scala 137:16]
  wire  _T_180 = _T_178 & _T_122; // @[lsu_stbuf.scala 137:27]
  wire  _T_182 = _T_178 & dual_stbuf_write_r; // @[lsu_stbuf.scala 138:29]
  wire  _T_184 = _T_182 & _T_126; // @[lsu_stbuf.scala 138:50]
  wire  _T_185 = _T_180 | _T_184; // @[lsu_stbuf.scala 137:51]
  wire  _T_186 = 2'h3 == WrPtrPlus1; // @[lsu_stbuf.scala 139:18]
  wire  _T_187 = _T_186 & dual_stbuf_write_r; // @[lsu_stbuf.scala 139:34]
  wire  _T_190 = _T_187 & _T_132; // @[lsu_stbuf.scala 139:55]
  wire  _T_191 = _T_185 | _T_190; // @[lsu_stbuf.scala 138:74]
  wire  _T_193 = _T_191 | store_matchvec_lo_r[3]; // @[lsu_stbuf.scala 139:103]
  wire  _T_195 = _T_193 | store_matchvec_hi_r[3]; // @[lsu_stbuf.scala 140:30]
  wire  _T_196 = io_ldst_stbuf_reqvld_r & _T_195; // @[lsu_stbuf.scala 136:76]
  wire [3:0] stbuf_wr_en = {_T_196,_T_177,_T_158,_T_139}; // @[Cat.scala 29:58]
  wire  _T_219 = ~ldst_dual_r; // @[lsu_stbuf.scala 142:53]
  wire  _T_220 = _T_219 | io_store_stbuf_reqvld_r; // @[lsu_stbuf.scala 142:66]
  wire  _T_223 = _T_220 & _T_121; // @[lsu_stbuf.scala 142:93]
  wire  _T_225 = _T_223 & _T_122; // @[lsu_stbuf.scala 142:123]
  wire  _T_227 = _T_225 | store_matchvec_lo_r[0]; // @[lsu_stbuf.scala 142:147]
  wire  _T_232 = _T_220 & _T_140; // @[lsu_stbuf.scala 142:93]
  wire  _T_234 = _T_232 & _T_122; // @[lsu_stbuf.scala 142:123]
  wire  _T_236 = _T_234 | store_matchvec_lo_r[1]; // @[lsu_stbuf.scala 142:147]
  wire  _T_241 = _T_220 & _T_159; // @[lsu_stbuf.scala 142:93]
  wire  _T_243 = _T_241 & _T_122; // @[lsu_stbuf.scala 142:123]
  wire  _T_245 = _T_243 | store_matchvec_lo_r[2]; // @[lsu_stbuf.scala 142:147]
  wire  _T_250 = _T_220 & _T_178; // @[lsu_stbuf.scala 142:93]
  wire  _T_252 = _T_250 & _T_122; // @[lsu_stbuf.scala 142:123]
  wire  _T_254 = _T_252 | store_matchvec_lo_r[3]; // @[lsu_stbuf.scala 142:147]
  wire [3:0] sel_lo = {_T_254,_T_245,_T_236,_T_227}; // @[Cat.scala 29:58]
  reg [3:0] stbuf_byteen_0; // @[lsu_stbuf.scala 165:92]
  wire [3:0] _T_274 = stbuf_byteen_0 | store_byteen_lo_r; // @[lsu_stbuf.scala 145:86]
  wire [3:0] _T_275 = stbuf_byteen_0 | store_byteen_hi_r; // @[lsu_stbuf.scala 145:123]
  wire [3:0] stbuf_byteenin_0 = sel_lo[0] ? _T_274 : _T_275; // @[lsu_stbuf.scala 145:58]
  reg [3:0] stbuf_byteen_1; // @[lsu_stbuf.scala 165:92]
  wire [3:0] _T_278 = stbuf_byteen_1 | store_byteen_lo_r; // @[lsu_stbuf.scala 145:86]
  wire [3:0] _T_279 = stbuf_byteen_1 | store_byteen_hi_r; // @[lsu_stbuf.scala 145:123]
  wire [3:0] stbuf_byteenin_1 = sel_lo[1] ? _T_278 : _T_279; // @[lsu_stbuf.scala 145:58]
  reg [3:0] stbuf_byteen_2; // @[lsu_stbuf.scala 165:92]
  wire [3:0] _T_282 = stbuf_byteen_2 | store_byteen_lo_r; // @[lsu_stbuf.scala 145:86]
  wire [3:0] _T_283 = stbuf_byteen_2 | store_byteen_hi_r; // @[lsu_stbuf.scala 145:123]
  wire [3:0] stbuf_byteenin_2 = sel_lo[2] ? _T_282 : _T_283; // @[lsu_stbuf.scala 145:58]
  reg [3:0] stbuf_byteen_3; // @[lsu_stbuf.scala 165:92]
  wire [3:0] _T_286 = stbuf_byteen_3 | store_byteen_lo_r; // @[lsu_stbuf.scala 145:86]
  wire [3:0] _T_287 = stbuf_byteen_3 | store_byteen_hi_r; // @[lsu_stbuf.scala 145:123]
  wire [3:0] stbuf_byteenin_3 = sel_lo[3] ? _T_286 : _T_287; // @[lsu_stbuf.scala 145:58]
  wire  _T_291 = ~stbuf_byteen_0[0]; // @[lsu_stbuf.scala 147:67]
  wire  _T_293 = _T_291 | store_byteen_lo_r[0]; // @[lsu_stbuf.scala 147:87]
  reg [31:0] stbuf_data_0; // @[lib.scala 374:16]
  wire [7:0] _T_296 = _T_293 ? io_store_datafn_lo_r[7:0] : stbuf_data_0[7:0]; // @[lsu_stbuf.scala 147:66]
  wire  _T_300 = _T_291 | store_byteen_hi_r[0]; // @[lsu_stbuf.scala 148:29]
  wire [7:0] _T_303 = _T_300 ? io_store_datafn_hi_r[7:0] : stbuf_data_0[7:0]; // @[lsu_stbuf.scala 148:8]
  wire [7:0] datain1_0 = sel_lo[0] ? _T_296 : _T_303; // @[lsu_stbuf.scala 147:51]
  wire  _T_307 = ~stbuf_byteen_1[0]; // @[lsu_stbuf.scala 147:67]
  wire  _T_309 = _T_307 | store_byteen_lo_r[0]; // @[lsu_stbuf.scala 147:87]
  reg [31:0] stbuf_data_1; // @[lib.scala 374:16]
  wire [7:0] _T_312 = _T_309 ? io_store_datafn_lo_r[7:0] : stbuf_data_1[7:0]; // @[lsu_stbuf.scala 147:66]
  wire  _T_316 = _T_307 | store_byteen_hi_r[0]; // @[lsu_stbuf.scala 148:29]
  wire [7:0] _T_319 = _T_316 ? io_store_datafn_hi_r[7:0] : stbuf_data_1[7:0]; // @[lsu_stbuf.scala 148:8]
  wire [7:0] datain1_1 = sel_lo[1] ? _T_312 : _T_319; // @[lsu_stbuf.scala 147:51]
  wire  _T_323 = ~stbuf_byteen_2[0]; // @[lsu_stbuf.scala 147:67]
  wire  _T_325 = _T_323 | store_byteen_lo_r[0]; // @[lsu_stbuf.scala 147:87]
  reg [31:0] stbuf_data_2; // @[lib.scala 374:16]
  wire [7:0] _T_328 = _T_325 ? io_store_datafn_lo_r[7:0] : stbuf_data_2[7:0]; // @[lsu_stbuf.scala 147:66]
  wire  _T_332 = _T_323 | store_byteen_hi_r[0]; // @[lsu_stbuf.scala 148:29]
  wire [7:0] _T_335 = _T_332 ? io_store_datafn_hi_r[7:0] : stbuf_data_2[7:0]; // @[lsu_stbuf.scala 148:8]
  wire [7:0] datain1_2 = sel_lo[2] ? _T_328 : _T_335; // @[lsu_stbuf.scala 147:51]
  wire  _T_339 = ~stbuf_byteen_3[0]; // @[lsu_stbuf.scala 147:67]
  wire  _T_341 = _T_339 | store_byteen_lo_r[0]; // @[lsu_stbuf.scala 147:87]
  reg [31:0] stbuf_data_3; // @[lib.scala 374:16]
  wire [7:0] _T_344 = _T_341 ? io_store_datafn_lo_r[7:0] : stbuf_data_3[7:0]; // @[lsu_stbuf.scala 147:66]
  wire  _T_348 = _T_339 | store_byteen_hi_r[0]; // @[lsu_stbuf.scala 148:29]
  wire [7:0] _T_351 = _T_348 ? io_store_datafn_hi_r[7:0] : stbuf_data_3[7:0]; // @[lsu_stbuf.scala 148:8]
  wire [7:0] datain1_3 = sel_lo[3] ? _T_344 : _T_351; // @[lsu_stbuf.scala 147:51]
  wire  _T_355 = ~stbuf_byteen_0[1]; // @[lsu_stbuf.scala 150:68]
  wire  _T_357 = _T_355 | store_byteen_lo_r[1]; // @[lsu_stbuf.scala 150:88]
  wire [7:0] _T_360 = _T_357 ? io_store_datafn_lo_r[15:8] : stbuf_data_0[15:8]; // @[lsu_stbuf.scala 150:67]
  wire  _T_364 = _T_355 | store_byteen_hi_r[1]; // @[lsu_stbuf.scala 151:29]
  wire [7:0] _T_367 = _T_364 ? io_store_datafn_hi_r[15:8] : stbuf_data_0[15:8]; // @[lsu_stbuf.scala 151:8]
  wire [7:0] datain2_0 = sel_lo[0] ? _T_360 : _T_367; // @[lsu_stbuf.scala 150:52]
  wire  _T_371 = ~stbuf_byteen_1[1]; // @[lsu_stbuf.scala 150:68]
  wire  _T_373 = _T_371 | store_byteen_lo_r[1]; // @[lsu_stbuf.scala 150:88]
  wire [7:0] _T_376 = _T_373 ? io_store_datafn_lo_r[15:8] : stbuf_data_1[15:8]; // @[lsu_stbuf.scala 150:67]
  wire  _T_380 = _T_371 | store_byteen_hi_r[1]; // @[lsu_stbuf.scala 151:29]
  wire [7:0] _T_383 = _T_380 ? io_store_datafn_hi_r[15:8] : stbuf_data_1[15:8]; // @[lsu_stbuf.scala 151:8]
  wire [7:0] datain2_1 = sel_lo[1] ? _T_376 : _T_383; // @[lsu_stbuf.scala 150:52]
  wire  _T_387 = ~stbuf_byteen_2[1]; // @[lsu_stbuf.scala 150:68]
  wire  _T_389 = _T_387 | store_byteen_lo_r[1]; // @[lsu_stbuf.scala 150:88]
  wire [7:0] _T_392 = _T_389 ? io_store_datafn_lo_r[15:8] : stbuf_data_2[15:8]; // @[lsu_stbuf.scala 150:67]
  wire  _T_396 = _T_387 | store_byteen_hi_r[1]; // @[lsu_stbuf.scala 151:29]
  wire [7:0] _T_399 = _T_396 ? io_store_datafn_hi_r[15:8] : stbuf_data_2[15:8]; // @[lsu_stbuf.scala 151:8]
  wire [7:0] datain2_2 = sel_lo[2] ? _T_392 : _T_399; // @[lsu_stbuf.scala 150:52]
  wire  _T_403 = ~stbuf_byteen_3[1]; // @[lsu_stbuf.scala 150:68]
  wire  _T_405 = _T_403 | store_byteen_lo_r[1]; // @[lsu_stbuf.scala 150:88]
  wire [7:0] _T_408 = _T_405 ? io_store_datafn_lo_r[15:8] : stbuf_data_3[15:8]; // @[lsu_stbuf.scala 150:67]
  wire  _T_412 = _T_403 | store_byteen_hi_r[1]; // @[lsu_stbuf.scala 151:29]
  wire [7:0] _T_415 = _T_412 ? io_store_datafn_hi_r[15:8] : stbuf_data_3[15:8]; // @[lsu_stbuf.scala 151:8]
  wire [7:0] datain2_3 = sel_lo[3] ? _T_408 : _T_415; // @[lsu_stbuf.scala 150:52]
  wire  _T_419 = ~stbuf_byteen_0[2]; // @[lsu_stbuf.scala 153:68]
  wire  _T_421 = _T_419 | store_byteen_lo_r[2]; // @[lsu_stbuf.scala 153:88]
  wire [7:0] _T_424 = _T_421 ? io_store_datafn_lo_r[23:16] : stbuf_data_0[23:16]; // @[lsu_stbuf.scala 153:67]
  wire  _T_428 = _T_419 | store_byteen_hi_r[2]; // @[lsu_stbuf.scala 154:29]
  wire [7:0] _T_431 = _T_428 ? io_store_datafn_hi_r[23:16] : stbuf_data_0[23:16]; // @[lsu_stbuf.scala 154:8]
  wire [7:0] datain3_0 = sel_lo[0] ? _T_424 : _T_431; // @[lsu_stbuf.scala 153:52]
  wire  _T_435 = ~stbuf_byteen_1[2]; // @[lsu_stbuf.scala 153:68]
  wire  _T_437 = _T_435 | store_byteen_lo_r[2]; // @[lsu_stbuf.scala 153:88]
  wire [7:0] _T_440 = _T_437 ? io_store_datafn_lo_r[23:16] : stbuf_data_1[23:16]; // @[lsu_stbuf.scala 153:67]
  wire  _T_444 = _T_435 | store_byteen_hi_r[2]; // @[lsu_stbuf.scala 154:29]
  wire [7:0] _T_447 = _T_444 ? io_store_datafn_hi_r[23:16] : stbuf_data_1[23:16]; // @[lsu_stbuf.scala 154:8]
  wire [7:0] datain3_1 = sel_lo[1] ? _T_440 : _T_447; // @[lsu_stbuf.scala 153:52]
  wire  _T_451 = ~stbuf_byteen_2[2]; // @[lsu_stbuf.scala 153:68]
  wire  _T_453 = _T_451 | store_byteen_lo_r[2]; // @[lsu_stbuf.scala 153:88]
  wire [7:0] _T_456 = _T_453 ? io_store_datafn_lo_r[23:16] : stbuf_data_2[23:16]; // @[lsu_stbuf.scala 153:67]
  wire  _T_460 = _T_451 | store_byteen_hi_r[2]; // @[lsu_stbuf.scala 154:29]
  wire [7:0] _T_463 = _T_460 ? io_store_datafn_hi_r[23:16] : stbuf_data_2[23:16]; // @[lsu_stbuf.scala 154:8]
  wire [7:0] datain3_2 = sel_lo[2] ? _T_456 : _T_463; // @[lsu_stbuf.scala 153:52]
  wire  _T_467 = ~stbuf_byteen_3[2]; // @[lsu_stbuf.scala 153:68]
  wire  _T_469 = _T_467 | store_byteen_lo_r[2]; // @[lsu_stbuf.scala 153:88]
  wire [7:0] _T_472 = _T_469 ? io_store_datafn_lo_r[23:16] : stbuf_data_3[23:16]; // @[lsu_stbuf.scala 153:67]
  wire  _T_476 = _T_467 | store_byteen_hi_r[2]; // @[lsu_stbuf.scala 154:29]
  wire [7:0] _T_479 = _T_476 ? io_store_datafn_hi_r[23:16] : stbuf_data_3[23:16]; // @[lsu_stbuf.scala 154:8]
  wire [7:0] datain3_3 = sel_lo[3] ? _T_472 : _T_479; // @[lsu_stbuf.scala 153:52]
  wire  _T_483 = ~stbuf_byteen_0[3]; // @[lsu_stbuf.scala 156:68]
  wire  _T_485 = _T_483 | store_byteen_lo_r[3]; // @[lsu_stbuf.scala 156:88]
  wire [7:0] _T_488 = _T_485 ? io_store_datafn_lo_r[31:24] : stbuf_data_0[31:24]; // @[lsu_stbuf.scala 156:67]
  wire  _T_492 = _T_483 | store_byteen_hi_r[3]; // @[lsu_stbuf.scala 157:29]
  wire [7:0] _T_495 = _T_492 ? io_store_datafn_hi_r[31:24] : stbuf_data_0[31:24]; // @[lsu_stbuf.scala 157:8]
  wire [7:0] datain4_0 = sel_lo[0] ? _T_488 : _T_495; // @[lsu_stbuf.scala 156:52]
  wire  _T_499 = ~stbuf_byteen_1[3]; // @[lsu_stbuf.scala 156:68]
  wire  _T_501 = _T_499 | store_byteen_lo_r[3]; // @[lsu_stbuf.scala 156:88]
  wire [7:0] _T_504 = _T_501 ? io_store_datafn_lo_r[31:24] : stbuf_data_1[31:24]; // @[lsu_stbuf.scala 156:67]
  wire  _T_508 = _T_499 | store_byteen_hi_r[3]; // @[lsu_stbuf.scala 157:29]
  wire [7:0] _T_511 = _T_508 ? io_store_datafn_hi_r[31:24] : stbuf_data_1[31:24]; // @[lsu_stbuf.scala 157:8]
  wire [7:0] datain4_1 = sel_lo[1] ? _T_504 : _T_511; // @[lsu_stbuf.scala 156:52]
  wire  _T_515 = ~stbuf_byteen_2[3]; // @[lsu_stbuf.scala 156:68]
  wire  _T_517 = _T_515 | store_byteen_lo_r[3]; // @[lsu_stbuf.scala 156:88]
  wire [7:0] _T_520 = _T_517 ? io_store_datafn_lo_r[31:24] : stbuf_data_2[31:24]; // @[lsu_stbuf.scala 156:67]
  wire  _T_524 = _T_515 | store_byteen_hi_r[3]; // @[lsu_stbuf.scala 157:29]
  wire [7:0] _T_527 = _T_524 ? io_store_datafn_hi_r[31:24] : stbuf_data_2[31:24]; // @[lsu_stbuf.scala 157:8]
  wire [7:0] datain4_2 = sel_lo[2] ? _T_520 : _T_527; // @[lsu_stbuf.scala 156:52]
  wire  _T_531 = ~stbuf_byteen_3[3]; // @[lsu_stbuf.scala 156:68]
  wire  _T_533 = _T_531 | store_byteen_lo_r[3]; // @[lsu_stbuf.scala 156:88]
  wire [7:0] _T_536 = _T_533 ? io_store_datafn_lo_r[31:24] : stbuf_data_3[31:24]; // @[lsu_stbuf.scala 156:67]
  wire  _T_540 = _T_531 | store_byteen_hi_r[3]; // @[lsu_stbuf.scala 157:29]
  wire [7:0] _T_543 = _T_540 ? io_store_datafn_hi_r[31:24] : stbuf_data_3[31:24]; // @[lsu_stbuf.scala 157:8]
  wire [7:0] datain4_3 = sel_lo[3] ? _T_536 : _T_543; // @[lsu_stbuf.scala 156:52]
  wire [15:0] _T_545 = {datain2_0,datain1_0}; // @[Cat.scala 29:58]
  wire [15:0] _T_546 = {datain4_0,datain3_0}; // @[Cat.scala 29:58]
  wire [15:0] _T_548 = {datain2_1,datain1_1}; // @[Cat.scala 29:58]
  wire [15:0] _T_549 = {datain4_1,datain3_1}; // @[Cat.scala 29:58]
  wire [15:0] _T_551 = {datain2_2,datain1_2}; // @[Cat.scala 29:58]
  wire [15:0] _T_552 = {datain4_2,datain3_2}; // @[Cat.scala 29:58]
  wire [15:0] _T_554 = {datain2_3,datain1_3}; // @[Cat.scala 29:58]
  wire [15:0] _T_555 = {datain4_3,datain3_3}; // @[Cat.scala 29:58]
  wire  _T_560 = stbuf_wr_en[0] | stbuf_vld[0]; // @[lsu_stbuf.scala 163:92]
  wire  _T_568 = stbuf_wr_en[1] | stbuf_vld[1]; // @[lsu_stbuf.scala 163:92]
  wire  _T_576 = stbuf_wr_en[2] | stbuf_vld[2]; // @[lsu_stbuf.scala 163:92]
  wire  _T_584 = stbuf_wr_en[3] | stbuf_vld[3]; // @[lsu_stbuf.scala 163:92]
  wire [15:0] cmpaddr_hi_m = {{2'd0}, io_end_addr_m[15:2]}; // @[lsu_stbuf.scala 200:16]
  wire  _T_789 = stbuf_addr_3[15:2] == cmpaddr_hi_m[13:0]; // @[lsu_stbuf.scala 206:115]
  wire  _T_791 = _T_789 & stbuf_vld[3]; // @[lsu_stbuf.scala 206:139]
  wire  _T_794 = _T_791 & _T_64; // @[lsu_stbuf.scala 206:154]
  wire  _T_795 = _T_794 & io_addr_in_dccm_m; // @[lsu_stbuf.scala 206:175]
  wire  _T_780 = stbuf_addr_2[15:2] == cmpaddr_hi_m[13:0]; // @[lsu_stbuf.scala 206:115]
  wire  _T_782 = _T_780 & stbuf_vld[2]; // @[lsu_stbuf.scala 206:139]
  wire  _T_785 = _T_782 & _T_53; // @[lsu_stbuf.scala 206:154]
  wire  _T_786 = _T_785 & io_addr_in_dccm_m; // @[lsu_stbuf.scala 206:175]
  wire  _T_771 = stbuf_addr_1[15:2] == cmpaddr_hi_m[13:0]; // @[lsu_stbuf.scala 206:115]
  wire  _T_773 = _T_771 & stbuf_vld[1]; // @[lsu_stbuf.scala 206:139]
  wire  _T_776 = _T_773 & _T_42; // @[lsu_stbuf.scala 206:154]
  wire  _T_777 = _T_776 & io_addr_in_dccm_m; // @[lsu_stbuf.scala 206:175]
  wire  _T_762 = stbuf_addr_0[15:2] == cmpaddr_hi_m[13:0]; // @[lsu_stbuf.scala 206:115]
  wire  _T_764 = _T_762 & stbuf_vld[0]; // @[lsu_stbuf.scala 206:139]
  wire  _T_767 = _T_764 & _T_31; // @[lsu_stbuf.scala 206:154]
  wire  _T_768 = _T_767 & io_addr_in_dccm_m; // @[lsu_stbuf.scala 206:175]
  wire [3:0] stbuf_match_hi = {_T_795,_T_786,_T_777,_T_768}; // @[Cat.scala 29:58]
  wire [15:0] cmpaddr_lo_m = {{2'd0}, io_lsu_addr_m[15:2]}; // @[lsu_stbuf.scala 203:17]
  wire  _T_827 = stbuf_addr_3[15:2] == cmpaddr_lo_m[13:0]; // @[lsu_stbuf.scala 207:115]
  wire  _T_829 = _T_827 & stbuf_vld[3]; // @[lsu_stbuf.scala 207:139]
  wire  _T_832 = _T_829 & _T_64; // @[lsu_stbuf.scala 207:154]
  wire  _T_833 = _T_832 & io_addr_in_dccm_m; // @[lsu_stbuf.scala 207:175]
  wire  _T_818 = stbuf_addr_2[15:2] == cmpaddr_lo_m[13:0]; // @[lsu_stbuf.scala 207:115]
  wire  _T_820 = _T_818 & stbuf_vld[2]; // @[lsu_stbuf.scala 207:139]
  wire  _T_823 = _T_820 & _T_53; // @[lsu_stbuf.scala 207:154]
  wire  _T_824 = _T_823 & io_addr_in_dccm_m; // @[lsu_stbuf.scala 207:175]
  wire  _T_809 = stbuf_addr_1[15:2] == cmpaddr_lo_m[13:0]; // @[lsu_stbuf.scala 207:115]
  wire  _T_811 = _T_809 & stbuf_vld[1]; // @[lsu_stbuf.scala 207:139]
  wire  _T_814 = _T_811 & _T_42; // @[lsu_stbuf.scala 207:154]
  wire  _T_815 = _T_814 & io_addr_in_dccm_m; // @[lsu_stbuf.scala 207:175]
  wire  _T_800 = stbuf_addr_0[15:2] == cmpaddr_lo_m[13:0]; // @[lsu_stbuf.scala 207:115]
  wire  _T_802 = _T_800 & stbuf_vld[0]; // @[lsu_stbuf.scala 207:139]
  wire  _T_805 = _T_802 & _T_31; // @[lsu_stbuf.scala 207:154]
  wire  _T_806 = _T_805 & io_addr_in_dccm_m; // @[lsu_stbuf.scala 207:175]
  wire [3:0] stbuf_match_lo = {_T_833,_T_824,_T_815,_T_806}; // @[Cat.scala 29:58]
  wire  _T_856 = stbuf_match_hi[3] | stbuf_match_lo[3]; // @[lsu_stbuf.scala 208:78]
  wire  _T_857 = _T_856 & io_lsu_pkt_m_valid; // @[lsu_stbuf.scala 208:99]
  wire  _T_858 = _T_857 & io_lsu_pkt_m_bits_dma; // @[lsu_stbuf.scala 208:120]
  wire  _T_859 = _T_858 & io_lsu_pkt_m_bits_store; // @[lsu_stbuf.scala 208:144]
  wire  _T_850 = stbuf_match_hi[2] | stbuf_match_lo[2]; // @[lsu_stbuf.scala 208:78]
  wire  _T_851 = _T_850 & io_lsu_pkt_m_valid; // @[lsu_stbuf.scala 208:99]
  wire  _T_852 = _T_851 & io_lsu_pkt_m_bits_dma; // @[lsu_stbuf.scala 208:120]
  wire  _T_853 = _T_852 & io_lsu_pkt_m_bits_store; // @[lsu_stbuf.scala 208:144]
  wire  _T_844 = stbuf_match_hi[1] | stbuf_match_lo[1]; // @[lsu_stbuf.scala 208:78]
  wire  _T_845 = _T_844 & io_lsu_pkt_m_valid; // @[lsu_stbuf.scala 208:99]
  wire  _T_846 = _T_845 & io_lsu_pkt_m_bits_dma; // @[lsu_stbuf.scala 208:120]
  wire  _T_847 = _T_846 & io_lsu_pkt_m_bits_store; // @[lsu_stbuf.scala 208:144]
  wire  _T_838 = stbuf_match_hi[0] | stbuf_match_lo[0]; // @[lsu_stbuf.scala 208:78]
  wire  _T_839 = _T_838 & io_lsu_pkt_m_valid; // @[lsu_stbuf.scala 208:99]
  wire  _T_840 = _T_839 & io_lsu_pkt_m_bits_dma; // @[lsu_stbuf.scala 208:120]
  wire  _T_841 = _T_840 & io_lsu_pkt_m_bits_store; // @[lsu_stbuf.scala 208:144]
  wire [3:0] stbuf_dma_kill_en = {_T_859,_T_853,_T_847,_T_841}; // @[Cat.scala 29:58]
  wire  _T_595 = stbuf_dma_kill_en[0] | stbuf_dma_kill[0]; // @[lsu_stbuf.scala 164:96]
  wire  _T_603 = stbuf_dma_kill_en[1] | stbuf_dma_kill[1]; // @[lsu_stbuf.scala 164:96]
  wire  _T_611 = stbuf_dma_kill_en[2] | stbuf_dma_kill[2]; // @[lsu_stbuf.scala 164:96]
  wire  _T_619 = stbuf_dma_kill_en[3] | stbuf_dma_kill[3]; // @[lsu_stbuf.scala 164:96]
  wire [3:0] _T_629 = stbuf_wr_en[0] ? stbuf_byteenin_0 : stbuf_byteen_0; // @[lsu_stbuf.scala 165:96]
  wire [3:0] _T_633 = _T_34 ? 4'hf : 4'h0; // @[Bitwise.scala 72:12]
  wire [3:0] _T_638 = stbuf_wr_en[1] ? stbuf_byteenin_1 : stbuf_byteen_1; // @[lsu_stbuf.scala 165:96]
  wire [3:0] _T_642 = _T_45 ? 4'hf : 4'h0; // @[Bitwise.scala 72:12]
  wire [3:0] _T_647 = stbuf_wr_en[2] ? stbuf_byteenin_2 : stbuf_byteen_2; // @[lsu_stbuf.scala 165:96]
  wire [3:0] _T_651 = _T_56 ? 4'hf : 4'h0; // @[Bitwise.scala 72:12]
  wire [3:0] _T_656 = stbuf_wr_en[3] ? stbuf_byteenin_3 : stbuf_byteen_3; // @[lsu_stbuf.scala 165:96]
  wire [3:0] _T_660 = _T_67 ? 4'hf : 4'h0; // @[Bitwise.scala 72:12]
  reg  ldst_dual_m; // @[lsu_stbuf.scala 170:52]
  wire [3:0] _T_689 = stbuf_vld >> RdPtr; // @[lsu_stbuf.scala 174:43]
  wire [3:0] _T_691 = stbuf_dma_kill >> RdPtr; // @[lsu_stbuf.scala 174:67]
  wire  _T_698 = ~_T_691[0]; // @[lsu_stbuf.scala 175:46]
  wire  _T_699 = _T_689[0] & _T_698; // @[lsu_stbuf.scala 175:44]
  wire  _T_700 = |stbuf_dma_kill_en; // @[lsu_stbuf.scala 175:91]
  wire  _T_701 = ~_T_700; // @[lsu_stbuf.scala 175:71]
  wire [15:0] _GEN_1 = 2'h1 == RdPtr ? stbuf_addr_1 : stbuf_addr_0; // @[lsu_stbuf.scala 176:22]
  wire [15:0] _GEN_2 = 2'h2 == RdPtr ? stbuf_addr_2 : _GEN_1; // @[lsu_stbuf.scala 176:22]
  wire [31:0] _GEN_5 = 2'h1 == RdPtr ? stbuf_data_1 : stbuf_data_0; // @[lsu_stbuf.scala 177:22]
  wire [31:0] _GEN_6 = 2'h2 == RdPtr ? stbuf_data_2 : _GEN_5; // @[lsu_stbuf.scala 177:22]
  wire  _T_703 = ~dual_stbuf_write_r; // @[lsu_stbuf.scala 179:44]
  wire  _T_704 = io_ldst_stbuf_reqvld_r & _T_703; // @[lsu_stbuf.scala 179:42]
  wire  _T_705 = store_coalesce_hi_r | store_coalesce_lo_r; // @[lsu_stbuf.scala 179:88]
  wire  _T_706 = ~_T_705; // @[lsu_stbuf.scala 179:66]
  wire  _T_707 = _T_704 & _T_706; // @[lsu_stbuf.scala 179:64]
  wire  _T_708 = io_ldst_stbuf_reqvld_r & dual_stbuf_write_r; // @[lsu_stbuf.scala 180:30]
  wire  _T_709 = store_coalesce_hi_r & store_coalesce_lo_r; // @[lsu_stbuf.scala 180:76]
  wire  _T_710 = ~_T_709; // @[lsu_stbuf.scala 180:54]
  wire  _T_711 = _T_708 & _T_710; // @[lsu_stbuf.scala 180:52]
  wire  WrPtrEn = _T_707 | _T_711; // @[lsu_stbuf.scala 179:113]
  wire  _T_716 = _T_708 & _T_706; // @[lsu_stbuf.scala 181:67]
  wire [3:0] _T_721 = {3'h0,stbuf_vld[0]}; // @[Cat.scala 29:58]
  wire [3:0] _T_723 = {3'h0,stbuf_vld[1]}; // @[Cat.scala 29:58]
  wire [3:0] _T_725 = {3'h0,stbuf_vld[2]}; // @[Cat.scala 29:58]
  wire [3:0] _T_727 = {3'h0,stbuf_vld[3]}; // @[Cat.scala 29:58]
  wire [3:0] _T_730 = _T_721 + _T_723; // @[lsu_stbuf.scala 188:101]
  wire [3:0] _T_732 = _T_730 + _T_725; // @[lsu_stbuf.scala 188:101]
  wire [3:0] stbuf_numvld_any = _T_732 + _T_727; // @[lsu_stbuf.scala 188:101]
  wire  _T_734 = io_lsu_pkt_m_valid & io_lsu_pkt_m_bits_store; // @[lsu_stbuf.scala 189:39]
  wire  _T_735 = _T_734 & io_addr_in_dccm_m; // @[lsu_stbuf.scala 189:65]
  wire  _T_736 = ~io_lsu_pkt_m_bits_dma; // @[lsu_stbuf.scala 189:87]
  wire  isdccmst_m = _T_735 & _T_736; // @[lsu_stbuf.scala 189:85]
  wire  _T_737 = io_lsu_pkt_r_valid & io_lsu_pkt_r_bits_store; // @[lsu_stbuf.scala 190:39]
  wire  _T_738 = _T_737 & io_addr_in_dccm_r; // @[lsu_stbuf.scala 190:65]
  wire  _T_739 = ~io_lsu_pkt_r_bits_dma; // @[lsu_stbuf.scala 190:87]
  wire  isdccmst_r = _T_738 & _T_739; // @[lsu_stbuf.scala 190:85]
  wire [1:0] _T_740 = {1'h0,isdccmst_m}; // @[Cat.scala 29:58]
  wire  _T_741 = isdccmst_m & ldst_dual_m; // @[lsu_stbuf.scala 192:62]
  wire [2:0] _GEN_14 = {{1'd0}, _T_740}; // @[lsu_stbuf.scala 192:47]
  wire [2:0] _T_742 = _GEN_14 << _T_741; // @[lsu_stbuf.scala 192:47]
  wire [1:0] _T_743 = {1'h0,isdccmst_r}; // @[Cat.scala 29:58]
  wire  _T_744 = isdccmst_r & ldst_dual_r; // @[lsu_stbuf.scala 193:62]
  wire [2:0] _GEN_15 = {{1'd0}, _T_743}; // @[lsu_stbuf.scala 193:47]
  wire [2:0] _T_745 = _GEN_15 << _T_744; // @[lsu_stbuf.scala 193:47]
  wire [1:0] stbuf_specvld_m = _T_742[1:0]; // @[lsu_stbuf.scala 192:19]
  wire [3:0] _T_746 = {2'h0,stbuf_specvld_m}; // @[Cat.scala 29:58]
  wire [3:0] _T_748 = stbuf_numvld_any + _T_746; // @[lsu_stbuf.scala 194:44]
  wire [1:0] stbuf_specvld_r = _T_745[1:0]; // @[lsu_stbuf.scala 193:19]
  wire [3:0] _T_749 = {2'h0,stbuf_specvld_r}; // @[Cat.scala 29:58]
  wire [3:0] stbuf_specvld_any = _T_748 + _T_749; // @[lsu_stbuf.scala 194:78]
  wire  _T_751 = ~ldst_dual_d; // @[lsu_stbuf.scala 196:34]
  wire  _T_752 = _T_751 & io_dec_lsu_valid_raw_d; // @[lsu_stbuf.scala 196:47]
  wire  _T_754 = stbuf_specvld_any >= 4'h4; // @[lsu_stbuf.scala 196:99]
  wire  _T_755 = stbuf_specvld_any >= 4'h3; // @[lsu_stbuf.scala 196:140]
  wire  _T_865 = stbuf_match_hi[0] & stbuf_byteen_0[0]; // @[lsu_stbuf.scala 211:116]
  wire  stbuf_fwdbyteenvec_hi_0_0 = _T_865 & stbuf_vld[0]; // @[lsu_stbuf.scala 211:137]
  wire  _T_869 = stbuf_match_hi[0] & stbuf_byteen_0[1]; // @[lsu_stbuf.scala 211:116]
  wire  stbuf_fwdbyteenvec_hi_0_1 = _T_869 & stbuf_vld[0]; // @[lsu_stbuf.scala 211:137]
  wire  _T_873 = stbuf_match_hi[0] & stbuf_byteen_0[2]; // @[lsu_stbuf.scala 211:116]
  wire  stbuf_fwdbyteenvec_hi_0_2 = _T_873 & stbuf_vld[0]; // @[lsu_stbuf.scala 211:137]
  wire  _T_877 = stbuf_match_hi[0] & stbuf_byteen_0[3]; // @[lsu_stbuf.scala 211:116]
  wire  stbuf_fwdbyteenvec_hi_0_3 = _T_877 & stbuf_vld[0]; // @[lsu_stbuf.scala 211:137]
  wire  _T_881 = stbuf_match_hi[1] & stbuf_byteen_1[0]; // @[lsu_stbuf.scala 211:116]
  wire  stbuf_fwdbyteenvec_hi_1_0 = _T_881 & stbuf_vld[1]; // @[lsu_stbuf.scala 211:137]
  wire  _T_885 = stbuf_match_hi[1] & stbuf_byteen_1[1]; // @[lsu_stbuf.scala 211:116]
  wire  stbuf_fwdbyteenvec_hi_1_1 = _T_885 & stbuf_vld[1]; // @[lsu_stbuf.scala 211:137]
  wire  _T_889 = stbuf_match_hi[1] & stbuf_byteen_1[2]; // @[lsu_stbuf.scala 211:116]
  wire  stbuf_fwdbyteenvec_hi_1_2 = _T_889 & stbuf_vld[1]; // @[lsu_stbuf.scala 211:137]
  wire  _T_893 = stbuf_match_hi[1] & stbuf_byteen_1[3]; // @[lsu_stbuf.scala 211:116]
  wire  stbuf_fwdbyteenvec_hi_1_3 = _T_893 & stbuf_vld[1]; // @[lsu_stbuf.scala 211:137]
  wire  _T_897 = stbuf_match_hi[2] & stbuf_byteen_2[0]; // @[lsu_stbuf.scala 211:116]
  wire  stbuf_fwdbyteenvec_hi_2_0 = _T_897 & stbuf_vld[2]; // @[lsu_stbuf.scala 211:137]
  wire  _T_901 = stbuf_match_hi[2] & stbuf_byteen_2[1]; // @[lsu_stbuf.scala 211:116]
  wire  stbuf_fwdbyteenvec_hi_2_1 = _T_901 & stbuf_vld[2]; // @[lsu_stbuf.scala 211:137]
  wire  _T_905 = stbuf_match_hi[2] & stbuf_byteen_2[2]; // @[lsu_stbuf.scala 211:116]
  wire  stbuf_fwdbyteenvec_hi_2_2 = _T_905 & stbuf_vld[2]; // @[lsu_stbuf.scala 211:137]
  wire  _T_909 = stbuf_match_hi[2] & stbuf_byteen_2[3]; // @[lsu_stbuf.scala 211:116]
  wire  stbuf_fwdbyteenvec_hi_2_3 = _T_909 & stbuf_vld[2]; // @[lsu_stbuf.scala 211:137]
  wire  _T_913 = stbuf_match_hi[3] & stbuf_byteen_3[0]; // @[lsu_stbuf.scala 211:116]
  wire  stbuf_fwdbyteenvec_hi_3_0 = _T_913 & stbuf_vld[3]; // @[lsu_stbuf.scala 211:137]
  wire  _T_917 = stbuf_match_hi[3] & stbuf_byteen_3[1]; // @[lsu_stbuf.scala 211:116]
  wire  stbuf_fwdbyteenvec_hi_3_1 = _T_917 & stbuf_vld[3]; // @[lsu_stbuf.scala 211:137]
  wire  _T_921 = stbuf_match_hi[3] & stbuf_byteen_3[2]; // @[lsu_stbuf.scala 211:116]
  wire  stbuf_fwdbyteenvec_hi_3_2 = _T_921 & stbuf_vld[3]; // @[lsu_stbuf.scala 211:137]
  wire  _T_925 = stbuf_match_hi[3] & stbuf_byteen_3[3]; // @[lsu_stbuf.scala 211:116]
  wire  stbuf_fwdbyteenvec_hi_3_3 = _T_925 & stbuf_vld[3]; // @[lsu_stbuf.scala 211:137]
  wire  _T_929 = stbuf_match_lo[0] & stbuf_byteen_0[0]; // @[lsu_stbuf.scala 212:116]
  wire  stbuf_fwdbyteenvec_lo_0_0 = _T_929 & stbuf_vld[0]; // @[lsu_stbuf.scala 212:137]
  wire  _T_933 = stbuf_match_lo[0] & stbuf_byteen_0[1]; // @[lsu_stbuf.scala 212:116]
  wire  stbuf_fwdbyteenvec_lo_0_1 = _T_933 & stbuf_vld[0]; // @[lsu_stbuf.scala 212:137]
  wire  _T_937 = stbuf_match_lo[0] & stbuf_byteen_0[2]; // @[lsu_stbuf.scala 212:116]
  wire  stbuf_fwdbyteenvec_lo_0_2 = _T_937 & stbuf_vld[0]; // @[lsu_stbuf.scala 212:137]
  wire  _T_941 = stbuf_match_lo[0] & stbuf_byteen_0[3]; // @[lsu_stbuf.scala 212:116]
  wire  stbuf_fwdbyteenvec_lo_0_3 = _T_941 & stbuf_vld[0]; // @[lsu_stbuf.scala 212:137]
  wire  _T_945 = stbuf_match_lo[1] & stbuf_byteen_1[0]; // @[lsu_stbuf.scala 212:116]
  wire  stbuf_fwdbyteenvec_lo_1_0 = _T_945 & stbuf_vld[1]; // @[lsu_stbuf.scala 212:137]
  wire  _T_949 = stbuf_match_lo[1] & stbuf_byteen_1[1]; // @[lsu_stbuf.scala 212:116]
  wire  stbuf_fwdbyteenvec_lo_1_1 = _T_949 & stbuf_vld[1]; // @[lsu_stbuf.scala 212:137]
  wire  _T_953 = stbuf_match_lo[1] & stbuf_byteen_1[2]; // @[lsu_stbuf.scala 212:116]
  wire  stbuf_fwdbyteenvec_lo_1_2 = _T_953 & stbuf_vld[1]; // @[lsu_stbuf.scala 212:137]
  wire  _T_957 = stbuf_match_lo[1] & stbuf_byteen_1[3]; // @[lsu_stbuf.scala 212:116]
  wire  stbuf_fwdbyteenvec_lo_1_3 = _T_957 & stbuf_vld[1]; // @[lsu_stbuf.scala 212:137]
  wire  _T_961 = stbuf_match_lo[2] & stbuf_byteen_2[0]; // @[lsu_stbuf.scala 212:116]
  wire  stbuf_fwdbyteenvec_lo_2_0 = _T_961 & stbuf_vld[2]; // @[lsu_stbuf.scala 212:137]
  wire  _T_965 = stbuf_match_lo[2] & stbuf_byteen_2[1]; // @[lsu_stbuf.scala 212:116]
  wire  stbuf_fwdbyteenvec_lo_2_1 = _T_965 & stbuf_vld[2]; // @[lsu_stbuf.scala 212:137]
  wire  _T_969 = stbuf_match_lo[2] & stbuf_byteen_2[2]; // @[lsu_stbuf.scala 212:116]
  wire  stbuf_fwdbyteenvec_lo_2_2 = _T_969 & stbuf_vld[2]; // @[lsu_stbuf.scala 212:137]
  wire  _T_973 = stbuf_match_lo[2] & stbuf_byteen_2[3]; // @[lsu_stbuf.scala 212:116]
  wire  stbuf_fwdbyteenvec_lo_2_3 = _T_973 & stbuf_vld[2]; // @[lsu_stbuf.scala 212:137]
  wire  _T_977 = stbuf_match_lo[3] & stbuf_byteen_3[0]; // @[lsu_stbuf.scala 212:116]
  wire  stbuf_fwdbyteenvec_lo_3_0 = _T_977 & stbuf_vld[3]; // @[lsu_stbuf.scala 212:137]
  wire  _T_981 = stbuf_match_lo[3] & stbuf_byteen_3[1]; // @[lsu_stbuf.scala 212:116]
  wire  stbuf_fwdbyteenvec_lo_3_1 = _T_981 & stbuf_vld[3]; // @[lsu_stbuf.scala 212:137]
  wire  _T_985 = stbuf_match_lo[3] & stbuf_byteen_3[2]; // @[lsu_stbuf.scala 212:116]
  wire  stbuf_fwdbyteenvec_lo_3_2 = _T_985 & stbuf_vld[3]; // @[lsu_stbuf.scala 212:137]
  wire  _T_989 = stbuf_match_lo[3] & stbuf_byteen_3[3]; // @[lsu_stbuf.scala 212:116]
  wire  stbuf_fwdbyteenvec_lo_3_3 = _T_989 & stbuf_vld[3]; // @[lsu_stbuf.scala 212:137]
  wire  _T_991 = stbuf_fwdbyteenvec_hi_0_0 | stbuf_fwdbyteenvec_hi_1_0; // @[lsu_stbuf.scala 213:147]
  wire  _T_992 = _T_991 | stbuf_fwdbyteenvec_hi_2_0; // @[lsu_stbuf.scala 213:147]
  wire  stbuf_fwdbyteen_hi_pre_m_0 = _T_992 | stbuf_fwdbyteenvec_hi_3_0; // @[lsu_stbuf.scala 213:147]
  wire  _T_993 = stbuf_fwdbyteenvec_hi_0_1 | stbuf_fwdbyteenvec_hi_1_1; // @[lsu_stbuf.scala 213:147]
  wire  _T_994 = _T_993 | stbuf_fwdbyteenvec_hi_2_1; // @[lsu_stbuf.scala 213:147]
  wire  stbuf_fwdbyteen_hi_pre_m_1 = _T_994 | stbuf_fwdbyteenvec_hi_3_1; // @[lsu_stbuf.scala 213:147]
  wire  _T_995 = stbuf_fwdbyteenvec_hi_0_2 | stbuf_fwdbyteenvec_hi_1_2; // @[lsu_stbuf.scala 213:147]
  wire  _T_996 = _T_995 | stbuf_fwdbyteenvec_hi_2_2; // @[lsu_stbuf.scala 213:147]
  wire  stbuf_fwdbyteen_hi_pre_m_2 = _T_996 | stbuf_fwdbyteenvec_hi_3_2; // @[lsu_stbuf.scala 213:147]
  wire  _T_997 = stbuf_fwdbyteenvec_hi_0_3 | stbuf_fwdbyteenvec_hi_1_3; // @[lsu_stbuf.scala 213:147]
  wire  _T_998 = _T_997 | stbuf_fwdbyteenvec_hi_2_3; // @[lsu_stbuf.scala 213:147]
  wire  stbuf_fwdbyteen_hi_pre_m_3 = _T_998 | stbuf_fwdbyteenvec_hi_3_3; // @[lsu_stbuf.scala 213:147]
  wire  _T_999 = stbuf_fwdbyteenvec_lo_0_0 | stbuf_fwdbyteenvec_lo_1_0; // @[lsu_stbuf.scala 214:147]
  wire  _T_1000 = _T_999 | stbuf_fwdbyteenvec_lo_2_0; // @[lsu_stbuf.scala 214:147]
  wire  stbuf_fwdbyteen_lo_pre_m_0 = _T_1000 | stbuf_fwdbyteenvec_lo_3_0; // @[lsu_stbuf.scala 214:147]
  wire  _T_1001 = stbuf_fwdbyteenvec_lo_0_1 | stbuf_fwdbyteenvec_lo_1_1; // @[lsu_stbuf.scala 214:147]
  wire  _T_1002 = _T_1001 | stbuf_fwdbyteenvec_lo_2_1; // @[lsu_stbuf.scala 214:147]
  wire  stbuf_fwdbyteen_lo_pre_m_1 = _T_1002 | stbuf_fwdbyteenvec_lo_3_1; // @[lsu_stbuf.scala 214:147]
  wire  _T_1003 = stbuf_fwdbyteenvec_lo_0_2 | stbuf_fwdbyteenvec_lo_1_2; // @[lsu_stbuf.scala 214:147]
  wire  _T_1004 = _T_1003 | stbuf_fwdbyteenvec_lo_2_2; // @[lsu_stbuf.scala 214:147]
  wire  stbuf_fwdbyteen_lo_pre_m_2 = _T_1004 | stbuf_fwdbyteenvec_lo_3_2; // @[lsu_stbuf.scala 214:147]
  wire  _T_1005 = stbuf_fwdbyteenvec_lo_0_3 | stbuf_fwdbyteenvec_lo_1_3; // @[lsu_stbuf.scala 214:147]
  wire  _T_1006 = _T_1005 | stbuf_fwdbyteenvec_lo_2_3; // @[lsu_stbuf.scala 214:147]
  wire  stbuf_fwdbyteen_lo_pre_m_3 = _T_1006 | stbuf_fwdbyteenvec_lo_3_3; // @[lsu_stbuf.scala 214:147]
  wire [31:0] _T_1009 = stbuf_match_hi[0] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_1010 = _T_1009 & stbuf_data_0; // @[lsu_stbuf.scala 216:97]
  wire [31:0] _T_1013 = stbuf_match_hi[1] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_1014 = _T_1013 & stbuf_data_1; // @[lsu_stbuf.scala 216:97]
  wire [31:0] _T_1017 = stbuf_match_hi[2] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_1018 = _T_1017 & stbuf_data_2; // @[lsu_stbuf.scala 216:97]
  wire [31:0] _T_1021 = stbuf_match_hi[3] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_1022 = _T_1021 & stbuf_data_3; // @[lsu_stbuf.scala 216:97]
  wire [31:0] _T_1024 = _T_1022 | _T_1018; // @[lsu_stbuf.scala 216:130]
  wire [31:0] _T_1025 = _T_1024 | _T_1014; // @[lsu_stbuf.scala 216:130]
  wire [31:0] stbuf_fwddata_hi_pre_m = _T_1025 | _T_1010; // @[lsu_stbuf.scala 216:130]
  wire [31:0] _T_1028 = stbuf_match_lo[0] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_1029 = _T_1028 & stbuf_data_0; // @[lsu_stbuf.scala 217:97]
  wire [31:0] _T_1032 = stbuf_match_lo[1] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_1033 = _T_1032 & stbuf_data_1; // @[lsu_stbuf.scala 217:97]
  wire [31:0] _T_1036 = stbuf_match_lo[2] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_1037 = _T_1036 & stbuf_data_2; // @[lsu_stbuf.scala 217:97]
  wire [31:0] _T_1040 = stbuf_match_lo[3] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_1041 = _T_1040 & stbuf_data_3; // @[lsu_stbuf.scala 217:97]
  wire [31:0] _T_1043 = _T_1041 | _T_1037; // @[lsu_stbuf.scala 217:130]
  wire [31:0] _T_1044 = _T_1043 | _T_1033; // @[lsu_stbuf.scala 217:130]
  wire [31:0] stbuf_fwddata_lo_pre_m = _T_1044 | _T_1029; // @[lsu_stbuf.scala 217:130]
  wire  _T_1049 = io_lsu_addr_m[31:2] == io_lsu_addr_r[31:2]; // @[lsu_stbuf.scala 224:49]
  wire  _T_1050 = _T_1049 & io_lsu_pkt_r_valid; // @[lsu_stbuf.scala 224:74]
  wire  _T_1051 = _T_1050 & io_lsu_pkt_r_bits_store; // @[lsu_stbuf.scala 224:95]
  wire  ld_addr_rhit_lo_lo = _T_1051 & _T_739; // @[lsu_stbuf.scala 224:121]
  wire  _T_1055 = io_end_addr_m[31:2] == io_lsu_addr_r[31:2]; // @[lsu_stbuf.scala 225:49]
  wire  _T_1056 = _T_1055 & io_lsu_pkt_r_valid; // @[lsu_stbuf.scala 225:74]
  wire  _T_1057 = _T_1056 & io_lsu_pkt_r_bits_store; // @[lsu_stbuf.scala 225:95]
  wire  ld_addr_rhit_lo_hi = _T_1057 & _T_739; // @[lsu_stbuf.scala 225:121]
  wire  _T_1061 = io_lsu_addr_m[31:2] == io_end_addr_r[31:2]; // @[lsu_stbuf.scala 226:49]
  wire  _T_1062 = _T_1061 & io_lsu_pkt_r_valid; // @[lsu_stbuf.scala 226:74]
  wire  _T_1063 = _T_1062 & io_lsu_pkt_r_bits_store; // @[lsu_stbuf.scala 226:95]
  wire  _T_1065 = _T_1063 & _T_739; // @[lsu_stbuf.scala 226:121]
  wire  ld_addr_rhit_hi_lo = _T_1065 & dual_stbuf_write_r; // @[lsu_stbuf.scala 226:146]
  wire  _T_1068 = io_end_addr_m[31:2] == io_end_addr_r[31:2]; // @[lsu_stbuf.scala 227:49]
  wire  _T_1069 = _T_1068 & io_lsu_pkt_r_valid; // @[lsu_stbuf.scala 227:74]
  wire  _T_1070 = _T_1069 & io_lsu_pkt_r_bits_store; // @[lsu_stbuf.scala 227:95]
  wire  _T_1072 = _T_1070 & _T_739; // @[lsu_stbuf.scala 227:121]
  wire  ld_addr_rhit_hi_hi = _T_1072 & dual_stbuf_write_r; // @[lsu_stbuf.scala 227:146]
  wire  _T_1074 = ld_addr_rhit_lo_lo & store_byteen_ext_r[0]; // @[lsu_stbuf.scala 229:79]
  wire  _T_1076 = ld_addr_rhit_lo_lo & store_byteen_ext_r[1]; // @[lsu_stbuf.scala 229:79]
  wire  _T_1078 = ld_addr_rhit_lo_lo & store_byteen_ext_r[2]; // @[lsu_stbuf.scala 229:79]
  wire  _T_1080 = ld_addr_rhit_lo_lo & store_byteen_ext_r[3]; // @[lsu_stbuf.scala 229:79]
  wire [3:0] ld_byte_rhit_lo_lo = {_T_1080,_T_1078,_T_1076,_T_1074}; // @[Cat.scala 29:58]
  wire  _T_1085 = ld_addr_rhit_lo_hi & store_byteen_ext_r[0]; // @[lsu_stbuf.scala 230:79]
  wire  _T_1087 = ld_addr_rhit_lo_hi & store_byteen_ext_r[1]; // @[lsu_stbuf.scala 230:79]
  wire  _T_1089 = ld_addr_rhit_lo_hi & store_byteen_ext_r[2]; // @[lsu_stbuf.scala 230:79]
  wire  _T_1091 = ld_addr_rhit_lo_hi & store_byteen_ext_r[3]; // @[lsu_stbuf.scala 230:79]
  wire [3:0] ld_byte_rhit_lo_hi = {_T_1091,_T_1089,_T_1087,_T_1085}; // @[Cat.scala 29:58]
  wire  _T_1096 = ld_addr_rhit_hi_lo & store_byteen_ext_r[4]; // @[lsu_stbuf.scala 231:79]
  wire  _T_1098 = ld_addr_rhit_hi_lo & store_byteen_ext_r[5]; // @[lsu_stbuf.scala 231:79]
  wire  _T_1100 = ld_addr_rhit_hi_lo & store_byteen_ext_r[6]; // @[lsu_stbuf.scala 231:79]
  wire  _T_1102 = ld_addr_rhit_hi_lo & store_byteen_ext_r[7]; // @[lsu_stbuf.scala 231:79]
  wire [3:0] ld_byte_rhit_hi_lo = {_T_1102,_T_1100,_T_1098,_T_1096}; // @[Cat.scala 29:58]
  wire  _T_1107 = ld_addr_rhit_hi_hi & store_byteen_ext_r[4]; // @[lsu_stbuf.scala 232:79]
  wire  _T_1109 = ld_addr_rhit_hi_hi & store_byteen_ext_r[5]; // @[lsu_stbuf.scala 232:79]
  wire  _T_1111 = ld_addr_rhit_hi_hi & store_byteen_ext_r[6]; // @[lsu_stbuf.scala 232:79]
  wire  _T_1113 = ld_addr_rhit_hi_hi & store_byteen_ext_r[7]; // @[lsu_stbuf.scala 232:79]
  wire [3:0] ld_byte_rhit_hi_hi = {_T_1113,_T_1111,_T_1109,_T_1107}; // @[Cat.scala 29:58]
  wire  _T_1119 = ld_byte_rhit_lo_lo[0] | ld_byte_rhit_hi_lo[0]; // @[lsu_stbuf.scala 234:79]
  wire  _T_1122 = ld_byte_rhit_lo_lo[1] | ld_byte_rhit_hi_lo[1]; // @[lsu_stbuf.scala 234:79]
  wire  _T_1125 = ld_byte_rhit_lo_lo[2] | ld_byte_rhit_hi_lo[2]; // @[lsu_stbuf.scala 234:79]
  wire  _T_1128 = ld_byte_rhit_lo_lo[3] | ld_byte_rhit_hi_lo[3]; // @[lsu_stbuf.scala 234:79]
  wire [3:0] ld_byte_rhit_lo = {_T_1128,_T_1125,_T_1122,_T_1119}; // @[Cat.scala 29:58]
  wire  _T_1134 = ld_byte_rhit_lo_hi[0] | ld_byte_rhit_hi_hi[0]; // @[lsu_stbuf.scala 235:79]
  wire  _T_1137 = ld_byte_rhit_lo_hi[1] | ld_byte_rhit_hi_hi[1]; // @[lsu_stbuf.scala 235:79]
  wire  _T_1140 = ld_byte_rhit_lo_hi[2] | ld_byte_rhit_hi_hi[2]; // @[lsu_stbuf.scala 235:79]
  wire  _T_1143 = ld_byte_rhit_lo_hi[3] | ld_byte_rhit_hi_hi[3]; // @[lsu_stbuf.scala 235:79]
  wire [3:0] ld_byte_rhit_hi = {_T_1143,_T_1140,_T_1137,_T_1134}; // @[Cat.scala 29:58]
  wire [7:0] _T_1149 = ld_byte_rhit_lo_lo[0] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_1151 = _T_1149 & io_store_data_lo_r[7:0]; // @[lsu_stbuf.scala 237:53]
  wire [7:0] _T_1154 = ld_byte_rhit_hi_lo[0] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_1156 = _T_1154 & io_store_data_hi_r[7:0]; // @[lsu_stbuf.scala 237:114]
  wire [7:0] fwdpipe1_lo = _T_1151 | _T_1156; // @[lsu_stbuf.scala 237:80]
  wire [7:0] _T_1159 = ld_byte_rhit_lo_lo[1] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_1161 = _T_1159 & io_store_data_lo_r[15:8]; // @[lsu_stbuf.scala 238:53]
  wire [7:0] _T_1164 = ld_byte_rhit_hi_lo[1] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_1166 = _T_1164 & io_store_data_hi_r[15:8]; // @[lsu_stbuf.scala 238:115]
  wire [7:0] fwdpipe2_lo = _T_1161 | _T_1166; // @[lsu_stbuf.scala 238:81]
  wire [7:0] _T_1169 = ld_byte_rhit_lo_lo[2] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_1171 = _T_1169 & io_store_data_lo_r[23:16]; // @[lsu_stbuf.scala 239:53]
  wire [7:0] _T_1174 = ld_byte_rhit_hi_lo[2] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_1176 = _T_1174 & io_store_data_hi_r[23:16]; // @[lsu_stbuf.scala 239:116]
  wire [7:0] fwdpipe3_lo = _T_1171 | _T_1176; // @[lsu_stbuf.scala 239:82]
  wire [7:0] _T_1179 = ld_byte_rhit_lo_lo[3] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_1181 = _T_1179 & io_store_data_lo_r[31:24]; // @[lsu_stbuf.scala 240:53]
  wire [7:0] _T_1184 = ld_byte_rhit_hi_lo[3] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_1186 = _T_1184 & io_store_data_hi_r[31:24]; // @[lsu_stbuf.scala 240:116]
  wire [7:0] fwdpipe4_lo = _T_1181 | _T_1186; // @[lsu_stbuf.scala 240:82]
  wire [31:0] ld_fwddata_rpipe_lo = {fwdpipe4_lo,fwdpipe3_lo,fwdpipe2_lo,fwdpipe1_lo}; // @[Cat.scala 29:58]
  wire [7:0] _T_1192 = ld_byte_rhit_lo_hi[0] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_1194 = _T_1192 & io_store_data_lo_r[7:0]; // @[lsu_stbuf.scala 243:53]
  wire [7:0] _T_1197 = ld_byte_rhit_hi_hi[0] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_1199 = _T_1197 & io_store_data_hi_r[7:0]; // @[lsu_stbuf.scala 243:114]
  wire [7:0] fwdpipe1_hi = _T_1194 | _T_1199; // @[lsu_stbuf.scala 243:80]
  wire [7:0] _T_1202 = ld_byte_rhit_lo_hi[1] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_1204 = _T_1202 & io_store_data_lo_r[15:8]; // @[lsu_stbuf.scala 244:53]
  wire [7:0] _T_1207 = ld_byte_rhit_hi_hi[1] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_1209 = _T_1207 & io_store_data_hi_r[15:8]; // @[lsu_stbuf.scala 244:115]
  wire [7:0] fwdpipe2_hi = _T_1204 | _T_1209; // @[lsu_stbuf.scala 244:81]
  wire [7:0] _T_1212 = ld_byte_rhit_lo_hi[2] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_1214 = _T_1212 & io_store_data_lo_r[23:16]; // @[lsu_stbuf.scala 245:53]
  wire [7:0] _T_1217 = ld_byte_rhit_hi_hi[2] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_1219 = _T_1217 & io_store_data_hi_r[23:16]; // @[lsu_stbuf.scala 245:116]
  wire [7:0] fwdpipe3_hi = _T_1214 | _T_1219; // @[lsu_stbuf.scala 245:82]
  wire [7:0] _T_1222 = ld_byte_rhit_lo_hi[3] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_1224 = _T_1222 & io_store_data_lo_r[31:24]; // @[lsu_stbuf.scala 246:53]
  wire [7:0] _T_1227 = ld_byte_rhit_hi_hi[3] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_1229 = _T_1227 & io_store_data_hi_r[31:24]; // @[lsu_stbuf.scala 246:116]
  wire [7:0] fwdpipe4_hi = _T_1224 | _T_1229; // @[lsu_stbuf.scala 246:82]
  wire [31:0] ld_fwddata_rpipe_hi = {fwdpipe4_hi,fwdpipe3_hi,fwdpipe2_hi,fwdpipe1_hi}; // @[Cat.scala 29:58]
  wire  _T_1264 = ld_byte_rhit_hi[0] | stbuf_fwdbyteen_hi_pre_m_0; // @[lsu_stbuf.scala 252:83]
  wire  _T_1266 = ld_byte_rhit_hi[1] | stbuf_fwdbyteen_hi_pre_m_1; // @[lsu_stbuf.scala 252:83]
  wire  _T_1268 = ld_byte_rhit_hi[2] | stbuf_fwdbyteen_hi_pre_m_2; // @[lsu_stbuf.scala 252:83]
  wire  _T_1270 = ld_byte_rhit_hi[3] | stbuf_fwdbyteen_hi_pre_m_3; // @[lsu_stbuf.scala 252:83]
  wire [2:0] _T_1272 = {_T_1270,_T_1268,_T_1266}; // @[Cat.scala 29:58]
  wire  _T_1275 = ld_byte_rhit_lo[0] | stbuf_fwdbyteen_lo_pre_m_0; // @[lsu_stbuf.scala 253:83]
  wire  _T_1277 = ld_byte_rhit_lo[1] | stbuf_fwdbyteen_lo_pre_m_1; // @[lsu_stbuf.scala 253:83]
  wire  _T_1279 = ld_byte_rhit_lo[2] | stbuf_fwdbyteen_lo_pre_m_2; // @[lsu_stbuf.scala 253:83]
  wire  _T_1281 = ld_byte_rhit_lo[3] | stbuf_fwdbyteen_lo_pre_m_3; // @[lsu_stbuf.scala 253:83]
  wire [2:0] _T_1283 = {_T_1281,_T_1279,_T_1277}; // @[Cat.scala 29:58]
  wire [7:0] stbuf_fwdpipe1_lo = ld_byte_rhit_lo[0] ? ld_fwddata_rpipe_lo[7:0] : stbuf_fwddata_lo_pre_m[7:0]; // @[lsu_stbuf.scala 256:30]
  wire [7:0] stbuf_fwdpipe2_lo = ld_byte_rhit_lo[1] ? ld_fwddata_rpipe_lo[15:8] : stbuf_fwddata_lo_pre_m[15:8]; // @[lsu_stbuf.scala 257:30]
  wire [7:0] stbuf_fwdpipe3_lo = ld_byte_rhit_lo[2] ? ld_fwddata_rpipe_lo[23:16] : stbuf_fwddata_lo_pre_m[23:16]; // @[lsu_stbuf.scala 258:30]
  wire [7:0] stbuf_fwdpipe4_lo = ld_byte_rhit_lo[3] ? ld_fwddata_rpipe_lo[31:24] : stbuf_fwddata_lo_pre_m[31:24]; // @[lsu_stbuf.scala 259:30]
  wire [15:0] _T_1297 = {stbuf_fwdpipe2_lo,stbuf_fwdpipe1_lo}; // @[Cat.scala 29:58]
  wire [15:0] _T_1298 = {stbuf_fwdpipe4_lo,stbuf_fwdpipe3_lo}; // @[Cat.scala 29:58]
  wire [7:0] stbuf_fwdpipe1_hi = ld_byte_rhit_hi[0] ? ld_fwddata_rpipe_hi[7:0] : stbuf_fwddata_hi_pre_m[7:0]; // @[lsu_stbuf.scala 262:30]
  wire [7:0] stbuf_fwdpipe2_hi = ld_byte_rhit_hi[1] ? ld_fwddata_rpipe_hi[15:8] : stbuf_fwddata_hi_pre_m[15:8]; // @[lsu_stbuf.scala 263:30]
  wire [7:0] stbuf_fwdpipe3_hi = ld_byte_rhit_hi[2] ? ld_fwddata_rpipe_hi[23:16] : stbuf_fwddata_hi_pre_m[23:16]; // @[lsu_stbuf.scala 264:30]
  wire [7:0] stbuf_fwdpipe4_hi = ld_byte_rhit_hi[3] ? ld_fwddata_rpipe_hi[31:24] : stbuf_fwddata_hi_pre_m[31:24]; // @[lsu_stbuf.scala 265:30]
  wire [15:0] _T_1312 = {stbuf_fwdpipe2_hi,stbuf_fwdpipe1_hi}; // @[Cat.scala 29:58]
  wire [15:0] _T_1313 = {stbuf_fwdpipe4_hi,stbuf_fwdpipe3_hi}; // @[Cat.scala 29:58]
  rvclkhdr rvclkhdr ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_io_l1clk),
    .io_clk(rvclkhdr_io_clk),
    .io_en(rvclkhdr_io_en),
    .io_scan_mode(rvclkhdr_io_scan_mode)
  );
  rvclkhdr rvclkhdr_1 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_1_io_l1clk),
    .io_clk(rvclkhdr_1_io_clk),
    .io_en(rvclkhdr_1_io_en),
    .io_scan_mode(rvclkhdr_1_io_scan_mode)
  );
  rvclkhdr rvclkhdr_2 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_2_io_l1clk),
    .io_clk(rvclkhdr_2_io_clk),
    .io_en(rvclkhdr_2_io_en),
    .io_scan_mode(rvclkhdr_2_io_scan_mode)
  );
  rvclkhdr rvclkhdr_3 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_3_io_l1clk),
    .io_clk(rvclkhdr_3_io_clk),
    .io_en(rvclkhdr_3_io_en),
    .io_scan_mode(rvclkhdr_3_io_scan_mode)
  );
  rvclkhdr rvclkhdr_4 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_4_io_l1clk),
    .io_clk(rvclkhdr_4_io_clk),
    .io_en(rvclkhdr_4_io_en),
    .io_scan_mode(rvclkhdr_4_io_scan_mode)
  );
  rvclkhdr rvclkhdr_5 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_5_io_l1clk),
    .io_clk(rvclkhdr_5_io_clk),
    .io_en(rvclkhdr_5_io_en),
    .io_scan_mode(rvclkhdr_5_io_scan_mode)
  );
  rvclkhdr rvclkhdr_6 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_6_io_l1clk),
    .io_clk(rvclkhdr_6_io_clk),
    .io_en(rvclkhdr_6_io_en),
    .io_scan_mode(rvclkhdr_6_io_scan_mode)
  );
  rvclkhdr rvclkhdr_7 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_7_io_l1clk),
    .io_clk(rvclkhdr_7_io_clk),
    .io_en(rvclkhdr_7_io_en),
    .io_scan_mode(rvclkhdr_7_io_scan_mode)
  );
  assign io_stbuf_reqvld_any = _T_699 & _T_701; // @[lsu_stbuf.scala 51:47 lsu_stbuf.scala 175:24]
  assign io_stbuf_reqvld_flushed_any = _T_689[0] & _T_691[0]; // @[lsu_stbuf.scala 52:35 lsu_stbuf.scala 174:31]
  assign io_stbuf_addr_any = 2'h3 == RdPtr ? stbuf_addr_3 : _GEN_2; // @[lsu_stbuf.scala 53:35 lsu_stbuf.scala 176:22]
  assign io_stbuf_data_any = 2'h3 == RdPtr ? stbuf_data_3 : _GEN_6; // @[lsu_stbuf.scala 54:35 lsu_stbuf.scala 177:22]
  assign io_lsu_stbuf_full_any = _T_752 ? _T_754 : _T_755; // @[lsu_stbuf.scala 55:43 lsu_stbuf.scala 196:26]
  assign io_lsu_stbuf_empty_any = stbuf_numvld_any == 4'h0; // @[lsu_stbuf.scala 56:43 lsu_stbuf.scala 197:26]
  assign io_ldst_stbuf_reqvld_r = io_lsu_commit_r & io_store_stbuf_reqvld_r; // @[lsu_stbuf.scala 57:43 lsu_stbuf.scala 128:26]
  assign io_stbuf_fwddata_hi_m = {_T_1313,_T_1312}; // @[lsu_stbuf.scala 58:43 lsu_stbuf.scala 266:25]
  assign io_stbuf_fwddata_lo_m = {_T_1298,_T_1297}; // @[lsu_stbuf.scala 59:43 lsu_stbuf.scala 260:25]
  assign io_stbuf_fwdbyteen_hi_m = {_T_1272,_T_1264}; // @[lsu_stbuf.scala 60:37 lsu_stbuf.scala 252:27]
  assign io_stbuf_fwdbyteen_lo_m = {_T_1283,_T_1275}; // @[lsu_stbuf.scala 61:37 lsu_stbuf.scala 253:27]
  assign rvclkhdr_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_io_en = stbuf_wr_en[0]; // @[lib.scala 371:17]
  assign rvclkhdr_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_1_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_1_io_en = stbuf_wr_en[0]; // @[lib.scala 371:17]
  assign rvclkhdr_1_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_2_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_2_io_en = stbuf_wr_en[1]; // @[lib.scala 371:17]
  assign rvclkhdr_2_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_3_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_3_io_en = stbuf_wr_en[1]; // @[lib.scala 371:17]
  assign rvclkhdr_3_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_4_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_4_io_en = stbuf_wr_en[2]; // @[lib.scala 371:17]
  assign rvclkhdr_4_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_5_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_5_io_en = stbuf_wr_en[2]; // @[lib.scala 371:17]
  assign rvclkhdr_5_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_6_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_6_io_en = stbuf_wr_en[3]; // @[lib.scala 371:17]
  assign rvclkhdr_6_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_7_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_7_io_en = stbuf_wr_en[3]; // @[lib.scala 371:17]
  assign rvclkhdr_7_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ldst_dual_r = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  RdPtr = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  WrPtr = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  stbuf_addr_0 = _RAND_3[15:0];
  _RAND_4 = {1{`RANDOM}};
  _T_588 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  _T_580 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  _T_572 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  _T_564 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  _T_623 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  _T_615 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  _T_607 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  _T_599 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  stbuf_addr_1 = _RAND_12[15:0];
  _RAND_13 = {1{`RANDOM}};
  stbuf_addr_2 = _RAND_13[15:0];
  _RAND_14 = {1{`RANDOM}};
  stbuf_addr_3 = _RAND_14[15:0];
  _RAND_15 = {1{`RANDOM}};
  stbuf_byteen_0 = _RAND_15[3:0];
  _RAND_16 = {1{`RANDOM}};
  stbuf_byteen_1 = _RAND_16[3:0];
  _RAND_17 = {1{`RANDOM}};
  stbuf_byteen_2 = _RAND_17[3:0];
  _RAND_18 = {1{`RANDOM}};
  stbuf_byteen_3 = _RAND_18[3:0];
  _RAND_19 = {1{`RANDOM}};
  stbuf_data_0 = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  stbuf_data_1 = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  stbuf_data_2 = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  stbuf_data_3 = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  ldst_dual_m = _RAND_23[0:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    ldst_dual_r = 1'h0;
  end
  if (reset) begin
    RdPtr = 2'h0;
  end
  if (reset) begin
    WrPtr = 2'h0;
  end
  if (reset) begin
    stbuf_addr_0 = 16'h0;
  end
  if (reset) begin
    _T_588 = 1'h0;
  end
  if (reset) begin
    _T_580 = 1'h0;
  end
  if (reset) begin
    _T_572 = 1'h0;
  end
  if (reset) begin
    _T_564 = 1'h0;
  end
  if (reset) begin
    _T_623 = 1'h0;
  end
  if (reset) begin
    _T_615 = 1'h0;
  end
  if (reset) begin
    _T_607 = 1'h0;
  end
  if (reset) begin
    _T_599 = 1'h0;
  end
  if (reset) begin
    stbuf_addr_1 = 16'h0;
  end
  if (reset) begin
    stbuf_addr_2 = 16'h0;
  end
  if (reset) begin
    stbuf_addr_3 = 16'h0;
  end
  if (reset) begin
    stbuf_byteen_0 = 4'h0;
  end
  if (reset) begin
    stbuf_byteen_1 = 4'h0;
  end
  if (reset) begin
    stbuf_byteen_2 = 4'h0;
  end
  if (reset) begin
    stbuf_byteen_3 = 4'h0;
  end
  if (reset) begin
    stbuf_data_0 = 32'h0;
  end
  if (reset) begin
    stbuf_data_1 = 32'h0;
  end
  if (reset) begin
    stbuf_data_2 = 32'h0;
  end
  if (reset) begin
    stbuf_data_3 = 32'h0;
  end
  if (reset) begin
    ldst_dual_m = 1'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge io_lsu_c1_r_clk or posedge reset) begin
    if (reset) begin
      ldst_dual_r <= 1'h0;
    end else begin
      ldst_dual_r <= ldst_dual_m;
    end
  end
  always @(posedge io_lsu_stbuf_c1_clk or posedge reset) begin
    if (reset) begin
      RdPtr <= 2'h0;
    end else if (_T_212) begin
      RdPtr <= RdPtrPlus1;
    end
  end
  always @(posedge io_lsu_stbuf_c1_clk or posedge reset) begin
    if (reset) begin
      WrPtr <= 2'h0;
    end else if (WrPtrEn) begin
      if (_T_716) begin
        WrPtr <= WrPtrPlus2;
      end else begin
        WrPtr <= WrPtrPlus1;
      end
    end
  end
  always @(posedge rvclkhdr_io_l1clk or posedge reset) begin
    if (reset) begin
      stbuf_addr_0 <= 16'h0;
    end else if (sel_lo[0]) begin
      stbuf_addr_0 <= io_lsu_addr_r[15:0];
    end else begin
      stbuf_addr_0 <= io_end_addr_r[15:0];
    end
  end
  always @(posedge io_lsu_free_c2_clk or posedge reset) begin
    if (reset) begin
      _T_588 <= 1'h0;
    end else begin
      _T_588 <= _T_584 & _T_67;
    end
  end
  always @(posedge io_lsu_free_c2_clk or posedge reset) begin
    if (reset) begin
      _T_580 <= 1'h0;
    end else begin
      _T_580 <= _T_576 & _T_56;
    end
  end
  always @(posedge io_lsu_free_c2_clk or posedge reset) begin
    if (reset) begin
      _T_572 <= 1'h0;
    end else begin
      _T_572 <= _T_568 & _T_45;
    end
  end
  always @(posedge io_lsu_free_c2_clk or posedge reset) begin
    if (reset) begin
      _T_564 <= 1'h0;
    end else begin
      _T_564 <= _T_560 & _T_34;
    end
  end
  always @(posedge io_lsu_free_c2_clk or posedge reset) begin
    if (reset) begin
      _T_623 <= 1'h0;
    end else begin
      _T_623 <= _T_619 & _T_67;
    end
  end
  always @(posedge io_lsu_free_c2_clk or posedge reset) begin
    if (reset) begin
      _T_615 <= 1'h0;
    end else begin
      _T_615 <= _T_611 & _T_56;
    end
  end
  always @(posedge io_lsu_free_c2_clk or posedge reset) begin
    if (reset) begin
      _T_607 <= 1'h0;
    end else begin
      _T_607 <= _T_603 & _T_45;
    end
  end
  always @(posedge io_lsu_free_c2_clk or posedge reset) begin
    if (reset) begin
      _T_599 <= 1'h0;
    end else begin
      _T_599 <= _T_595 & _T_34;
    end
  end
  always @(posedge rvclkhdr_2_io_l1clk or posedge reset) begin
    if (reset) begin
      stbuf_addr_1 <= 16'h0;
    end else if (sel_lo[1]) begin
      stbuf_addr_1 <= io_lsu_addr_r[15:0];
    end else begin
      stbuf_addr_1 <= io_end_addr_r[15:0];
    end
  end
  always @(posedge rvclkhdr_4_io_l1clk or posedge reset) begin
    if (reset) begin
      stbuf_addr_2 <= 16'h0;
    end else if (sel_lo[2]) begin
      stbuf_addr_2 <= io_lsu_addr_r[15:0];
    end else begin
      stbuf_addr_2 <= io_end_addr_r[15:0];
    end
  end
  always @(posedge rvclkhdr_6_io_l1clk or posedge reset) begin
    if (reset) begin
      stbuf_addr_3 <= 16'h0;
    end else if (sel_lo[3]) begin
      stbuf_addr_3 <= io_lsu_addr_r[15:0];
    end else begin
      stbuf_addr_3 <= io_end_addr_r[15:0];
    end
  end
  always @(posedge io_lsu_stbuf_c1_clk or posedge reset) begin
    if (reset) begin
      stbuf_byteen_0 <= 4'h0;
    end else begin
      stbuf_byteen_0 <= _T_629 & _T_633;
    end
  end
  always @(posedge io_lsu_stbuf_c1_clk or posedge reset) begin
    if (reset) begin
      stbuf_byteen_1 <= 4'h0;
    end else begin
      stbuf_byteen_1 <= _T_638 & _T_642;
    end
  end
  always @(posedge io_lsu_stbuf_c1_clk or posedge reset) begin
    if (reset) begin
      stbuf_byteen_2 <= 4'h0;
    end else begin
      stbuf_byteen_2 <= _T_647 & _T_651;
    end
  end
  always @(posedge io_lsu_stbuf_c1_clk or posedge reset) begin
    if (reset) begin
      stbuf_byteen_3 <= 4'h0;
    end else begin
      stbuf_byteen_3 <= _T_656 & _T_660;
    end
  end
  always @(posedge rvclkhdr_1_io_l1clk or posedge reset) begin
    if (reset) begin
      stbuf_data_0 <= 32'h0;
    end else begin
      stbuf_data_0 <= {_T_546,_T_545};
    end
  end
  always @(posedge rvclkhdr_3_io_l1clk or posedge reset) begin
    if (reset) begin
      stbuf_data_1 <= 32'h0;
    end else begin
      stbuf_data_1 <= {_T_549,_T_548};
    end
  end
  always @(posedge rvclkhdr_5_io_l1clk or posedge reset) begin
    if (reset) begin
      stbuf_data_2 <= 32'h0;
    end else begin
      stbuf_data_2 <= {_T_552,_T_551};
    end
  end
  always @(posedge rvclkhdr_7_io_l1clk or posedge reset) begin
    if (reset) begin
      stbuf_data_3 <= 32'h0;
    end else begin
      stbuf_data_3 <= {_T_555,_T_554};
    end
  end
  always @(posedge io_lsu_c1_m_clk or posedge reset) begin
    if (reset) begin
      ldst_dual_m <= 1'h0;
    end else begin
      ldst_dual_m <= io_lsu_addr_d[2] != io_end_addr_d[2];
    end
  end
endmodule
module lsu_ecc(
  input         clock,
  input         reset,
  input         io_lsu_c2_r_clk,
  input         io_lsu_pkt_m_valid,
  input         io_lsu_pkt_m_bits_load,
  input         io_lsu_pkt_m_bits_store,
  input         io_lsu_pkt_m_bits_dma,
  input  [31:0] io_stbuf_data_any,
  input         io_dec_tlu_core_ecc_disable,
  input  [15:0] io_lsu_addr_m,
  input  [15:0] io_end_addr_m,
  input  [31:0] io_dccm_rdata_hi_m,
  input  [31:0] io_dccm_rdata_lo_m,
  input  [6:0]  io_dccm_data_ecc_hi_m,
  input  [6:0]  io_dccm_data_ecc_lo_m,
  input         io_ld_single_ecc_error_r,
  input         io_ld_single_ecc_error_r_ff,
  input         io_lsu_dccm_rden_m,
  input         io_addr_in_dccm_m,
  input         io_dma_dccm_wen,
  input  [31:0] io_dma_dccm_wdata_lo,
  input  [31:0] io_dma_dccm_wdata_hi,
  input         io_scan_mode,
  output [31:0] io_sec_data_hi_r,
  output [31:0] io_sec_data_lo_r,
  output [31:0] io_sec_data_hi_m,
  output [31:0] io_sec_data_lo_m,
  output [31:0] io_sec_data_hi_r_ff,
  output [31:0] io_sec_data_lo_r_ff,
  output [6:0]  io_dma_dccm_wdata_ecc_hi,
  output [6:0]  io_dma_dccm_wdata_ecc_lo,
  output [6:0]  io_stbuf_ecc_any,
  output [6:0]  io_sec_data_ecc_hi_r_ff,
  output [6:0]  io_sec_data_ecc_lo_r_ff,
  output        io_single_ecc_error_hi_r,
  output        io_single_ecc_error_lo_r,
  output        io_lsu_single_ecc_error_r,
  output        io_lsu_double_ecc_error_r,
  output        io_lsu_single_ecc_error_m,
  output        io_lsu_double_ecc_error_m
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  wire  rvclkhdr_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_1_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_1_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_1_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_1_io_scan_mode; // @[lib.scala 368:23]
  wire  _T_96 = ^io_dccm_rdata_hi_m; // @[lib.scala 193:30]
  wire  _T_97 = ^io_dccm_data_ecc_hi_m; // @[lib.scala 193:44]
  wire  _T_98 = _T_96 ^ _T_97; // @[lib.scala 193:35]
  wire [5:0] _T_106 = {io_dccm_rdata_hi_m[31],io_dccm_rdata_hi_m[30],io_dccm_rdata_hi_m[29],io_dccm_rdata_hi_m[28],io_dccm_rdata_hi_m[27],io_dccm_rdata_hi_m[26]}; // @[lib.scala 193:76]
  wire  _T_107 = ^_T_106; // @[lib.scala 193:83]
  wire  _T_108 = io_dccm_data_ecc_hi_m[5] ^ _T_107; // @[lib.scala 193:71]
  wire [6:0] _T_115 = {io_dccm_rdata_hi_m[17],io_dccm_rdata_hi_m[16],io_dccm_rdata_hi_m[15],io_dccm_rdata_hi_m[14],io_dccm_rdata_hi_m[13],io_dccm_rdata_hi_m[12],io_dccm_rdata_hi_m[11]}; // @[lib.scala 193:103]
  wire [14:0] _T_123 = {io_dccm_rdata_hi_m[25],io_dccm_rdata_hi_m[24],io_dccm_rdata_hi_m[23],io_dccm_rdata_hi_m[22],io_dccm_rdata_hi_m[21],io_dccm_rdata_hi_m[20],io_dccm_rdata_hi_m[19],io_dccm_rdata_hi_m[18],_T_115}; // @[lib.scala 193:103]
  wire  _T_124 = ^_T_123; // @[lib.scala 193:110]
  wire  _T_125 = io_dccm_data_ecc_hi_m[4] ^ _T_124; // @[lib.scala 193:98]
  wire [6:0] _T_132 = {io_dccm_rdata_hi_m[10],io_dccm_rdata_hi_m[9],io_dccm_rdata_hi_m[8],io_dccm_rdata_hi_m[7],io_dccm_rdata_hi_m[6],io_dccm_rdata_hi_m[5],io_dccm_rdata_hi_m[4]}; // @[lib.scala 193:130]
  wire [14:0] _T_140 = {io_dccm_rdata_hi_m[25],io_dccm_rdata_hi_m[24],io_dccm_rdata_hi_m[23],io_dccm_rdata_hi_m[22],io_dccm_rdata_hi_m[21],io_dccm_rdata_hi_m[20],io_dccm_rdata_hi_m[19],io_dccm_rdata_hi_m[18],_T_132}; // @[lib.scala 193:130]
  wire  _T_141 = ^_T_140; // @[lib.scala 193:137]
  wire  _T_142 = io_dccm_data_ecc_hi_m[3] ^ _T_141; // @[lib.scala 193:125]
  wire [8:0] _T_151 = {io_dccm_rdata_hi_m[15],io_dccm_rdata_hi_m[14],io_dccm_rdata_hi_m[10],io_dccm_rdata_hi_m[9],io_dccm_rdata_hi_m[8],io_dccm_rdata_hi_m[7],io_dccm_rdata_hi_m[3],io_dccm_rdata_hi_m[2],io_dccm_rdata_hi_m[1]}; // @[lib.scala 193:157]
  wire [17:0] _T_160 = {io_dccm_rdata_hi_m[31],io_dccm_rdata_hi_m[30],io_dccm_rdata_hi_m[29],io_dccm_rdata_hi_m[25],io_dccm_rdata_hi_m[24],io_dccm_rdata_hi_m[23],io_dccm_rdata_hi_m[22],io_dccm_rdata_hi_m[17],io_dccm_rdata_hi_m[16],_T_151}; // @[lib.scala 193:157]
  wire  _T_161 = ^_T_160; // @[lib.scala 193:164]
  wire  _T_162 = io_dccm_data_ecc_hi_m[2] ^ _T_161; // @[lib.scala 193:152]
  wire [8:0] _T_171 = {io_dccm_rdata_hi_m[13],io_dccm_rdata_hi_m[12],io_dccm_rdata_hi_m[10],io_dccm_rdata_hi_m[9],io_dccm_rdata_hi_m[6],io_dccm_rdata_hi_m[5],io_dccm_rdata_hi_m[3],io_dccm_rdata_hi_m[2],io_dccm_rdata_hi_m[0]}; // @[lib.scala 193:184]
  wire [17:0] _T_180 = {io_dccm_rdata_hi_m[31],io_dccm_rdata_hi_m[28],io_dccm_rdata_hi_m[27],io_dccm_rdata_hi_m[25],io_dccm_rdata_hi_m[24],io_dccm_rdata_hi_m[21],io_dccm_rdata_hi_m[20],io_dccm_rdata_hi_m[17],io_dccm_rdata_hi_m[16],_T_171}; // @[lib.scala 193:184]
  wire  _T_181 = ^_T_180; // @[lib.scala 193:191]
  wire  _T_182 = io_dccm_data_ecc_hi_m[1] ^ _T_181; // @[lib.scala 193:179]
  wire [8:0] _T_191 = {io_dccm_rdata_hi_m[13],io_dccm_rdata_hi_m[11],io_dccm_rdata_hi_m[10],io_dccm_rdata_hi_m[8],io_dccm_rdata_hi_m[6],io_dccm_rdata_hi_m[4],io_dccm_rdata_hi_m[3],io_dccm_rdata_hi_m[1],io_dccm_rdata_hi_m[0]}; // @[lib.scala 193:211]
  wire [17:0] _T_200 = {io_dccm_rdata_hi_m[30],io_dccm_rdata_hi_m[28],io_dccm_rdata_hi_m[26],io_dccm_rdata_hi_m[25],io_dccm_rdata_hi_m[23],io_dccm_rdata_hi_m[21],io_dccm_rdata_hi_m[19],io_dccm_rdata_hi_m[17],io_dccm_rdata_hi_m[15],_T_191}; // @[lib.scala 193:211]
  wire  _T_201 = ^_T_200; // @[lib.scala 193:218]
  wire  _T_202 = io_dccm_data_ecc_hi_m[0] ^ _T_201; // @[lib.scala 193:206]
  wire [6:0] _T_208 = {_T_98,_T_108,_T_125,_T_142,_T_162,_T_182,_T_202}; // @[Cat.scala 29:58]
  wire  _T_209 = _T_208 != 7'h0; // @[lib.scala 194:44]
  wire  _T_1131 = ~io_dec_tlu_core_ecc_disable; // @[lsu_ecc.scala 107:73]
  wire  _T_1138 = io_lsu_pkt_m_bits_load | io_lsu_pkt_m_bits_store; // @[lsu_ecc.scala 125:65]
  wire  _T_1139 = io_lsu_pkt_m_valid & _T_1138; // @[lsu_ecc.scala 125:39]
  wire  _T_1140 = _T_1139 & io_addr_in_dccm_m; // @[lsu_ecc.scala 125:92]
  wire  is_ldst_m = _T_1140 & io_lsu_dccm_rden_m; // @[lsu_ecc.scala 125:112]
  wire  ldst_dual_m = io_lsu_addr_m[2] != io_end_addr_m[2]; // @[lsu_ecc.scala 124:39]
  wire  _T_1144 = ldst_dual_m | io_lsu_pkt_m_bits_dma; // @[lsu_ecc.scala 127:48]
  wire  _T_1145 = is_ldst_m & _T_1144; // @[lsu_ecc.scala 127:33]
  wire  is_ldst_hi_m = _T_1145 & _T_1131; // @[lsu_ecc.scala 127:73]
  wire  _T_210 = is_ldst_hi_m & _T_209; // @[lib.scala 194:32]
  wire  single_ecc_error_hi_any = _T_210 & _T_208[6]; // @[lib.scala 194:53]
  wire  _T_215 = ~_T_208[6]; // @[lib.scala 195:55]
  wire  double_ecc_error_hi_any = _T_210 & _T_215; // @[lib.scala 195:53]
  wire  _T_218 = _T_208[5:0] == 6'h1; // @[lib.scala 199:41]
  wire  _T_220 = _T_208[5:0] == 6'h2; // @[lib.scala 199:41]
  wire  _T_222 = _T_208[5:0] == 6'h3; // @[lib.scala 199:41]
  wire  _T_224 = _T_208[5:0] == 6'h4; // @[lib.scala 199:41]
  wire  _T_226 = _T_208[5:0] == 6'h5; // @[lib.scala 199:41]
  wire  _T_228 = _T_208[5:0] == 6'h6; // @[lib.scala 199:41]
  wire  _T_230 = _T_208[5:0] == 6'h7; // @[lib.scala 199:41]
  wire  _T_232 = _T_208[5:0] == 6'h8; // @[lib.scala 199:41]
  wire  _T_234 = _T_208[5:0] == 6'h9; // @[lib.scala 199:41]
  wire  _T_236 = _T_208[5:0] == 6'ha; // @[lib.scala 199:41]
  wire  _T_238 = _T_208[5:0] == 6'hb; // @[lib.scala 199:41]
  wire  _T_240 = _T_208[5:0] == 6'hc; // @[lib.scala 199:41]
  wire  _T_242 = _T_208[5:0] == 6'hd; // @[lib.scala 199:41]
  wire  _T_244 = _T_208[5:0] == 6'he; // @[lib.scala 199:41]
  wire  _T_246 = _T_208[5:0] == 6'hf; // @[lib.scala 199:41]
  wire  _T_248 = _T_208[5:0] == 6'h10; // @[lib.scala 199:41]
  wire  _T_250 = _T_208[5:0] == 6'h11; // @[lib.scala 199:41]
  wire  _T_252 = _T_208[5:0] == 6'h12; // @[lib.scala 199:41]
  wire  _T_254 = _T_208[5:0] == 6'h13; // @[lib.scala 199:41]
  wire  _T_256 = _T_208[5:0] == 6'h14; // @[lib.scala 199:41]
  wire  _T_258 = _T_208[5:0] == 6'h15; // @[lib.scala 199:41]
  wire  _T_260 = _T_208[5:0] == 6'h16; // @[lib.scala 199:41]
  wire  _T_262 = _T_208[5:0] == 6'h17; // @[lib.scala 199:41]
  wire  _T_264 = _T_208[5:0] == 6'h18; // @[lib.scala 199:41]
  wire  _T_266 = _T_208[5:0] == 6'h19; // @[lib.scala 199:41]
  wire  _T_268 = _T_208[5:0] == 6'h1a; // @[lib.scala 199:41]
  wire  _T_270 = _T_208[5:0] == 6'h1b; // @[lib.scala 199:41]
  wire  _T_272 = _T_208[5:0] == 6'h1c; // @[lib.scala 199:41]
  wire  _T_274 = _T_208[5:0] == 6'h1d; // @[lib.scala 199:41]
  wire  _T_276 = _T_208[5:0] == 6'h1e; // @[lib.scala 199:41]
  wire  _T_278 = _T_208[5:0] == 6'h1f; // @[lib.scala 199:41]
  wire  _T_280 = _T_208[5:0] == 6'h20; // @[lib.scala 199:41]
  wire  _T_282 = _T_208[5:0] == 6'h21; // @[lib.scala 199:41]
  wire  _T_284 = _T_208[5:0] == 6'h22; // @[lib.scala 199:41]
  wire  _T_286 = _T_208[5:0] == 6'h23; // @[lib.scala 199:41]
  wire  _T_288 = _T_208[5:0] == 6'h24; // @[lib.scala 199:41]
  wire  _T_290 = _T_208[5:0] == 6'h25; // @[lib.scala 199:41]
  wire  _T_292 = _T_208[5:0] == 6'h26; // @[lib.scala 199:41]
  wire  _T_294 = _T_208[5:0] == 6'h27; // @[lib.scala 199:41]
  wire [7:0] _T_309 = {io_dccm_data_ecc_hi_m[3],io_dccm_rdata_hi_m[3:1],io_dccm_data_ecc_hi_m[2],io_dccm_rdata_hi_m[0],io_dccm_data_ecc_hi_m[1:0]}; // @[Cat.scala 29:58]
  wire [38:0] _T_315 = {io_dccm_data_ecc_hi_m[6],io_dccm_rdata_hi_m[31:26],io_dccm_data_ecc_hi_m[5],io_dccm_rdata_hi_m[25:11],io_dccm_data_ecc_hi_m[4],io_dccm_rdata_hi_m[10:4],_T_309}; // @[Cat.scala 29:58]
  wire [9:0] _T_333 = {_T_254,_T_252,_T_250,_T_248,_T_246,_T_244,_T_242,_T_240,_T_238,_T_236}; // @[lib.scala 202:69]
  wire [18:0] _T_334 = {_T_333,_T_234,_T_232,_T_230,_T_228,_T_226,_T_224,_T_222,_T_220,_T_218}; // @[lib.scala 202:69]
  wire [9:0] _T_343 = {_T_274,_T_272,_T_270,_T_268,_T_266,_T_264,_T_262,_T_260,_T_258,_T_256}; // @[lib.scala 202:69]
  wire [9:0] _T_352 = {_T_294,_T_292,_T_290,_T_288,_T_286,_T_284,_T_282,_T_280,_T_278,_T_276}; // @[lib.scala 202:69]
  wire [38:0] _T_354 = {_T_352,_T_343,_T_334}; // @[lib.scala 202:69]
  wire [38:0] _T_355 = _T_354 ^ _T_315; // @[lib.scala 202:76]
  wire [38:0] _T_356 = single_ecc_error_hi_any ? _T_355 : _T_315; // @[lib.scala 202:31]
  wire [3:0] _T_362 = {_T_356[6:4],_T_356[2]}; // @[Cat.scala 29:58]
  wire [27:0] _T_364 = {_T_356[37:32],_T_356[30:16],_T_356[14:8]}; // @[Cat.scala 29:58]
  wire  _T_474 = ^io_dccm_rdata_lo_m; // @[lib.scala 193:30]
  wire  _T_475 = ^io_dccm_data_ecc_lo_m; // @[lib.scala 193:44]
  wire  _T_476 = _T_474 ^ _T_475; // @[lib.scala 193:35]
  wire [5:0] _T_484 = {io_dccm_rdata_lo_m[31],io_dccm_rdata_lo_m[30],io_dccm_rdata_lo_m[29],io_dccm_rdata_lo_m[28],io_dccm_rdata_lo_m[27],io_dccm_rdata_lo_m[26]}; // @[lib.scala 193:76]
  wire  _T_485 = ^_T_484; // @[lib.scala 193:83]
  wire  _T_486 = io_dccm_data_ecc_lo_m[5] ^ _T_485; // @[lib.scala 193:71]
  wire [6:0] _T_493 = {io_dccm_rdata_lo_m[17],io_dccm_rdata_lo_m[16],io_dccm_rdata_lo_m[15],io_dccm_rdata_lo_m[14],io_dccm_rdata_lo_m[13],io_dccm_rdata_lo_m[12],io_dccm_rdata_lo_m[11]}; // @[lib.scala 193:103]
  wire [14:0] _T_501 = {io_dccm_rdata_lo_m[25],io_dccm_rdata_lo_m[24],io_dccm_rdata_lo_m[23],io_dccm_rdata_lo_m[22],io_dccm_rdata_lo_m[21],io_dccm_rdata_lo_m[20],io_dccm_rdata_lo_m[19],io_dccm_rdata_lo_m[18],_T_493}; // @[lib.scala 193:103]
  wire  _T_502 = ^_T_501; // @[lib.scala 193:110]
  wire  _T_503 = io_dccm_data_ecc_lo_m[4] ^ _T_502; // @[lib.scala 193:98]
  wire [6:0] _T_510 = {io_dccm_rdata_lo_m[10],io_dccm_rdata_lo_m[9],io_dccm_rdata_lo_m[8],io_dccm_rdata_lo_m[7],io_dccm_rdata_lo_m[6],io_dccm_rdata_lo_m[5],io_dccm_rdata_lo_m[4]}; // @[lib.scala 193:130]
  wire [14:0] _T_518 = {io_dccm_rdata_lo_m[25],io_dccm_rdata_lo_m[24],io_dccm_rdata_lo_m[23],io_dccm_rdata_lo_m[22],io_dccm_rdata_lo_m[21],io_dccm_rdata_lo_m[20],io_dccm_rdata_lo_m[19],io_dccm_rdata_lo_m[18],_T_510}; // @[lib.scala 193:130]
  wire  _T_519 = ^_T_518; // @[lib.scala 193:137]
  wire  _T_520 = io_dccm_data_ecc_lo_m[3] ^ _T_519; // @[lib.scala 193:125]
  wire [8:0] _T_529 = {io_dccm_rdata_lo_m[15],io_dccm_rdata_lo_m[14],io_dccm_rdata_lo_m[10],io_dccm_rdata_lo_m[9],io_dccm_rdata_lo_m[8],io_dccm_rdata_lo_m[7],io_dccm_rdata_lo_m[3],io_dccm_rdata_lo_m[2],io_dccm_rdata_lo_m[1]}; // @[lib.scala 193:157]
  wire [17:0] _T_538 = {io_dccm_rdata_lo_m[31],io_dccm_rdata_lo_m[30],io_dccm_rdata_lo_m[29],io_dccm_rdata_lo_m[25],io_dccm_rdata_lo_m[24],io_dccm_rdata_lo_m[23],io_dccm_rdata_lo_m[22],io_dccm_rdata_lo_m[17],io_dccm_rdata_lo_m[16],_T_529}; // @[lib.scala 193:157]
  wire  _T_539 = ^_T_538; // @[lib.scala 193:164]
  wire  _T_540 = io_dccm_data_ecc_lo_m[2] ^ _T_539; // @[lib.scala 193:152]
  wire [8:0] _T_549 = {io_dccm_rdata_lo_m[13],io_dccm_rdata_lo_m[12],io_dccm_rdata_lo_m[10],io_dccm_rdata_lo_m[9],io_dccm_rdata_lo_m[6],io_dccm_rdata_lo_m[5],io_dccm_rdata_lo_m[3],io_dccm_rdata_lo_m[2],io_dccm_rdata_lo_m[0]}; // @[lib.scala 193:184]
  wire [17:0] _T_558 = {io_dccm_rdata_lo_m[31],io_dccm_rdata_lo_m[28],io_dccm_rdata_lo_m[27],io_dccm_rdata_lo_m[25],io_dccm_rdata_lo_m[24],io_dccm_rdata_lo_m[21],io_dccm_rdata_lo_m[20],io_dccm_rdata_lo_m[17],io_dccm_rdata_lo_m[16],_T_549}; // @[lib.scala 193:184]
  wire  _T_559 = ^_T_558; // @[lib.scala 193:191]
  wire  _T_560 = io_dccm_data_ecc_lo_m[1] ^ _T_559; // @[lib.scala 193:179]
  wire [8:0] _T_569 = {io_dccm_rdata_lo_m[13],io_dccm_rdata_lo_m[11],io_dccm_rdata_lo_m[10],io_dccm_rdata_lo_m[8],io_dccm_rdata_lo_m[6],io_dccm_rdata_lo_m[4],io_dccm_rdata_lo_m[3],io_dccm_rdata_lo_m[1],io_dccm_rdata_lo_m[0]}; // @[lib.scala 193:211]
  wire [17:0] _T_578 = {io_dccm_rdata_lo_m[30],io_dccm_rdata_lo_m[28],io_dccm_rdata_lo_m[26],io_dccm_rdata_lo_m[25],io_dccm_rdata_lo_m[23],io_dccm_rdata_lo_m[21],io_dccm_rdata_lo_m[19],io_dccm_rdata_lo_m[17],io_dccm_rdata_lo_m[15],_T_569}; // @[lib.scala 193:211]
  wire  _T_579 = ^_T_578; // @[lib.scala 193:218]
  wire  _T_580 = io_dccm_data_ecc_lo_m[0] ^ _T_579; // @[lib.scala 193:206]
  wire [6:0] _T_586 = {_T_476,_T_486,_T_503,_T_520,_T_540,_T_560,_T_580}; // @[Cat.scala 29:58]
  wire  _T_587 = _T_586 != 7'h0; // @[lib.scala 194:44]
  wire  is_ldst_lo_m = is_ldst_m & _T_1131; // @[lsu_ecc.scala 126:33]
  wire  _T_588 = is_ldst_lo_m & _T_587; // @[lib.scala 194:32]
  wire  single_ecc_error_lo_any = _T_588 & _T_586[6]; // @[lib.scala 194:53]
  wire  _T_593 = ~_T_586[6]; // @[lib.scala 195:55]
  wire  double_ecc_error_lo_any = _T_588 & _T_593; // @[lib.scala 195:53]
  wire  _T_596 = _T_586[5:0] == 6'h1; // @[lib.scala 199:41]
  wire  _T_598 = _T_586[5:0] == 6'h2; // @[lib.scala 199:41]
  wire  _T_600 = _T_586[5:0] == 6'h3; // @[lib.scala 199:41]
  wire  _T_602 = _T_586[5:0] == 6'h4; // @[lib.scala 199:41]
  wire  _T_604 = _T_586[5:0] == 6'h5; // @[lib.scala 199:41]
  wire  _T_606 = _T_586[5:0] == 6'h6; // @[lib.scala 199:41]
  wire  _T_608 = _T_586[5:0] == 6'h7; // @[lib.scala 199:41]
  wire  _T_610 = _T_586[5:0] == 6'h8; // @[lib.scala 199:41]
  wire  _T_612 = _T_586[5:0] == 6'h9; // @[lib.scala 199:41]
  wire  _T_614 = _T_586[5:0] == 6'ha; // @[lib.scala 199:41]
  wire  _T_616 = _T_586[5:0] == 6'hb; // @[lib.scala 199:41]
  wire  _T_618 = _T_586[5:0] == 6'hc; // @[lib.scala 199:41]
  wire  _T_620 = _T_586[5:0] == 6'hd; // @[lib.scala 199:41]
  wire  _T_622 = _T_586[5:0] == 6'he; // @[lib.scala 199:41]
  wire  _T_624 = _T_586[5:0] == 6'hf; // @[lib.scala 199:41]
  wire  _T_626 = _T_586[5:0] == 6'h10; // @[lib.scala 199:41]
  wire  _T_628 = _T_586[5:0] == 6'h11; // @[lib.scala 199:41]
  wire  _T_630 = _T_586[5:0] == 6'h12; // @[lib.scala 199:41]
  wire  _T_632 = _T_586[5:0] == 6'h13; // @[lib.scala 199:41]
  wire  _T_634 = _T_586[5:0] == 6'h14; // @[lib.scala 199:41]
  wire  _T_636 = _T_586[5:0] == 6'h15; // @[lib.scala 199:41]
  wire  _T_638 = _T_586[5:0] == 6'h16; // @[lib.scala 199:41]
  wire  _T_640 = _T_586[5:0] == 6'h17; // @[lib.scala 199:41]
  wire  _T_642 = _T_586[5:0] == 6'h18; // @[lib.scala 199:41]
  wire  _T_644 = _T_586[5:0] == 6'h19; // @[lib.scala 199:41]
  wire  _T_646 = _T_586[5:0] == 6'h1a; // @[lib.scala 199:41]
  wire  _T_648 = _T_586[5:0] == 6'h1b; // @[lib.scala 199:41]
  wire  _T_650 = _T_586[5:0] == 6'h1c; // @[lib.scala 199:41]
  wire  _T_652 = _T_586[5:0] == 6'h1d; // @[lib.scala 199:41]
  wire  _T_654 = _T_586[5:0] == 6'h1e; // @[lib.scala 199:41]
  wire  _T_656 = _T_586[5:0] == 6'h1f; // @[lib.scala 199:41]
  wire  _T_658 = _T_586[5:0] == 6'h20; // @[lib.scala 199:41]
  wire  _T_660 = _T_586[5:0] == 6'h21; // @[lib.scala 199:41]
  wire  _T_662 = _T_586[5:0] == 6'h22; // @[lib.scala 199:41]
  wire  _T_664 = _T_586[5:0] == 6'h23; // @[lib.scala 199:41]
  wire  _T_666 = _T_586[5:0] == 6'h24; // @[lib.scala 199:41]
  wire  _T_668 = _T_586[5:0] == 6'h25; // @[lib.scala 199:41]
  wire  _T_670 = _T_586[5:0] == 6'h26; // @[lib.scala 199:41]
  wire  _T_672 = _T_586[5:0] == 6'h27; // @[lib.scala 199:41]
  wire [7:0] _T_687 = {io_dccm_data_ecc_lo_m[3],io_dccm_rdata_lo_m[3:1],io_dccm_data_ecc_lo_m[2],io_dccm_rdata_lo_m[0],io_dccm_data_ecc_lo_m[1:0]}; // @[Cat.scala 29:58]
  wire [38:0] _T_693 = {io_dccm_data_ecc_lo_m[6],io_dccm_rdata_lo_m[31:26],io_dccm_data_ecc_lo_m[5],io_dccm_rdata_lo_m[25:11],io_dccm_data_ecc_lo_m[4],io_dccm_rdata_lo_m[10:4],_T_687}; // @[Cat.scala 29:58]
  wire [9:0] _T_711 = {_T_632,_T_630,_T_628,_T_626,_T_624,_T_622,_T_620,_T_618,_T_616,_T_614}; // @[lib.scala 202:69]
  wire [18:0] _T_712 = {_T_711,_T_612,_T_610,_T_608,_T_606,_T_604,_T_602,_T_600,_T_598,_T_596}; // @[lib.scala 202:69]
  wire [9:0] _T_721 = {_T_652,_T_650,_T_648,_T_646,_T_644,_T_642,_T_640,_T_638,_T_636,_T_634}; // @[lib.scala 202:69]
  wire [9:0] _T_730 = {_T_672,_T_670,_T_668,_T_666,_T_664,_T_662,_T_660,_T_658,_T_656,_T_654}; // @[lib.scala 202:69]
  wire [38:0] _T_732 = {_T_730,_T_721,_T_712}; // @[lib.scala 202:69]
  wire [38:0] _T_733 = _T_732 ^ _T_693; // @[lib.scala 202:76]
  wire [38:0] _T_734 = single_ecc_error_lo_any ? _T_733 : _T_693; // @[lib.scala 202:31]
  wire [3:0] _T_740 = {_T_734[6:4],_T_734[2]}; // @[Cat.scala 29:58]
  wire [27:0] _T_742 = {_T_734[37:32],_T_734[30:16],_T_734[14:8]}; // @[Cat.scala 29:58]
  wire [31:0] _T_1158 = io_dma_dccm_wen ? io_dma_dccm_wdata_lo : io_stbuf_data_any; // @[lsu_ecc.scala 149:87]
  wire [31:0] dccm_wdata_lo_any = io_ld_single_ecc_error_r_ff ? io_sec_data_lo_r_ff : _T_1158; // @[lsu_ecc.scala 149:27]
  wire  _T_774 = dccm_wdata_lo_any[0] ^ dccm_wdata_lo_any[1]; // @[lib.scala 119:74]
  wire  _T_775 = _T_774 ^ dccm_wdata_lo_any[3]; // @[lib.scala 119:74]
  wire  _T_776 = _T_775 ^ dccm_wdata_lo_any[4]; // @[lib.scala 119:74]
  wire  _T_777 = _T_776 ^ dccm_wdata_lo_any[6]; // @[lib.scala 119:74]
  wire  _T_778 = _T_777 ^ dccm_wdata_lo_any[8]; // @[lib.scala 119:74]
  wire  _T_779 = _T_778 ^ dccm_wdata_lo_any[10]; // @[lib.scala 119:74]
  wire  _T_780 = _T_779 ^ dccm_wdata_lo_any[11]; // @[lib.scala 119:74]
  wire  _T_781 = _T_780 ^ dccm_wdata_lo_any[13]; // @[lib.scala 119:74]
  wire  _T_782 = _T_781 ^ dccm_wdata_lo_any[15]; // @[lib.scala 119:74]
  wire  _T_783 = _T_782 ^ dccm_wdata_lo_any[17]; // @[lib.scala 119:74]
  wire  _T_784 = _T_783 ^ dccm_wdata_lo_any[19]; // @[lib.scala 119:74]
  wire  _T_785 = _T_784 ^ dccm_wdata_lo_any[21]; // @[lib.scala 119:74]
  wire  _T_786 = _T_785 ^ dccm_wdata_lo_any[23]; // @[lib.scala 119:74]
  wire  _T_787 = _T_786 ^ dccm_wdata_lo_any[25]; // @[lib.scala 119:74]
  wire  _T_788 = _T_787 ^ dccm_wdata_lo_any[26]; // @[lib.scala 119:74]
  wire  _T_789 = _T_788 ^ dccm_wdata_lo_any[28]; // @[lib.scala 119:74]
  wire  _T_790 = _T_789 ^ dccm_wdata_lo_any[30]; // @[lib.scala 119:74]
  wire  _T_809 = dccm_wdata_lo_any[0] ^ dccm_wdata_lo_any[2]; // @[lib.scala 119:74]
  wire  _T_810 = _T_809 ^ dccm_wdata_lo_any[3]; // @[lib.scala 119:74]
  wire  _T_811 = _T_810 ^ dccm_wdata_lo_any[5]; // @[lib.scala 119:74]
  wire  _T_812 = _T_811 ^ dccm_wdata_lo_any[6]; // @[lib.scala 119:74]
  wire  _T_813 = _T_812 ^ dccm_wdata_lo_any[9]; // @[lib.scala 119:74]
  wire  _T_814 = _T_813 ^ dccm_wdata_lo_any[10]; // @[lib.scala 119:74]
  wire  _T_815 = _T_814 ^ dccm_wdata_lo_any[12]; // @[lib.scala 119:74]
  wire  _T_816 = _T_815 ^ dccm_wdata_lo_any[13]; // @[lib.scala 119:74]
  wire  _T_817 = _T_816 ^ dccm_wdata_lo_any[16]; // @[lib.scala 119:74]
  wire  _T_818 = _T_817 ^ dccm_wdata_lo_any[17]; // @[lib.scala 119:74]
  wire  _T_819 = _T_818 ^ dccm_wdata_lo_any[20]; // @[lib.scala 119:74]
  wire  _T_820 = _T_819 ^ dccm_wdata_lo_any[21]; // @[lib.scala 119:74]
  wire  _T_821 = _T_820 ^ dccm_wdata_lo_any[24]; // @[lib.scala 119:74]
  wire  _T_822 = _T_821 ^ dccm_wdata_lo_any[25]; // @[lib.scala 119:74]
  wire  _T_823 = _T_822 ^ dccm_wdata_lo_any[27]; // @[lib.scala 119:74]
  wire  _T_824 = _T_823 ^ dccm_wdata_lo_any[28]; // @[lib.scala 119:74]
  wire  _T_825 = _T_824 ^ dccm_wdata_lo_any[31]; // @[lib.scala 119:74]
  wire  _T_844 = dccm_wdata_lo_any[1] ^ dccm_wdata_lo_any[2]; // @[lib.scala 119:74]
  wire  _T_845 = _T_844 ^ dccm_wdata_lo_any[3]; // @[lib.scala 119:74]
  wire  _T_846 = _T_845 ^ dccm_wdata_lo_any[7]; // @[lib.scala 119:74]
  wire  _T_847 = _T_846 ^ dccm_wdata_lo_any[8]; // @[lib.scala 119:74]
  wire  _T_848 = _T_847 ^ dccm_wdata_lo_any[9]; // @[lib.scala 119:74]
  wire  _T_849 = _T_848 ^ dccm_wdata_lo_any[10]; // @[lib.scala 119:74]
  wire  _T_850 = _T_849 ^ dccm_wdata_lo_any[14]; // @[lib.scala 119:74]
  wire  _T_851 = _T_850 ^ dccm_wdata_lo_any[15]; // @[lib.scala 119:74]
  wire  _T_852 = _T_851 ^ dccm_wdata_lo_any[16]; // @[lib.scala 119:74]
  wire  _T_853 = _T_852 ^ dccm_wdata_lo_any[17]; // @[lib.scala 119:74]
  wire  _T_854 = _T_853 ^ dccm_wdata_lo_any[22]; // @[lib.scala 119:74]
  wire  _T_855 = _T_854 ^ dccm_wdata_lo_any[23]; // @[lib.scala 119:74]
  wire  _T_856 = _T_855 ^ dccm_wdata_lo_any[24]; // @[lib.scala 119:74]
  wire  _T_857 = _T_856 ^ dccm_wdata_lo_any[25]; // @[lib.scala 119:74]
  wire  _T_858 = _T_857 ^ dccm_wdata_lo_any[29]; // @[lib.scala 119:74]
  wire  _T_859 = _T_858 ^ dccm_wdata_lo_any[30]; // @[lib.scala 119:74]
  wire  _T_860 = _T_859 ^ dccm_wdata_lo_any[31]; // @[lib.scala 119:74]
  wire  _T_876 = dccm_wdata_lo_any[4] ^ dccm_wdata_lo_any[5]; // @[lib.scala 119:74]
  wire  _T_877 = _T_876 ^ dccm_wdata_lo_any[6]; // @[lib.scala 119:74]
  wire  _T_878 = _T_877 ^ dccm_wdata_lo_any[7]; // @[lib.scala 119:74]
  wire  _T_879 = _T_878 ^ dccm_wdata_lo_any[8]; // @[lib.scala 119:74]
  wire  _T_880 = _T_879 ^ dccm_wdata_lo_any[9]; // @[lib.scala 119:74]
  wire  _T_881 = _T_880 ^ dccm_wdata_lo_any[10]; // @[lib.scala 119:74]
  wire  _T_882 = _T_881 ^ dccm_wdata_lo_any[18]; // @[lib.scala 119:74]
  wire  _T_883 = _T_882 ^ dccm_wdata_lo_any[19]; // @[lib.scala 119:74]
  wire  _T_884 = _T_883 ^ dccm_wdata_lo_any[20]; // @[lib.scala 119:74]
  wire  _T_885 = _T_884 ^ dccm_wdata_lo_any[21]; // @[lib.scala 119:74]
  wire  _T_886 = _T_885 ^ dccm_wdata_lo_any[22]; // @[lib.scala 119:74]
  wire  _T_887 = _T_886 ^ dccm_wdata_lo_any[23]; // @[lib.scala 119:74]
  wire  _T_888 = _T_887 ^ dccm_wdata_lo_any[24]; // @[lib.scala 119:74]
  wire  _T_889 = _T_888 ^ dccm_wdata_lo_any[25]; // @[lib.scala 119:74]
  wire  _T_905 = dccm_wdata_lo_any[11] ^ dccm_wdata_lo_any[12]; // @[lib.scala 119:74]
  wire  _T_906 = _T_905 ^ dccm_wdata_lo_any[13]; // @[lib.scala 119:74]
  wire  _T_907 = _T_906 ^ dccm_wdata_lo_any[14]; // @[lib.scala 119:74]
  wire  _T_908 = _T_907 ^ dccm_wdata_lo_any[15]; // @[lib.scala 119:74]
  wire  _T_909 = _T_908 ^ dccm_wdata_lo_any[16]; // @[lib.scala 119:74]
  wire  _T_910 = _T_909 ^ dccm_wdata_lo_any[17]; // @[lib.scala 119:74]
  wire  _T_911 = _T_910 ^ dccm_wdata_lo_any[18]; // @[lib.scala 119:74]
  wire  _T_912 = _T_911 ^ dccm_wdata_lo_any[19]; // @[lib.scala 119:74]
  wire  _T_913 = _T_912 ^ dccm_wdata_lo_any[20]; // @[lib.scala 119:74]
  wire  _T_914 = _T_913 ^ dccm_wdata_lo_any[21]; // @[lib.scala 119:74]
  wire  _T_915 = _T_914 ^ dccm_wdata_lo_any[22]; // @[lib.scala 119:74]
  wire  _T_916 = _T_915 ^ dccm_wdata_lo_any[23]; // @[lib.scala 119:74]
  wire  _T_917 = _T_916 ^ dccm_wdata_lo_any[24]; // @[lib.scala 119:74]
  wire  _T_918 = _T_917 ^ dccm_wdata_lo_any[25]; // @[lib.scala 119:74]
  wire  _T_925 = dccm_wdata_lo_any[26] ^ dccm_wdata_lo_any[27]; // @[lib.scala 119:74]
  wire  _T_926 = _T_925 ^ dccm_wdata_lo_any[28]; // @[lib.scala 119:74]
  wire  _T_927 = _T_926 ^ dccm_wdata_lo_any[29]; // @[lib.scala 119:74]
  wire  _T_928 = _T_927 ^ dccm_wdata_lo_any[30]; // @[lib.scala 119:74]
  wire  _T_929 = _T_928 ^ dccm_wdata_lo_any[31]; // @[lib.scala 119:74]
  wire [5:0] _T_934 = {_T_929,_T_918,_T_889,_T_860,_T_825,_T_790}; // @[Cat.scala 29:58]
  wire  _T_935 = ^dccm_wdata_lo_any; // @[lib.scala 127:13]
  wire  _T_936 = ^_T_934; // @[lib.scala 127:23]
  wire  _T_937 = _T_935 ^ _T_936; // @[lib.scala 127:18]
  wire [31:0] _T_1162 = io_dma_dccm_wen ? io_dma_dccm_wdata_hi : io_stbuf_data_any; // @[lsu_ecc.scala 150:87]
  wire [31:0] dccm_wdata_hi_any = io_ld_single_ecc_error_r_ff ? io_sec_data_hi_r_ff : _T_1162; // @[lsu_ecc.scala 150:27]
  wire  _T_956 = dccm_wdata_hi_any[0] ^ dccm_wdata_hi_any[1]; // @[lib.scala 119:74]
  wire  _T_957 = _T_956 ^ dccm_wdata_hi_any[3]; // @[lib.scala 119:74]
  wire  _T_958 = _T_957 ^ dccm_wdata_hi_any[4]; // @[lib.scala 119:74]
  wire  _T_959 = _T_958 ^ dccm_wdata_hi_any[6]; // @[lib.scala 119:74]
  wire  _T_960 = _T_959 ^ dccm_wdata_hi_any[8]; // @[lib.scala 119:74]
  wire  _T_961 = _T_960 ^ dccm_wdata_hi_any[10]; // @[lib.scala 119:74]
  wire  _T_962 = _T_961 ^ dccm_wdata_hi_any[11]; // @[lib.scala 119:74]
  wire  _T_963 = _T_962 ^ dccm_wdata_hi_any[13]; // @[lib.scala 119:74]
  wire  _T_964 = _T_963 ^ dccm_wdata_hi_any[15]; // @[lib.scala 119:74]
  wire  _T_965 = _T_964 ^ dccm_wdata_hi_any[17]; // @[lib.scala 119:74]
  wire  _T_966 = _T_965 ^ dccm_wdata_hi_any[19]; // @[lib.scala 119:74]
  wire  _T_967 = _T_966 ^ dccm_wdata_hi_any[21]; // @[lib.scala 119:74]
  wire  _T_968 = _T_967 ^ dccm_wdata_hi_any[23]; // @[lib.scala 119:74]
  wire  _T_969 = _T_968 ^ dccm_wdata_hi_any[25]; // @[lib.scala 119:74]
  wire  _T_970 = _T_969 ^ dccm_wdata_hi_any[26]; // @[lib.scala 119:74]
  wire  _T_971 = _T_970 ^ dccm_wdata_hi_any[28]; // @[lib.scala 119:74]
  wire  _T_972 = _T_971 ^ dccm_wdata_hi_any[30]; // @[lib.scala 119:74]
  wire  _T_991 = dccm_wdata_hi_any[0] ^ dccm_wdata_hi_any[2]; // @[lib.scala 119:74]
  wire  _T_992 = _T_991 ^ dccm_wdata_hi_any[3]; // @[lib.scala 119:74]
  wire  _T_993 = _T_992 ^ dccm_wdata_hi_any[5]; // @[lib.scala 119:74]
  wire  _T_994 = _T_993 ^ dccm_wdata_hi_any[6]; // @[lib.scala 119:74]
  wire  _T_995 = _T_994 ^ dccm_wdata_hi_any[9]; // @[lib.scala 119:74]
  wire  _T_996 = _T_995 ^ dccm_wdata_hi_any[10]; // @[lib.scala 119:74]
  wire  _T_997 = _T_996 ^ dccm_wdata_hi_any[12]; // @[lib.scala 119:74]
  wire  _T_998 = _T_997 ^ dccm_wdata_hi_any[13]; // @[lib.scala 119:74]
  wire  _T_999 = _T_998 ^ dccm_wdata_hi_any[16]; // @[lib.scala 119:74]
  wire  _T_1000 = _T_999 ^ dccm_wdata_hi_any[17]; // @[lib.scala 119:74]
  wire  _T_1001 = _T_1000 ^ dccm_wdata_hi_any[20]; // @[lib.scala 119:74]
  wire  _T_1002 = _T_1001 ^ dccm_wdata_hi_any[21]; // @[lib.scala 119:74]
  wire  _T_1003 = _T_1002 ^ dccm_wdata_hi_any[24]; // @[lib.scala 119:74]
  wire  _T_1004 = _T_1003 ^ dccm_wdata_hi_any[25]; // @[lib.scala 119:74]
  wire  _T_1005 = _T_1004 ^ dccm_wdata_hi_any[27]; // @[lib.scala 119:74]
  wire  _T_1006 = _T_1005 ^ dccm_wdata_hi_any[28]; // @[lib.scala 119:74]
  wire  _T_1007 = _T_1006 ^ dccm_wdata_hi_any[31]; // @[lib.scala 119:74]
  wire  _T_1026 = dccm_wdata_hi_any[1] ^ dccm_wdata_hi_any[2]; // @[lib.scala 119:74]
  wire  _T_1027 = _T_1026 ^ dccm_wdata_hi_any[3]; // @[lib.scala 119:74]
  wire  _T_1028 = _T_1027 ^ dccm_wdata_hi_any[7]; // @[lib.scala 119:74]
  wire  _T_1029 = _T_1028 ^ dccm_wdata_hi_any[8]; // @[lib.scala 119:74]
  wire  _T_1030 = _T_1029 ^ dccm_wdata_hi_any[9]; // @[lib.scala 119:74]
  wire  _T_1031 = _T_1030 ^ dccm_wdata_hi_any[10]; // @[lib.scala 119:74]
  wire  _T_1032 = _T_1031 ^ dccm_wdata_hi_any[14]; // @[lib.scala 119:74]
  wire  _T_1033 = _T_1032 ^ dccm_wdata_hi_any[15]; // @[lib.scala 119:74]
  wire  _T_1034 = _T_1033 ^ dccm_wdata_hi_any[16]; // @[lib.scala 119:74]
  wire  _T_1035 = _T_1034 ^ dccm_wdata_hi_any[17]; // @[lib.scala 119:74]
  wire  _T_1036 = _T_1035 ^ dccm_wdata_hi_any[22]; // @[lib.scala 119:74]
  wire  _T_1037 = _T_1036 ^ dccm_wdata_hi_any[23]; // @[lib.scala 119:74]
  wire  _T_1038 = _T_1037 ^ dccm_wdata_hi_any[24]; // @[lib.scala 119:74]
  wire  _T_1039 = _T_1038 ^ dccm_wdata_hi_any[25]; // @[lib.scala 119:74]
  wire  _T_1040 = _T_1039 ^ dccm_wdata_hi_any[29]; // @[lib.scala 119:74]
  wire  _T_1041 = _T_1040 ^ dccm_wdata_hi_any[30]; // @[lib.scala 119:74]
  wire  _T_1042 = _T_1041 ^ dccm_wdata_hi_any[31]; // @[lib.scala 119:74]
  wire  _T_1058 = dccm_wdata_hi_any[4] ^ dccm_wdata_hi_any[5]; // @[lib.scala 119:74]
  wire  _T_1059 = _T_1058 ^ dccm_wdata_hi_any[6]; // @[lib.scala 119:74]
  wire  _T_1060 = _T_1059 ^ dccm_wdata_hi_any[7]; // @[lib.scala 119:74]
  wire  _T_1061 = _T_1060 ^ dccm_wdata_hi_any[8]; // @[lib.scala 119:74]
  wire  _T_1062 = _T_1061 ^ dccm_wdata_hi_any[9]; // @[lib.scala 119:74]
  wire  _T_1063 = _T_1062 ^ dccm_wdata_hi_any[10]; // @[lib.scala 119:74]
  wire  _T_1064 = _T_1063 ^ dccm_wdata_hi_any[18]; // @[lib.scala 119:74]
  wire  _T_1065 = _T_1064 ^ dccm_wdata_hi_any[19]; // @[lib.scala 119:74]
  wire  _T_1066 = _T_1065 ^ dccm_wdata_hi_any[20]; // @[lib.scala 119:74]
  wire  _T_1067 = _T_1066 ^ dccm_wdata_hi_any[21]; // @[lib.scala 119:74]
  wire  _T_1068 = _T_1067 ^ dccm_wdata_hi_any[22]; // @[lib.scala 119:74]
  wire  _T_1069 = _T_1068 ^ dccm_wdata_hi_any[23]; // @[lib.scala 119:74]
  wire  _T_1070 = _T_1069 ^ dccm_wdata_hi_any[24]; // @[lib.scala 119:74]
  wire  _T_1071 = _T_1070 ^ dccm_wdata_hi_any[25]; // @[lib.scala 119:74]
  wire  _T_1087 = dccm_wdata_hi_any[11] ^ dccm_wdata_hi_any[12]; // @[lib.scala 119:74]
  wire  _T_1088 = _T_1087 ^ dccm_wdata_hi_any[13]; // @[lib.scala 119:74]
  wire  _T_1089 = _T_1088 ^ dccm_wdata_hi_any[14]; // @[lib.scala 119:74]
  wire  _T_1090 = _T_1089 ^ dccm_wdata_hi_any[15]; // @[lib.scala 119:74]
  wire  _T_1091 = _T_1090 ^ dccm_wdata_hi_any[16]; // @[lib.scala 119:74]
  wire  _T_1092 = _T_1091 ^ dccm_wdata_hi_any[17]; // @[lib.scala 119:74]
  wire  _T_1093 = _T_1092 ^ dccm_wdata_hi_any[18]; // @[lib.scala 119:74]
  wire  _T_1094 = _T_1093 ^ dccm_wdata_hi_any[19]; // @[lib.scala 119:74]
  wire  _T_1095 = _T_1094 ^ dccm_wdata_hi_any[20]; // @[lib.scala 119:74]
  wire  _T_1096 = _T_1095 ^ dccm_wdata_hi_any[21]; // @[lib.scala 119:74]
  wire  _T_1097 = _T_1096 ^ dccm_wdata_hi_any[22]; // @[lib.scala 119:74]
  wire  _T_1098 = _T_1097 ^ dccm_wdata_hi_any[23]; // @[lib.scala 119:74]
  wire  _T_1099 = _T_1098 ^ dccm_wdata_hi_any[24]; // @[lib.scala 119:74]
  wire  _T_1100 = _T_1099 ^ dccm_wdata_hi_any[25]; // @[lib.scala 119:74]
  wire  _T_1107 = dccm_wdata_hi_any[26] ^ dccm_wdata_hi_any[27]; // @[lib.scala 119:74]
  wire  _T_1108 = _T_1107 ^ dccm_wdata_hi_any[28]; // @[lib.scala 119:74]
  wire  _T_1109 = _T_1108 ^ dccm_wdata_hi_any[29]; // @[lib.scala 119:74]
  wire  _T_1110 = _T_1109 ^ dccm_wdata_hi_any[30]; // @[lib.scala 119:74]
  wire  _T_1111 = _T_1110 ^ dccm_wdata_hi_any[31]; // @[lib.scala 119:74]
  wire [5:0] _T_1116 = {_T_1111,_T_1100,_T_1071,_T_1042,_T_1007,_T_972}; // @[Cat.scala 29:58]
  wire  _T_1117 = ^dccm_wdata_hi_any; // @[lib.scala 127:13]
  wire  _T_1118 = ^_T_1116; // @[lib.scala 127:23]
  wire  _T_1119 = _T_1117 ^ _T_1118; // @[lib.scala 127:18]
  reg  _T_1150; // @[lsu_ecc.scala 141:72]
  reg  _T_1151; // @[lsu_ecc.scala 142:72]
  reg  _T_1152; // @[lsu_ecc.scala 143:72]
  reg  _T_1153; // @[lsu_ecc.scala 144:72]
  reg [31:0] _T_1154; // @[lsu_ecc.scala 145:72]
  reg [31:0] _T_1155; // @[lsu_ecc.scala 146:72]
  reg [31:0] _T_1164; // @[lib.scala 374:16]
  reg [31:0] _T_1165; // @[lib.scala 374:16]
  rvclkhdr rvclkhdr ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_io_l1clk),
    .io_clk(rvclkhdr_io_clk),
    .io_en(rvclkhdr_io_en),
    .io_scan_mode(rvclkhdr_io_scan_mode)
  );
  rvclkhdr rvclkhdr_1 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_1_io_l1clk),
    .io_clk(rvclkhdr_1_io_clk),
    .io_en(rvclkhdr_1_io_en),
    .io_scan_mode(rvclkhdr_1_io_scan_mode)
  );
  assign io_sec_data_hi_r = _T_1154; // @[lsu_ecc.scala 114:22 lsu_ecc.scala 145:62]
  assign io_sec_data_lo_r = _T_1155; // @[lsu_ecc.scala 117:25 lsu_ecc.scala 146:62]
  assign io_sec_data_hi_m = {_T_364,_T_362}; // @[lsu_ecc.scala 90:32 lsu_ecc.scala 134:27]
  assign io_sec_data_lo_m = {_T_742,_T_740}; // @[lsu_ecc.scala 91:32 lsu_ecc.scala 136:27]
  assign io_sec_data_hi_r_ff = _T_1164; // @[lsu_ecc.scala 157:23]
  assign io_sec_data_lo_r_ff = _T_1165; // @[lsu_ecc.scala 158:23]
  assign io_dma_dccm_wdata_ecc_hi = {_T_1119,_T_1116}; // @[lsu_ecc.scala 154:28]
  assign io_dma_dccm_wdata_ecc_lo = {_T_937,_T_934}; // @[lsu_ecc.scala 155:28]
  assign io_stbuf_ecc_any = {_T_937,_T_934}; // @[lsu_ecc.scala 153:28]
  assign io_sec_data_ecc_hi_r_ff = {_T_1119,_T_1116}; // @[lsu_ecc.scala 151:28]
  assign io_sec_data_ecc_lo_r_ff = {_T_937,_T_934}; // @[lsu_ecc.scala 152:28]
  assign io_single_ecc_error_hi_r = _T_1153; // @[lsu_ecc.scala 115:31 lsu_ecc.scala 144:62]
  assign io_single_ecc_error_lo_r = _T_1152; // @[lsu_ecc.scala 118:31 lsu_ecc.scala 143:62]
  assign io_lsu_single_ecc_error_r = _T_1150; // @[lsu_ecc.scala 120:31 lsu_ecc.scala 141:62]
  assign io_lsu_double_ecc_error_r = _T_1151; // @[lsu_ecc.scala 121:31 lsu_ecc.scala 142:62]
  assign io_lsu_single_ecc_error_m = single_ecc_error_hi_any | single_ecc_error_lo_any; // @[lsu_ecc.scala 92:30 lsu_ecc.scala 138:33]
  assign io_lsu_double_ecc_error_m = double_ecc_error_hi_any | double_ecc_error_lo_any; // @[lsu_ecc.scala 93:30 lsu_ecc.scala 139:33]
  assign rvclkhdr_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_io_en = io_ld_single_ecc_error_r; // @[lib.scala 371:17]
  assign rvclkhdr_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_1_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_1_io_en = io_ld_single_ecc_error_r; // @[lib.scala 371:17]
  assign rvclkhdr_1_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_1150 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  _T_1151 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  _T_1152 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  _T_1153 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  _T_1154 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  _T_1155 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  _T_1164 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  _T_1165 = _RAND_7[31:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    _T_1150 = 1'h0;
  end
  if (reset) begin
    _T_1151 = 1'h0;
  end
  if (reset) begin
    _T_1152 = 1'h0;
  end
  if (reset) begin
    _T_1153 = 1'h0;
  end
  if (reset) begin
    _T_1154 = 32'h0;
  end
  if (reset) begin
    _T_1155 = 32'h0;
  end
  if (reset) begin
    _T_1164 = 32'h0;
  end
  if (reset) begin
    _T_1165 = 32'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge io_lsu_c2_r_clk or posedge reset) begin
    if (reset) begin
      _T_1150 <= 1'h0;
    end else begin
      _T_1150 <= io_lsu_single_ecc_error_m;
    end
  end
  always @(posedge io_lsu_c2_r_clk or posedge reset) begin
    if (reset) begin
      _T_1151 <= 1'h0;
    end else begin
      _T_1151 <= io_lsu_double_ecc_error_m;
    end
  end
  always @(posedge io_lsu_c2_r_clk or posedge reset) begin
    if (reset) begin
      _T_1152 <= 1'h0;
    end else begin
      _T_1152 <= _T_588 & _T_586[6];
    end
  end
  always @(posedge io_lsu_c2_r_clk or posedge reset) begin
    if (reset) begin
      _T_1153 <= 1'h0;
    end else begin
      _T_1153 <= _T_210 & _T_208[6];
    end
  end
  always @(posedge io_lsu_c2_r_clk or posedge reset) begin
    if (reset) begin
      _T_1154 <= 32'h0;
    end else begin
      _T_1154 <= io_sec_data_hi_m;
    end
  end
  always @(posedge io_lsu_c2_r_clk or posedge reset) begin
    if (reset) begin
      _T_1155 <= 32'h0;
    end else begin
      _T_1155 <= io_sec_data_lo_m;
    end
  end
  always @(posedge rvclkhdr_io_l1clk or posedge reset) begin
    if (reset) begin
      _T_1164 <= 32'h0;
    end else begin
      _T_1164 <= io_sec_data_hi_r;
    end
  end
  always @(posedge rvclkhdr_1_io_l1clk or posedge reset) begin
    if (reset) begin
      _T_1165 <= 32'h0;
    end else begin
      _T_1165 <= io_sec_data_lo_r;
    end
  end
endmodule
module lsu_trigger(
  input         io_trigger_pkt_any_0_select,
  input         io_trigger_pkt_any_0_match_pkt,
  input         io_trigger_pkt_any_0_store,
  input         io_trigger_pkt_any_0_load,
  input  [31:0] io_trigger_pkt_any_0_tdata2,
  input         io_trigger_pkt_any_1_select,
  input         io_trigger_pkt_any_1_match_pkt,
  input         io_trigger_pkt_any_1_store,
  input         io_trigger_pkt_any_1_load,
  input  [31:0] io_trigger_pkt_any_1_tdata2,
  input         io_trigger_pkt_any_2_select,
  input         io_trigger_pkt_any_2_match_pkt,
  input         io_trigger_pkt_any_2_store,
  input         io_trigger_pkt_any_2_load,
  input  [31:0] io_trigger_pkt_any_2_tdata2,
  input         io_trigger_pkt_any_3_select,
  input         io_trigger_pkt_any_3_match_pkt,
  input         io_trigger_pkt_any_3_store,
  input         io_trigger_pkt_any_3_load,
  input  [31:0] io_trigger_pkt_any_3_tdata2,
  input         io_lsu_pkt_m_valid,
  input         io_lsu_pkt_m_bits_half,
  input         io_lsu_pkt_m_bits_word,
  input         io_lsu_pkt_m_bits_load,
  input         io_lsu_pkt_m_bits_store,
  input         io_lsu_pkt_m_bits_dma,
  input  [31:0] io_lsu_addr_m,
  input  [31:0] io_store_data_m,
  output [3:0]  io_lsu_trigger_match_m
);
  wire [15:0] _T_1 = io_lsu_pkt_m_bits_word ? 16'hffff : 16'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _T_3 = _T_1 & io_store_data_m[31:16]; // @[lsu_trigger.scala 16:66]
  wire  _T_4 = io_lsu_pkt_m_bits_half | io_lsu_pkt_m_bits_word; // @[lsu_trigger.scala 16:124]
  wire [7:0] _T_6 = _T_4 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_8 = _T_6 & io_store_data_m[15:8]; // @[lsu_trigger.scala 16:151]
  wire [31:0] store_data_trigger_m = {_T_3,_T_8,io_store_data_m[7:0]}; // @[Cat.scala 29:58]
  wire  _T_12 = ~io_trigger_pkt_any_0_select; // @[lsu_trigger.scala 17:53]
  wire  _T_13 = io_trigger_pkt_any_0_select & io_trigger_pkt_any_0_store; // @[lsu_trigger.scala 17:136]
  wire [31:0] _T_15 = _T_12 ? io_lsu_addr_m : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_16 = _T_13 ? store_data_trigger_m : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] lsu_match_data_0 = _T_15 | _T_16; // @[Mux.scala 27:72]
  wire  _T_19 = ~io_trigger_pkt_any_1_select; // @[lsu_trigger.scala 17:53]
  wire  _T_20 = io_trigger_pkt_any_1_select & io_trigger_pkt_any_1_store; // @[lsu_trigger.scala 17:136]
  wire [31:0] _T_22 = _T_19 ? io_lsu_addr_m : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_23 = _T_20 ? store_data_trigger_m : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] lsu_match_data_1 = _T_22 | _T_23; // @[Mux.scala 27:72]
  wire  _T_26 = ~io_trigger_pkt_any_2_select; // @[lsu_trigger.scala 17:53]
  wire  _T_27 = io_trigger_pkt_any_2_select & io_trigger_pkt_any_2_store; // @[lsu_trigger.scala 17:136]
  wire [31:0] _T_29 = _T_26 ? io_lsu_addr_m : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_30 = _T_27 ? store_data_trigger_m : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] lsu_match_data_2 = _T_29 | _T_30; // @[Mux.scala 27:72]
  wire  _T_33 = ~io_trigger_pkt_any_3_select; // @[lsu_trigger.scala 17:53]
  wire  _T_34 = io_trigger_pkt_any_3_select & io_trigger_pkt_any_3_store; // @[lsu_trigger.scala 17:136]
  wire [31:0] _T_36 = _T_33 ? io_lsu_addr_m : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_37 = _T_34 ? store_data_trigger_m : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] lsu_match_data_3 = _T_36 | _T_37; // @[Mux.scala 27:72]
  wire  _T_39 = ~io_lsu_pkt_m_bits_dma; // @[lsu_trigger.scala 18:71]
  wire  _T_40 = io_lsu_pkt_m_valid & _T_39; // @[lsu_trigger.scala 18:69]
  wire  _T_41 = io_trigger_pkt_any_0_store & io_lsu_pkt_m_bits_store; // @[lsu_trigger.scala 18:126]
  wire  _T_42 = io_trigger_pkt_any_0_load & io_lsu_pkt_m_bits_load; // @[lsu_trigger.scala 19:33]
  wire  _T_44 = _T_42 & _T_12; // @[lsu_trigger.scala 19:58]
  wire  _T_45 = _T_41 | _T_44; // @[lsu_trigger.scala 18:152]
  wire  _T_46 = _T_40 & _T_45; // @[lsu_trigger.scala 18:94]
  wire  _T_49 = &io_trigger_pkt_any_0_tdata2; // @[lib.scala 101:45]
  wire  _T_50 = ~_T_49; // @[lib.scala 101:39]
  wire  _T_51 = io_trigger_pkt_any_0_match_pkt & _T_50; // @[lib.scala 101:37]
  wire  _T_54 = io_trigger_pkt_any_0_tdata2[0] == lsu_match_data_0[0]; // @[lib.scala 102:52]
  wire  _T_55 = _T_51 | _T_54; // @[lib.scala 102:41]
  wire  _T_57 = &io_trigger_pkt_any_0_tdata2[0]; // @[lib.scala 104:36]
  wire  _T_58 = _T_57 & _T_51; // @[lib.scala 104:41]
  wire  _T_61 = io_trigger_pkt_any_0_tdata2[1] == lsu_match_data_0[1]; // @[lib.scala 104:78]
  wire  _T_62 = _T_58 | _T_61; // @[lib.scala 104:23]
  wire  _T_64 = &io_trigger_pkt_any_0_tdata2[1:0]; // @[lib.scala 104:36]
  wire  _T_65 = _T_64 & _T_51; // @[lib.scala 104:41]
  wire  _T_68 = io_trigger_pkt_any_0_tdata2[2] == lsu_match_data_0[2]; // @[lib.scala 104:78]
  wire  _T_69 = _T_65 | _T_68; // @[lib.scala 104:23]
  wire  _T_71 = &io_trigger_pkt_any_0_tdata2[2:0]; // @[lib.scala 104:36]
  wire  _T_72 = _T_71 & _T_51; // @[lib.scala 104:41]
  wire  _T_75 = io_trigger_pkt_any_0_tdata2[3] == lsu_match_data_0[3]; // @[lib.scala 104:78]
  wire  _T_76 = _T_72 | _T_75; // @[lib.scala 104:23]
  wire  _T_78 = &io_trigger_pkt_any_0_tdata2[3:0]; // @[lib.scala 104:36]
  wire  _T_79 = _T_78 & _T_51; // @[lib.scala 104:41]
  wire  _T_82 = io_trigger_pkt_any_0_tdata2[4] == lsu_match_data_0[4]; // @[lib.scala 104:78]
  wire  _T_83 = _T_79 | _T_82; // @[lib.scala 104:23]
  wire  _T_85 = &io_trigger_pkt_any_0_tdata2[4:0]; // @[lib.scala 104:36]
  wire  _T_86 = _T_85 & _T_51; // @[lib.scala 104:41]
  wire  _T_89 = io_trigger_pkt_any_0_tdata2[5] == lsu_match_data_0[5]; // @[lib.scala 104:78]
  wire  _T_90 = _T_86 | _T_89; // @[lib.scala 104:23]
  wire  _T_92 = &io_trigger_pkt_any_0_tdata2[5:0]; // @[lib.scala 104:36]
  wire  _T_93 = _T_92 & _T_51; // @[lib.scala 104:41]
  wire  _T_96 = io_trigger_pkt_any_0_tdata2[6] == lsu_match_data_0[6]; // @[lib.scala 104:78]
  wire  _T_97 = _T_93 | _T_96; // @[lib.scala 104:23]
  wire  _T_99 = &io_trigger_pkt_any_0_tdata2[6:0]; // @[lib.scala 104:36]
  wire  _T_100 = _T_99 & _T_51; // @[lib.scala 104:41]
  wire  _T_103 = io_trigger_pkt_any_0_tdata2[7] == lsu_match_data_0[7]; // @[lib.scala 104:78]
  wire  _T_104 = _T_100 | _T_103; // @[lib.scala 104:23]
  wire  _T_106 = &io_trigger_pkt_any_0_tdata2[7:0]; // @[lib.scala 104:36]
  wire  _T_107 = _T_106 & _T_51; // @[lib.scala 104:41]
  wire  _T_110 = io_trigger_pkt_any_0_tdata2[8] == lsu_match_data_0[8]; // @[lib.scala 104:78]
  wire  _T_111 = _T_107 | _T_110; // @[lib.scala 104:23]
  wire  _T_113 = &io_trigger_pkt_any_0_tdata2[8:0]; // @[lib.scala 104:36]
  wire  _T_114 = _T_113 & _T_51; // @[lib.scala 104:41]
  wire  _T_117 = io_trigger_pkt_any_0_tdata2[9] == lsu_match_data_0[9]; // @[lib.scala 104:78]
  wire  _T_118 = _T_114 | _T_117; // @[lib.scala 104:23]
  wire  _T_120 = &io_trigger_pkt_any_0_tdata2[9:0]; // @[lib.scala 104:36]
  wire  _T_121 = _T_120 & _T_51; // @[lib.scala 104:41]
  wire  _T_124 = io_trigger_pkt_any_0_tdata2[10] == lsu_match_data_0[10]; // @[lib.scala 104:78]
  wire  _T_125 = _T_121 | _T_124; // @[lib.scala 104:23]
  wire  _T_127 = &io_trigger_pkt_any_0_tdata2[10:0]; // @[lib.scala 104:36]
  wire  _T_128 = _T_127 & _T_51; // @[lib.scala 104:41]
  wire  _T_131 = io_trigger_pkt_any_0_tdata2[11] == lsu_match_data_0[11]; // @[lib.scala 104:78]
  wire  _T_132 = _T_128 | _T_131; // @[lib.scala 104:23]
  wire  _T_134 = &io_trigger_pkt_any_0_tdata2[11:0]; // @[lib.scala 104:36]
  wire  _T_135 = _T_134 & _T_51; // @[lib.scala 104:41]
  wire  _T_138 = io_trigger_pkt_any_0_tdata2[12] == lsu_match_data_0[12]; // @[lib.scala 104:78]
  wire  _T_139 = _T_135 | _T_138; // @[lib.scala 104:23]
  wire  _T_141 = &io_trigger_pkt_any_0_tdata2[12:0]; // @[lib.scala 104:36]
  wire  _T_142 = _T_141 & _T_51; // @[lib.scala 104:41]
  wire  _T_145 = io_trigger_pkt_any_0_tdata2[13] == lsu_match_data_0[13]; // @[lib.scala 104:78]
  wire  _T_146 = _T_142 | _T_145; // @[lib.scala 104:23]
  wire  _T_148 = &io_trigger_pkt_any_0_tdata2[13:0]; // @[lib.scala 104:36]
  wire  _T_149 = _T_148 & _T_51; // @[lib.scala 104:41]
  wire  _T_152 = io_trigger_pkt_any_0_tdata2[14] == lsu_match_data_0[14]; // @[lib.scala 104:78]
  wire  _T_153 = _T_149 | _T_152; // @[lib.scala 104:23]
  wire  _T_155 = &io_trigger_pkt_any_0_tdata2[14:0]; // @[lib.scala 104:36]
  wire  _T_156 = _T_155 & _T_51; // @[lib.scala 104:41]
  wire  _T_159 = io_trigger_pkt_any_0_tdata2[15] == lsu_match_data_0[15]; // @[lib.scala 104:78]
  wire  _T_160 = _T_156 | _T_159; // @[lib.scala 104:23]
  wire  _T_162 = &io_trigger_pkt_any_0_tdata2[15:0]; // @[lib.scala 104:36]
  wire  _T_163 = _T_162 & _T_51; // @[lib.scala 104:41]
  wire  _T_166 = io_trigger_pkt_any_0_tdata2[16] == lsu_match_data_0[16]; // @[lib.scala 104:78]
  wire  _T_167 = _T_163 | _T_166; // @[lib.scala 104:23]
  wire  _T_169 = &io_trigger_pkt_any_0_tdata2[16:0]; // @[lib.scala 104:36]
  wire  _T_170 = _T_169 & _T_51; // @[lib.scala 104:41]
  wire  _T_173 = io_trigger_pkt_any_0_tdata2[17] == lsu_match_data_0[17]; // @[lib.scala 104:78]
  wire  _T_174 = _T_170 | _T_173; // @[lib.scala 104:23]
  wire  _T_176 = &io_trigger_pkt_any_0_tdata2[17:0]; // @[lib.scala 104:36]
  wire  _T_177 = _T_176 & _T_51; // @[lib.scala 104:41]
  wire  _T_180 = io_trigger_pkt_any_0_tdata2[18] == lsu_match_data_0[18]; // @[lib.scala 104:78]
  wire  _T_181 = _T_177 | _T_180; // @[lib.scala 104:23]
  wire  _T_183 = &io_trigger_pkt_any_0_tdata2[18:0]; // @[lib.scala 104:36]
  wire  _T_184 = _T_183 & _T_51; // @[lib.scala 104:41]
  wire  _T_187 = io_trigger_pkt_any_0_tdata2[19] == lsu_match_data_0[19]; // @[lib.scala 104:78]
  wire  _T_188 = _T_184 | _T_187; // @[lib.scala 104:23]
  wire  _T_190 = &io_trigger_pkt_any_0_tdata2[19:0]; // @[lib.scala 104:36]
  wire  _T_191 = _T_190 & _T_51; // @[lib.scala 104:41]
  wire  _T_194 = io_trigger_pkt_any_0_tdata2[20] == lsu_match_data_0[20]; // @[lib.scala 104:78]
  wire  _T_195 = _T_191 | _T_194; // @[lib.scala 104:23]
  wire  _T_197 = &io_trigger_pkt_any_0_tdata2[20:0]; // @[lib.scala 104:36]
  wire  _T_198 = _T_197 & _T_51; // @[lib.scala 104:41]
  wire  _T_201 = io_trigger_pkt_any_0_tdata2[21] == lsu_match_data_0[21]; // @[lib.scala 104:78]
  wire  _T_202 = _T_198 | _T_201; // @[lib.scala 104:23]
  wire  _T_204 = &io_trigger_pkt_any_0_tdata2[21:0]; // @[lib.scala 104:36]
  wire  _T_205 = _T_204 & _T_51; // @[lib.scala 104:41]
  wire  _T_208 = io_trigger_pkt_any_0_tdata2[22] == lsu_match_data_0[22]; // @[lib.scala 104:78]
  wire  _T_209 = _T_205 | _T_208; // @[lib.scala 104:23]
  wire  _T_211 = &io_trigger_pkt_any_0_tdata2[22:0]; // @[lib.scala 104:36]
  wire  _T_212 = _T_211 & _T_51; // @[lib.scala 104:41]
  wire  _T_215 = io_trigger_pkt_any_0_tdata2[23] == lsu_match_data_0[23]; // @[lib.scala 104:78]
  wire  _T_216 = _T_212 | _T_215; // @[lib.scala 104:23]
  wire  _T_218 = &io_trigger_pkt_any_0_tdata2[23:0]; // @[lib.scala 104:36]
  wire  _T_219 = _T_218 & _T_51; // @[lib.scala 104:41]
  wire  _T_222 = io_trigger_pkt_any_0_tdata2[24] == lsu_match_data_0[24]; // @[lib.scala 104:78]
  wire  _T_223 = _T_219 | _T_222; // @[lib.scala 104:23]
  wire  _T_225 = &io_trigger_pkt_any_0_tdata2[24:0]; // @[lib.scala 104:36]
  wire  _T_226 = _T_225 & _T_51; // @[lib.scala 104:41]
  wire  _T_229 = io_trigger_pkt_any_0_tdata2[25] == lsu_match_data_0[25]; // @[lib.scala 104:78]
  wire  _T_230 = _T_226 | _T_229; // @[lib.scala 104:23]
  wire  _T_232 = &io_trigger_pkt_any_0_tdata2[25:0]; // @[lib.scala 104:36]
  wire  _T_233 = _T_232 & _T_51; // @[lib.scala 104:41]
  wire  _T_236 = io_trigger_pkt_any_0_tdata2[26] == lsu_match_data_0[26]; // @[lib.scala 104:78]
  wire  _T_237 = _T_233 | _T_236; // @[lib.scala 104:23]
  wire  _T_239 = &io_trigger_pkt_any_0_tdata2[26:0]; // @[lib.scala 104:36]
  wire  _T_240 = _T_239 & _T_51; // @[lib.scala 104:41]
  wire  _T_243 = io_trigger_pkt_any_0_tdata2[27] == lsu_match_data_0[27]; // @[lib.scala 104:78]
  wire  _T_244 = _T_240 | _T_243; // @[lib.scala 104:23]
  wire  _T_246 = &io_trigger_pkt_any_0_tdata2[27:0]; // @[lib.scala 104:36]
  wire  _T_247 = _T_246 & _T_51; // @[lib.scala 104:41]
  wire  _T_250 = io_trigger_pkt_any_0_tdata2[28] == lsu_match_data_0[28]; // @[lib.scala 104:78]
  wire  _T_251 = _T_247 | _T_250; // @[lib.scala 104:23]
  wire  _T_253 = &io_trigger_pkt_any_0_tdata2[28:0]; // @[lib.scala 104:36]
  wire  _T_254 = _T_253 & _T_51; // @[lib.scala 104:41]
  wire  _T_257 = io_trigger_pkt_any_0_tdata2[29] == lsu_match_data_0[29]; // @[lib.scala 104:78]
  wire  _T_258 = _T_254 | _T_257; // @[lib.scala 104:23]
  wire  _T_260 = &io_trigger_pkt_any_0_tdata2[29:0]; // @[lib.scala 104:36]
  wire  _T_261 = _T_260 & _T_51; // @[lib.scala 104:41]
  wire  _T_264 = io_trigger_pkt_any_0_tdata2[30] == lsu_match_data_0[30]; // @[lib.scala 104:78]
  wire  _T_265 = _T_261 | _T_264; // @[lib.scala 104:23]
  wire  _T_267 = &io_trigger_pkt_any_0_tdata2[30:0]; // @[lib.scala 104:36]
  wire  _T_268 = _T_267 & _T_51; // @[lib.scala 104:41]
  wire  _T_271 = io_trigger_pkt_any_0_tdata2[31] == lsu_match_data_0[31]; // @[lib.scala 104:78]
  wire  _T_272 = _T_268 | _T_271; // @[lib.scala 104:23]
  wire [7:0] _T_279 = {_T_104,_T_97,_T_90,_T_83,_T_76,_T_69,_T_62,_T_55}; // @[lib.scala 105:14]
  wire [15:0] _T_287 = {_T_160,_T_153,_T_146,_T_139,_T_132,_T_125,_T_118,_T_111,_T_279}; // @[lib.scala 105:14]
  wire [7:0] _T_294 = {_T_216,_T_209,_T_202,_T_195,_T_188,_T_181,_T_174,_T_167}; // @[lib.scala 105:14]
  wire [31:0] _T_303 = {_T_272,_T_265,_T_258,_T_251,_T_244,_T_237,_T_230,_T_223,_T_294,_T_287}; // @[lib.scala 105:14]
  wire  _T_304 = &_T_303; // @[lib.scala 105:25]
  wire  _T_305 = _T_46 & _T_304; // @[lsu_trigger.scala 19:92]
  wire  _T_308 = io_trigger_pkt_any_1_store & io_lsu_pkt_m_bits_store; // @[lsu_trigger.scala 18:126]
  wire  _T_309 = io_trigger_pkt_any_1_load & io_lsu_pkt_m_bits_load; // @[lsu_trigger.scala 19:33]
  wire  _T_311 = _T_309 & _T_19; // @[lsu_trigger.scala 19:58]
  wire  _T_312 = _T_308 | _T_311; // @[lsu_trigger.scala 18:152]
  wire  _T_313 = _T_40 & _T_312; // @[lsu_trigger.scala 18:94]
  wire  _T_316 = &io_trigger_pkt_any_1_tdata2; // @[lib.scala 101:45]
  wire  _T_317 = ~_T_316; // @[lib.scala 101:39]
  wire  _T_318 = io_trigger_pkt_any_1_match_pkt & _T_317; // @[lib.scala 101:37]
  wire  _T_321 = io_trigger_pkt_any_1_tdata2[0] == lsu_match_data_1[0]; // @[lib.scala 102:52]
  wire  _T_322 = _T_318 | _T_321; // @[lib.scala 102:41]
  wire  _T_324 = &io_trigger_pkt_any_1_tdata2[0]; // @[lib.scala 104:36]
  wire  _T_325 = _T_324 & _T_318; // @[lib.scala 104:41]
  wire  _T_328 = io_trigger_pkt_any_1_tdata2[1] == lsu_match_data_1[1]; // @[lib.scala 104:78]
  wire  _T_329 = _T_325 | _T_328; // @[lib.scala 104:23]
  wire  _T_331 = &io_trigger_pkt_any_1_tdata2[1:0]; // @[lib.scala 104:36]
  wire  _T_332 = _T_331 & _T_318; // @[lib.scala 104:41]
  wire  _T_335 = io_trigger_pkt_any_1_tdata2[2] == lsu_match_data_1[2]; // @[lib.scala 104:78]
  wire  _T_336 = _T_332 | _T_335; // @[lib.scala 104:23]
  wire  _T_338 = &io_trigger_pkt_any_1_tdata2[2:0]; // @[lib.scala 104:36]
  wire  _T_339 = _T_338 & _T_318; // @[lib.scala 104:41]
  wire  _T_342 = io_trigger_pkt_any_1_tdata2[3] == lsu_match_data_1[3]; // @[lib.scala 104:78]
  wire  _T_343 = _T_339 | _T_342; // @[lib.scala 104:23]
  wire  _T_345 = &io_trigger_pkt_any_1_tdata2[3:0]; // @[lib.scala 104:36]
  wire  _T_346 = _T_345 & _T_318; // @[lib.scala 104:41]
  wire  _T_349 = io_trigger_pkt_any_1_tdata2[4] == lsu_match_data_1[4]; // @[lib.scala 104:78]
  wire  _T_350 = _T_346 | _T_349; // @[lib.scala 104:23]
  wire  _T_352 = &io_trigger_pkt_any_1_tdata2[4:0]; // @[lib.scala 104:36]
  wire  _T_353 = _T_352 & _T_318; // @[lib.scala 104:41]
  wire  _T_356 = io_trigger_pkt_any_1_tdata2[5] == lsu_match_data_1[5]; // @[lib.scala 104:78]
  wire  _T_357 = _T_353 | _T_356; // @[lib.scala 104:23]
  wire  _T_359 = &io_trigger_pkt_any_1_tdata2[5:0]; // @[lib.scala 104:36]
  wire  _T_360 = _T_359 & _T_318; // @[lib.scala 104:41]
  wire  _T_363 = io_trigger_pkt_any_1_tdata2[6] == lsu_match_data_1[6]; // @[lib.scala 104:78]
  wire  _T_364 = _T_360 | _T_363; // @[lib.scala 104:23]
  wire  _T_366 = &io_trigger_pkt_any_1_tdata2[6:0]; // @[lib.scala 104:36]
  wire  _T_367 = _T_366 & _T_318; // @[lib.scala 104:41]
  wire  _T_370 = io_trigger_pkt_any_1_tdata2[7] == lsu_match_data_1[7]; // @[lib.scala 104:78]
  wire  _T_371 = _T_367 | _T_370; // @[lib.scala 104:23]
  wire  _T_373 = &io_trigger_pkt_any_1_tdata2[7:0]; // @[lib.scala 104:36]
  wire  _T_374 = _T_373 & _T_318; // @[lib.scala 104:41]
  wire  _T_377 = io_trigger_pkt_any_1_tdata2[8] == lsu_match_data_1[8]; // @[lib.scala 104:78]
  wire  _T_378 = _T_374 | _T_377; // @[lib.scala 104:23]
  wire  _T_380 = &io_trigger_pkt_any_1_tdata2[8:0]; // @[lib.scala 104:36]
  wire  _T_381 = _T_380 & _T_318; // @[lib.scala 104:41]
  wire  _T_384 = io_trigger_pkt_any_1_tdata2[9] == lsu_match_data_1[9]; // @[lib.scala 104:78]
  wire  _T_385 = _T_381 | _T_384; // @[lib.scala 104:23]
  wire  _T_387 = &io_trigger_pkt_any_1_tdata2[9:0]; // @[lib.scala 104:36]
  wire  _T_388 = _T_387 & _T_318; // @[lib.scala 104:41]
  wire  _T_391 = io_trigger_pkt_any_1_tdata2[10] == lsu_match_data_1[10]; // @[lib.scala 104:78]
  wire  _T_392 = _T_388 | _T_391; // @[lib.scala 104:23]
  wire  _T_394 = &io_trigger_pkt_any_1_tdata2[10:0]; // @[lib.scala 104:36]
  wire  _T_395 = _T_394 & _T_318; // @[lib.scala 104:41]
  wire  _T_398 = io_trigger_pkt_any_1_tdata2[11] == lsu_match_data_1[11]; // @[lib.scala 104:78]
  wire  _T_399 = _T_395 | _T_398; // @[lib.scala 104:23]
  wire  _T_401 = &io_trigger_pkt_any_1_tdata2[11:0]; // @[lib.scala 104:36]
  wire  _T_402 = _T_401 & _T_318; // @[lib.scala 104:41]
  wire  _T_405 = io_trigger_pkt_any_1_tdata2[12] == lsu_match_data_1[12]; // @[lib.scala 104:78]
  wire  _T_406 = _T_402 | _T_405; // @[lib.scala 104:23]
  wire  _T_408 = &io_trigger_pkt_any_1_tdata2[12:0]; // @[lib.scala 104:36]
  wire  _T_409 = _T_408 & _T_318; // @[lib.scala 104:41]
  wire  _T_412 = io_trigger_pkt_any_1_tdata2[13] == lsu_match_data_1[13]; // @[lib.scala 104:78]
  wire  _T_413 = _T_409 | _T_412; // @[lib.scala 104:23]
  wire  _T_415 = &io_trigger_pkt_any_1_tdata2[13:0]; // @[lib.scala 104:36]
  wire  _T_416 = _T_415 & _T_318; // @[lib.scala 104:41]
  wire  _T_419 = io_trigger_pkt_any_1_tdata2[14] == lsu_match_data_1[14]; // @[lib.scala 104:78]
  wire  _T_420 = _T_416 | _T_419; // @[lib.scala 104:23]
  wire  _T_422 = &io_trigger_pkt_any_1_tdata2[14:0]; // @[lib.scala 104:36]
  wire  _T_423 = _T_422 & _T_318; // @[lib.scala 104:41]
  wire  _T_426 = io_trigger_pkt_any_1_tdata2[15] == lsu_match_data_1[15]; // @[lib.scala 104:78]
  wire  _T_427 = _T_423 | _T_426; // @[lib.scala 104:23]
  wire  _T_429 = &io_trigger_pkt_any_1_tdata2[15:0]; // @[lib.scala 104:36]
  wire  _T_430 = _T_429 & _T_318; // @[lib.scala 104:41]
  wire  _T_433 = io_trigger_pkt_any_1_tdata2[16] == lsu_match_data_1[16]; // @[lib.scala 104:78]
  wire  _T_434 = _T_430 | _T_433; // @[lib.scala 104:23]
  wire  _T_436 = &io_trigger_pkt_any_1_tdata2[16:0]; // @[lib.scala 104:36]
  wire  _T_437 = _T_436 & _T_318; // @[lib.scala 104:41]
  wire  _T_440 = io_trigger_pkt_any_1_tdata2[17] == lsu_match_data_1[17]; // @[lib.scala 104:78]
  wire  _T_441 = _T_437 | _T_440; // @[lib.scala 104:23]
  wire  _T_443 = &io_trigger_pkt_any_1_tdata2[17:0]; // @[lib.scala 104:36]
  wire  _T_444 = _T_443 & _T_318; // @[lib.scala 104:41]
  wire  _T_447 = io_trigger_pkt_any_1_tdata2[18] == lsu_match_data_1[18]; // @[lib.scala 104:78]
  wire  _T_448 = _T_444 | _T_447; // @[lib.scala 104:23]
  wire  _T_450 = &io_trigger_pkt_any_1_tdata2[18:0]; // @[lib.scala 104:36]
  wire  _T_451 = _T_450 & _T_318; // @[lib.scala 104:41]
  wire  _T_454 = io_trigger_pkt_any_1_tdata2[19] == lsu_match_data_1[19]; // @[lib.scala 104:78]
  wire  _T_455 = _T_451 | _T_454; // @[lib.scala 104:23]
  wire  _T_457 = &io_trigger_pkt_any_1_tdata2[19:0]; // @[lib.scala 104:36]
  wire  _T_458 = _T_457 & _T_318; // @[lib.scala 104:41]
  wire  _T_461 = io_trigger_pkt_any_1_tdata2[20] == lsu_match_data_1[20]; // @[lib.scala 104:78]
  wire  _T_462 = _T_458 | _T_461; // @[lib.scala 104:23]
  wire  _T_464 = &io_trigger_pkt_any_1_tdata2[20:0]; // @[lib.scala 104:36]
  wire  _T_465 = _T_464 & _T_318; // @[lib.scala 104:41]
  wire  _T_468 = io_trigger_pkt_any_1_tdata2[21] == lsu_match_data_1[21]; // @[lib.scala 104:78]
  wire  _T_469 = _T_465 | _T_468; // @[lib.scala 104:23]
  wire  _T_471 = &io_trigger_pkt_any_1_tdata2[21:0]; // @[lib.scala 104:36]
  wire  _T_472 = _T_471 & _T_318; // @[lib.scala 104:41]
  wire  _T_475 = io_trigger_pkt_any_1_tdata2[22] == lsu_match_data_1[22]; // @[lib.scala 104:78]
  wire  _T_476 = _T_472 | _T_475; // @[lib.scala 104:23]
  wire  _T_478 = &io_trigger_pkt_any_1_tdata2[22:0]; // @[lib.scala 104:36]
  wire  _T_479 = _T_478 & _T_318; // @[lib.scala 104:41]
  wire  _T_482 = io_trigger_pkt_any_1_tdata2[23] == lsu_match_data_1[23]; // @[lib.scala 104:78]
  wire  _T_483 = _T_479 | _T_482; // @[lib.scala 104:23]
  wire  _T_485 = &io_trigger_pkt_any_1_tdata2[23:0]; // @[lib.scala 104:36]
  wire  _T_486 = _T_485 & _T_318; // @[lib.scala 104:41]
  wire  _T_489 = io_trigger_pkt_any_1_tdata2[24] == lsu_match_data_1[24]; // @[lib.scala 104:78]
  wire  _T_490 = _T_486 | _T_489; // @[lib.scala 104:23]
  wire  _T_492 = &io_trigger_pkt_any_1_tdata2[24:0]; // @[lib.scala 104:36]
  wire  _T_493 = _T_492 & _T_318; // @[lib.scala 104:41]
  wire  _T_496 = io_trigger_pkt_any_1_tdata2[25] == lsu_match_data_1[25]; // @[lib.scala 104:78]
  wire  _T_497 = _T_493 | _T_496; // @[lib.scala 104:23]
  wire  _T_499 = &io_trigger_pkt_any_1_tdata2[25:0]; // @[lib.scala 104:36]
  wire  _T_500 = _T_499 & _T_318; // @[lib.scala 104:41]
  wire  _T_503 = io_trigger_pkt_any_1_tdata2[26] == lsu_match_data_1[26]; // @[lib.scala 104:78]
  wire  _T_504 = _T_500 | _T_503; // @[lib.scala 104:23]
  wire  _T_506 = &io_trigger_pkt_any_1_tdata2[26:0]; // @[lib.scala 104:36]
  wire  _T_507 = _T_506 & _T_318; // @[lib.scala 104:41]
  wire  _T_510 = io_trigger_pkt_any_1_tdata2[27] == lsu_match_data_1[27]; // @[lib.scala 104:78]
  wire  _T_511 = _T_507 | _T_510; // @[lib.scala 104:23]
  wire  _T_513 = &io_trigger_pkt_any_1_tdata2[27:0]; // @[lib.scala 104:36]
  wire  _T_514 = _T_513 & _T_318; // @[lib.scala 104:41]
  wire  _T_517 = io_trigger_pkt_any_1_tdata2[28] == lsu_match_data_1[28]; // @[lib.scala 104:78]
  wire  _T_518 = _T_514 | _T_517; // @[lib.scala 104:23]
  wire  _T_520 = &io_trigger_pkt_any_1_tdata2[28:0]; // @[lib.scala 104:36]
  wire  _T_521 = _T_520 & _T_318; // @[lib.scala 104:41]
  wire  _T_524 = io_trigger_pkt_any_1_tdata2[29] == lsu_match_data_1[29]; // @[lib.scala 104:78]
  wire  _T_525 = _T_521 | _T_524; // @[lib.scala 104:23]
  wire  _T_527 = &io_trigger_pkt_any_1_tdata2[29:0]; // @[lib.scala 104:36]
  wire  _T_528 = _T_527 & _T_318; // @[lib.scala 104:41]
  wire  _T_531 = io_trigger_pkt_any_1_tdata2[30] == lsu_match_data_1[30]; // @[lib.scala 104:78]
  wire  _T_532 = _T_528 | _T_531; // @[lib.scala 104:23]
  wire  _T_534 = &io_trigger_pkt_any_1_tdata2[30:0]; // @[lib.scala 104:36]
  wire  _T_535 = _T_534 & _T_318; // @[lib.scala 104:41]
  wire  _T_538 = io_trigger_pkt_any_1_tdata2[31] == lsu_match_data_1[31]; // @[lib.scala 104:78]
  wire  _T_539 = _T_535 | _T_538; // @[lib.scala 104:23]
  wire [7:0] _T_546 = {_T_371,_T_364,_T_357,_T_350,_T_343,_T_336,_T_329,_T_322}; // @[lib.scala 105:14]
  wire [15:0] _T_554 = {_T_427,_T_420,_T_413,_T_406,_T_399,_T_392,_T_385,_T_378,_T_546}; // @[lib.scala 105:14]
  wire [7:0] _T_561 = {_T_483,_T_476,_T_469,_T_462,_T_455,_T_448,_T_441,_T_434}; // @[lib.scala 105:14]
  wire [31:0] _T_570 = {_T_539,_T_532,_T_525,_T_518,_T_511,_T_504,_T_497,_T_490,_T_561,_T_554}; // @[lib.scala 105:14]
  wire  _T_571 = &_T_570; // @[lib.scala 105:25]
  wire  _T_572 = _T_313 & _T_571; // @[lsu_trigger.scala 19:92]
  wire  _T_575 = io_trigger_pkt_any_2_store & io_lsu_pkt_m_bits_store; // @[lsu_trigger.scala 18:126]
  wire  _T_576 = io_trigger_pkt_any_2_load & io_lsu_pkt_m_bits_load; // @[lsu_trigger.scala 19:33]
  wire  _T_578 = _T_576 & _T_26; // @[lsu_trigger.scala 19:58]
  wire  _T_579 = _T_575 | _T_578; // @[lsu_trigger.scala 18:152]
  wire  _T_580 = _T_40 & _T_579; // @[lsu_trigger.scala 18:94]
  wire  _T_583 = &io_trigger_pkt_any_2_tdata2; // @[lib.scala 101:45]
  wire  _T_584 = ~_T_583; // @[lib.scala 101:39]
  wire  _T_585 = io_trigger_pkt_any_2_match_pkt & _T_584; // @[lib.scala 101:37]
  wire  _T_588 = io_trigger_pkt_any_2_tdata2[0] == lsu_match_data_2[0]; // @[lib.scala 102:52]
  wire  _T_589 = _T_585 | _T_588; // @[lib.scala 102:41]
  wire  _T_591 = &io_trigger_pkt_any_2_tdata2[0]; // @[lib.scala 104:36]
  wire  _T_592 = _T_591 & _T_585; // @[lib.scala 104:41]
  wire  _T_595 = io_trigger_pkt_any_2_tdata2[1] == lsu_match_data_2[1]; // @[lib.scala 104:78]
  wire  _T_596 = _T_592 | _T_595; // @[lib.scala 104:23]
  wire  _T_598 = &io_trigger_pkt_any_2_tdata2[1:0]; // @[lib.scala 104:36]
  wire  _T_599 = _T_598 & _T_585; // @[lib.scala 104:41]
  wire  _T_602 = io_trigger_pkt_any_2_tdata2[2] == lsu_match_data_2[2]; // @[lib.scala 104:78]
  wire  _T_603 = _T_599 | _T_602; // @[lib.scala 104:23]
  wire  _T_605 = &io_trigger_pkt_any_2_tdata2[2:0]; // @[lib.scala 104:36]
  wire  _T_606 = _T_605 & _T_585; // @[lib.scala 104:41]
  wire  _T_609 = io_trigger_pkt_any_2_tdata2[3] == lsu_match_data_2[3]; // @[lib.scala 104:78]
  wire  _T_610 = _T_606 | _T_609; // @[lib.scala 104:23]
  wire  _T_612 = &io_trigger_pkt_any_2_tdata2[3:0]; // @[lib.scala 104:36]
  wire  _T_613 = _T_612 & _T_585; // @[lib.scala 104:41]
  wire  _T_616 = io_trigger_pkt_any_2_tdata2[4] == lsu_match_data_2[4]; // @[lib.scala 104:78]
  wire  _T_617 = _T_613 | _T_616; // @[lib.scala 104:23]
  wire  _T_619 = &io_trigger_pkt_any_2_tdata2[4:0]; // @[lib.scala 104:36]
  wire  _T_620 = _T_619 & _T_585; // @[lib.scala 104:41]
  wire  _T_623 = io_trigger_pkt_any_2_tdata2[5] == lsu_match_data_2[5]; // @[lib.scala 104:78]
  wire  _T_624 = _T_620 | _T_623; // @[lib.scala 104:23]
  wire  _T_626 = &io_trigger_pkt_any_2_tdata2[5:0]; // @[lib.scala 104:36]
  wire  _T_627 = _T_626 & _T_585; // @[lib.scala 104:41]
  wire  _T_630 = io_trigger_pkt_any_2_tdata2[6] == lsu_match_data_2[6]; // @[lib.scala 104:78]
  wire  _T_631 = _T_627 | _T_630; // @[lib.scala 104:23]
  wire  _T_633 = &io_trigger_pkt_any_2_tdata2[6:0]; // @[lib.scala 104:36]
  wire  _T_634 = _T_633 & _T_585; // @[lib.scala 104:41]
  wire  _T_637 = io_trigger_pkt_any_2_tdata2[7] == lsu_match_data_2[7]; // @[lib.scala 104:78]
  wire  _T_638 = _T_634 | _T_637; // @[lib.scala 104:23]
  wire  _T_640 = &io_trigger_pkt_any_2_tdata2[7:0]; // @[lib.scala 104:36]
  wire  _T_641 = _T_640 & _T_585; // @[lib.scala 104:41]
  wire  _T_644 = io_trigger_pkt_any_2_tdata2[8] == lsu_match_data_2[8]; // @[lib.scala 104:78]
  wire  _T_645 = _T_641 | _T_644; // @[lib.scala 104:23]
  wire  _T_647 = &io_trigger_pkt_any_2_tdata2[8:0]; // @[lib.scala 104:36]
  wire  _T_648 = _T_647 & _T_585; // @[lib.scala 104:41]
  wire  _T_651 = io_trigger_pkt_any_2_tdata2[9] == lsu_match_data_2[9]; // @[lib.scala 104:78]
  wire  _T_652 = _T_648 | _T_651; // @[lib.scala 104:23]
  wire  _T_654 = &io_trigger_pkt_any_2_tdata2[9:0]; // @[lib.scala 104:36]
  wire  _T_655 = _T_654 & _T_585; // @[lib.scala 104:41]
  wire  _T_658 = io_trigger_pkt_any_2_tdata2[10] == lsu_match_data_2[10]; // @[lib.scala 104:78]
  wire  _T_659 = _T_655 | _T_658; // @[lib.scala 104:23]
  wire  _T_661 = &io_trigger_pkt_any_2_tdata2[10:0]; // @[lib.scala 104:36]
  wire  _T_662 = _T_661 & _T_585; // @[lib.scala 104:41]
  wire  _T_665 = io_trigger_pkt_any_2_tdata2[11] == lsu_match_data_2[11]; // @[lib.scala 104:78]
  wire  _T_666 = _T_662 | _T_665; // @[lib.scala 104:23]
  wire  _T_668 = &io_trigger_pkt_any_2_tdata2[11:0]; // @[lib.scala 104:36]
  wire  _T_669 = _T_668 & _T_585; // @[lib.scala 104:41]
  wire  _T_672 = io_trigger_pkt_any_2_tdata2[12] == lsu_match_data_2[12]; // @[lib.scala 104:78]
  wire  _T_673 = _T_669 | _T_672; // @[lib.scala 104:23]
  wire  _T_675 = &io_trigger_pkt_any_2_tdata2[12:0]; // @[lib.scala 104:36]
  wire  _T_676 = _T_675 & _T_585; // @[lib.scala 104:41]
  wire  _T_679 = io_trigger_pkt_any_2_tdata2[13] == lsu_match_data_2[13]; // @[lib.scala 104:78]
  wire  _T_680 = _T_676 | _T_679; // @[lib.scala 104:23]
  wire  _T_682 = &io_trigger_pkt_any_2_tdata2[13:0]; // @[lib.scala 104:36]
  wire  _T_683 = _T_682 & _T_585; // @[lib.scala 104:41]
  wire  _T_686 = io_trigger_pkt_any_2_tdata2[14] == lsu_match_data_2[14]; // @[lib.scala 104:78]
  wire  _T_687 = _T_683 | _T_686; // @[lib.scala 104:23]
  wire  _T_689 = &io_trigger_pkt_any_2_tdata2[14:0]; // @[lib.scala 104:36]
  wire  _T_690 = _T_689 & _T_585; // @[lib.scala 104:41]
  wire  _T_693 = io_trigger_pkt_any_2_tdata2[15] == lsu_match_data_2[15]; // @[lib.scala 104:78]
  wire  _T_694 = _T_690 | _T_693; // @[lib.scala 104:23]
  wire  _T_696 = &io_trigger_pkt_any_2_tdata2[15:0]; // @[lib.scala 104:36]
  wire  _T_697 = _T_696 & _T_585; // @[lib.scala 104:41]
  wire  _T_700 = io_trigger_pkt_any_2_tdata2[16] == lsu_match_data_2[16]; // @[lib.scala 104:78]
  wire  _T_701 = _T_697 | _T_700; // @[lib.scala 104:23]
  wire  _T_703 = &io_trigger_pkt_any_2_tdata2[16:0]; // @[lib.scala 104:36]
  wire  _T_704 = _T_703 & _T_585; // @[lib.scala 104:41]
  wire  _T_707 = io_trigger_pkt_any_2_tdata2[17] == lsu_match_data_2[17]; // @[lib.scala 104:78]
  wire  _T_708 = _T_704 | _T_707; // @[lib.scala 104:23]
  wire  _T_710 = &io_trigger_pkt_any_2_tdata2[17:0]; // @[lib.scala 104:36]
  wire  _T_711 = _T_710 & _T_585; // @[lib.scala 104:41]
  wire  _T_714 = io_trigger_pkt_any_2_tdata2[18] == lsu_match_data_2[18]; // @[lib.scala 104:78]
  wire  _T_715 = _T_711 | _T_714; // @[lib.scala 104:23]
  wire  _T_717 = &io_trigger_pkt_any_2_tdata2[18:0]; // @[lib.scala 104:36]
  wire  _T_718 = _T_717 & _T_585; // @[lib.scala 104:41]
  wire  _T_721 = io_trigger_pkt_any_2_tdata2[19] == lsu_match_data_2[19]; // @[lib.scala 104:78]
  wire  _T_722 = _T_718 | _T_721; // @[lib.scala 104:23]
  wire  _T_724 = &io_trigger_pkt_any_2_tdata2[19:0]; // @[lib.scala 104:36]
  wire  _T_725 = _T_724 & _T_585; // @[lib.scala 104:41]
  wire  _T_728 = io_trigger_pkt_any_2_tdata2[20] == lsu_match_data_2[20]; // @[lib.scala 104:78]
  wire  _T_729 = _T_725 | _T_728; // @[lib.scala 104:23]
  wire  _T_731 = &io_trigger_pkt_any_2_tdata2[20:0]; // @[lib.scala 104:36]
  wire  _T_732 = _T_731 & _T_585; // @[lib.scala 104:41]
  wire  _T_735 = io_trigger_pkt_any_2_tdata2[21] == lsu_match_data_2[21]; // @[lib.scala 104:78]
  wire  _T_736 = _T_732 | _T_735; // @[lib.scala 104:23]
  wire  _T_738 = &io_trigger_pkt_any_2_tdata2[21:0]; // @[lib.scala 104:36]
  wire  _T_739 = _T_738 & _T_585; // @[lib.scala 104:41]
  wire  _T_742 = io_trigger_pkt_any_2_tdata2[22] == lsu_match_data_2[22]; // @[lib.scala 104:78]
  wire  _T_743 = _T_739 | _T_742; // @[lib.scala 104:23]
  wire  _T_745 = &io_trigger_pkt_any_2_tdata2[22:0]; // @[lib.scala 104:36]
  wire  _T_746 = _T_745 & _T_585; // @[lib.scala 104:41]
  wire  _T_749 = io_trigger_pkt_any_2_tdata2[23] == lsu_match_data_2[23]; // @[lib.scala 104:78]
  wire  _T_750 = _T_746 | _T_749; // @[lib.scala 104:23]
  wire  _T_752 = &io_trigger_pkt_any_2_tdata2[23:0]; // @[lib.scala 104:36]
  wire  _T_753 = _T_752 & _T_585; // @[lib.scala 104:41]
  wire  _T_756 = io_trigger_pkt_any_2_tdata2[24] == lsu_match_data_2[24]; // @[lib.scala 104:78]
  wire  _T_757 = _T_753 | _T_756; // @[lib.scala 104:23]
  wire  _T_759 = &io_trigger_pkt_any_2_tdata2[24:0]; // @[lib.scala 104:36]
  wire  _T_760 = _T_759 & _T_585; // @[lib.scala 104:41]
  wire  _T_763 = io_trigger_pkt_any_2_tdata2[25] == lsu_match_data_2[25]; // @[lib.scala 104:78]
  wire  _T_764 = _T_760 | _T_763; // @[lib.scala 104:23]
  wire  _T_766 = &io_trigger_pkt_any_2_tdata2[25:0]; // @[lib.scala 104:36]
  wire  _T_767 = _T_766 & _T_585; // @[lib.scala 104:41]
  wire  _T_770 = io_trigger_pkt_any_2_tdata2[26] == lsu_match_data_2[26]; // @[lib.scala 104:78]
  wire  _T_771 = _T_767 | _T_770; // @[lib.scala 104:23]
  wire  _T_773 = &io_trigger_pkt_any_2_tdata2[26:0]; // @[lib.scala 104:36]
  wire  _T_774 = _T_773 & _T_585; // @[lib.scala 104:41]
  wire  _T_777 = io_trigger_pkt_any_2_tdata2[27] == lsu_match_data_2[27]; // @[lib.scala 104:78]
  wire  _T_778 = _T_774 | _T_777; // @[lib.scala 104:23]
  wire  _T_780 = &io_trigger_pkt_any_2_tdata2[27:0]; // @[lib.scala 104:36]
  wire  _T_781 = _T_780 & _T_585; // @[lib.scala 104:41]
  wire  _T_784 = io_trigger_pkt_any_2_tdata2[28] == lsu_match_data_2[28]; // @[lib.scala 104:78]
  wire  _T_785 = _T_781 | _T_784; // @[lib.scala 104:23]
  wire  _T_787 = &io_trigger_pkt_any_2_tdata2[28:0]; // @[lib.scala 104:36]
  wire  _T_788 = _T_787 & _T_585; // @[lib.scala 104:41]
  wire  _T_791 = io_trigger_pkt_any_2_tdata2[29] == lsu_match_data_2[29]; // @[lib.scala 104:78]
  wire  _T_792 = _T_788 | _T_791; // @[lib.scala 104:23]
  wire  _T_794 = &io_trigger_pkt_any_2_tdata2[29:0]; // @[lib.scala 104:36]
  wire  _T_795 = _T_794 & _T_585; // @[lib.scala 104:41]
  wire  _T_798 = io_trigger_pkt_any_2_tdata2[30] == lsu_match_data_2[30]; // @[lib.scala 104:78]
  wire  _T_799 = _T_795 | _T_798; // @[lib.scala 104:23]
  wire  _T_801 = &io_trigger_pkt_any_2_tdata2[30:0]; // @[lib.scala 104:36]
  wire  _T_802 = _T_801 & _T_585; // @[lib.scala 104:41]
  wire  _T_805 = io_trigger_pkt_any_2_tdata2[31] == lsu_match_data_2[31]; // @[lib.scala 104:78]
  wire  _T_806 = _T_802 | _T_805; // @[lib.scala 104:23]
  wire [7:0] _T_813 = {_T_638,_T_631,_T_624,_T_617,_T_610,_T_603,_T_596,_T_589}; // @[lib.scala 105:14]
  wire [15:0] _T_821 = {_T_694,_T_687,_T_680,_T_673,_T_666,_T_659,_T_652,_T_645,_T_813}; // @[lib.scala 105:14]
  wire [7:0] _T_828 = {_T_750,_T_743,_T_736,_T_729,_T_722,_T_715,_T_708,_T_701}; // @[lib.scala 105:14]
  wire [31:0] _T_837 = {_T_806,_T_799,_T_792,_T_785,_T_778,_T_771,_T_764,_T_757,_T_828,_T_821}; // @[lib.scala 105:14]
  wire  _T_838 = &_T_837; // @[lib.scala 105:25]
  wire  _T_839 = _T_580 & _T_838; // @[lsu_trigger.scala 19:92]
  wire  _T_842 = io_trigger_pkt_any_3_store & io_lsu_pkt_m_bits_store; // @[lsu_trigger.scala 18:126]
  wire  _T_843 = io_trigger_pkt_any_3_load & io_lsu_pkt_m_bits_load; // @[lsu_trigger.scala 19:33]
  wire  _T_845 = _T_843 & _T_33; // @[lsu_trigger.scala 19:58]
  wire  _T_846 = _T_842 | _T_845; // @[lsu_trigger.scala 18:152]
  wire  _T_847 = _T_40 & _T_846; // @[lsu_trigger.scala 18:94]
  wire  _T_850 = &io_trigger_pkt_any_3_tdata2; // @[lib.scala 101:45]
  wire  _T_851 = ~_T_850; // @[lib.scala 101:39]
  wire  _T_852 = io_trigger_pkt_any_3_match_pkt & _T_851; // @[lib.scala 101:37]
  wire  _T_855 = io_trigger_pkt_any_3_tdata2[0] == lsu_match_data_3[0]; // @[lib.scala 102:52]
  wire  _T_856 = _T_852 | _T_855; // @[lib.scala 102:41]
  wire  _T_858 = &io_trigger_pkt_any_3_tdata2[0]; // @[lib.scala 104:36]
  wire  _T_859 = _T_858 & _T_852; // @[lib.scala 104:41]
  wire  _T_862 = io_trigger_pkt_any_3_tdata2[1] == lsu_match_data_3[1]; // @[lib.scala 104:78]
  wire  _T_863 = _T_859 | _T_862; // @[lib.scala 104:23]
  wire  _T_865 = &io_trigger_pkt_any_3_tdata2[1:0]; // @[lib.scala 104:36]
  wire  _T_866 = _T_865 & _T_852; // @[lib.scala 104:41]
  wire  _T_869 = io_trigger_pkt_any_3_tdata2[2] == lsu_match_data_3[2]; // @[lib.scala 104:78]
  wire  _T_870 = _T_866 | _T_869; // @[lib.scala 104:23]
  wire  _T_872 = &io_trigger_pkt_any_3_tdata2[2:0]; // @[lib.scala 104:36]
  wire  _T_873 = _T_872 & _T_852; // @[lib.scala 104:41]
  wire  _T_876 = io_trigger_pkt_any_3_tdata2[3] == lsu_match_data_3[3]; // @[lib.scala 104:78]
  wire  _T_877 = _T_873 | _T_876; // @[lib.scala 104:23]
  wire  _T_879 = &io_trigger_pkt_any_3_tdata2[3:0]; // @[lib.scala 104:36]
  wire  _T_880 = _T_879 & _T_852; // @[lib.scala 104:41]
  wire  _T_883 = io_trigger_pkt_any_3_tdata2[4] == lsu_match_data_3[4]; // @[lib.scala 104:78]
  wire  _T_884 = _T_880 | _T_883; // @[lib.scala 104:23]
  wire  _T_886 = &io_trigger_pkt_any_3_tdata2[4:0]; // @[lib.scala 104:36]
  wire  _T_887 = _T_886 & _T_852; // @[lib.scala 104:41]
  wire  _T_890 = io_trigger_pkt_any_3_tdata2[5] == lsu_match_data_3[5]; // @[lib.scala 104:78]
  wire  _T_891 = _T_887 | _T_890; // @[lib.scala 104:23]
  wire  _T_893 = &io_trigger_pkt_any_3_tdata2[5:0]; // @[lib.scala 104:36]
  wire  _T_894 = _T_893 & _T_852; // @[lib.scala 104:41]
  wire  _T_897 = io_trigger_pkt_any_3_tdata2[6] == lsu_match_data_3[6]; // @[lib.scala 104:78]
  wire  _T_898 = _T_894 | _T_897; // @[lib.scala 104:23]
  wire  _T_900 = &io_trigger_pkt_any_3_tdata2[6:0]; // @[lib.scala 104:36]
  wire  _T_901 = _T_900 & _T_852; // @[lib.scala 104:41]
  wire  _T_904 = io_trigger_pkt_any_3_tdata2[7] == lsu_match_data_3[7]; // @[lib.scala 104:78]
  wire  _T_905 = _T_901 | _T_904; // @[lib.scala 104:23]
  wire  _T_907 = &io_trigger_pkt_any_3_tdata2[7:0]; // @[lib.scala 104:36]
  wire  _T_908 = _T_907 & _T_852; // @[lib.scala 104:41]
  wire  _T_911 = io_trigger_pkt_any_3_tdata2[8] == lsu_match_data_3[8]; // @[lib.scala 104:78]
  wire  _T_912 = _T_908 | _T_911; // @[lib.scala 104:23]
  wire  _T_914 = &io_trigger_pkt_any_3_tdata2[8:0]; // @[lib.scala 104:36]
  wire  _T_915 = _T_914 & _T_852; // @[lib.scala 104:41]
  wire  _T_918 = io_trigger_pkt_any_3_tdata2[9] == lsu_match_data_3[9]; // @[lib.scala 104:78]
  wire  _T_919 = _T_915 | _T_918; // @[lib.scala 104:23]
  wire  _T_921 = &io_trigger_pkt_any_3_tdata2[9:0]; // @[lib.scala 104:36]
  wire  _T_922 = _T_921 & _T_852; // @[lib.scala 104:41]
  wire  _T_925 = io_trigger_pkt_any_3_tdata2[10] == lsu_match_data_3[10]; // @[lib.scala 104:78]
  wire  _T_926 = _T_922 | _T_925; // @[lib.scala 104:23]
  wire  _T_928 = &io_trigger_pkt_any_3_tdata2[10:0]; // @[lib.scala 104:36]
  wire  _T_929 = _T_928 & _T_852; // @[lib.scala 104:41]
  wire  _T_932 = io_trigger_pkt_any_3_tdata2[11] == lsu_match_data_3[11]; // @[lib.scala 104:78]
  wire  _T_933 = _T_929 | _T_932; // @[lib.scala 104:23]
  wire  _T_935 = &io_trigger_pkt_any_3_tdata2[11:0]; // @[lib.scala 104:36]
  wire  _T_936 = _T_935 & _T_852; // @[lib.scala 104:41]
  wire  _T_939 = io_trigger_pkt_any_3_tdata2[12] == lsu_match_data_3[12]; // @[lib.scala 104:78]
  wire  _T_940 = _T_936 | _T_939; // @[lib.scala 104:23]
  wire  _T_942 = &io_trigger_pkt_any_3_tdata2[12:0]; // @[lib.scala 104:36]
  wire  _T_943 = _T_942 & _T_852; // @[lib.scala 104:41]
  wire  _T_946 = io_trigger_pkt_any_3_tdata2[13] == lsu_match_data_3[13]; // @[lib.scala 104:78]
  wire  _T_947 = _T_943 | _T_946; // @[lib.scala 104:23]
  wire  _T_949 = &io_trigger_pkt_any_3_tdata2[13:0]; // @[lib.scala 104:36]
  wire  _T_950 = _T_949 & _T_852; // @[lib.scala 104:41]
  wire  _T_953 = io_trigger_pkt_any_3_tdata2[14] == lsu_match_data_3[14]; // @[lib.scala 104:78]
  wire  _T_954 = _T_950 | _T_953; // @[lib.scala 104:23]
  wire  _T_956 = &io_trigger_pkt_any_3_tdata2[14:0]; // @[lib.scala 104:36]
  wire  _T_957 = _T_956 & _T_852; // @[lib.scala 104:41]
  wire  _T_960 = io_trigger_pkt_any_3_tdata2[15] == lsu_match_data_3[15]; // @[lib.scala 104:78]
  wire  _T_961 = _T_957 | _T_960; // @[lib.scala 104:23]
  wire  _T_963 = &io_trigger_pkt_any_3_tdata2[15:0]; // @[lib.scala 104:36]
  wire  _T_964 = _T_963 & _T_852; // @[lib.scala 104:41]
  wire  _T_967 = io_trigger_pkt_any_3_tdata2[16] == lsu_match_data_3[16]; // @[lib.scala 104:78]
  wire  _T_968 = _T_964 | _T_967; // @[lib.scala 104:23]
  wire  _T_970 = &io_trigger_pkt_any_3_tdata2[16:0]; // @[lib.scala 104:36]
  wire  _T_971 = _T_970 & _T_852; // @[lib.scala 104:41]
  wire  _T_974 = io_trigger_pkt_any_3_tdata2[17] == lsu_match_data_3[17]; // @[lib.scala 104:78]
  wire  _T_975 = _T_971 | _T_974; // @[lib.scala 104:23]
  wire  _T_977 = &io_trigger_pkt_any_3_tdata2[17:0]; // @[lib.scala 104:36]
  wire  _T_978 = _T_977 & _T_852; // @[lib.scala 104:41]
  wire  _T_981 = io_trigger_pkt_any_3_tdata2[18] == lsu_match_data_3[18]; // @[lib.scala 104:78]
  wire  _T_982 = _T_978 | _T_981; // @[lib.scala 104:23]
  wire  _T_984 = &io_trigger_pkt_any_3_tdata2[18:0]; // @[lib.scala 104:36]
  wire  _T_985 = _T_984 & _T_852; // @[lib.scala 104:41]
  wire  _T_988 = io_trigger_pkt_any_3_tdata2[19] == lsu_match_data_3[19]; // @[lib.scala 104:78]
  wire  _T_989 = _T_985 | _T_988; // @[lib.scala 104:23]
  wire  _T_991 = &io_trigger_pkt_any_3_tdata2[19:0]; // @[lib.scala 104:36]
  wire  _T_992 = _T_991 & _T_852; // @[lib.scala 104:41]
  wire  _T_995 = io_trigger_pkt_any_3_tdata2[20] == lsu_match_data_3[20]; // @[lib.scala 104:78]
  wire  _T_996 = _T_992 | _T_995; // @[lib.scala 104:23]
  wire  _T_998 = &io_trigger_pkt_any_3_tdata2[20:0]; // @[lib.scala 104:36]
  wire  _T_999 = _T_998 & _T_852; // @[lib.scala 104:41]
  wire  _T_1002 = io_trigger_pkt_any_3_tdata2[21] == lsu_match_data_3[21]; // @[lib.scala 104:78]
  wire  _T_1003 = _T_999 | _T_1002; // @[lib.scala 104:23]
  wire  _T_1005 = &io_trigger_pkt_any_3_tdata2[21:0]; // @[lib.scala 104:36]
  wire  _T_1006 = _T_1005 & _T_852; // @[lib.scala 104:41]
  wire  _T_1009 = io_trigger_pkt_any_3_tdata2[22] == lsu_match_data_3[22]; // @[lib.scala 104:78]
  wire  _T_1010 = _T_1006 | _T_1009; // @[lib.scala 104:23]
  wire  _T_1012 = &io_trigger_pkt_any_3_tdata2[22:0]; // @[lib.scala 104:36]
  wire  _T_1013 = _T_1012 & _T_852; // @[lib.scala 104:41]
  wire  _T_1016 = io_trigger_pkt_any_3_tdata2[23] == lsu_match_data_3[23]; // @[lib.scala 104:78]
  wire  _T_1017 = _T_1013 | _T_1016; // @[lib.scala 104:23]
  wire  _T_1019 = &io_trigger_pkt_any_3_tdata2[23:0]; // @[lib.scala 104:36]
  wire  _T_1020 = _T_1019 & _T_852; // @[lib.scala 104:41]
  wire  _T_1023 = io_trigger_pkt_any_3_tdata2[24] == lsu_match_data_3[24]; // @[lib.scala 104:78]
  wire  _T_1024 = _T_1020 | _T_1023; // @[lib.scala 104:23]
  wire  _T_1026 = &io_trigger_pkt_any_3_tdata2[24:0]; // @[lib.scala 104:36]
  wire  _T_1027 = _T_1026 & _T_852; // @[lib.scala 104:41]
  wire  _T_1030 = io_trigger_pkt_any_3_tdata2[25] == lsu_match_data_3[25]; // @[lib.scala 104:78]
  wire  _T_1031 = _T_1027 | _T_1030; // @[lib.scala 104:23]
  wire  _T_1033 = &io_trigger_pkt_any_3_tdata2[25:0]; // @[lib.scala 104:36]
  wire  _T_1034 = _T_1033 & _T_852; // @[lib.scala 104:41]
  wire  _T_1037 = io_trigger_pkt_any_3_tdata2[26] == lsu_match_data_3[26]; // @[lib.scala 104:78]
  wire  _T_1038 = _T_1034 | _T_1037; // @[lib.scala 104:23]
  wire  _T_1040 = &io_trigger_pkt_any_3_tdata2[26:0]; // @[lib.scala 104:36]
  wire  _T_1041 = _T_1040 & _T_852; // @[lib.scala 104:41]
  wire  _T_1044 = io_trigger_pkt_any_3_tdata2[27] == lsu_match_data_3[27]; // @[lib.scala 104:78]
  wire  _T_1045 = _T_1041 | _T_1044; // @[lib.scala 104:23]
  wire  _T_1047 = &io_trigger_pkt_any_3_tdata2[27:0]; // @[lib.scala 104:36]
  wire  _T_1048 = _T_1047 & _T_852; // @[lib.scala 104:41]
  wire  _T_1051 = io_trigger_pkt_any_3_tdata2[28] == lsu_match_data_3[28]; // @[lib.scala 104:78]
  wire  _T_1052 = _T_1048 | _T_1051; // @[lib.scala 104:23]
  wire  _T_1054 = &io_trigger_pkt_any_3_tdata2[28:0]; // @[lib.scala 104:36]
  wire  _T_1055 = _T_1054 & _T_852; // @[lib.scala 104:41]
  wire  _T_1058 = io_trigger_pkt_any_3_tdata2[29] == lsu_match_data_3[29]; // @[lib.scala 104:78]
  wire  _T_1059 = _T_1055 | _T_1058; // @[lib.scala 104:23]
  wire  _T_1061 = &io_trigger_pkt_any_3_tdata2[29:0]; // @[lib.scala 104:36]
  wire  _T_1062 = _T_1061 & _T_852; // @[lib.scala 104:41]
  wire  _T_1065 = io_trigger_pkt_any_3_tdata2[30] == lsu_match_data_3[30]; // @[lib.scala 104:78]
  wire  _T_1066 = _T_1062 | _T_1065; // @[lib.scala 104:23]
  wire  _T_1068 = &io_trigger_pkt_any_3_tdata2[30:0]; // @[lib.scala 104:36]
  wire  _T_1069 = _T_1068 & _T_852; // @[lib.scala 104:41]
  wire  _T_1072 = io_trigger_pkt_any_3_tdata2[31] == lsu_match_data_3[31]; // @[lib.scala 104:78]
  wire  _T_1073 = _T_1069 | _T_1072; // @[lib.scala 104:23]
  wire [7:0] _T_1080 = {_T_905,_T_898,_T_891,_T_884,_T_877,_T_870,_T_863,_T_856}; // @[lib.scala 105:14]
  wire [15:0] _T_1088 = {_T_961,_T_954,_T_947,_T_940,_T_933,_T_926,_T_919,_T_912,_T_1080}; // @[lib.scala 105:14]
  wire [7:0] _T_1095 = {_T_1017,_T_1010,_T_1003,_T_996,_T_989,_T_982,_T_975,_T_968}; // @[lib.scala 105:14]
  wire [31:0] _T_1104 = {_T_1073,_T_1066,_T_1059,_T_1052,_T_1045,_T_1038,_T_1031,_T_1024,_T_1095,_T_1088}; // @[lib.scala 105:14]
  wire  _T_1105 = &_T_1104; // @[lib.scala 105:25]
  wire  _T_1106 = _T_847 & _T_1105; // @[lsu_trigger.scala 19:92]
  wire [2:0] _T_1108 = {_T_1106,_T_839,_T_572}; // @[Cat.scala 29:58]
  assign io_lsu_trigger_match_m = {_T_1108,_T_305}; // @[lsu_trigger.scala 18:26]
endmodule
module lsu_clkdomain(
  input   clock,
  input   reset,
  input   io_free_clk,
  input   io_clk_override,
  input   io_dma_dccm_req,
  input   io_ldst_stbuf_reqvld_r,
  input   io_stbuf_reqvld_any,
  input   io_stbuf_reqvld_flushed_any,
  input   io_lsu_busreq_r,
  input   io_lsu_bus_buffer_pend_any,
  input   io_lsu_bus_buffer_empty_any,
  input   io_lsu_stbuf_empty_any,
  input   io_lsu_bus_clk_en,
  input   io_lsu_p_valid,
  input   io_lsu_pkt_d_valid,
  input   io_lsu_pkt_d_bits_store,
  input   io_lsu_pkt_m_valid,
  input   io_lsu_pkt_m_bits_store,
  input   io_lsu_pkt_r_valid,
  output  io_lsu_c1_m_clk,
  output  io_lsu_c1_r_clk,
  output  io_lsu_c2_m_clk,
  output  io_lsu_c2_r_clk,
  output  io_lsu_store_c1_m_clk,
  output  io_lsu_store_c1_r_clk,
  output  io_lsu_stbuf_c1_clk,
  output  io_lsu_bus_obuf_c1_clk,
  output  io_lsu_bus_ibuf_c1_clk,
  output  io_lsu_bus_buf_c1_clk,
  output  io_lsu_busm_clk,
  output  io_lsu_free_c2_clk,
  input   io_scan_mode
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire  rvclkhdr_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_1_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_1_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_1_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_1_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_2_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_2_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_2_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_2_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_3_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_3_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_3_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_3_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_4_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_4_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_4_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_4_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_5_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_5_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_5_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_5_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_6_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_6_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_6_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_6_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_7_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_7_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_7_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_7_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_8_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_8_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_8_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_8_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_9_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_9_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_9_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_9_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_10_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_10_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_10_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_10_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_11_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_11_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_11_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_11_io_scan_mode; // @[lib.scala 343:22]
  wire  _T = io_lsu_p_valid | io_dma_dccm_req; // @[lsu_clkdomain.scala 62:51]
  reg  lsu_c1_d_clken_q; // @[lsu_clkdomain.scala 81:67]
  wire  _T_1 = io_lsu_pkt_d_valid | lsu_c1_d_clken_q; // @[lsu_clkdomain.scala 63:51]
  wire  lsu_c1_m_clken = _T_1 | io_clk_override; // @[lsu_clkdomain.scala 63:70]
  reg  lsu_c1_m_clken_q; // @[lsu_clkdomain.scala 82:67]
  wire  _T_2 = io_lsu_pkt_m_valid | lsu_c1_m_clken_q; // @[lsu_clkdomain.scala 64:51]
  wire  lsu_c1_r_clken = _T_2 | io_clk_override; // @[lsu_clkdomain.scala 64:70]
  wire  _T_3 = lsu_c1_m_clken | lsu_c1_m_clken_q; // @[lsu_clkdomain.scala 66:47]
  reg  lsu_c1_r_clken_q; // @[lsu_clkdomain.scala 83:67]
  wire  _T_4 = lsu_c1_r_clken | lsu_c1_r_clken_q; // @[lsu_clkdomain.scala 67:47]
  wire  _T_5 = lsu_c1_m_clken & io_lsu_pkt_d_bits_store; // @[lsu_clkdomain.scala 69:49]
  wire  _T_6 = lsu_c1_r_clken & io_lsu_pkt_m_bits_store; // @[lsu_clkdomain.scala 70:49]
  wire  _T_7 = io_ldst_stbuf_reqvld_r | io_stbuf_reqvld_any; // @[lsu_clkdomain.scala 71:55]
  wire  _T_8 = _T_7 | io_stbuf_reqvld_flushed_any; // @[lsu_clkdomain.scala 71:77]
  wire  _T_9 = io_lsu_bus_buffer_pend_any | io_lsu_busreq_r; // @[lsu_clkdomain.scala 73:61]
  wire  _T_10 = _T_9 | io_clk_override; // @[lsu_clkdomain.scala 73:79]
  wire  _T_11 = ~io_lsu_bus_buffer_empty_any; // @[lsu_clkdomain.scala 74:32]
  wire  _T_12 = _T_11 | io_lsu_busreq_r; // @[lsu_clkdomain.scala 74:61]
  wire  _T_13 = io_lsu_p_valid | io_lsu_pkt_d_valid; // @[lsu_clkdomain.scala 76:48]
  wire  _T_14 = _T_13 | io_lsu_pkt_m_valid; // @[lsu_clkdomain.scala 76:69]
  wire  _T_15 = _T_14 | io_lsu_pkt_r_valid; // @[lsu_clkdomain.scala 76:90]
  wire  _T_17 = _T_15 | _T_11; // @[lsu_clkdomain.scala 76:112]
  wire  _T_18 = ~io_lsu_stbuf_empty_any; // @[lsu_clkdomain.scala 76:145]
  wire  _T_19 = _T_17 | _T_18; // @[lsu_clkdomain.scala 76:143]
  wire  lsu_free_c1_clken = _T_19 | io_clk_override; // @[lsu_clkdomain.scala 76:169]
  reg  lsu_free_c1_clken_q; // @[lsu_clkdomain.scala 80:60]
  wire  _T_20 = lsu_free_c1_clken | lsu_free_c1_clken_q; // @[lsu_clkdomain.scala 77:50]
  rvclkhdr rvclkhdr ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_io_l1clk),
    .io_clk(rvclkhdr_io_clk),
    .io_en(rvclkhdr_io_en),
    .io_scan_mode(rvclkhdr_io_scan_mode)
  );
  rvclkhdr rvclkhdr_1 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_1_io_l1clk),
    .io_clk(rvclkhdr_1_io_clk),
    .io_en(rvclkhdr_1_io_en),
    .io_scan_mode(rvclkhdr_1_io_scan_mode)
  );
  rvclkhdr rvclkhdr_2 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_2_io_l1clk),
    .io_clk(rvclkhdr_2_io_clk),
    .io_en(rvclkhdr_2_io_en),
    .io_scan_mode(rvclkhdr_2_io_scan_mode)
  );
  rvclkhdr rvclkhdr_3 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_3_io_l1clk),
    .io_clk(rvclkhdr_3_io_clk),
    .io_en(rvclkhdr_3_io_en),
    .io_scan_mode(rvclkhdr_3_io_scan_mode)
  );
  rvclkhdr rvclkhdr_4 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_4_io_l1clk),
    .io_clk(rvclkhdr_4_io_clk),
    .io_en(rvclkhdr_4_io_en),
    .io_scan_mode(rvclkhdr_4_io_scan_mode)
  );
  rvclkhdr rvclkhdr_5 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_5_io_l1clk),
    .io_clk(rvclkhdr_5_io_clk),
    .io_en(rvclkhdr_5_io_en),
    .io_scan_mode(rvclkhdr_5_io_scan_mode)
  );
  rvclkhdr rvclkhdr_6 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_6_io_l1clk),
    .io_clk(rvclkhdr_6_io_clk),
    .io_en(rvclkhdr_6_io_en),
    .io_scan_mode(rvclkhdr_6_io_scan_mode)
  );
  rvclkhdr rvclkhdr_7 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_7_io_l1clk),
    .io_clk(rvclkhdr_7_io_clk),
    .io_en(rvclkhdr_7_io_en),
    .io_scan_mode(rvclkhdr_7_io_scan_mode)
  );
  rvclkhdr rvclkhdr_8 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_8_io_l1clk),
    .io_clk(rvclkhdr_8_io_clk),
    .io_en(rvclkhdr_8_io_en),
    .io_scan_mode(rvclkhdr_8_io_scan_mode)
  );
  rvclkhdr rvclkhdr_9 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_9_io_l1clk),
    .io_clk(rvclkhdr_9_io_clk),
    .io_en(rvclkhdr_9_io_en),
    .io_scan_mode(rvclkhdr_9_io_scan_mode)
  );
  rvclkhdr rvclkhdr_10 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_10_io_l1clk),
    .io_clk(rvclkhdr_10_io_clk),
    .io_en(rvclkhdr_10_io_en),
    .io_scan_mode(rvclkhdr_10_io_scan_mode)
  );
  rvclkhdr rvclkhdr_11 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_11_io_l1clk),
    .io_clk(rvclkhdr_11_io_clk),
    .io_en(rvclkhdr_11_io_en),
    .io_scan_mode(rvclkhdr_11_io_scan_mode)
  );
  assign io_lsu_c1_m_clk = rvclkhdr_io_l1clk; // @[lsu_clkdomain.scala 85:26]
  assign io_lsu_c1_r_clk = rvclkhdr_1_io_l1clk; // @[lsu_clkdomain.scala 86:26]
  assign io_lsu_c2_m_clk = rvclkhdr_2_io_l1clk; // @[lsu_clkdomain.scala 87:26]
  assign io_lsu_c2_r_clk = rvclkhdr_3_io_l1clk; // @[lsu_clkdomain.scala 88:26]
  assign io_lsu_store_c1_m_clk = rvclkhdr_4_io_l1clk; // @[lsu_clkdomain.scala 89:26]
  assign io_lsu_store_c1_r_clk = rvclkhdr_5_io_l1clk; // @[lsu_clkdomain.scala 90:26]
  assign io_lsu_stbuf_c1_clk = rvclkhdr_6_io_l1clk; // @[lsu_clkdomain.scala 91:26]
  assign io_lsu_bus_obuf_c1_clk = rvclkhdr_8_io_l1clk; // @[lsu_clkdomain.scala 93:26]
  assign io_lsu_bus_ibuf_c1_clk = rvclkhdr_7_io_l1clk; // @[lsu_clkdomain.scala 92:26]
  assign io_lsu_bus_buf_c1_clk = rvclkhdr_9_io_l1clk; // @[lsu_clkdomain.scala 94:26]
  assign io_lsu_busm_clk = rvclkhdr_10_io_l1clk; // @[lsu_clkdomain.scala 95:26]
  assign io_lsu_free_c2_clk = rvclkhdr_11_io_l1clk; // @[lsu_clkdomain.scala 96:26]
  assign rvclkhdr_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_io_en = _T_1 | io_clk_override; // @[lib.scala 345:16]
  assign rvclkhdr_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_1_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_1_io_en = _T_2 | io_clk_override; // @[lib.scala 345:16]
  assign rvclkhdr_1_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_2_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_2_io_en = _T_3 | io_clk_override; // @[lib.scala 345:16]
  assign rvclkhdr_2_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_3_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_3_io_en = _T_4 | io_clk_override; // @[lib.scala 345:16]
  assign rvclkhdr_3_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_4_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_4_io_en = _T_5 | io_clk_override; // @[lib.scala 345:16]
  assign rvclkhdr_4_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_5_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_5_io_en = _T_6 | io_clk_override; // @[lib.scala 345:16]
  assign rvclkhdr_5_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_6_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_6_io_en = _T_8 | io_clk_override; // @[lib.scala 345:16]
  assign rvclkhdr_6_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_7_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_7_io_en = io_lsu_busreq_r | io_clk_override; // @[lib.scala 345:16]
  assign rvclkhdr_7_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_8_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_8_io_en = _T_10 & io_lsu_bus_clk_en; // @[lib.scala 345:16]
  assign rvclkhdr_8_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_9_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_9_io_en = _T_12 | io_clk_override; // @[lib.scala 345:16]
  assign rvclkhdr_9_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_10_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_10_io_en = io_lsu_bus_clk_en; // @[lib.scala 345:16]
  assign rvclkhdr_10_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_11_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_11_io_en = _T_20 | io_clk_override; // @[lib.scala 345:16]
  assign rvclkhdr_11_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  lsu_c1_d_clken_q = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  lsu_c1_m_clken_q = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  lsu_c1_r_clken_q = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  lsu_free_c1_clken_q = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    lsu_c1_d_clken_q = 1'h0;
  end
  if (reset) begin
    lsu_c1_m_clken_q = 1'h0;
  end
  if (reset) begin
    lsu_c1_r_clken_q = 1'h0;
  end
  if (reset) begin
    lsu_free_c1_clken_q = 1'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge io_lsu_free_c2_clk or posedge reset) begin
    if (reset) begin
      lsu_c1_d_clken_q <= 1'h0;
    end else begin
      lsu_c1_d_clken_q <= _T | io_clk_override;
    end
  end
  always @(posedge io_lsu_free_c2_clk or posedge reset) begin
    if (reset) begin
      lsu_c1_m_clken_q <= 1'h0;
    end else begin
      lsu_c1_m_clken_q <= _T_1 | io_clk_override;
    end
  end
  always @(posedge io_lsu_free_c2_clk or posedge reset) begin
    if (reset) begin
      lsu_c1_r_clken_q <= 1'h0;
    end else begin
      lsu_c1_r_clken_q <= _T_2 | io_clk_override;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      lsu_free_c1_clken_q <= 1'h0;
    end else begin
      lsu_free_c1_clken_q <= _T_19 | io_clk_override;
    end
  end
endmodule
module lsu_bus_buffer(
  input         clock,
  input         reset,
  input         io_scan_mode,
  output        io_tlu_busbuff_lsu_pmu_bus_misaligned,
  output        io_tlu_busbuff_lsu_pmu_bus_error,
  output        io_tlu_busbuff_lsu_pmu_bus_busy,
  input         io_tlu_busbuff_dec_tlu_external_ldfwd_disable,
  input         io_tlu_busbuff_dec_tlu_wb_coalescing_disable,
  input         io_tlu_busbuff_dec_tlu_sideeffect_posted_disable,
  output        io_tlu_busbuff_lsu_imprecise_error_load_any,
  output        io_tlu_busbuff_lsu_imprecise_error_store_any,
  output [31:0] io_tlu_busbuff_lsu_imprecise_error_addr_any,
  output        io_dctl_busbuff_lsu_nonblock_load_valid_m,
  output [1:0]  io_dctl_busbuff_lsu_nonblock_load_tag_m,
  output        io_dctl_busbuff_lsu_nonblock_load_inv_r,
  output [1:0]  io_dctl_busbuff_lsu_nonblock_load_inv_tag_r,
  output        io_dctl_busbuff_lsu_nonblock_load_data_valid,
  output        io_dctl_busbuff_lsu_nonblock_load_data_error,
  output [1:0]  io_dctl_busbuff_lsu_nonblock_load_data_tag,
  output [31:0] io_dctl_busbuff_lsu_nonblock_load_data,
  input         io_dec_tlu_force_halt,
  input         io_lsu_c2_r_clk,
  input         io_lsu_bus_ibuf_c1_clk,
  input         io_lsu_bus_obuf_c1_clk,
  input         io_lsu_bus_buf_c1_clk,
  input         io_lsu_free_c2_clk,
  input         io_lsu_busm_clk,
  input         io_dec_lsu_valid_raw_d,
  input         io_lsu_pkt_m_valid,
  input         io_lsu_pkt_m_bits_load,
  input         io_lsu_pkt_r_bits_by,
  input         io_lsu_pkt_r_bits_half,
  input         io_lsu_pkt_r_bits_word,
  input         io_lsu_pkt_r_bits_load,
  input         io_lsu_pkt_r_bits_store,
  input         io_lsu_pkt_r_bits_unsign,
  input  [31:0] io_lsu_addr_m,
  input  [31:0] io_end_addr_m,
  input  [31:0] io_lsu_addr_r,
  input  [31:0] io_end_addr_r,
  input  [31:0] io_store_data_r,
  input         io_no_word_merge_r,
  input         io_no_dword_merge_r,
  input         io_lsu_busreq_m,
  input         io_ld_full_hit_m,
  input         io_flush_m_up,
  input         io_flush_r,
  input         io_lsu_commit_r,
  input         io_is_sideeffects_r,
  input         io_ldst_dual_d,
  input         io_ldst_dual_m,
  input         io_ldst_dual_r,
  input  [7:0]  io_ldst_byteen_ext_m,
  output        io_lsu_axi_aw_valid,
  output [31:0] io_lsu_axi_aw_bits_addr,
  output [2:0]  io_lsu_axi_aw_bits_size,
  output        io_lsu_axi_w_valid,
  output [7:0]  io_lsu_axi_w_bits_strb,
  output        io_lsu_axi_ar_valid,
  output [31:0] io_lsu_axi_ar_bits_addr,
  output [2:0]  io_lsu_axi_ar_bits_size,
  input         io_lsu_bus_clk_en,
  input         io_lsu_bus_clk_en_q,
  output        io_lsu_busreq_r,
  output        io_lsu_bus_buffer_pend_any,
  output        io_lsu_bus_buffer_full_any,
  output        io_lsu_bus_buffer_empty_any,
  output [3:0]  io_ld_byte_hit_buf_lo,
  output [3:0]  io_ld_byte_hit_buf_hi,
  output [31:0] io_ld_fwddata_buf_lo,
  output [31:0] io_ld_fwddata_buf_hi
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
`endif // RANDOMIZE_REG_INIT
  wire  rvclkhdr_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_1_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_1_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_1_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_1_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_2_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_2_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_2_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_2_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_3_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_3_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_3_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_3_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_4_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_4_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_4_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_4_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_5_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_5_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_5_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_5_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_6_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_6_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_6_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_6_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_7_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_7_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_7_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_7_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_8_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_8_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_8_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_8_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_9_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_9_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_9_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_9_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_10_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_10_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_10_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_10_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_11_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_11_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_11_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_11_io_scan_mode; // @[lib.scala 368:23]
  wire [3:0] ldst_byteen_hi_m = io_ldst_byteen_ext_m[7:4]; // @[lsu_bus_buffer.scala 72:46]
  wire [3:0] ldst_byteen_lo_m = io_ldst_byteen_ext_m[3:0]; // @[lsu_bus_buffer.scala 73:46]
  reg [31:0] buf_addr_0; // @[lib.scala 374:16]
  wire  _T_2 = io_lsu_addr_m[31:2] == buf_addr_0[31:2]; // @[lsu_bus_buffer.scala 75:74]
  reg  _T_4360; // @[Reg.scala 27:20]
  reg  _T_4357; // @[Reg.scala 27:20]
  reg  _T_4354; // @[Reg.scala 27:20]
  reg  _T_4351; // @[Reg.scala 27:20]
  wire [3:0] buf_write = {_T_4360,_T_4357,_T_4354,_T_4351}; // @[Cat.scala 29:58]
  wire  _T_4 = _T_2 & buf_write[0]; // @[lsu_bus_buffer.scala 75:98]
  reg [2:0] buf_state_0; // @[Reg.scala 27:20]
  wire  _T_5 = buf_state_0 != 3'h0; // @[lsu_bus_buffer.scala 75:129]
  wire  _T_6 = _T_4 & _T_5; // @[lsu_bus_buffer.scala 75:113]
  wire  ld_addr_hitvec_lo_0 = _T_6 & io_lsu_busreq_m; // @[lsu_bus_buffer.scala 75:141]
  reg [31:0] buf_addr_1; // @[lib.scala 374:16]
  wire  _T_9 = io_lsu_addr_m[31:2] == buf_addr_1[31:2]; // @[lsu_bus_buffer.scala 75:74]
  wire  _T_11 = _T_9 & buf_write[1]; // @[lsu_bus_buffer.scala 75:98]
  reg [2:0] buf_state_1; // @[Reg.scala 27:20]
  wire  _T_12 = buf_state_1 != 3'h0; // @[lsu_bus_buffer.scala 75:129]
  wire  _T_13 = _T_11 & _T_12; // @[lsu_bus_buffer.scala 75:113]
  wire  ld_addr_hitvec_lo_1 = _T_13 & io_lsu_busreq_m; // @[lsu_bus_buffer.scala 75:141]
  reg [31:0] buf_addr_2; // @[lib.scala 374:16]
  wire  _T_16 = io_lsu_addr_m[31:2] == buf_addr_2[31:2]; // @[lsu_bus_buffer.scala 75:74]
  wire  _T_18 = _T_16 & buf_write[2]; // @[lsu_bus_buffer.scala 75:98]
  reg [2:0] buf_state_2; // @[Reg.scala 27:20]
  wire  _T_19 = buf_state_2 != 3'h0; // @[lsu_bus_buffer.scala 75:129]
  wire  _T_20 = _T_18 & _T_19; // @[lsu_bus_buffer.scala 75:113]
  wire  ld_addr_hitvec_lo_2 = _T_20 & io_lsu_busreq_m; // @[lsu_bus_buffer.scala 75:141]
  reg [31:0] buf_addr_3; // @[lib.scala 374:16]
  wire  _T_23 = io_lsu_addr_m[31:2] == buf_addr_3[31:2]; // @[lsu_bus_buffer.scala 75:74]
  wire  _T_25 = _T_23 & buf_write[3]; // @[lsu_bus_buffer.scala 75:98]
  reg [2:0] buf_state_3; // @[Reg.scala 27:20]
  wire  _T_26 = buf_state_3 != 3'h0; // @[lsu_bus_buffer.scala 75:129]
  wire  _T_27 = _T_25 & _T_26; // @[lsu_bus_buffer.scala 75:113]
  wire  ld_addr_hitvec_lo_3 = _T_27 & io_lsu_busreq_m; // @[lsu_bus_buffer.scala 75:141]
  wire  _T_30 = io_end_addr_m[31:2] == buf_addr_0[31:2]; // @[lsu_bus_buffer.scala 76:74]
  wire  _T_32 = _T_30 & buf_write[0]; // @[lsu_bus_buffer.scala 76:98]
  wire  _T_34 = _T_32 & _T_5; // @[lsu_bus_buffer.scala 76:113]
  wire  ld_addr_hitvec_hi_0 = _T_34 & io_lsu_busreq_m; // @[lsu_bus_buffer.scala 76:141]
  wire  _T_37 = io_end_addr_m[31:2] == buf_addr_1[31:2]; // @[lsu_bus_buffer.scala 76:74]
  wire  _T_39 = _T_37 & buf_write[1]; // @[lsu_bus_buffer.scala 76:98]
  wire  _T_41 = _T_39 & _T_12; // @[lsu_bus_buffer.scala 76:113]
  wire  ld_addr_hitvec_hi_1 = _T_41 & io_lsu_busreq_m; // @[lsu_bus_buffer.scala 76:141]
  wire  _T_44 = io_end_addr_m[31:2] == buf_addr_2[31:2]; // @[lsu_bus_buffer.scala 76:74]
  wire  _T_46 = _T_44 & buf_write[2]; // @[lsu_bus_buffer.scala 76:98]
  wire  _T_48 = _T_46 & _T_19; // @[lsu_bus_buffer.scala 76:113]
  wire  ld_addr_hitvec_hi_2 = _T_48 & io_lsu_busreq_m; // @[lsu_bus_buffer.scala 76:141]
  wire  _T_51 = io_end_addr_m[31:2] == buf_addr_3[31:2]; // @[lsu_bus_buffer.scala 76:74]
  wire  _T_53 = _T_51 & buf_write[3]; // @[lsu_bus_buffer.scala 76:98]
  wire  _T_55 = _T_53 & _T_26; // @[lsu_bus_buffer.scala 76:113]
  wire  ld_addr_hitvec_hi_3 = _T_55 & io_lsu_busreq_m; // @[lsu_bus_buffer.scala 76:141]
  reg [3:0] buf_byteen_3; // @[Reg.scala 27:20]
  wire  _T_99 = ld_addr_hitvec_lo_3 & buf_byteen_3[0]; // @[lsu_bus_buffer.scala 140:95]
  wire  _T_101 = _T_99 & ldst_byteen_lo_m[0]; // @[lsu_bus_buffer.scala 140:114]
  reg [3:0] buf_byteen_2; // @[Reg.scala 27:20]
  wire  _T_95 = ld_addr_hitvec_lo_2 & buf_byteen_2[0]; // @[lsu_bus_buffer.scala 140:95]
  wire  _T_97 = _T_95 & ldst_byteen_lo_m[0]; // @[lsu_bus_buffer.scala 140:114]
  reg [3:0] buf_byteen_1; // @[Reg.scala 27:20]
  wire  _T_91 = ld_addr_hitvec_lo_1 & buf_byteen_1[0]; // @[lsu_bus_buffer.scala 140:95]
  wire  _T_93 = _T_91 & ldst_byteen_lo_m[0]; // @[lsu_bus_buffer.scala 140:114]
  reg [3:0] buf_byteen_0; // @[Reg.scala 27:20]
  wire  _T_87 = ld_addr_hitvec_lo_0 & buf_byteen_0[0]; // @[lsu_bus_buffer.scala 140:95]
  wire  _T_89 = _T_87 & ldst_byteen_lo_m[0]; // @[lsu_bus_buffer.scala 140:114]
  wire [3:0] ld_byte_hitvec_lo_0 = {_T_101,_T_97,_T_93,_T_89}; // @[Cat.scala 29:58]
  reg [3:0] buf_ageQ_3; // @[lsu_bus_buffer.scala 499:60]
  wire  _T_2621 = buf_state_3 == 3'h2; // @[lsu_bus_buffer.scala 411:93]
  wire  _T_4107 = 3'h0 == buf_state_3; // @[Conditional.scala 37:30]
  wire  _T_4130 = 3'h1 == buf_state_3; // @[Conditional.scala 37:30]
  wire  _T_4134 = 3'h2 == buf_state_3; // @[Conditional.scala 37:30]
  reg [1:0] _T_1848; // @[Reg.scala 27:20]
  wire [2:0] obuf_tag0 = {{1'd0}, _T_1848}; // @[lsu_bus_buffer.scala 351:13]
  wire  _T_4141 = obuf_tag0 == 3'h3; // @[lsu_bus_buffer.scala 454:48]
  reg  obuf_merge; // @[Reg.scala 27:20]
  reg [1:0] obuf_tag1; // @[Reg.scala 27:20]
  wire [2:0] _GEN_358 = {{1'd0}, obuf_tag1}; // @[lsu_bus_buffer.scala 454:104]
  wire  _T_4142 = _GEN_358 == 3'h3; // @[lsu_bus_buffer.scala 454:104]
  wire  _T_4143 = obuf_merge & _T_4142; // @[lsu_bus_buffer.scala 454:91]
  wire  _T_4144 = _T_4141 | _T_4143; // @[lsu_bus_buffer.scala 454:77]
  reg  obuf_valid; // @[lsu_bus_buffer.scala 345:54]
  wire  _T_4145 = _T_4144 & obuf_valid; // @[lsu_bus_buffer.scala 454:135]
  reg  obuf_wr_enQ; // @[lsu_bus_buffer.scala 344:55]
  wire  _T_4146 = _T_4145 & obuf_wr_enQ; // @[lsu_bus_buffer.scala 454:148]
  wire  _GEN_280 = _T_4134 & _T_4146; // @[Conditional.scala 39:67]
  wire  _GEN_293 = _T_4130 ? 1'h0 : _GEN_280; // @[Conditional.scala 39:67]
  wire  buf_cmd_state_bus_en_3 = _T_4107 ? 1'h0 : _GEN_293; // @[Conditional.scala 40:58]
  wire  _T_2622 = _T_2621 & buf_cmd_state_bus_en_3; // @[lsu_bus_buffer.scala 411:103]
  wire  _T_2623 = ~_T_2622; // @[lsu_bus_buffer.scala 411:78]
  wire  _T_2624 = buf_ageQ_3[3] & _T_2623; // @[lsu_bus_buffer.scala 411:76]
  wire  _T_2616 = buf_state_2 == 3'h2; // @[lsu_bus_buffer.scala 411:93]
  wire  _T_3914 = 3'h0 == buf_state_2; // @[Conditional.scala 37:30]
  wire  _T_3937 = 3'h1 == buf_state_2; // @[Conditional.scala 37:30]
  wire  _T_3941 = 3'h2 == buf_state_2; // @[Conditional.scala 37:30]
  wire  _T_3948 = obuf_tag0 == 3'h2; // @[lsu_bus_buffer.scala 454:48]
  wire  _T_3949 = _GEN_358 == 3'h2; // @[lsu_bus_buffer.scala 454:104]
  wire  _T_3950 = obuf_merge & _T_3949; // @[lsu_bus_buffer.scala 454:91]
  wire  _T_3951 = _T_3948 | _T_3950; // @[lsu_bus_buffer.scala 454:77]
  wire  _T_3952 = _T_3951 & obuf_valid; // @[lsu_bus_buffer.scala 454:135]
  wire  _T_3953 = _T_3952 & obuf_wr_enQ; // @[lsu_bus_buffer.scala 454:148]
  wire  _GEN_204 = _T_3941 & _T_3953; // @[Conditional.scala 39:67]
  wire  _GEN_217 = _T_3937 ? 1'h0 : _GEN_204; // @[Conditional.scala 39:67]
  wire  buf_cmd_state_bus_en_2 = _T_3914 ? 1'h0 : _GEN_217; // @[Conditional.scala 40:58]
  wire  _T_2617 = _T_2616 & buf_cmd_state_bus_en_2; // @[lsu_bus_buffer.scala 411:103]
  wire  _T_2618 = ~_T_2617; // @[lsu_bus_buffer.scala 411:78]
  wire  _T_2619 = buf_ageQ_3[2] & _T_2618; // @[lsu_bus_buffer.scala 411:76]
  wire  _T_2611 = buf_state_1 == 3'h2; // @[lsu_bus_buffer.scala 411:93]
  wire  _T_3721 = 3'h0 == buf_state_1; // @[Conditional.scala 37:30]
  wire  _T_3744 = 3'h1 == buf_state_1; // @[Conditional.scala 37:30]
  wire  _T_3748 = 3'h2 == buf_state_1; // @[Conditional.scala 37:30]
  wire  _T_3755 = obuf_tag0 == 3'h1; // @[lsu_bus_buffer.scala 454:48]
  wire  _T_3756 = _GEN_358 == 3'h1; // @[lsu_bus_buffer.scala 454:104]
  wire  _T_3757 = obuf_merge & _T_3756; // @[lsu_bus_buffer.scala 454:91]
  wire  _T_3758 = _T_3755 | _T_3757; // @[lsu_bus_buffer.scala 454:77]
  wire  _T_3759 = _T_3758 & obuf_valid; // @[lsu_bus_buffer.scala 454:135]
  wire  _T_3760 = _T_3759 & obuf_wr_enQ; // @[lsu_bus_buffer.scala 454:148]
  wire  _GEN_128 = _T_3748 & _T_3760; // @[Conditional.scala 39:67]
  wire  _GEN_141 = _T_3744 ? 1'h0 : _GEN_128; // @[Conditional.scala 39:67]
  wire  buf_cmd_state_bus_en_1 = _T_3721 ? 1'h0 : _GEN_141; // @[Conditional.scala 40:58]
  wire  _T_2612 = _T_2611 & buf_cmd_state_bus_en_1; // @[lsu_bus_buffer.scala 411:103]
  wire  _T_2613 = ~_T_2612; // @[lsu_bus_buffer.scala 411:78]
  wire  _T_2614 = buf_ageQ_3[1] & _T_2613; // @[lsu_bus_buffer.scala 411:76]
  wire  _T_2606 = buf_state_0 == 3'h2; // @[lsu_bus_buffer.scala 411:93]
  wire  _T_3528 = 3'h0 == buf_state_0; // @[Conditional.scala 37:30]
  wire  _T_3551 = 3'h1 == buf_state_0; // @[Conditional.scala 37:30]
  wire  _T_3555 = 3'h2 == buf_state_0; // @[Conditional.scala 37:30]
  wire  _T_3562 = obuf_tag0 == 3'h0; // @[lsu_bus_buffer.scala 454:48]
  wire  _T_3563 = _GEN_358 == 3'h0; // @[lsu_bus_buffer.scala 454:104]
  wire  _T_3564 = obuf_merge & _T_3563; // @[lsu_bus_buffer.scala 454:91]
  wire  _T_3565 = _T_3562 | _T_3564; // @[lsu_bus_buffer.scala 454:77]
  wire  _T_3566 = _T_3565 & obuf_valid; // @[lsu_bus_buffer.scala 454:135]
  wire  _T_3567 = _T_3566 & obuf_wr_enQ; // @[lsu_bus_buffer.scala 454:148]
  wire  _GEN_52 = _T_3555 & _T_3567; // @[Conditional.scala 39:67]
  wire  _GEN_65 = _T_3551 ? 1'h0 : _GEN_52; // @[Conditional.scala 39:67]
  wire  buf_cmd_state_bus_en_0 = _T_3528 ? 1'h0 : _GEN_65; // @[Conditional.scala 40:58]
  wire  _T_2607 = _T_2606 & buf_cmd_state_bus_en_0; // @[lsu_bus_buffer.scala 411:103]
  wire  _T_2608 = ~_T_2607; // @[lsu_bus_buffer.scala 411:78]
  wire  _T_2609 = buf_ageQ_3[0] & _T_2608; // @[lsu_bus_buffer.scala 411:76]
  wire [3:0] buf_age_3 = {_T_2624,_T_2619,_T_2614,_T_2609}; // @[Cat.scala 29:58]
  wire  _T_2723 = ~buf_age_3[2]; // @[lsu_bus_buffer.scala 412:89]
  wire  _T_2725 = _T_2723 & _T_19; // @[lsu_bus_buffer.scala 412:104]
  wire  _T_2717 = ~buf_age_3[1]; // @[lsu_bus_buffer.scala 412:89]
  wire  _T_2719 = _T_2717 & _T_12; // @[lsu_bus_buffer.scala 412:104]
  wire  _T_2711 = ~buf_age_3[0]; // @[lsu_bus_buffer.scala 412:89]
  wire  _T_2713 = _T_2711 & _T_5; // @[lsu_bus_buffer.scala 412:104]
  wire [3:0] buf_age_younger_3 = {1'h0,_T_2725,_T_2719,_T_2713}; // @[Cat.scala 29:58]
  wire [3:0] _T_255 = ld_byte_hitvec_lo_0 & buf_age_younger_3; // @[lsu_bus_buffer.scala 145:122]
  wire  _T_256 = |_T_255; // @[lsu_bus_buffer.scala 145:144]
  wire  _T_257 = ~_T_256; // @[lsu_bus_buffer.scala 145:99]
  wire  _T_258 = ld_byte_hitvec_lo_0[3] & _T_257; // @[lsu_bus_buffer.scala 145:97]
  reg [31:0] ibuf_addr; // @[lib.scala 374:16]
  wire  _T_512 = io_lsu_addr_m[31:2] == ibuf_addr[31:2]; // @[lsu_bus_buffer.scala 151:51]
  reg  ibuf_write; // @[Reg.scala 27:20]
  wire  _T_513 = _T_512 & ibuf_write; // @[lsu_bus_buffer.scala 151:73]
  reg  ibuf_valid; // @[lsu_bus_buffer.scala 238:54]
  wire  _T_514 = _T_513 & ibuf_valid; // @[lsu_bus_buffer.scala 151:86]
  wire  ld_addr_ibuf_hit_lo = _T_514 & io_lsu_busreq_m; // @[lsu_bus_buffer.scala 151:99]
  wire [3:0] _T_521 = ld_addr_ibuf_hit_lo ? 4'hf : 4'h0; // @[Bitwise.scala 72:12]
  reg [3:0] ibuf_byteen; // @[Reg.scala 27:20]
  wire [3:0] _T_522 = _T_521 & ibuf_byteen; // @[lsu_bus_buffer.scala 156:55]
  wire [3:0] ld_byte_ibuf_hit_lo = _T_522 & ldst_byteen_lo_m; // @[lsu_bus_buffer.scala 156:69]
  wire  _T_260 = ~ld_byte_ibuf_hit_lo[0]; // @[lsu_bus_buffer.scala 145:150]
  wire  _T_261 = _T_258 & _T_260; // @[lsu_bus_buffer.scala 145:148]
  reg [3:0] buf_ageQ_2; // @[lsu_bus_buffer.scala 499:60]
  wire  _T_2601 = buf_ageQ_2[3] & _T_2623; // @[lsu_bus_buffer.scala 411:76]
  wire  _T_2596 = buf_ageQ_2[2] & _T_2618; // @[lsu_bus_buffer.scala 411:76]
  wire  _T_2591 = buf_ageQ_2[1] & _T_2613; // @[lsu_bus_buffer.scala 411:76]
  wire  _T_2586 = buf_ageQ_2[0] & _T_2608; // @[lsu_bus_buffer.scala 411:76]
  wire [3:0] buf_age_2 = {_T_2601,_T_2596,_T_2591,_T_2586}; // @[Cat.scala 29:58]
  wire  _T_2702 = ~buf_age_2[3]; // @[lsu_bus_buffer.scala 412:89]
  wire  _T_2704 = _T_2702 & _T_26; // @[lsu_bus_buffer.scala 412:104]
  wire  _T_2690 = ~buf_age_2[1]; // @[lsu_bus_buffer.scala 412:89]
  wire  _T_2692 = _T_2690 & _T_12; // @[lsu_bus_buffer.scala 412:104]
  wire  _T_2684 = ~buf_age_2[0]; // @[lsu_bus_buffer.scala 412:89]
  wire  _T_2686 = _T_2684 & _T_5; // @[lsu_bus_buffer.scala 412:104]
  wire [3:0] buf_age_younger_2 = {_T_2704,1'h0,_T_2692,_T_2686}; // @[Cat.scala 29:58]
  wire [3:0] _T_247 = ld_byte_hitvec_lo_0 & buf_age_younger_2; // @[lsu_bus_buffer.scala 145:122]
  wire  _T_248 = |_T_247; // @[lsu_bus_buffer.scala 145:144]
  wire  _T_249 = ~_T_248; // @[lsu_bus_buffer.scala 145:99]
  wire  _T_250 = ld_byte_hitvec_lo_0[2] & _T_249; // @[lsu_bus_buffer.scala 145:97]
  wire  _T_253 = _T_250 & _T_260; // @[lsu_bus_buffer.scala 145:148]
  reg [3:0] buf_ageQ_1; // @[lsu_bus_buffer.scala 499:60]
  wire  _T_2578 = buf_ageQ_1[3] & _T_2623; // @[lsu_bus_buffer.scala 411:76]
  wire  _T_2573 = buf_ageQ_1[2] & _T_2618; // @[lsu_bus_buffer.scala 411:76]
  wire  _T_2568 = buf_ageQ_1[1] & _T_2613; // @[lsu_bus_buffer.scala 411:76]
  wire  _T_2563 = buf_ageQ_1[0] & _T_2608; // @[lsu_bus_buffer.scala 411:76]
  wire [3:0] buf_age_1 = {_T_2578,_T_2573,_T_2568,_T_2563}; // @[Cat.scala 29:58]
  wire  _T_2675 = ~buf_age_1[3]; // @[lsu_bus_buffer.scala 412:89]
  wire  _T_2677 = _T_2675 & _T_26; // @[lsu_bus_buffer.scala 412:104]
  wire  _T_2669 = ~buf_age_1[2]; // @[lsu_bus_buffer.scala 412:89]
  wire  _T_2671 = _T_2669 & _T_19; // @[lsu_bus_buffer.scala 412:104]
  wire  _T_2657 = ~buf_age_1[0]; // @[lsu_bus_buffer.scala 412:89]
  wire  _T_2659 = _T_2657 & _T_5; // @[lsu_bus_buffer.scala 412:104]
  wire [3:0] buf_age_younger_1 = {_T_2677,_T_2671,1'h0,_T_2659}; // @[Cat.scala 29:58]
  wire [3:0] _T_239 = ld_byte_hitvec_lo_0 & buf_age_younger_1; // @[lsu_bus_buffer.scala 145:122]
  wire  _T_240 = |_T_239; // @[lsu_bus_buffer.scala 145:144]
  wire  _T_241 = ~_T_240; // @[lsu_bus_buffer.scala 145:99]
  wire  _T_242 = ld_byte_hitvec_lo_0[1] & _T_241; // @[lsu_bus_buffer.scala 145:97]
  wire  _T_245 = _T_242 & _T_260; // @[lsu_bus_buffer.scala 145:148]
  reg [3:0] buf_ageQ_0; // @[lsu_bus_buffer.scala 499:60]
  wire  _T_2555 = buf_ageQ_0[3] & _T_2623; // @[lsu_bus_buffer.scala 411:76]
  wire  _T_2550 = buf_ageQ_0[2] & _T_2618; // @[lsu_bus_buffer.scala 411:76]
  wire  _T_2545 = buf_ageQ_0[1] & _T_2613; // @[lsu_bus_buffer.scala 411:76]
  wire  _T_2540 = buf_ageQ_0[0] & _T_2608; // @[lsu_bus_buffer.scala 411:76]
  wire [3:0] buf_age_0 = {_T_2555,_T_2550,_T_2545,_T_2540}; // @[Cat.scala 29:58]
  wire  _T_2648 = ~buf_age_0[3]; // @[lsu_bus_buffer.scala 412:89]
  wire  _T_2650 = _T_2648 & _T_26; // @[lsu_bus_buffer.scala 412:104]
  wire  _T_2642 = ~buf_age_0[2]; // @[lsu_bus_buffer.scala 412:89]
  wire  _T_2644 = _T_2642 & _T_19; // @[lsu_bus_buffer.scala 412:104]
  wire  _T_2636 = ~buf_age_0[1]; // @[lsu_bus_buffer.scala 412:89]
  wire  _T_2638 = _T_2636 & _T_12; // @[lsu_bus_buffer.scala 412:104]
  wire [3:0] buf_age_younger_0 = {_T_2650,_T_2644,_T_2638,1'h0}; // @[Cat.scala 29:58]
  wire [3:0] _T_231 = ld_byte_hitvec_lo_0 & buf_age_younger_0; // @[lsu_bus_buffer.scala 145:122]
  wire  _T_232 = |_T_231; // @[lsu_bus_buffer.scala 145:144]
  wire  _T_233 = ~_T_232; // @[lsu_bus_buffer.scala 145:99]
  wire  _T_234 = ld_byte_hitvec_lo_0[0] & _T_233; // @[lsu_bus_buffer.scala 145:97]
  wire  _T_237 = _T_234 & _T_260; // @[lsu_bus_buffer.scala 145:148]
  wire [3:0] ld_byte_hitvecfn_lo_0 = {_T_261,_T_253,_T_245,_T_237}; // @[Cat.scala 29:58]
  wire  _T_56 = |ld_byte_hitvecfn_lo_0; // @[lsu_bus_buffer.scala 137:73]
  wire  _T_58 = _T_56 | ld_byte_ibuf_hit_lo[0]; // @[lsu_bus_buffer.scala 137:77]
  wire  _T_117 = ld_addr_hitvec_lo_3 & buf_byteen_3[1]; // @[lsu_bus_buffer.scala 140:95]
  wire  _T_119 = _T_117 & ldst_byteen_lo_m[1]; // @[lsu_bus_buffer.scala 140:114]
  wire  _T_113 = ld_addr_hitvec_lo_2 & buf_byteen_2[1]; // @[lsu_bus_buffer.scala 140:95]
  wire  _T_115 = _T_113 & ldst_byteen_lo_m[1]; // @[lsu_bus_buffer.scala 140:114]
  wire  _T_109 = ld_addr_hitvec_lo_1 & buf_byteen_1[1]; // @[lsu_bus_buffer.scala 140:95]
  wire  _T_111 = _T_109 & ldst_byteen_lo_m[1]; // @[lsu_bus_buffer.scala 140:114]
  wire  _T_105 = ld_addr_hitvec_lo_0 & buf_byteen_0[1]; // @[lsu_bus_buffer.scala 140:95]
  wire  _T_107 = _T_105 & ldst_byteen_lo_m[1]; // @[lsu_bus_buffer.scala 140:114]
  wire [3:0] ld_byte_hitvec_lo_1 = {_T_119,_T_115,_T_111,_T_107}; // @[Cat.scala 29:58]
  wire [3:0] _T_290 = ld_byte_hitvec_lo_1 & buf_age_younger_3; // @[lsu_bus_buffer.scala 145:122]
  wire  _T_291 = |_T_290; // @[lsu_bus_buffer.scala 145:144]
  wire  _T_292 = ~_T_291; // @[lsu_bus_buffer.scala 145:99]
  wire  _T_293 = ld_byte_hitvec_lo_1[3] & _T_292; // @[lsu_bus_buffer.scala 145:97]
  wire  _T_295 = ~ld_byte_ibuf_hit_lo[1]; // @[lsu_bus_buffer.scala 145:150]
  wire  _T_296 = _T_293 & _T_295; // @[lsu_bus_buffer.scala 145:148]
  wire [3:0] _T_282 = ld_byte_hitvec_lo_1 & buf_age_younger_2; // @[lsu_bus_buffer.scala 145:122]
  wire  _T_283 = |_T_282; // @[lsu_bus_buffer.scala 145:144]
  wire  _T_284 = ~_T_283; // @[lsu_bus_buffer.scala 145:99]
  wire  _T_285 = ld_byte_hitvec_lo_1[2] & _T_284; // @[lsu_bus_buffer.scala 145:97]
  wire  _T_288 = _T_285 & _T_295; // @[lsu_bus_buffer.scala 145:148]
  wire [3:0] _T_274 = ld_byte_hitvec_lo_1 & buf_age_younger_1; // @[lsu_bus_buffer.scala 145:122]
  wire  _T_275 = |_T_274; // @[lsu_bus_buffer.scala 145:144]
  wire  _T_276 = ~_T_275; // @[lsu_bus_buffer.scala 145:99]
  wire  _T_277 = ld_byte_hitvec_lo_1[1] & _T_276; // @[lsu_bus_buffer.scala 145:97]
  wire  _T_280 = _T_277 & _T_295; // @[lsu_bus_buffer.scala 145:148]
  wire [3:0] _T_266 = ld_byte_hitvec_lo_1 & buf_age_younger_0; // @[lsu_bus_buffer.scala 145:122]
  wire  _T_267 = |_T_266; // @[lsu_bus_buffer.scala 145:144]
  wire  _T_268 = ~_T_267; // @[lsu_bus_buffer.scala 145:99]
  wire  _T_269 = ld_byte_hitvec_lo_1[0] & _T_268; // @[lsu_bus_buffer.scala 145:97]
  wire  _T_272 = _T_269 & _T_295; // @[lsu_bus_buffer.scala 145:148]
  wire [3:0] ld_byte_hitvecfn_lo_1 = {_T_296,_T_288,_T_280,_T_272}; // @[Cat.scala 29:58]
  wire  _T_59 = |ld_byte_hitvecfn_lo_1; // @[lsu_bus_buffer.scala 137:73]
  wire  _T_61 = _T_59 | ld_byte_ibuf_hit_lo[1]; // @[lsu_bus_buffer.scala 137:77]
  wire  _T_135 = ld_addr_hitvec_lo_3 & buf_byteen_3[2]; // @[lsu_bus_buffer.scala 140:95]
  wire  _T_137 = _T_135 & ldst_byteen_lo_m[2]; // @[lsu_bus_buffer.scala 140:114]
  wire  _T_131 = ld_addr_hitvec_lo_2 & buf_byteen_2[2]; // @[lsu_bus_buffer.scala 140:95]
  wire  _T_133 = _T_131 & ldst_byteen_lo_m[2]; // @[lsu_bus_buffer.scala 140:114]
  wire  _T_127 = ld_addr_hitvec_lo_1 & buf_byteen_1[2]; // @[lsu_bus_buffer.scala 140:95]
  wire  _T_129 = _T_127 & ldst_byteen_lo_m[2]; // @[lsu_bus_buffer.scala 140:114]
  wire  _T_123 = ld_addr_hitvec_lo_0 & buf_byteen_0[2]; // @[lsu_bus_buffer.scala 140:95]
  wire  _T_125 = _T_123 & ldst_byteen_lo_m[2]; // @[lsu_bus_buffer.scala 140:114]
  wire [3:0] ld_byte_hitvec_lo_2 = {_T_137,_T_133,_T_129,_T_125}; // @[Cat.scala 29:58]
  wire [3:0] _T_325 = ld_byte_hitvec_lo_2 & buf_age_younger_3; // @[lsu_bus_buffer.scala 145:122]
  wire  _T_326 = |_T_325; // @[lsu_bus_buffer.scala 145:144]
  wire  _T_327 = ~_T_326; // @[lsu_bus_buffer.scala 145:99]
  wire  _T_328 = ld_byte_hitvec_lo_2[3] & _T_327; // @[lsu_bus_buffer.scala 145:97]
  wire  _T_330 = ~ld_byte_ibuf_hit_lo[2]; // @[lsu_bus_buffer.scala 145:150]
  wire  _T_331 = _T_328 & _T_330; // @[lsu_bus_buffer.scala 145:148]
  wire [3:0] _T_317 = ld_byte_hitvec_lo_2 & buf_age_younger_2; // @[lsu_bus_buffer.scala 145:122]
  wire  _T_318 = |_T_317; // @[lsu_bus_buffer.scala 145:144]
  wire  _T_319 = ~_T_318; // @[lsu_bus_buffer.scala 145:99]
  wire  _T_320 = ld_byte_hitvec_lo_2[2] & _T_319; // @[lsu_bus_buffer.scala 145:97]
  wire  _T_323 = _T_320 & _T_330; // @[lsu_bus_buffer.scala 145:148]
  wire [3:0] _T_309 = ld_byte_hitvec_lo_2 & buf_age_younger_1; // @[lsu_bus_buffer.scala 145:122]
  wire  _T_310 = |_T_309; // @[lsu_bus_buffer.scala 145:144]
  wire  _T_311 = ~_T_310; // @[lsu_bus_buffer.scala 145:99]
  wire  _T_312 = ld_byte_hitvec_lo_2[1] & _T_311; // @[lsu_bus_buffer.scala 145:97]
  wire  _T_315 = _T_312 & _T_330; // @[lsu_bus_buffer.scala 145:148]
  wire [3:0] _T_301 = ld_byte_hitvec_lo_2 & buf_age_younger_0; // @[lsu_bus_buffer.scala 145:122]
  wire  _T_302 = |_T_301; // @[lsu_bus_buffer.scala 145:144]
  wire  _T_303 = ~_T_302; // @[lsu_bus_buffer.scala 145:99]
  wire  _T_304 = ld_byte_hitvec_lo_2[0] & _T_303; // @[lsu_bus_buffer.scala 145:97]
  wire  _T_307 = _T_304 & _T_330; // @[lsu_bus_buffer.scala 145:148]
  wire [3:0] ld_byte_hitvecfn_lo_2 = {_T_331,_T_323,_T_315,_T_307}; // @[Cat.scala 29:58]
  wire  _T_62 = |ld_byte_hitvecfn_lo_2; // @[lsu_bus_buffer.scala 137:73]
  wire  _T_64 = _T_62 | ld_byte_ibuf_hit_lo[2]; // @[lsu_bus_buffer.scala 137:77]
  wire  _T_153 = ld_addr_hitvec_lo_3 & buf_byteen_3[3]; // @[lsu_bus_buffer.scala 140:95]
  wire  _T_155 = _T_153 & ldst_byteen_lo_m[3]; // @[lsu_bus_buffer.scala 140:114]
  wire  _T_149 = ld_addr_hitvec_lo_2 & buf_byteen_2[3]; // @[lsu_bus_buffer.scala 140:95]
  wire  _T_151 = _T_149 & ldst_byteen_lo_m[3]; // @[lsu_bus_buffer.scala 140:114]
  wire  _T_145 = ld_addr_hitvec_lo_1 & buf_byteen_1[3]; // @[lsu_bus_buffer.scala 140:95]
  wire  _T_147 = _T_145 & ldst_byteen_lo_m[3]; // @[lsu_bus_buffer.scala 140:114]
  wire  _T_141 = ld_addr_hitvec_lo_0 & buf_byteen_0[3]; // @[lsu_bus_buffer.scala 140:95]
  wire  _T_143 = _T_141 & ldst_byteen_lo_m[3]; // @[lsu_bus_buffer.scala 140:114]
  wire [3:0] ld_byte_hitvec_lo_3 = {_T_155,_T_151,_T_147,_T_143}; // @[Cat.scala 29:58]
  wire [3:0] _T_360 = ld_byte_hitvec_lo_3 & buf_age_younger_3; // @[lsu_bus_buffer.scala 145:122]
  wire  _T_361 = |_T_360; // @[lsu_bus_buffer.scala 145:144]
  wire  _T_362 = ~_T_361; // @[lsu_bus_buffer.scala 145:99]
  wire  _T_363 = ld_byte_hitvec_lo_3[3] & _T_362; // @[lsu_bus_buffer.scala 145:97]
  wire  _T_365 = ~ld_byte_ibuf_hit_lo[3]; // @[lsu_bus_buffer.scala 145:150]
  wire  _T_366 = _T_363 & _T_365; // @[lsu_bus_buffer.scala 145:148]
  wire [3:0] _T_352 = ld_byte_hitvec_lo_3 & buf_age_younger_2; // @[lsu_bus_buffer.scala 145:122]
  wire  _T_353 = |_T_352; // @[lsu_bus_buffer.scala 145:144]
  wire  _T_354 = ~_T_353; // @[lsu_bus_buffer.scala 145:99]
  wire  _T_355 = ld_byte_hitvec_lo_3[2] & _T_354; // @[lsu_bus_buffer.scala 145:97]
  wire  _T_358 = _T_355 & _T_365; // @[lsu_bus_buffer.scala 145:148]
  wire [3:0] _T_344 = ld_byte_hitvec_lo_3 & buf_age_younger_1; // @[lsu_bus_buffer.scala 145:122]
  wire  _T_345 = |_T_344; // @[lsu_bus_buffer.scala 145:144]
  wire  _T_346 = ~_T_345; // @[lsu_bus_buffer.scala 145:99]
  wire  _T_347 = ld_byte_hitvec_lo_3[1] & _T_346; // @[lsu_bus_buffer.scala 145:97]
  wire  _T_350 = _T_347 & _T_365; // @[lsu_bus_buffer.scala 145:148]
  wire [3:0] _T_336 = ld_byte_hitvec_lo_3 & buf_age_younger_0; // @[lsu_bus_buffer.scala 145:122]
  wire  _T_337 = |_T_336; // @[lsu_bus_buffer.scala 145:144]
  wire  _T_338 = ~_T_337; // @[lsu_bus_buffer.scala 145:99]
  wire  _T_339 = ld_byte_hitvec_lo_3[0] & _T_338; // @[lsu_bus_buffer.scala 145:97]
  wire  _T_342 = _T_339 & _T_365; // @[lsu_bus_buffer.scala 145:148]
  wire [3:0] ld_byte_hitvecfn_lo_3 = {_T_366,_T_358,_T_350,_T_342}; // @[Cat.scala 29:58]
  wire  _T_65 = |ld_byte_hitvecfn_lo_3; // @[lsu_bus_buffer.scala 137:73]
  wire  _T_67 = _T_65 | ld_byte_ibuf_hit_lo[3]; // @[lsu_bus_buffer.scala 137:77]
  wire [2:0] _T_69 = {_T_67,_T_64,_T_61}; // @[Cat.scala 29:58]
  wire  _T_171 = ld_addr_hitvec_hi_3 & buf_byteen_3[0]; // @[lsu_bus_buffer.scala 141:95]
  wire  _T_173 = _T_171 & ldst_byteen_hi_m[0]; // @[lsu_bus_buffer.scala 141:114]
  wire  _T_167 = ld_addr_hitvec_hi_2 & buf_byteen_2[0]; // @[lsu_bus_buffer.scala 141:95]
  wire  _T_169 = _T_167 & ldst_byteen_hi_m[0]; // @[lsu_bus_buffer.scala 141:114]
  wire  _T_163 = ld_addr_hitvec_hi_1 & buf_byteen_1[0]; // @[lsu_bus_buffer.scala 141:95]
  wire  _T_165 = _T_163 & ldst_byteen_hi_m[0]; // @[lsu_bus_buffer.scala 141:114]
  wire  _T_159 = ld_addr_hitvec_hi_0 & buf_byteen_0[0]; // @[lsu_bus_buffer.scala 141:95]
  wire  _T_161 = _T_159 & ldst_byteen_hi_m[0]; // @[lsu_bus_buffer.scala 141:114]
  wire [3:0] ld_byte_hitvec_hi_0 = {_T_173,_T_169,_T_165,_T_161}; // @[Cat.scala 29:58]
  wire [3:0] _T_395 = ld_byte_hitvec_hi_0 & buf_age_younger_3; // @[lsu_bus_buffer.scala 146:122]
  wire  _T_396 = |_T_395; // @[lsu_bus_buffer.scala 146:144]
  wire  _T_397 = ~_T_396; // @[lsu_bus_buffer.scala 146:99]
  wire  _T_398 = ld_byte_hitvec_hi_0[3] & _T_397; // @[lsu_bus_buffer.scala 146:97]
  wire  _T_517 = io_end_addr_m[31:2] == ibuf_addr[31:2]; // @[lsu_bus_buffer.scala 152:51]
  wire  _T_518 = _T_517 & ibuf_write; // @[lsu_bus_buffer.scala 152:73]
  wire  _T_519 = _T_518 & ibuf_valid; // @[lsu_bus_buffer.scala 152:86]
  wire  ld_addr_ibuf_hit_hi = _T_519 & io_lsu_busreq_m; // @[lsu_bus_buffer.scala 152:99]
  wire [3:0] _T_525 = ld_addr_ibuf_hit_hi ? 4'hf : 4'h0; // @[Bitwise.scala 72:12]
  wire [3:0] _T_526 = _T_525 & ibuf_byteen; // @[lsu_bus_buffer.scala 157:55]
  wire [3:0] ld_byte_ibuf_hit_hi = _T_526 & ldst_byteen_hi_m; // @[lsu_bus_buffer.scala 157:69]
  wire  _T_400 = ~ld_byte_ibuf_hit_hi[0]; // @[lsu_bus_buffer.scala 146:150]
  wire  _T_401 = _T_398 & _T_400; // @[lsu_bus_buffer.scala 146:148]
  wire [3:0] _T_387 = ld_byte_hitvec_hi_0 & buf_age_younger_2; // @[lsu_bus_buffer.scala 146:122]
  wire  _T_388 = |_T_387; // @[lsu_bus_buffer.scala 146:144]
  wire  _T_389 = ~_T_388; // @[lsu_bus_buffer.scala 146:99]
  wire  _T_390 = ld_byte_hitvec_hi_0[2] & _T_389; // @[lsu_bus_buffer.scala 146:97]
  wire  _T_393 = _T_390 & _T_400; // @[lsu_bus_buffer.scala 146:148]
  wire [3:0] _T_379 = ld_byte_hitvec_hi_0 & buf_age_younger_1; // @[lsu_bus_buffer.scala 146:122]
  wire  _T_380 = |_T_379; // @[lsu_bus_buffer.scala 146:144]
  wire  _T_381 = ~_T_380; // @[lsu_bus_buffer.scala 146:99]
  wire  _T_382 = ld_byte_hitvec_hi_0[1] & _T_381; // @[lsu_bus_buffer.scala 146:97]
  wire  _T_385 = _T_382 & _T_400; // @[lsu_bus_buffer.scala 146:148]
  wire [3:0] _T_371 = ld_byte_hitvec_hi_0 & buf_age_younger_0; // @[lsu_bus_buffer.scala 146:122]
  wire  _T_372 = |_T_371; // @[lsu_bus_buffer.scala 146:144]
  wire  _T_373 = ~_T_372; // @[lsu_bus_buffer.scala 146:99]
  wire  _T_374 = ld_byte_hitvec_hi_0[0] & _T_373; // @[lsu_bus_buffer.scala 146:97]
  wire  _T_377 = _T_374 & _T_400; // @[lsu_bus_buffer.scala 146:148]
  wire [3:0] ld_byte_hitvecfn_hi_0 = {_T_401,_T_393,_T_385,_T_377}; // @[Cat.scala 29:58]
  wire  _T_71 = |ld_byte_hitvecfn_hi_0; // @[lsu_bus_buffer.scala 138:73]
  wire  _T_73 = _T_71 | ld_byte_ibuf_hit_hi[0]; // @[lsu_bus_buffer.scala 138:77]
  wire  _T_189 = ld_addr_hitvec_hi_3 & buf_byteen_3[1]; // @[lsu_bus_buffer.scala 141:95]
  wire  _T_191 = _T_189 & ldst_byteen_hi_m[1]; // @[lsu_bus_buffer.scala 141:114]
  wire  _T_185 = ld_addr_hitvec_hi_2 & buf_byteen_2[1]; // @[lsu_bus_buffer.scala 141:95]
  wire  _T_187 = _T_185 & ldst_byteen_hi_m[1]; // @[lsu_bus_buffer.scala 141:114]
  wire  _T_181 = ld_addr_hitvec_hi_1 & buf_byteen_1[1]; // @[lsu_bus_buffer.scala 141:95]
  wire  _T_183 = _T_181 & ldst_byteen_hi_m[1]; // @[lsu_bus_buffer.scala 141:114]
  wire  _T_177 = ld_addr_hitvec_hi_0 & buf_byteen_0[1]; // @[lsu_bus_buffer.scala 141:95]
  wire  _T_179 = _T_177 & ldst_byteen_hi_m[1]; // @[lsu_bus_buffer.scala 141:114]
  wire [3:0] ld_byte_hitvec_hi_1 = {_T_191,_T_187,_T_183,_T_179}; // @[Cat.scala 29:58]
  wire [3:0] _T_430 = ld_byte_hitvec_hi_1 & buf_age_younger_3; // @[lsu_bus_buffer.scala 146:122]
  wire  _T_431 = |_T_430; // @[lsu_bus_buffer.scala 146:144]
  wire  _T_432 = ~_T_431; // @[lsu_bus_buffer.scala 146:99]
  wire  _T_433 = ld_byte_hitvec_hi_1[3] & _T_432; // @[lsu_bus_buffer.scala 146:97]
  wire  _T_435 = ~ld_byte_ibuf_hit_hi[1]; // @[lsu_bus_buffer.scala 146:150]
  wire  _T_436 = _T_433 & _T_435; // @[lsu_bus_buffer.scala 146:148]
  wire [3:0] _T_422 = ld_byte_hitvec_hi_1 & buf_age_younger_2; // @[lsu_bus_buffer.scala 146:122]
  wire  _T_423 = |_T_422; // @[lsu_bus_buffer.scala 146:144]
  wire  _T_424 = ~_T_423; // @[lsu_bus_buffer.scala 146:99]
  wire  _T_425 = ld_byte_hitvec_hi_1[2] & _T_424; // @[lsu_bus_buffer.scala 146:97]
  wire  _T_428 = _T_425 & _T_435; // @[lsu_bus_buffer.scala 146:148]
  wire [3:0] _T_414 = ld_byte_hitvec_hi_1 & buf_age_younger_1; // @[lsu_bus_buffer.scala 146:122]
  wire  _T_415 = |_T_414; // @[lsu_bus_buffer.scala 146:144]
  wire  _T_416 = ~_T_415; // @[lsu_bus_buffer.scala 146:99]
  wire  _T_417 = ld_byte_hitvec_hi_1[1] & _T_416; // @[lsu_bus_buffer.scala 146:97]
  wire  _T_420 = _T_417 & _T_435; // @[lsu_bus_buffer.scala 146:148]
  wire [3:0] _T_406 = ld_byte_hitvec_hi_1 & buf_age_younger_0; // @[lsu_bus_buffer.scala 146:122]
  wire  _T_407 = |_T_406; // @[lsu_bus_buffer.scala 146:144]
  wire  _T_408 = ~_T_407; // @[lsu_bus_buffer.scala 146:99]
  wire  _T_409 = ld_byte_hitvec_hi_1[0] & _T_408; // @[lsu_bus_buffer.scala 146:97]
  wire  _T_412 = _T_409 & _T_435; // @[lsu_bus_buffer.scala 146:148]
  wire [3:0] ld_byte_hitvecfn_hi_1 = {_T_436,_T_428,_T_420,_T_412}; // @[Cat.scala 29:58]
  wire  _T_74 = |ld_byte_hitvecfn_hi_1; // @[lsu_bus_buffer.scala 138:73]
  wire  _T_76 = _T_74 | ld_byte_ibuf_hit_hi[1]; // @[lsu_bus_buffer.scala 138:77]
  wire  _T_207 = ld_addr_hitvec_hi_3 & buf_byteen_3[2]; // @[lsu_bus_buffer.scala 141:95]
  wire  _T_209 = _T_207 & ldst_byteen_hi_m[2]; // @[lsu_bus_buffer.scala 141:114]
  wire  _T_203 = ld_addr_hitvec_hi_2 & buf_byteen_2[2]; // @[lsu_bus_buffer.scala 141:95]
  wire  _T_205 = _T_203 & ldst_byteen_hi_m[2]; // @[lsu_bus_buffer.scala 141:114]
  wire  _T_199 = ld_addr_hitvec_hi_1 & buf_byteen_1[2]; // @[lsu_bus_buffer.scala 141:95]
  wire  _T_201 = _T_199 & ldst_byteen_hi_m[2]; // @[lsu_bus_buffer.scala 141:114]
  wire  _T_195 = ld_addr_hitvec_hi_0 & buf_byteen_0[2]; // @[lsu_bus_buffer.scala 141:95]
  wire  _T_197 = _T_195 & ldst_byteen_hi_m[2]; // @[lsu_bus_buffer.scala 141:114]
  wire [3:0] ld_byte_hitvec_hi_2 = {_T_209,_T_205,_T_201,_T_197}; // @[Cat.scala 29:58]
  wire [3:0] _T_465 = ld_byte_hitvec_hi_2 & buf_age_younger_3; // @[lsu_bus_buffer.scala 146:122]
  wire  _T_466 = |_T_465; // @[lsu_bus_buffer.scala 146:144]
  wire  _T_467 = ~_T_466; // @[lsu_bus_buffer.scala 146:99]
  wire  _T_468 = ld_byte_hitvec_hi_2[3] & _T_467; // @[lsu_bus_buffer.scala 146:97]
  wire  _T_470 = ~ld_byte_ibuf_hit_hi[2]; // @[lsu_bus_buffer.scala 146:150]
  wire  _T_471 = _T_468 & _T_470; // @[lsu_bus_buffer.scala 146:148]
  wire [3:0] _T_457 = ld_byte_hitvec_hi_2 & buf_age_younger_2; // @[lsu_bus_buffer.scala 146:122]
  wire  _T_458 = |_T_457; // @[lsu_bus_buffer.scala 146:144]
  wire  _T_459 = ~_T_458; // @[lsu_bus_buffer.scala 146:99]
  wire  _T_460 = ld_byte_hitvec_hi_2[2] & _T_459; // @[lsu_bus_buffer.scala 146:97]
  wire  _T_463 = _T_460 & _T_470; // @[lsu_bus_buffer.scala 146:148]
  wire [3:0] _T_449 = ld_byte_hitvec_hi_2 & buf_age_younger_1; // @[lsu_bus_buffer.scala 146:122]
  wire  _T_450 = |_T_449; // @[lsu_bus_buffer.scala 146:144]
  wire  _T_451 = ~_T_450; // @[lsu_bus_buffer.scala 146:99]
  wire  _T_452 = ld_byte_hitvec_hi_2[1] & _T_451; // @[lsu_bus_buffer.scala 146:97]
  wire  _T_455 = _T_452 & _T_470; // @[lsu_bus_buffer.scala 146:148]
  wire [3:0] _T_441 = ld_byte_hitvec_hi_2 & buf_age_younger_0; // @[lsu_bus_buffer.scala 146:122]
  wire  _T_442 = |_T_441; // @[lsu_bus_buffer.scala 146:144]
  wire  _T_443 = ~_T_442; // @[lsu_bus_buffer.scala 146:99]
  wire  _T_444 = ld_byte_hitvec_hi_2[0] & _T_443; // @[lsu_bus_buffer.scala 146:97]
  wire  _T_447 = _T_444 & _T_470; // @[lsu_bus_buffer.scala 146:148]
  wire [3:0] ld_byte_hitvecfn_hi_2 = {_T_471,_T_463,_T_455,_T_447}; // @[Cat.scala 29:58]
  wire  _T_77 = |ld_byte_hitvecfn_hi_2; // @[lsu_bus_buffer.scala 138:73]
  wire  _T_79 = _T_77 | ld_byte_ibuf_hit_hi[2]; // @[lsu_bus_buffer.scala 138:77]
  wire  _T_225 = ld_addr_hitvec_hi_3 & buf_byteen_3[3]; // @[lsu_bus_buffer.scala 141:95]
  wire  _T_227 = _T_225 & ldst_byteen_hi_m[3]; // @[lsu_bus_buffer.scala 141:114]
  wire  _T_221 = ld_addr_hitvec_hi_2 & buf_byteen_2[3]; // @[lsu_bus_buffer.scala 141:95]
  wire  _T_223 = _T_221 & ldst_byteen_hi_m[3]; // @[lsu_bus_buffer.scala 141:114]
  wire  _T_217 = ld_addr_hitvec_hi_1 & buf_byteen_1[3]; // @[lsu_bus_buffer.scala 141:95]
  wire  _T_219 = _T_217 & ldst_byteen_hi_m[3]; // @[lsu_bus_buffer.scala 141:114]
  wire  _T_213 = ld_addr_hitvec_hi_0 & buf_byteen_0[3]; // @[lsu_bus_buffer.scala 141:95]
  wire  _T_215 = _T_213 & ldst_byteen_hi_m[3]; // @[lsu_bus_buffer.scala 141:114]
  wire [3:0] ld_byte_hitvec_hi_3 = {_T_227,_T_223,_T_219,_T_215}; // @[Cat.scala 29:58]
  wire [3:0] _T_500 = ld_byte_hitvec_hi_3 & buf_age_younger_3; // @[lsu_bus_buffer.scala 146:122]
  wire  _T_501 = |_T_500; // @[lsu_bus_buffer.scala 146:144]
  wire  _T_502 = ~_T_501; // @[lsu_bus_buffer.scala 146:99]
  wire  _T_503 = ld_byte_hitvec_hi_3[3] & _T_502; // @[lsu_bus_buffer.scala 146:97]
  wire  _T_505 = ~ld_byte_ibuf_hit_hi[3]; // @[lsu_bus_buffer.scala 146:150]
  wire  _T_506 = _T_503 & _T_505; // @[lsu_bus_buffer.scala 146:148]
  wire [3:0] _T_492 = ld_byte_hitvec_hi_3 & buf_age_younger_2; // @[lsu_bus_buffer.scala 146:122]
  wire  _T_493 = |_T_492; // @[lsu_bus_buffer.scala 146:144]
  wire  _T_494 = ~_T_493; // @[lsu_bus_buffer.scala 146:99]
  wire  _T_495 = ld_byte_hitvec_hi_3[2] & _T_494; // @[lsu_bus_buffer.scala 146:97]
  wire  _T_498 = _T_495 & _T_505; // @[lsu_bus_buffer.scala 146:148]
  wire [3:0] _T_484 = ld_byte_hitvec_hi_3 & buf_age_younger_1; // @[lsu_bus_buffer.scala 146:122]
  wire  _T_485 = |_T_484; // @[lsu_bus_buffer.scala 146:144]
  wire  _T_486 = ~_T_485; // @[lsu_bus_buffer.scala 146:99]
  wire  _T_487 = ld_byte_hitvec_hi_3[1] & _T_486; // @[lsu_bus_buffer.scala 146:97]
  wire  _T_490 = _T_487 & _T_505; // @[lsu_bus_buffer.scala 146:148]
  wire [3:0] _T_476 = ld_byte_hitvec_hi_3 & buf_age_younger_0; // @[lsu_bus_buffer.scala 146:122]
  wire  _T_477 = |_T_476; // @[lsu_bus_buffer.scala 146:144]
  wire  _T_478 = ~_T_477; // @[lsu_bus_buffer.scala 146:99]
  wire  _T_479 = ld_byte_hitvec_hi_3[0] & _T_478; // @[lsu_bus_buffer.scala 146:97]
  wire  _T_482 = _T_479 & _T_505; // @[lsu_bus_buffer.scala 146:148]
  wire [3:0] ld_byte_hitvecfn_hi_3 = {_T_506,_T_498,_T_490,_T_482}; // @[Cat.scala 29:58]
  wire  _T_80 = |ld_byte_hitvecfn_hi_3; // @[lsu_bus_buffer.scala 138:73]
  wire  _T_82 = _T_80 | ld_byte_ibuf_hit_hi[3]; // @[lsu_bus_buffer.scala 138:77]
  wire [2:0] _T_84 = {_T_82,_T_79,_T_76}; // @[Cat.scala 29:58]
  wire [7:0] _T_530 = ld_byte_ibuf_hit_lo[0] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_533 = ld_byte_ibuf_hit_lo[1] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_536 = ld_byte_ibuf_hit_lo[2] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_539 = ld_byte_ibuf_hit_lo[3] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [31:0] ld_fwddata_buf_lo_initial = {_T_539,_T_536,_T_533,_T_530}; // @[Cat.scala 29:58]
  wire [7:0] _T_544 = ld_byte_ibuf_hit_hi[0] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_547 = ld_byte_ibuf_hit_hi[1] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_550 = ld_byte_ibuf_hit_hi[2] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_553 = ld_byte_ibuf_hit_hi[3] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [31:0] ld_fwddata_buf_hi_initial = {_T_553,_T_550,_T_547,_T_544}; // @[Cat.scala 29:58]
  wire [7:0] _T_558 = ld_byte_hitvecfn_lo_3[0] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  reg [31:0] buf_data_0; // @[lib.scala 374:16]
  wire [7:0] _T_560 = _T_558 & buf_data_0[31:24]; // @[lsu_bus_buffer.scala 164:91]
  wire [7:0] _T_563 = ld_byte_hitvecfn_lo_3[1] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  reg [31:0] buf_data_1; // @[lib.scala 374:16]
  wire [7:0] _T_565 = _T_563 & buf_data_1[31:24]; // @[lsu_bus_buffer.scala 164:91]
  wire [7:0] _T_568 = ld_byte_hitvecfn_lo_3[2] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  reg [31:0] buf_data_2; // @[lib.scala 374:16]
  wire [7:0] _T_570 = _T_568 & buf_data_2[31:24]; // @[lsu_bus_buffer.scala 164:91]
  wire [7:0] _T_573 = ld_byte_hitvecfn_lo_3[3] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  reg [31:0] buf_data_3; // @[lib.scala 374:16]
  wire [7:0] _T_575 = _T_573 & buf_data_3[31:24]; // @[lsu_bus_buffer.scala 164:91]
  wire [7:0] _T_576 = _T_560 | _T_565; // @[lsu_bus_buffer.scala 164:123]
  wire [7:0] _T_577 = _T_576 | _T_570; // @[lsu_bus_buffer.scala 164:123]
  wire [7:0] _T_578 = _T_577 | _T_575; // @[lsu_bus_buffer.scala 164:123]
  wire [7:0] _T_581 = ld_byte_hitvecfn_lo_2[0] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_583 = _T_581 & buf_data_0[23:16]; // @[lsu_bus_buffer.scala 165:65]
  wire [7:0] _T_586 = ld_byte_hitvecfn_lo_2[1] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_588 = _T_586 & buf_data_1[23:16]; // @[lsu_bus_buffer.scala 165:65]
  wire [7:0] _T_591 = ld_byte_hitvecfn_lo_2[2] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_593 = _T_591 & buf_data_2[23:16]; // @[lsu_bus_buffer.scala 165:65]
  wire [7:0] _T_596 = ld_byte_hitvecfn_lo_2[3] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_598 = _T_596 & buf_data_3[23:16]; // @[lsu_bus_buffer.scala 165:65]
  wire [7:0] _T_599 = _T_583 | _T_588; // @[lsu_bus_buffer.scala 165:97]
  wire [7:0] _T_600 = _T_599 | _T_593; // @[lsu_bus_buffer.scala 165:97]
  wire [7:0] _T_601 = _T_600 | _T_598; // @[lsu_bus_buffer.scala 165:97]
  wire [7:0] _T_604 = ld_byte_hitvecfn_lo_1[0] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_606 = _T_604 & buf_data_0[15:8]; // @[lsu_bus_buffer.scala 166:65]
  wire [7:0] _T_609 = ld_byte_hitvecfn_lo_1[1] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_611 = _T_609 & buf_data_1[15:8]; // @[lsu_bus_buffer.scala 166:65]
  wire [7:0] _T_614 = ld_byte_hitvecfn_lo_1[2] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_616 = _T_614 & buf_data_2[15:8]; // @[lsu_bus_buffer.scala 166:65]
  wire [7:0] _T_619 = ld_byte_hitvecfn_lo_1[3] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_621 = _T_619 & buf_data_3[15:8]; // @[lsu_bus_buffer.scala 166:65]
  wire [7:0] _T_622 = _T_606 | _T_611; // @[lsu_bus_buffer.scala 166:97]
  wire [7:0] _T_623 = _T_622 | _T_616; // @[lsu_bus_buffer.scala 166:97]
  wire [7:0] _T_624 = _T_623 | _T_621; // @[lsu_bus_buffer.scala 166:97]
  wire [7:0] _T_627 = ld_byte_hitvecfn_lo_0[0] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_629 = _T_627 & buf_data_0[7:0]; // @[lsu_bus_buffer.scala 167:65]
  wire [7:0] _T_632 = ld_byte_hitvecfn_lo_0[1] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_634 = _T_632 & buf_data_1[7:0]; // @[lsu_bus_buffer.scala 167:65]
  wire [7:0] _T_637 = ld_byte_hitvecfn_lo_0[2] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_639 = _T_637 & buf_data_2[7:0]; // @[lsu_bus_buffer.scala 167:65]
  wire [7:0] _T_642 = ld_byte_hitvecfn_lo_0[3] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_644 = _T_642 & buf_data_3[7:0]; // @[lsu_bus_buffer.scala 167:65]
  wire [7:0] _T_645 = _T_629 | _T_634; // @[lsu_bus_buffer.scala 167:97]
  wire [7:0] _T_646 = _T_645 | _T_639; // @[lsu_bus_buffer.scala 167:97]
  wire [7:0] _T_647 = _T_646 | _T_644; // @[lsu_bus_buffer.scala 167:97]
  wire [31:0] _T_650 = {_T_578,_T_601,_T_624,_T_647}; // @[Cat.scala 29:58]
  reg [31:0] ibuf_data; // @[lib.scala 374:16]
  wire [31:0] _T_651 = ld_fwddata_buf_lo_initial & ibuf_data; // @[lsu_bus_buffer.scala 168:32]
  wire [7:0] _T_655 = ld_byte_hitvecfn_hi_3[0] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_657 = _T_655 & buf_data_0[31:24]; // @[lsu_bus_buffer.scala 170:91]
  wire [7:0] _T_660 = ld_byte_hitvecfn_hi_3[1] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_662 = _T_660 & buf_data_1[31:24]; // @[lsu_bus_buffer.scala 170:91]
  wire [7:0] _T_665 = ld_byte_hitvecfn_hi_3[2] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_667 = _T_665 & buf_data_2[31:24]; // @[lsu_bus_buffer.scala 170:91]
  wire [7:0] _T_670 = ld_byte_hitvecfn_hi_3[3] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_672 = _T_670 & buf_data_3[31:24]; // @[lsu_bus_buffer.scala 170:91]
  wire [7:0] _T_673 = _T_657 | _T_662; // @[lsu_bus_buffer.scala 170:123]
  wire [7:0] _T_674 = _T_673 | _T_667; // @[lsu_bus_buffer.scala 170:123]
  wire [7:0] _T_675 = _T_674 | _T_672; // @[lsu_bus_buffer.scala 170:123]
  wire [7:0] _T_678 = ld_byte_hitvecfn_hi_2[0] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_680 = _T_678 & buf_data_0[23:16]; // @[lsu_bus_buffer.scala 171:65]
  wire [7:0] _T_683 = ld_byte_hitvecfn_hi_2[1] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_685 = _T_683 & buf_data_1[23:16]; // @[lsu_bus_buffer.scala 171:65]
  wire [7:0] _T_688 = ld_byte_hitvecfn_hi_2[2] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_690 = _T_688 & buf_data_2[23:16]; // @[lsu_bus_buffer.scala 171:65]
  wire [7:0] _T_693 = ld_byte_hitvecfn_hi_2[3] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_695 = _T_693 & buf_data_3[23:16]; // @[lsu_bus_buffer.scala 171:65]
  wire [7:0] _T_696 = _T_680 | _T_685; // @[lsu_bus_buffer.scala 171:97]
  wire [7:0] _T_697 = _T_696 | _T_690; // @[lsu_bus_buffer.scala 171:97]
  wire [7:0] _T_698 = _T_697 | _T_695; // @[lsu_bus_buffer.scala 171:97]
  wire [7:0] _T_701 = ld_byte_hitvecfn_hi_1[0] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_703 = _T_701 & buf_data_0[15:8]; // @[lsu_bus_buffer.scala 172:65]
  wire [7:0] _T_706 = ld_byte_hitvecfn_hi_1[1] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_708 = _T_706 & buf_data_1[15:8]; // @[lsu_bus_buffer.scala 172:65]
  wire [7:0] _T_711 = ld_byte_hitvecfn_hi_1[2] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_713 = _T_711 & buf_data_2[15:8]; // @[lsu_bus_buffer.scala 172:65]
  wire [7:0] _T_716 = ld_byte_hitvecfn_hi_1[3] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_718 = _T_716 & buf_data_3[15:8]; // @[lsu_bus_buffer.scala 172:65]
  wire [7:0] _T_719 = _T_703 | _T_708; // @[lsu_bus_buffer.scala 172:97]
  wire [7:0] _T_720 = _T_719 | _T_713; // @[lsu_bus_buffer.scala 172:97]
  wire [7:0] _T_721 = _T_720 | _T_718; // @[lsu_bus_buffer.scala 172:97]
  wire [7:0] _T_724 = ld_byte_hitvecfn_hi_0[0] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_726 = _T_724 & buf_data_0[7:0]; // @[lsu_bus_buffer.scala 173:65]
  wire [7:0] _T_729 = ld_byte_hitvecfn_hi_0[1] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_731 = _T_729 & buf_data_1[7:0]; // @[lsu_bus_buffer.scala 173:65]
  wire [7:0] _T_734 = ld_byte_hitvecfn_hi_0[2] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_736 = _T_734 & buf_data_2[7:0]; // @[lsu_bus_buffer.scala 173:65]
  wire [7:0] _T_739 = ld_byte_hitvecfn_hi_0[3] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_741 = _T_739 & buf_data_3[7:0]; // @[lsu_bus_buffer.scala 173:65]
  wire [7:0] _T_742 = _T_726 | _T_731; // @[lsu_bus_buffer.scala 173:97]
  wire [7:0] _T_743 = _T_742 | _T_736; // @[lsu_bus_buffer.scala 173:97]
  wire [7:0] _T_744 = _T_743 | _T_741; // @[lsu_bus_buffer.scala 173:97]
  wire [31:0] _T_747 = {_T_675,_T_698,_T_721,_T_744}; // @[Cat.scala 29:58]
  wire [31:0] _T_748 = ld_fwddata_buf_hi_initial & ibuf_data; // @[lsu_bus_buffer.scala 174:32]
  wire [3:0] _T_750 = io_lsu_pkt_r_bits_by ? 4'h1 : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_751 = io_lsu_pkt_r_bits_half ? 4'h3 : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_752 = io_lsu_pkt_r_bits_word ? 4'hf : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_753 = _T_750 | _T_751; // @[Mux.scala 27:72]
  wire [3:0] ldst_byteen_r = _T_753 | _T_752; // @[Mux.scala 27:72]
  wire  _T_756 = io_lsu_addr_r[1:0] == 2'h0; // @[lsu_bus_buffer.scala 181:55]
  wire  _T_758 = io_lsu_addr_r[1:0] == 2'h1; // @[lsu_bus_buffer.scala 182:24]
  wire [3:0] _T_760 = {3'h0,ldst_byteen_r[3]}; // @[Cat.scala 29:58]
  wire  _T_762 = io_lsu_addr_r[1:0] == 2'h2; // @[lsu_bus_buffer.scala 183:24]
  wire [3:0] _T_764 = {2'h0,ldst_byteen_r[3:2]}; // @[Cat.scala 29:58]
  wire  _T_766 = io_lsu_addr_r[1:0] == 2'h3; // @[lsu_bus_buffer.scala 184:24]
  wire [3:0] _T_768 = {1'h0,ldst_byteen_r[3:1]}; // @[Cat.scala 29:58]
  wire [3:0] _T_770 = _T_758 ? _T_760 : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_771 = _T_762 ? _T_764 : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_772 = _T_766 ? _T_768 : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_774 = _T_770 | _T_771; // @[Mux.scala 27:72]
  wire [3:0] ldst_byteen_hi_r = _T_774 | _T_772; // @[Mux.scala 27:72]
  wire [3:0] _T_781 = {ldst_byteen_r[2:0],1'h0}; // @[Cat.scala 29:58]
  wire [3:0] _T_785 = {ldst_byteen_r[1:0],2'h0}; // @[Cat.scala 29:58]
  wire [3:0] _T_789 = {ldst_byteen_r[0],3'h0}; // @[Cat.scala 29:58]
  wire [3:0] _T_790 = _T_756 ? ldst_byteen_r : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_791 = _T_758 ? _T_781 : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_792 = _T_762 ? _T_785 : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_793 = _T_766 ? _T_789 : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_794 = _T_790 | _T_791; // @[Mux.scala 27:72]
  wire [3:0] _T_795 = _T_794 | _T_792; // @[Mux.scala 27:72]
  wire [3:0] ldst_byteen_lo_r = _T_795 | _T_793; // @[Mux.scala 27:72]
  wire [31:0] _T_802 = {24'h0,io_store_data_r[31:24]}; // @[Cat.scala 29:58]
  wire [31:0] _T_806 = {16'h0,io_store_data_r[31:16]}; // @[Cat.scala 29:58]
  wire [31:0] _T_810 = {8'h0,io_store_data_r[31:8]}; // @[Cat.scala 29:58]
  wire [31:0] _T_812 = _T_758 ? _T_802 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_813 = _T_762 ? _T_806 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_814 = _T_766 ? _T_810 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_816 = _T_812 | _T_813; // @[Mux.scala 27:72]
  wire [31:0] store_data_hi_r = _T_816 | _T_814; // @[Mux.scala 27:72]
  wire [31:0] _T_823 = {io_store_data_r[23:0],8'h0}; // @[Cat.scala 29:58]
  wire [31:0] _T_827 = {io_store_data_r[15:0],16'h0}; // @[Cat.scala 29:58]
  wire [31:0] _T_831 = {io_store_data_r[7:0],24'h0}; // @[Cat.scala 29:58]
  wire [31:0] _T_832 = _T_756 ? io_store_data_r : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_833 = _T_758 ? _T_823 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_834 = _T_762 ? _T_827 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_835 = _T_766 ? _T_831 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_836 = _T_832 | _T_833; // @[Mux.scala 27:72]
  wire [31:0] _T_837 = _T_836 | _T_834; // @[Mux.scala 27:72]
  wire [31:0] store_data_lo_r = _T_837 | _T_835; // @[Mux.scala 27:72]
  wire  ldst_samedw_r = io_lsu_addr_r[3] == io_end_addr_r[3]; // @[lsu_bus_buffer.scala 201:40]
  wire  _T_844 = ~io_lsu_addr_r[0]; // @[lsu_bus_buffer.scala 203:31]
  wire  _T_845 = io_lsu_pkt_r_bits_word & _T_756; // @[Mux.scala 27:72]
  wire  _T_846 = io_lsu_pkt_r_bits_half & _T_844; // @[Mux.scala 27:72]
  wire  _T_848 = _T_845 | _T_846; // @[Mux.scala 27:72]
  wire  is_aligned_r = _T_848 | io_lsu_pkt_r_bits_by; // @[Mux.scala 27:72]
  wire  _T_850 = io_lsu_pkt_r_bits_load | io_no_word_merge_r; // @[lsu_bus_buffer.scala 205:60]
  wire  _T_851 = io_lsu_busreq_r & _T_850; // @[lsu_bus_buffer.scala 205:34]
  wire  _T_852 = ~ibuf_valid; // @[lsu_bus_buffer.scala 205:84]
  wire  ibuf_byp = _T_851 & _T_852; // @[lsu_bus_buffer.scala 205:82]
  wire  _T_853 = io_lsu_busreq_r & io_lsu_commit_r; // @[lsu_bus_buffer.scala 206:36]
  wire  _T_854 = ~ibuf_byp; // @[lsu_bus_buffer.scala 206:56]
  wire  ibuf_wr_en = _T_853 & _T_854; // @[lsu_bus_buffer.scala 206:54]
  wire  _T_855 = ~ibuf_wr_en; // @[lsu_bus_buffer.scala 208:36]
  reg [2:0] ibuf_timer; // @[lsu_bus_buffer.scala 251:55]
  wire  _T_864 = ibuf_timer == 3'h7; // @[lsu_bus_buffer.scala 214:62]
  wire  _T_865 = ibuf_wr_en | _T_864; // @[lsu_bus_buffer.scala 214:48]
  wire  _T_929 = _T_853 & io_lsu_pkt_r_bits_store; // @[lsu_bus_buffer.scala 233:54]
  wire  _T_930 = _T_929 & ibuf_valid; // @[lsu_bus_buffer.scala 233:80]
  wire  _T_931 = _T_930 & ibuf_write; // @[lsu_bus_buffer.scala 233:93]
  wire  _T_934 = io_lsu_addr_r[31:2] == ibuf_addr[31:2]; // @[lsu_bus_buffer.scala 233:129]
  wire  _T_935 = _T_931 & _T_934; // @[lsu_bus_buffer.scala 233:106]
  wire  _T_936 = ~io_is_sideeffects_r; // @[lsu_bus_buffer.scala 233:152]
  wire  _T_937 = _T_935 & _T_936; // @[lsu_bus_buffer.scala 233:150]
  wire  _T_938 = ~io_tlu_busbuff_dec_tlu_wb_coalescing_disable; // @[lsu_bus_buffer.scala 233:175]
  wire  ibuf_merge_en = _T_937 & _T_938; // @[lsu_bus_buffer.scala 233:173]
  wire  ibuf_merge_in = ~io_ldst_dual_r; // @[lsu_bus_buffer.scala 234:20]
  wire  _T_866 = ibuf_merge_en & ibuf_merge_in; // @[lsu_bus_buffer.scala 214:98]
  wire  _T_867 = ~_T_866; // @[lsu_bus_buffer.scala 214:82]
  wire  _T_868 = _T_865 & _T_867; // @[lsu_bus_buffer.scala 214:80]
  wire  _T_869 = _T_868 | ibuf_byp; // @[lsu_bus_buffer.scala 215:5]
  wire  _T_857 = ~io_lsu_busreq_r; // @[lsu_bus_buffer.scala 209:44]
  wire  _T_858 = io_lsu_busreq_m & _T_857; // @[lsu_bus_buffer.scala 209:42]
  wire  _T_859 = _T_858 & ibuf_valid; // @[lsu_bus_buffer.scala 209:61]
  wire  _T_862 = ibuf_addr[31:2] != io_lsu_addr_m[31:2]; // @[lsu_bus_buffer.scala 209:120]
  wire  _T_863 = io_lsu_pkt_m_bits_load | _T_862; // @[lsu_bus_buffer.scala 209:100]
  wire  ibuf_force_drain = _T_859 & _T_863; // @[lsu_bus_buffer.scala 209:74]
  wire  _T_870 = _T_869 | ibuf_force_drain; // @[lsu_bus_buffer.scala 215:16]
  reg  ibuf_sideeffect; // @[Reg.scala 27:20]
  wire  _T_871 = _T_870 | ibuf_sideeffect; // @[lsu_bus_buffer.scala 215:35]
  wire  _T_872 = ~ibuf_write; // @[lsu_bus_buffer.scala 215:55]
  wire  _T_873 = _T_871 | _T_872; // @[lsu_bus_buffer.scala 215:53]
  wire  _T_874 = _T_873 | io_tlu_busbuff_dec_tlu_wb_coalescing_disable; // @[lsu_bus_buffer.scala 215:67]
  wire  ibuf_drain_vld = ibuf_valid & _T_874; // @[lsu_bus_buffer.scala 214:32]
  wire  _T_856 = ibuf_drain_vld & _T_855; // @[lsu_bus_buffer.scala 208:34]
  wire  ibuf_rst = _T_856 | io_dec_tlu_force_halt; // @[lsu_bus_buffer.scala 208:49]
  reg [1:0] WrPtr1_r; // @[lsu_bus_buffer.scala 615:49]
  reg [1:0] WrPtr0_r; // @[lsu_bus_buffer.scala 614:49]
  reg [1:0] ibuf_tag; // @[Reg.scala 27:20]
  wire [1:0] ibuf_sz_in = {io_lsu_pkt_r_bits_word,io_lsu_pkt_r_bits_half}; // @[Cat.scala 29:58]
  wire [3:0] _T_881 = ibuf_byteen | ldst_byteen_lo_r; // @[lsu_bus_buffer.scala 224:77]
  wire [7:0] _T_889 = ldst_byteen_lo_r[0] ? store_data_lo_r[7:0] : ibuf_data[7:0]; // @[lsu_bus_buffer.scala 229:8]
  wire [7:0] _T_892 = io_ldst_dual_r ? store_data_hi_r[7:0] : store_data_lo_r[7:0]; // @[lsu_bus_buffer.scala 230:8]
  wire [7:0] _T_893 = _T_866 ? _T_889 : _T_892; // @[lsu_bus_buffer.scala 228:46]
  wire [7:0] _T_898 = ldst_byteen_lo_r[1] ? store_data_lo_r[15:8] : ibuf_data[15:8]; // @[lsu_bus_buffer.scala 229:8]
  wire [7:0] _T_901 = io_ldst_dual_r ? store_data_hi_r[15:8] : store_data_lo_r[15:8]; // @[lsu_bus_buffer.scala 230:8]
  wire [7:0] _T_902 = _T_866 ? _T_898 : _T_901; // @[lsu_bus_buffer.scala 228:46]
  wire [7:0] _T_907 = ldst_byteen_lo_r[2] ? store_data_lo_r[23:16] : ibuf_data[23:16]; // @[lsu_bus_buffer.scala 229:8]
  wire [7:0] _T_910 = io_ldst_dual_r ? store_data_hi_r[23:16] : store_data_lo_r[23:16]; // @[lsu_bus_buffer.scala 230:8]
  wire [7:0] _T_911 = _T_866 ? _T_907 : _T_910; // @[lsu_bus_buffer.scala 228:46]
  wire [7:0] _T_916 = ldst_byteen_lo_r[3] ? store_data_lo_r[31:24] : ibuf_data[31:24]; // @[lsu_bus_buffer.scala 229:8]
  wire [7:0] _T_919 = io_ldst_dual_r ? store_data_hi_r[31:24] : store_data_lo_r[31:24]; // @[lsu_bus_buffer.scala 230:8]
  wire [7:0] _T_920 = _T_866 ? _T_916 : _T_919; // @[lsu_bus_buffer.scala 228:46]
  wire [23:0] _T_922 = {_T_920,_T_911,_T_902}; // @[Cat.scala 29:58]
  wire  _T_923 = ibuf_timer < 3'h7; // @[lsu_bus_buffer.scala 231:59]
  wire [2:0] _T_926 = ibuf_timer + 3'h1; // @[lsu_bus_buffer.scala 231:93]
  wire  _T_941 = ~ibuf_merge_in; // @[lsu_bus_buffer.scala 235:65]
  wire  _T_942 = ibuf_merge_en & _T_941; // @[lsu_bus_buffer.scala 235:63]
  wire  _T_945 = ibuf_byteen[0] | ldst_byteen_lo_r[0]; // @[lsu_bus_buffer.scala 235:96]
  wire  _T_947 = _T_942 ? _T_945 : ibuf_byteen[0]; // @[lsu_bus_buffer.scala 235:48]
  wire  _T_952 = ibuf_byteen[1] | ldst_byteen_lo_r[1]; // @[lsu_bus_buffer.scala 235:96]
  wire  _T_954 = _T_942 ? _T_952 : ibuf_byteen[1]; // @[lsu_bus_buffer.scala 235:48]
  wire  _T_959 = ibuf_byteen[2] | ldst_byteen_lo_r[2]; // @[lsu_bus_buffer.scala 235:96]
  wire  _T_961 = _T_942 ? _T_959 : ibuf_byteen[2]; // @[lsu_bus_buffer.scala 235:48]
  wire  _T_966 = ibuf_byteen[3] | ldst_byteen_lo_r[3]; // @[lsu_bus_buffer.scala 235:96]
  wire  _T_968 = _T_942 ? _T_966 : ibuf_byteen[3]; // @[lsu_bus_buffer.scala 235:48]
  wire [3:0] ibuf_byteen_out = {_T_968,_T_961,_T_954,_T_947}; // @[Cat.scala 29:58]
  wire [7:0] _T_978 = _T_942 ? _T_889 : ibuf_data[7:0]; // @[lsu_bus_buffer.scala 236:45]
  wire [7:0] _T_986 = _T_942 ? _T_898 : ibuf_data[15:8]; // @[lsu_bus_buffer.scala 236:45]
  wire [7:0] _T_994 = _T_942 ? _T_907 : ibuf_data[23:16]; // @[lsu_bus_buffer.scala 236:45]
  wire [7:0] _T_1002 = _T_942 ? _T_916 : ibuf_data[31:24]; // @[lsu_bus_buffer.scala 236:45]
  wire [31:0] ibuf_data_out = {_T_1002,_T_994,_T_986,_T_978}; // @[Cat.scala 29:58]
  wire  _T_1005 = ibuf_wr_en | ibuf_valid; // @[lsu_bus_buffer.scala 238:58]
  wire  _T_1006 = ~ibuf_rst; // @[lsu_bus_buffer.scala 238:93]
  reg [1:0] ibuf_dualtag; // @[Reg.scala 27:20]
  reg  ibuf_dual; // @[Reg.scala 27:20]
  reg  ibuf_samedw; // @[Reg.scala 27:20]
  reg  ibuf_nomerge; // @[Reg.scala 27:20]
  reg  ibuf_unsign; // @[Reg.scala 27:20]
  reg [1:0] ibuf_sz; // @[Reg.scala 27:20]
  wire  _T_4446 = buf_write[3] & _T_2621; // @[lsu_bus_buffer.scala 521:64]
  wire  _T_4447 = ~buf_cmd_state_bus_en_3; // @[lsu_bus_buffer.scala 521:91]
  wire  _T_4448 = _T_4446 & _T_4447; // @[lsu_bus_buffer.scala 521:89]
  wire  _T_4441 = buf_write[2] & _T_2616; // @[lsu_bus_buffer.scala 521:64]
  wire  _T_4442 = ~buf_cmd_state_bus_en_2; // @[lsu_bus_buffer.scala 521:91]
  wire  _T_4443 = _T_4441 & _T_4442; // @[lsu_bus_buffer.scala 521:89]
  wire [1:0] _T_4449 = _T_4448 + _T_4443; // @[lsu_bus_buffer.scala 521:142]
  wire  _T_4436 = buf_write[1] & _T_2611; // @[lsu_bus_buffer.scala 521:64]
  wire  _T_4437 = ~buf_cmd_state_bus_en_1; // @[lsu_bus_buffer.scala 521:91]
  wire  _T_4438 = _T_4436 & _T_4437; // @[lsu_bus_buffer.scala 521:89]
  wire [1:0] _GEN_362 = {{1'd0}, _T_4438}; // @[lsu_bus_buffer.scala 521:142]
  wire [2:0] _T_4450 = _T_4449 + _GEN_362; // @[lsu_bus_buffer.scala 521:142]
  wire  _T_4431 = buf_write[0] & _T_2606; // @[lsu_bus_buffer.scala 521:64]
  wire  _T_4432 = ~buf_cmd_state_bus_en_0; // @[lsu_bus_buffer.scala 521:91]
  wire  _T_4433 = _T_4431 & _T_4432; // @[lsu_bus_buffer.scala 521:89]
  wire [2:0] _GEN_363 = {{2'd0}, _T_4433}; // @[lsu_bus_buffer.scala 521:142]
  wire [3:0] buf_numvld_wrcmd_any = _T_4450 + _GEN_363; // @[lsu_bus_buffer.scala 521:142]
  wire  _T_1016 = buf_numvld_wrcmd_any == 4'h1; // @[lsu_bus_buffer.scala 261:43]
  wire  _T_4463 = _T_2621 & _T_4447; // @[lsu_bus_buffer.scala 522:73]
  wire  _T_4460 = _T_2616 & _T_4442; // @[lsu_bus_buffer.scala 522:73]
  wire [1:0] _T_4464 = _T_4463 + _T_4460; // @[lsu_bus_buffer.scala 522:126]
  wire  _T_4457 = _T_2611 & _T_4437; // @[lsu_bus_buffer.scala 522:73]
  wire [1:0] _GEN_364 = {{1'd0}, _T_4457}; // @[lsu_bus_buffer.scala 522:126]
  wire [2:0] _T_4465 = _T_4464 + _GEN_364; // @[lsu_bus_buffer.scala 522:126]
  wire  _T_4454 = _T_2606 & _T_4432; // @[lsu_bus_buffer.scala 522:73]
  wire [2:0] _GEN_365 = {{2'd0}, _T_4454}; // @[lsu_bus_buffer.scala 522:126]
  wire [3:0] buf_numvld_cmd_any = _T_4465 + _GEN_365; // @[lsu_bus_buffer.scala 522:126]
  wire  _T_1017 = buf_numvld_cmd_any == 4'h1; // @[lsu_bus_buffer.scala 261:72]
  wire  _T_1018 = _T_1016 & _T_1017; // @[lsu_bus_buffer.scala 261:51]
  reg [2:0] obuf_wr_timer; // @[lsu_bus_buffer.scala 360:54]
  wire  _T_1019 = obuf_wr_timer != 3'h7; // @[lsu_bus_buffer.scala 261:97]
  wire  _T_1020 = _T_1018 & _T_1019; // @[lsu_bus_buffer.scala 261:80]
  wire  _T_1022 = _T_1020 & _T_938; // @[lsu_bus_buffer.scala 261:114]
  wire  _T_1979 = |buf_age_3; // @[lsu_bus_buffer.scala 377:58]
  wire  _T_1980 = ~_T_1979; // @[lsu_bus_buffer.scala 377:45]
  wire  _T_1982 = _T_1980 & _T_2621; // @[lsu_bus_buffer.scala 377:63]
  wire  _T_1984 = _T_1982 & _T_4447; // @[lsu_bus_buffer.scala 377:88]
  wire  _T_1973 = |buf_age_2; // @[lsu_bus_buffer.scala 377:58]
  wire  _T_1974 = ~_T_1973; // @[lsu_bus_buffer.scala 377:45]
  wire  _T_1976 = _T_1974 & _T_2616; // @[lsu_bus_buffer.scala 377:63]
  wire  _T_1978 = _T_1976 & _T_4442; // @[lsu_bus_buffer.scala 377:88]
  wire  _T_1967 = |buf_age_1; // @[lsu_bus_buffer.scala 377:58]
  wire  _T_1968 = ~_T_1967; // @[lsu_bus_buffer.scala 377:45]
  wire  _T_1970 = _T_1968 & _T_2611; // @[lsu_bus_buffer.scala 377:63]
  wire  _T_1972 = _T_1970 & _T_4437; // @[lsu_bus_buffer.scala 377:88]
  wire  _T_1961 = |buf_age_0; // @[lsu_bus_buffer.scala 377:58]
  wire  _T_1962 = ~_T_1961; // @[lsu_bus_buffer.scala 377:45]
  wire  _T_1964 = _T_1962 & _T_2606; // @[lsu_bus_buffer.scala 377:63]
  wire  _T_1966 = _T_1964 & _T_4432; // @[lsu_bus_buffer.scala 377:88]
  wire [3:0] CmdPtr0Dec = {_T_1984,_T_1978,_T_1972,_T_1966}; // @[Cat.scala 29:58]
  wire [7:0] _T_2054 = {4'h0,_T_1984,_T_1978,_T_1972,_T_1966}; // @[Cat.scala 29:58]
  wire  _T_2057 = _T_2054[4] | _T_2054[5]; // @[lsu_bus_buffer.scala 385:42]
  wire  _T_2059 = _T_2057 | _T_2054[6]; // @[lsu_bus_buffer.scala 385:48]
  wire  _T_2061 = _T_2059 | _T_2054[7]; // @[lsu_bus_buffer.scala 385:54]
  wire  _T_2064 = _T_2054[2] | _T_2054[3]; // @[lsu_bus_buffer.scala 385:67]
  wire  _T_2066 = _T_2064 | _T_2054[6]; // @[lsu_bus_buffer.scala 385:73]
  wire  _T_2068 = _T_2066 | _T_2054[7]; // @[lsu_bus_buffer.scala 385:79]
  wire  _T_2071 = _T_2054[1] | _T_2054[3]; // @[lsu_bus_buffer.scala 385:92]
  wire  _T_2073 = _T_2071 | _T_2054[5]; // @[lsu_bus_buffer.scala 385:98]
  wire  _T_2075 = _T_2073 | _T_2054[7]; // @[lsu_bus_buffer.scala 385:104]
  wire [2:0] _T_2077 = {_T_2061,_T_2068,_T_2075}; // @[Cat.scala 29:58]
  wire [1:0] CmdPtr0 = _T_2077[1:0]; // @[lsu_bus_buffer.scala 390:11]
  wire  _T_1023 = CmdPtr0 == 2'h0; // @[lsu_bus_buffer.scala 262:114]
  wire  _T_1024 = CmdPtr0 == 2'h1; // @[lsu_bus_buffer.scala 262:114]
  wire  _T_1025 = CmdPtr0 == 2'h2; // @[lsu_bus_buffer.scala 262:114]
  wire  _T_1026 = CmdPtr0 == 2'h3; // @[lsu_bus_buffer.scala 262:114]
  reg  buf_nomerge_0; // @[Reg.scala 27:20]
  wire  _T_1027 = _T_1023 & buf_nomerge_0; // @[Mux.scala 27:72]
  reg  buf_nomerge_1; // @[Reg.scala 27:20]
  wire  _T_1028 = _T_1024 & buf_nomerge_1; // @[Mux.scala 27:72]
  reg  buf_nomerge_2; // @[Reg.scala 27:20]
  wire  _T_1029 = _T_1025 & buf_nomerge_2; // @[Mux.scala 27:72]
  reg  buf_nomerge_3; // @[Reg.scala 27:20]
  wire  _T_1030 = _T_1026 & buf_nomerge_3; // @[Mux.scala 27:72]
  wire  _T_1031 = _T_1027 | _T_1028; // @[Mux.scala 27:72]
  wire  _T_1032 = _T_1031 | _T_1029; // @[Mux.scala 27:72]
  wire  _T_1033 = _T_1032 | _T_1030; // @[Mux.scala 27:72]
  wire  _T_1035 = ~_T_1033; // @[lsu_bus_buffer.scala 262:31]
  wire  _T_1036 = _T_1022 & _T_1035; // @[lsu_bus_buffer.scala 262:29]
  reg  _T_4330; // @[Reg.scala 27:20]
  reg  _T_4327; // @[Reg.scala 27:20]
  reg  _T_4324; // @[Reg.scala 27:20]
  reg  _T_4321; // @[Reg.scala 27:20]
  wire [3:0] buf_sideeffect = {_T_4330,_T_4327,_T_4324,_T_4321}; // @[Cat.scala 29:58]
  wire  _T_1045 = _T_1023 & buf_sideeffect[0]; // @[Mux.scala 27:72]
  wire  _T_1046 = _T_1024 & buf_sideeffect[1]; // @[Mux.scala 27:72]
  wire  _T_1047 = _T_1025 & buf_sideeffect[2]; // @[Mux.scala 27:72]
  wire  _T_1048 = _T_1026 & buf_sideeffect[3]; // @[Mux.scala 27:72]
  wire  _T_1049 = _T_1045 | _T_1046; // @[Mux.scala 27:72]
  wire  _T_1050 = _T_1049 | _T_1047; // @[Mux.scala 27:72]
  wire  _T_1051 = _T_1050 | _T_1048; // @[Mux.scala 27:72]
  wire  _T_1053 = ~_T_1051; // @[lsu_bus_buffer.scala 263:5]
  wire  _T_1054 = _T_1036 & _T_1053; // @[lsu_bus_buffer.scala 262:140]
  wire  _T_1065 = _T_858 & _T_852; // @[lsu_bus_buffer.scala 265:58]
  wire  _T_1067 = _T_1065 & _T_1017; // @[lsu_bus_buffer.scala 265:72]
  wire [29:0] _T_1077 = _T_1023 ? buf_addr_0[31:2] : 30'h0; // @[Mux.scala 27:72]
  wire [29:0] _T_1078 = _T_1024 ? buf_addr_1[31:2] : 30'h0; // @[Mux.scala 27:72]
  wire [29:0] _T_1081 = _T_1077 | _T_1078; // @[Mux.scala 27:72]
  wire [29:0] _T_1079 = _T_1025 ? buf_addr_2[31:2] : 30'h0; // @[Mux.scala 27:72]
  wire [29:0] _T_1082 = _T_1081 | _T_1079; // @[Mux.scala 27:72]
  wire [29:0] _T_1080 = _T_1026 ? buf_addr_3[31:2] : 30'h0; // @[Mux.scala 27:72]
  wire [29:0] _T_1083 = _T_1082 | _T_1080; // @[Mux.scala 27:72]
  wire  _T_1085 = io_lsu_addr_m[31:2] != _T_1083; // @[lsu_bus_buffer.scala 265:123]
  wire  obuf_force_wr_en = _T_1067 & _T_1085; // @[lsu_bus_buffer.scala 265:101]
  wire  _T_1055 = ~obuf_force_wr_en; // @[lsu_bus_buffer.scala 263:119]
  wire  obuf_wr_wait = _T_1054 & _T_1055; // @[lsu_bus_buffer.scala 263:117]
  wire  _T_1056 = |buf_numvld_cmd_any; // @[lsu_bus_buffer.scala 264:75]
  wire  _T_1057 = obuf_wr_timer < 3'h7; // @[lsu_bus_buffer.scala 264:95]
  wire  _T_1058 = _T_1056 & _T_1057; // @[lsu_bus_buffer.scala 264:79]
  wire [2:0] _T_1060 = obuf_wr_timer + 3'h1; // @[lsu_bus_buffer.scala 264:123]
  wire  _T_4482 = buf_state_3 == 3'h1; // @[lsu_bus_buffer.scala 523:63]
  wire  _T_4486 = _T_4482 | _T_4463; // @[lsu_bus_buffer.scala 523:74]
  wire  _T_4477 = buf_state_2 == 3'h1; // @[lsu_bus_buffer.scala 523:63]
  wire  _T_4481 = _T_4477 | _T_4460; // @[lsu_bus_buffer.scala 523:74]
  wire [1:0] _T_4487 = _T_4486 + _T_4481; // @[lsu_bus_buffer.scala 523:154]
  wire  _T_4472 = buf_state_1 == 3'h1; // @[lsu_bus_buffer.scala 523:63]
  wire  _T_4476 = _T_4472 | _T_4457; // @[lsu_bus_buffer.scala 523:74]
  wire [1:0] _GEN_366 = {{1'd0}, _T_4476}; // @[lsu_bus_buffer.scala 523:154]
  wire [2:0] _T_4488 = _T_4487 + _GEN_366; // @[lsu_bus_buffer.scala 523:154]
  wire  _T_4467 = buf_state_0 == 3'h1; // @[lsu_bus_buffer.scala 523:63]
  wire  _T_4471 = _T_4467 | _T_4454; // @[lsu_bus_buffer.scala 523:74]
  wire [2:0] _GEN_367 = {{2'd0}, _T_4471}; // @[lsu_bus_buffer.scala 523:154]
  wire [3:0] buf_numvld_pend_any = _T_4488 + _GEN_367; // @[lsu_bus_buffer.scala 523:154]
  wire  _T_1087 = buf_numvld_pend_any == 4'h0; // @[lsu_bus_buffer.scala 267:53]
  wire  _T_1088 = ibuf_byp & _T_1087; // @[lsu_bus_buffer.scala 267:31]
  wire  _T_1089 = ~io_lsu_pkt_r_bits_store; // @[lsu_bus_buffer.scala 267:64]
  wire  _T_1090 = _T_1089 | io_no_dword_merge_r; // @[lsu_bus_buffer.scala 267:89]
  wire  ibuf_buf_byp = _T_1088 & _T_1090; // @[lsu_bus_buffer.scala 267:61]
  wire  _T_1091 = ibuf_buf_byp & io_lsu_commit_r; // @[lsu_bus_buffer.scala 282:32]
  wire  _T_4778 = buf_state_0 == 3'h3; // @[lsu_bus_buffer.scala 551:62]
  wire  _T_4780 = _T_4778 & buf_sideeffect[0]; // @[lsu_bus_buffer.scala 551:73]
  wire  _T_4781 = _T_4780 & io_tlu_busbuff_dec_tlu_sideeffect_posted_disable; // @[lsu_bus_buffer.scala 551:93]
  wire  _T_4782 = buf_state_1 == 3'h3; // @[lsu_bus_buffer.scala 551:62]
  wire  _T_4784 = _T_4782 & buf_sideeffect[1]; // @[lsu_bus_buffer.scala 551:73]
  wire  _T_4785 = _T_4784 & io_tlu_busbuff_dec_tlu_sideeffect_posted_disable; // @[lsu_bus_buffer.scala 551:93]
  wire  _T_4794 = _T_4781 | _T_4785; // @[lsu_bus_buffer.scala 551:153]
  wire  _T_4786 = buf_state_2 == 3'h3; // @[lsu_bus_buffer.scala 551:62]
  wire  _T_4788 = _T_4786 & buf_sideeffect[2]; // @[lsu_bus_buffer.scala 551:73]
  wire  _T_4789 = _T_4788 & io_tlu_busbuff_dec_tlu_sideeffect_posted_disable; // @[lsu_bus_buffer.scala 551:93]
  wire  _T_4795 = _T_4794 | _T_4789; // @[lsu_bus_buffer.scala 551:153]
  wire  _T_4790 = buf_state_3 == 3'h3; // @[lsu_bus_buffer.scala 551:62]
  wire  _T_4792 = _T_4790 & buf_sideeffect[3]; // @[lsu_bus_buffer.scala 551:73]
  wire  _T_4793 = _T_4792 & io_tlu_busbuff_dec_tlu_sideeffect_posted_disable; // @[lsu_bus_buffer.scala 551:93]
  wire  _T_4796 = _T_4795 | _T_4793; // @[lsu_bus_buffer.scala 551:153]
  reg  obuf_sideeffect; // @[Reg.scala 27:20]
  wire  _T_4797 = obuf_valid & obuf_sideeffect; // @[lsu_bus_buffer.scala 551:171]
  wire  _T_4798 = _T_4797 & io_tlu_busbuff_dec_tlu_sideeffect_posted_disable; // @[lsu_bus_buffer.scala 551:189]
  wire  bus_sideeffect_pend = _T_4796 | _T_4798; // @[lsu_bus_buffer.scala 551:157]
  wire  _T_1092 = io_is_sideeffects_r & bus_sideeffect_pend; // @[lsu_bus_buffer.scala 282:74]
  wire  _T_1093 = ~_T_1092; // @[lsu_bus_buffer.scala 282:52]
  wire  _T_1094 = _T_1091 & _T_1093; // @[lsu_bus_buffer.scala 282:50]
  wire [2:0] _T_1099 = _T_1023 ? buf_state_0 : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_1100 = _T_1024 ? buf_state_1 : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_1103 = _T_1099 | _T_1100; // @[Mux.scala 27:72]
  wire [2:0] _T_1101 = _T_1025 ? buf_state_2 : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_1104 = _T_1103 | _T_1101; // @[Mux.scala 27:72]
  wire [2:0] _T_1102 = _T_1026 ? buf_state_3 : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_1105 = _T_1104 | _T_1102; // @[Mux.scala 27:72]
  wire  _T_1107 = _T_1105 == 3'h2; // @[lsu_bus_buffer.scala 283:36]
  wire  found_cmdptr0 = |CmdPtr0Dec; // @[lsu_bus_buffer.scala 382:31]
  wire  _T_1108 = _T_1107 & found_cmdptr0; // @[lsu_bus_buffer.scala 283:47]
  wire [3:0] _T_1111 = {buf_cmd_state_bus_en_3,buf_cmd_state_bus_en_2,buf_cmd_state_bus_en_1,buf_cmd_state_bus_en_0}; // @[Cat.scala 29:58]
  wire  _T_1120 = _T_1023 & _T_1111[0]; // @[Mux.scala 27:72]
  wire  _T_1121 = _T_1024 & _T_1111[1]; // @[Mux.scala 27:72]
  wire  _T_1124 = _T_1120 | _T_1121; // @[Mux.scala 27:72]
  wire  _T_1122 = _T_1025 & _T_1111[2]; // @[Mux.scala 27:72]
  wire  _T_1125 = _T_1124 | _T_1122; // @[Mux.scala 27:72]
  wire  _T_1123 = _T_1026 & _T_1111[3]; // @[Mux.scala 27:72]
  wire  _T_1126 = _T_1125 | _T_1123; // @[Mux.scala 27:72]
  wire  _T_1128 = ~_T_1126; // @[lsu_bus_buffer.scala 284:23]
  wire  _T_1129 = _T_1108 & _T_1128; // @[lsu_bus_buffer.scala 284:21]
  wire  _T_1146 = _T_1051 & bus_sideeffect_pend; // @[lsu_bus_buffer.scala 284:141]
  wire  _T_1147 = ~_T_1146; // @[lsu_bus_buffer.scala 284:105]
  wire  _T_1148 = _T_1129 & _T_1147; // @[lsu_bus_buffer.scala 284:103]
  reg  buf_dual_3; // @[Reg.scala 27:20]
  reg  buf_dual_2; // @[Reg.scala 27:20]
  reg  buf_dual_1; // @[Reg.scala 27:20]
  reg  buf_dual_0; // @[Reg.scala 27:20]
  wire [3:0] _T_1151 = {buf_dual_3,buf_dual_2,buf_dual_1,buf_dual_0}; // @[Cat.scala 29:58]
  wire  _T_1160 = _T_1023 & _T_1151[0]; // @[Mux.scala 27:72]
  wire  _T_1161 = _T_1024 & _T_1151[1]; // @[Mux.scala 27:72]
  wire  _T_1164 = _T_1160 | _T_1161; // @[Mux.scala 27:72]
  wire  _T_1162 = _T_1025 & _T_1151[2]; // @[Mux.scala 27:72]
  wire  _T_1165 = _T_1164 | _T_1162; // @[Mux.scala 27:72]
  wire  _T_1163 = _T_1026 & _T_1151[3]; // @[Mux.scala 27:72]
  wire  _T_1166 = _T_1165 | _T_1163; // @[Mux.scala 27:72]
  reg  buf_samedw_3; // @[Reg.scala 27:20]
  reg  buf_samedw_2; // @[Reg.scala 27:20]
  reg  buf_samedw_1; // @[Reg.scala 27:20]
  reg  buf_samedw_0; // @[Reg.scala 27:20]
  wire [3:0] _T_1170 = {buf_samedw_3,buf_samedw_2,buf_samedw_1,buf_samedw_0}; // @[Cat.scala 29:58]
  wire  _T_1179 = _T_1023 & _T_1170[0]; // @[Mux.scala 27:72]
  wire  _T_1180 = _T_1024 & _T_1170[1]; // @[Mux.scala 27:72]
  wire  _T_1183 = _T_1179 | _T_1180; // @[Mux.scala 27:72]
  wire  _T_1181 = _T_1025 & _T_1170[2]; // @[Mux.scala 27:72]
  wire  _T_1184 = _T_1183 | _T_1181; // @[Mux.scala 27:72]
  wire  _T_1182 = _T_1026 & _T_1170[3]; // @[Mux.scala 27:72]
  wire  _T_1185 = _T_1184 | _T_1182; // @[Mux.scala 27:72]
  wire  _T_1187 = _T_1166 & _T_1185; // @[lsu_bus_buffer.scala 285:77]
  wire  _T_1196 = _T_1023 & buf_write[0]; // @[Mux.scala 27:72]
  wire  _T_1197 = _T_1024 & buf_write[1]; // @[Mux.scala 27:72]
  wire  _T_1200 = _T_1196 | _T_1197; // @[Mux.scala 27:72]
  wire  _T_1198 = _T_1025 & buf_write[2]; // @[Mux.scala 27:72]
  wire  _T_1201 = _T_1200 | _T_1198; // @[Mux.scala 27:72]
  wire  _T_1199 = _T_1026 & buf_write[3]; // @[Mux.scala 27:72]
  wire  _T_1202 = _T_1201 | _T_1199; // @[Mux.scala 27:72]
  wire  _T_1204 = ~_T_1202; // @[lsu_bus_buffer.scala 285:150]
  wire  _T_1205 = _T_1187 & _T_1204; // @[lsu_bus_buffer.scala 285:148]
  wire  _T_1206 = ~_T_1205; // @[lsu_bus_buffer.scala 285:8]
  wire [3:0] _T_2020 = ~CmdPtr0Dec; // @[lsu_bus_buffer.scala 378:62]
  wire [3:0] _T_2021 = buf_age_3 & _T_2020; // @[lsu_bus_buffer.scala 378:59]
  wire  _T_2022 = |_T_2021; // @[lsu_bus_buffer.scala 378:76]
  wire  _T_2023 = ~_T_2022; // @[lsu_bus_buffer.scala 378:45]
  wire  _T_2025 = ~CmdPtr0Dec[3]; // @[lsu_bus_buffer.scala 378:83]
  wire  _T_2026 = _T_2023 & _T_2025; // @[lsu_bus_buffer.scala 378:81]
  wire  _T_2028 = _T_2026 & _T_2621; // @[lsu_bus_buffer.scala 378:98]
  wire  _T_2030 = _T_2028 & _T_4447; // @[lsu_bus_buffer.scala 378:123]
  wire [3:0] _T_2010 = buf_age_2 & _T_2020; // @[lsu_bus_buffer.scala 378:59]
  wire  _T_2011 = |_T_2010; // @[lsu_bus_buffer.scala 378:76]
  wire  _T_2012 = ~_T_2011; // @[lsu_bus_buffer.scala 378:45]
  wire  _T_2014 = ~CmdPtr0Dec[2]; // @[lsu_bus_buffer.scala 378:83]
  wire  _T_2015 = _T_2012 & _T_2014; // @[lsu_bus_buffer.scala 378:81]
  wire  _T_2017 = _T_2015 & _T_2616; // @[lsu_bus_buffer.scala 378:98]
  wire  _T_2019 = _T_2017 & _T_4442; // @[lsu_bus_buffer.scala 378:123]
  wire [3:0] _T_1999 = buf_age_1 & _T_2020; // @[lsu_bus_buffer.scala 378:59]
  wire  _T_2000 = |_T_1999; // @[lsu_bus_buffer.scala 378:76]
  wire  _T_2001 = ~_T_2000; // @[lsu_bus_buffer.scala 378:45]
  wire  _T_2003 = ~CmdPtr0Dec[1]; // @[lsu_bus_buffer.scala 378:83]
  wire  _T_2004 = _T_2001 & _T_2003; // @[lsu_bus_buffer.scala 378:81]
  wire  _T_2006 = _T_2004 & _T_2611; // @[lsu_bus_buffer.scala 378:98]
  wire  _T_2008 = _T_2006 & _T_4437; // @[lsu_bus_buffer.scala 378:123]
  wire [3:0] _T_1988 = buf_age_0 & _T_2020; // @[lsu_bus_buffer.scala 378:59]
  wire  _T_1989 = |_T_1988; // @[lsu_bus_buffer.scala 378:76]
  wire  _T_1990 = ~_T_1989; // @[lsu_bus_buffer.scala 378:45]
  wire  _T_1992 = ~CmdPtr0Dec[0]; // @[lsu_bus_buffer.scala 378:83]
  wire  _T_1993 = _T_1990 & _T_1992; // @[lsu_bus_buffer.scala 378:81]
  wire  _T_1995 = _T_1993 & _T_2606; // @[lsu_bus_buffer.scala 378:98]
  wire  _T_1997 = _T_1995 & _T_4432; // @[lsu_bus_buffer.scala 378:123]
  wire [3:0] CmdPtr1Dec = {_T_2030,_T_2019,_T_2008,_T_1997}; // @[Cat.scala 29:58]
  wire  found_cmdptr1 = |CmdPtr1Dec; // @[lsu_bus_buffer.scala 383:31]
  wire  _T_1207 = _T_1206 | found_cmdptr1; // @[lsu_bus_buffer.scala 285:181]
  wire [3:0] _T_1210 = {buf_nomerge_3,buf_nomerge_2,buf_nomerge_1,buf_nomerge_0}; // @[Cat.scala 29:58]
  wire  _T_1219 = _T_1023 & _T_1210[0]; // @[Mux.scala 27:72]
  wire  _T_1220 = _T_1024 & _T_1210[1]; // @[Mux.scala 27:72]
  wire  _T_1223 = _T_1219 | _T_1220; // @[Mux.scala 27:72]
  wire  _T_1221 = _T_1025 & _T_1210[2]; // @[Mux.scala 27:72]
  wire  _T_1224 = _T_1223 | _T_1221; // @[Mux.scala 27:72]
  wire  _T_1222 = _T_1026 & _T_1210[3]; // @[Mux.scala 27:72]
  wire  _T_1225 = _T_1224 | _T_1222; // @[Mux.scala 27:72]
  wire  _T_1227 = _T_1207 | _T_1225; // @[lsu_bus_buffer.scala 285:197]
  wire  _T_1228 = _T_1227 | obuf_force_wr_en; // @[lsu_bus_buffer.scala 285:269]
  wire  _T_1229 = _T_1148 & _T_1228; // @[lsu_bus_buffer.scala 284:164]
  wire  _T_1230 = _T_1094 | _T_1229; // @[lsu_bus_buffer.scala 282:98]
  reg  obuf_write; // @[Reg.scala 27:20]
  wire  _T_1231 = ~obuf_valid; // @[lsu_bus_buffer.scala 286:48]
  reg  obuf_nosend; // @[Reg.scala 27:20]
  wire  _T_1233 = _T_1231 | obuf_nosend; // @[lsu_bus_buffer.scala 286:60]
  wire  _T_1234 = _T_1230 & _T_1233; // @[lsu_bus_buffer.scala 286:29]
  wire  _T_1235 = ~obuf_wr_wait; // @[lsu_bus_buffer.scala 286:77]
  wire  _T_1236 = _T_1234 & _T_1235; // @[lsu_bus_buffer.scala 286:75]
  reg [31:0] obuf_addr; // @[lib.scala 374:16]
  wire  _T_4804 = obuf_addr[31:3] == buf_addr_0[31:3]; // @[lsu_bus_buffer.scala 553:56]
  wire  _T_4805 = obuf_valid & _T_4804; // @[lsu_bus_buffer.scala 553:38]
  wire  _T_4807 = obuf_tag1 == 2'h0; // @[lsu_bus_buffer.scala 553:126]
  wire  _T_4808 = obuf_merge & _T_4807; // @[lsu_bus_buffer.scala 553:114]
  wire  _T_4809 = _T_3562 | _T_4808; // @[lsu_bus_buffer.scala 553:100]
  wire  _T_4810 = ~_T_4809; // @[lsu_bus_buffer.scala 553:80]
  wire  _T_4811 = _T_4805 & _T_4810; // @[lsu_bus_buffer.scala 553:78]
  wire  _T_4848 = _T_4778 & _T_4811; // @[Mux.scala 27:72]
  wire  _T_4816 = obuf_addr[31:3] == buf_addr_1[31:3]; // @[lsu_bus_buffer.scala 553:56]
  wire  _T_4817 = obuf_valid & _T_4816; // @[lsu_bus_buffer.scala 553:38]
  wire  _T_4819 = obuf_tag1 == 2'h1; // @[lsu_bus_buffer.scala 553:126]
  wire  _T_4820 = obuf_merge & _T_4819; // @[lsu_bus_buffer.scala 553:114]
  wire  _T_4821 = _T_3755 | _T_4820; // @[lsu_bus_buffer.scala 553:100]
  wire  _T_4822 = ~_T_4821; // @[lsu_bus_buffer.scala 553:80]
  wire  _T_4823 = _T_4817 & _T_4822; // @[lsu_bus_buffer.scala 553:78]
  wire  _T_4849 = _T_4782 & _T_4823; // @[Mux.scala 27:72]
  wire  _T_4852 = _T_4848 | _T_4849; // @[Mux.scala 27:72]
  wire  _T_4828 = obuf_addr[31:3] == buf_addr_2[31:3]; // @[lsu_bus_buffer.scala 553:56]
  wire  _T_4829 = obuf_valid & _T_4828; // @[lsu_bus_buffer.scala 553:38]
  wire  _T_4831 = obuf_tag1 == 2'h2; // @[lsu_bus_buffer.scala 553:126]
  wire  _T_4832 = obuf_merge & _T_4831; // @[lsu_bus_buffer.scala 553:114]
  wire  _T_4833 = _T_3948 | _T_4832; // @[lsu_bus_buffer.scala 553:100]
  wire  _T_4834 = ~_T_4833; // @[lsu_bus_buffer.scala 553:80]
  wire  _T_4835 = _T_4829 & _T_4834; // @[lsu_bus_buffer.scala 553:78]
  wire  _T_4850 = _T_4786 & _T_4835; // @[Mux.scala 27:72]
  wire  _T_4853 = _T_4852 | _T_4850; // @[Mux.scala 27:72]
  wire  _T_4840 = obuf_addr[31:3] == buf_addr_3[31:3]; // @[lsu_bus_buffer.scala 553:56]
  wire  _T_4841 = obuf_valid & _T_4840; // @[lsu_bus_buffer.scala 553:38]
  wire  _T_4843 = obuf_tag1 == 2'h3; // @[lsu_bus_buffer.scala 553:126]
  wire  _T_4844 = obuf_merge & _T_4843; // @[lsu_bus_buffer.scala 553:114]
  wire  _T_4845 = _T_4141 | _T_4844; // @[lsu_bus_buffer.scala 553:100]
  wire  _T_4846 = ~_T_4845; // @[lsu_bus_buffer.scala 553:80]
  wire  _T_4847 = _T_4841 & _T_4846; // @[lsu_bus_buffer.scala 553:78]
  wire  _T_4851 = _T_4790 & _T_4847; // @[Mux.scala 27:72]
  wire  bus_addr_match_pending = _T_4853 | _T_4851; // @[Mux.scala 27:72]
  wire  _T_1239 = ~bus_addr_match_pending; // @[lsu_bus_buffer.scala 286:118]
  wire  _T_1240 = _T_1236 & _T_1239; // @[lsu_bus_buffer.scala 286:116]
  wire  obuf_wr_en = _T_1240 & io_lsu_bus_clk_en; // @[lsu_bus_buffer.scala 286:142]
  wire  _T_1242 = obuf_valid & obuf_nosend; // @[lsu_bus_buffer.scala 288:47]
  wire  _T_1244 = ~obuf_wr_en; // @[lsu_bus_buffer.scala 288:65]
  wire  _T_1245 = _T_1242 & _T_1244; // @[lsu_bus_buffer.scala 288:63]
  wire  _T_1246 = _T_1245 & io_lsu_bus_clk_en; // @[lsu_bus_buffer.scala 288:77]
  wire  obuf_rst = _T_1246 | io_dec_tlu_force_halt; // @[lsu_bus_buffer.scala 288:98]
  wire  obuf_write_in = ibuf_buf_byp ? io_lsu_pkt_r_bits_store : _T_1202; // @[lsu_bus_buffer.scala 289:26]
  wire [31:0] _T_1283 = _T_1023 ? buf_addr_0 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1284 = _T_1024 ? buf_addr_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1285 = _T_1025 ? buf_addr_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1286 = _T_1026 ? buf_addr_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1287 = _T_1283 | _T_1284; // @[Mux.scala 27:72]
  wire [31:0] _T_1288 = _T_1287 | _T_1285; // @[Mux.scala 27:72]
  wire [31:0] _T_1289 = _T_1288 | _T_1286; // @[Mux.scala 27:72]
  wire [31:0] obuf_addr_in = ibuf_buf_byp ? io_lsu_addr_r : _T_1289; // @[lsu_bus_buffer.scala 291:25]
  reg [1:0] buf_sz_0; // @[Reg.scala 27:20]
  wire [1:0] _T_1296 = _T_1023 ? buf_sz_0 : 2'h0; // @[Mux.scala 27:72]
  reg [1:0] buf_sz_1; // @[Reg.scala 27:20]
  wire [1:0] _T_1297 = _T_1024 ? buf_sz_1 : 2'h0; // @[Mux.scala 27:72]
  reg [1:0] buf_sz_2; // @[Reg.scala 27:20]
  wire [1:0] _T_1298 = _T_1025 ? buf_sz_2 : 2'h0; // @[Mux.scala 27:72]
  reg [1:0] buf_sz_3; // @[Reg.scala 27:20]
  wire [1:0] _T_1299 = _T_1026 ? buf_sz_3 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_1300 = _T_1296 | _T_1297; // @[Mux.scala 27:72]
  wire [1:0] _T_1301 = _T_1300 | _T_1298; // @[Mux.scala 27:72]
  wire [1:0] _T_1302 = _T_1301 | _T_1299; // @[Mux.scala 27:72]
  wire [1:0] obuf_sz_in = ibuf_buf_byp ? ibuf_sz_in : _T_1302; // @[lsu_bus_buffer.scala 294:23]
  wire [7:0] _T_2079 = {4'h0,_T_2030,_T_2019,_T_2008,_T_1997}; // @[Cat.scala 29:58]
  wire  _T_2082 = _T_2079[4] | _T_2079[5]; // @[lsu_bus_buffer.scala 385:42]
  wire  _T_2084 = _T_2082 | _T_2079[6]; // @[lsu_bus_buffer.scala 385:48]
  wire  _T_2086 = _T_2084 | _T_2079[7]; // @[lsu_bus_buffer.scala 385:54]
  wire  _T_2089 = _T_2079[2] | _T_2079[3]; // @[lsu_bus_buffer.scala 385:67]
  wire  _T_2091 = _T_2089 | _T_2079[6]; // @[lsu_bus_buffer.scala 385:73]
  wire  _T_2093 = _T_2091 | _T_2079[7]; // @[lsu_bus_buffer.scala 385:79]
  wire  _T_2096 = _T_2079[1] | _T_2079[3]; // @[lsu_bus_buffer.scala 385:92]
  wire  _T_2098 = _T_2096 | _T_2079[5]; // @[lsu_bus_buffer.scala 385:98]
  wire  _T_2100 = _T_2098 | _T_2079[7]; // @[lsu_bus_buffer.scala 385:104]
  wire [2:0] _T_2102 = {_T_2086,_T_2093,_T_2100}; // @[Cat.scala 29:58]
  wire [1:0] CmdPtr1 = _T_2102[1:0]; // @[lsu_bus_buffer.scala 392:11]
  wire  _T_1311 = obuf_sz_in == 2'h0; // @[lsu_bus_buffer.scala 307:72]
  wire  _T_1314 = ~obuf_addr_in[0]; // @[lsu_bus_buffer.scala 307:98]
  wire  _T_1315 = obuf_sz_in[0] & _T_1314; // @[lsu_bus_buffer.scala 307:96]
  wire  _T_1316 = _T_1311 | _T_1315; // @[lsu_bus_buffer.scala 307:79]
  wire  _T_1319 = |obuf_addr_in[1:0]; // @[lsu_bus_buffer.scala 307:153]
  wire  _T_1320 = ~_T_1319; // @[lsu_bus_buffer.scala 307:134]
  wire  _T_1321 = obuf_sz_in[1] & _T_1320; // @[lsu_bus_buffer.scala 307:132]
  wire  _T_1322 = _T_1316 | _T_1321; // @[lsu_bus_buffer.scala 307:116]
  wire  obuf_aligned_in = ibuf_buf_byp ? is_aligned_r : _T_1322; // @[lsu_bus_buffer.scala 307:28]
  wire  _T_1339 = obuf_addr_in[31:3] == obuf_addr[31:3]; // @[lsu_bus_buffer.scala 321:40]
  wire  _T_1340 = _T_1339 & obuf_aligned_in; // @[lsu_bus_buffer.scala 321:60]
  wire  _T_1341 = ~obuf_sideeffect; // @[lsu_bus_buffer.scala 321:80]
  wire  _T_1342 = _T_1340 & _T_1341; // @[lsu_bus_buffer.scala 321:78]
  wire  _T_1343 = ~obuf_write; // @[lsu_bus_buffer.scala 321:99]
  wire  _T_1344 = _T_1342 & _T_1343; // @[lsu_bus_buffer.scala 321:97]
  wire  _T_1345 = ~obuf_write_in; // @[lsu_bus_buffer.scala 321:113]
  wire  _T_1346 = _T_1344 & _T_1345; // @[lsu_bus_buffer.scala 321:111]
  wire  _T_1347 = ~io_tlu_busbuff_dec_tlu_external_ldfwd_disable; // @[lsu_bus_buffer.scala 321:130]
  wire  _T_1348 = _T_1346 & _T_1347; // @[lsu_bus_buffer.scala 321:128]
  wire  _T_1349 = ~obuf_nosend; // @[lsu_bus_buffer.scala 322:20]
  wire  _T_1350 = obuf_valid & _T_1349; // @[lsu_bus_buffer.scala 322:18]
  wire  obuf_nosend_in = _T_1348 & _T_1350; // @[lsu_bus_buffer.scala 321:177]
  wire  _T_1333 = ~io_dec_tlu_force_halt; // @[lsu_bus_buffer.scala 316:37]
  wire [7:0] _T_1358 = {ldst_byteen_lo_r,4'h0}; // @[Cat.scala 29:58]
  wire [7:0] _T_1359 = {4'h0,ldst_byteen_lo_r}; // @[Cat.scala 29:58]
  wire [7:0] _T_1360 = io_lsu_addr_r[2] ? _T_1358 : _T_1359; // @[lsu_bus_buffer.scala 323:46]
  wire [3:0] _T_1379 = _T_1023 ? buf_byteen_0 : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_1380 = _T_1024 ? buf_byteen_1 : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_1381 = _T_1025 ? buf_byteen_2 : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_1382 = _T_1026 ? buf_byteen_3 : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_1383 = _T_1379 | _T_1380; // @[Mux.scala 27:72]
  wire [3:0] _T_1384 = _T_1383 | _T_1381; // @[Mux.scala 27:72]
  wire [3:0] _T_1385 = _T_1384 | _T_1382; // @[Mux.scala 27:72]
  wire [7:0] _T_1387 = {_T_1385,4'h0}; // @[Cat.scala 29:58]
  wire [7:0] _T_1400 = {4'h0,_T_1385}; // @[Cat.scala 29:58]
  wire [7:0] _T_1401 = _T_1289[2] ? _T_1387 : _T_1400; // @[lsu_bus_buffer.scala 324:8]
  wire [7:0] obuf_byteen0_in = ibuf_buf_byp ? _T_1360 : _T_1401; // @[lsu_bus_buffer.scala 323:28]
  wire [7:0] _T_1403 = {ldst_byteen_hi_r,4'h0}; // @[Cat.scala 29:58]
  wire [7:0] _T_1404 = {4'h0,ldst_byteen_hi_r}; // @[Cat.scala 29:58]
  wire [7:0] _T_1405 = io_end_addr_r[2] ? _T_1403 : _T_1404; // @[lsu_bus_buffer.scala 325:46]
  wire  _T_1406 = CmdPtr1 == 2'h0; // @[lsu_bus_buffer.scala 57:123]
  wire  _T_1407 = CmdPtr1 == 2'h1; // @[lsu_bus_buffer.scala 57:123]
  wire  _T_1408 = CmdPtr1 == 2'h2; // @[lsu_bus_buffer.scala 57:123]
  wire  _T_1409 = CmdPtr1 == 2'h3; // @[lsu_bus_buffer.scala 57:123]
  wire [31:0] _T_1410 = _T_1406 ? buf_addr_0 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1411 = _T_1407 ? buf_addr_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1412 = _T_1408 ? buf_addr_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1413 = _T_1409 ? buf_addr_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1414 = _T_1410 | _T_1411; // @[Mux.scala 27:72]
  wire [31:0] _T_1415 = _T_1414 | _T_1412; // @[Mux.scala 27:72]
  wire [31:0] _T_1416 = _T_1415 | _T_1413; // @[Mux.scala 27:72]
  wire [3:0] _T_1424 = _T_1406 ? buf_byteen_0 : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_1425 = _T_1407 ? buf_byteen_1 : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_1426 = _T_1408 ? buf_byteen_2 : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_1427 = _T_1409 ? buf_byteen_3 : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_1428 = _T_1424 | _T_1425; // @[Mux.scala 27:72]
  wire [3:0] _T_1429 = _T_1428 | _T_1426; // @[Mux.scala 27:72]
  wire [3:0] _T_1430 = _T_1429 | _T_1427; // @[Mux.scala 27:72]
  wire [7:0] _T_1432 = {_T_1430,4'h0}; // @[Cat.scala 29:58]
  wire [7:0] _T_1445 = {4'h0,_T_1430}; // @[Cat.scala 29:58]
  wire [7:0] _T_1446 = _T_1416[2] ? _T_1432 : _T_1445; // @[lsu_bus_buffer.scala 326:8]
  wire [7:0] obuf_byteen1_in = ibuf_buf_byp ? _T_1405 : _T_1446; // @[lsu_bus_buffer.scala 325:28]
  wire  _T_1621 = CmdPtr0 != CmdPtr1; // @[lsu_bus_buffer.scala 337:30]
  wire  _T_1622 = _T_1621 & found_cmdptr0; // @[lsu_bus_buffer.scala 337:43]
  wire  _T_1623 = _T_1622 & found_cmdptr1; // @[lsu_bus_buffer.scala 337:59]
  wire  _T_1637 = _T_1623 & _T_1107; // @[lsu_bus_buffer.scala 337:75]
  wire [2:0] _T_1642 = _T_1406 ? buf_state_0 : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_1643 = _T_1407 ? buf_state_1 : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_1646 = _T_1642 | _T_1643; // @[Mux.scala 27:72]
  wire [2:0] _T_1644 = _T_1408 ? buf_state_2 : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_1647 = _T_1646 | _T_1644; // @[Mux.scala 27:72]
  wire [2:0] _T_1645 = _T_1409 ? buf_state_3 : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_1648 = _T_1647 | _T_1645; // @[Mux.scala 27:72]
  wire  _T_1650 = _T_1648 == 3'h2; // @[lsu_bus_buffer.scala 337:150]
  wire  _T_1651 = _T_1637 & _T_1650; // @[lsu_bus_buffer.scala 337:118]
  wire  _T_1672 = _T_1651 & _T_1128; // @[lsu_bus_buffer.scala 337:161]
  wire  _T_1690 = _T_1672 & _T_1053; // @[lsu_bus_buffer.scala 338:85]
  wire  _T_1792 = _T_1204 & _T_1166; // @[lsu_bus_buffer.scala 341:38]
  reg  buf_dualhi_3; // @[Reg.scala 27:20]
  reg  buf_dualhi_2; // @[Reg.scala 27:20]
  reg  buf_dualhi_1; // @[Reg.scala 27:20]
  reg  buf_dualhi_0; // @[Reg.scala 27:20]
  wire [3:0] _T_1795 = {buf_dualhi_3,buf_dualhi_2,buf_dualhi_1,buf_dualhi_0}; // @[Cat.scala 29:58]
  wire  _T_1804 = _T_1023 & _T_1795[0]; // @[Mux.scala 27:72]
  wire  _T_1805 = _T_1024 & _T_1795[1]; // @[Mux.scala 27:72]
  wire  _T_1808 = _T_1804 | _T_1805; // @[Mux.scala 27:72]
  wire  _T_1806 = _T_1025 & _T_1795[2]; // @[Mux.scala 27:72]
  wire  _T_1809 = _T_1808 | _T_1806; // @[Mux.scala 27:72]
  wire  _T_1807 = _T_1026 & _T_1795[3]; // @[Mux.scala 27:72]
  wire  _T_1810 = _T_1809 | _T_1807; // @[Mux.scala 27:72]
  wire  _T_1812 = ~_T_1810; // @[lsu_bus_buffer.scala 341:109]
  wire  _T_1813 = _T_1792 & _T_1812; // @[lsu_bus_buffer.scala 341:107]
  wire  _T_1833 = _T_1813 & _T_1185; // @[lsu_bus_buffer.scala 341:179]
  wire  _T_1835 = _T_1690 & _T_1833; // @[lsu_bus_buffer.scala 338:122]
  wire  _T_1836 = ibuf_buf_byp & ldst_samedw_r; // @[lsu_bus_buffer.scala 342:19]
  wire  _T_1837 = _T_1836 & io_ldst_dual_r; // @[lsu_bus_buffer.scala 342:35]
  wire  obuf_merge_en = _T_1835 | _T_1837; // @[lsu_bus_buffer.scala 341:253]
  wire  _T_1539 = obuf_merge_en & obuf_byteen1_in[0]; // @[lsu_bus_buffer.scala 332:80]
  wire  _T_1540 = obuf_byteen0_in[0] | _T_1539; // @[lsu_bus_buffer.scala 332:63]
  wire  _T_1543 = obuf_merge_en & obuf_byteen1_in[1]; // @[lsu_bus_buffer.scala 332:80]
  wire  _T_1544 = obuf_byteen0_in[1] | _T_1543; // @[lsu_bus_buffer.scala 332:63]
  wire  _T_1547 = obuf_merge_en & obuf_byteen1_in[2]; // @[lsu_bus_buffer.scala 332:80]
  wire  _T_1548 = obuf_byteen0_in[2] | _T_1547; // @[lsu_bus_buffer.scala 332:63]
  wire  _T_1551 = obuf_merge_en & obuf_byteen1_in[3]; // @[lsu_bus_buffer.scala 332:80]
  wire  _T_1552 = obuf_byteen0_in[3] | _T_1551; // @[lsu_bus_buffer.scala 332:63]
  wire  _T_1555 = obuf_merge_en & obuf_byteen1_in[4]; // @[lsu_bus_buffer.scala 332:80]
  wire  _T_1556 = obuf_byteen0_in[4] | _T_1555; // @[lsu_bus_buffer.scala 332:63]
  wire  _T_1559 = obuf_merge_en & obuf_byteen1_in[5]; // @[lsu_bus_buffer.scala 332:80]
  wire  _T_1560 = obuf_byteen0_in[5] | _T_1559; // @[lsu_bus_buffer.scala 332:63]
  wire  _T_1563 = obuf_merge_en & obuf_byteen1_in[6]; // @[lsu_bus_buffer.scala 332:80]
  wire  _T_1564 = obuf_byteen0_in[6] | _T_1563; // @[lsu_bus_buffer.scala 332:63]
  wire  _T_1567 = obuf_merge_en & obuf_byteen1_in[7]; // @[lsu_bus_buffer.scala 332:80]
  wire  _T_1568 = obuf_byteen0_in[7] | _T_1567; // @[lsu_bus_buffer.scala 332:63]
  wire [7:0] obuf_byteen_in = {_T_1568,_T_1564,_T_1560,_T_1556,_T_1552,_T_1548,_T_1544,_T_1540}; // @[Cat.scala 29:58]
  wire  _T_1839 = obuf_wr_en | obuf_valid; // @[lsu_bus_buffer.scala 345:58]
  wire  _T_1840 = ~obuf_rst; // @[lsu_bus_buffer.scala 345:93]
  reg [1:0] obuf_sz; // @[Reg.scala 27:20]
  reg [7:0] obuf_byteen; // @[Reg.scala 27:20]
  wire  _T_1853 = buf_state_0 == 3'h0; // @[lsu_bus_buffer.scala 363:65]
  wire  _T_1854 = ibuf_tag == 2'h0; // @[lsu_bus_buffer.scala 364:30]
  wire  _T_1855 = ibuf_valid & _T_1854; // @[lsu_bus_buffer.scala 364:19]
  wire  _T_1856 = WrPtr0_r == 2'h0; // @[lsu_bus_buffer.scala 365:18]
  wire  _T_1857 = WrPtr1_r == 2'h0; // @[lsu_bus_buffer.scala 365:57]
  wire  _T_1858 = io_ldst_dual_r & _T_1857; // @[lsu_bus_buffer.scala 365:45]
  wire  _T_1859 = _T_1856 | _T_1858; // @[lsu_bus_buffer.scala 365:27]
  wire  _T_1860 = io_lsu_busreq_r & _T_1859; // @[lsu_bus_buffer.scala 364:58]
  wire  _T_1861 = _T_1855 | _T_1860; // @[lsu_bus_buffer.scala 364:39]
  wire  _T_1862 = ~_T_1861; // @[lsu_bus_buffer.scala 364:5]
  wire  _T_1863 = _T_1853 & _T_1862; // @[lsu_bus_buffer.scala 363:76]
  wire  _T_1864 = buf_state_1 == 3'h0; // @[lsu_bus_buffer.scala 363:65]
  wire  _T_1865 = ibuf_tag == 2'h1; // @[lsu_bus_buffer.scala 364:30]
  wire  _T_1866 = ibuf_valid & _T_1865; // @[lsu_bus_buffer.scala 364:19]
  wire  _T_1867 = WrPtr0_r == 2'h1; // @[lsu_bus_buffer.scala 365:18]
  wire  _T_1868 = WrPtr1_r == 2'h1; // @[lsu_bus_buffer.scala 365:57]
  wire  _T_1869 = io_ldst_dual_r & _T_1868; // @[lsu_bus_buffer.scala 365:45]
  wire  _T_1870 = _T_1867 | _T_1869; // @[lsu_bus_buffer.scala 365:27]
  wire  _T_1871 = io_lsu_busreq_r & _T_1870; // @[lsu_bus_buffer.scala 364:58]
  wire  _T_1872 = _T_1866 | _T_1871; // @[lsu_bus_buffer.scala 364:39]
  wire  _T_1873 = ~_T_1872; // @[lsu_bus_buffer.scala 364:5]
  wire  _T_1874 = _T_1864 & _T_1873; // @[lsu_bus_buffer.scala 363:76]
  wire  _T_1875 = buf_state_2 == 3'h0; // @[lsu_bus_buffer.scala 363:65]
  wire  _T_1876 = ibuf_tag == 2'h2; // @[lsu_bus_buffer.scala 364:30]
  wire  _T_1877 = ibuf_valid & _T_1876; // @[lsu_bus_buffer.scala 364:19]
  wire  _T_1878 = WrPtr0_r == 2'h2; // @[lsu_bus_buffer.scala 365:18]
  wire  _T_1879 = WrPtr1_r == 2'h2; // @[lsu_bus_buffer.scala 365:57]
  wire  _T_1880 = io_ldst_dual_r & _T_1879; // @[lsu_bus_buffer.scala 365:45]
  wire  _T_1881 = _T_1878 | _T_1880; // @[lsu_bus_buffer.scala 365:27]
  wire  _T_1882 = io_lsu_busreq_r & _T_1881; // @[lsu_bus_buffer.scala 364:58]
  wire  _T_1883 = _T_1877 | _T_1882; // @[lsu_bus_buffer.scala 364:39]
  wire  _T_1884 = ~_T_1883; // @[lsu_bus_buffer.scala 364:5]
  wire  _T_1885 = _T_1875 & _T_1884; // @[lsu_bus_buffer.scala 363:76]
  wire  _T_1886 = buf_state_3 == 3'h0; // @[lsu_bus_buffer.scala 363:65]
  wire  _T_1887 = ibuf_tag == 2'h3; // @[lsu_bus_buffer.scala 364:30]
  wire  _T_1889 = WrPtr0_r == 2'h3; // @[lsu_bus_buffer.scala 365:18]
  wire  _T_1890 = WrPtr1_r == 2'h3; // @[lsu_bus_buffer.scala 365:57]
  wire [1:0] _T_1898 = _T_1885 ? 2'h2 : 2'h3; // @[Mux.scala 98:16]
  wire [1:0] _T_1899 = _T_1874 ? 2'h1 : _T_1898; // @[Mux.scala 98:16]
  wire [1:0] WrPtr0_m = _T_1863 ? 2'h0 : _T_1899; // @[Mux.scala 98:16]
  wire  _T_1904 = WrPtr0_m == 2'h0; // @[lsu_bus_buffer.scala 370:33]
  wire  _T_1905 = io_lsu_busreq_m & _T_1904; // @[lsu_bus_buffer.scala 370:22]
  wire  _T_1906 = _T_1855 | _T_1905; // @[lsu_bus_buffer.scala 369:112]
  wire  _T_1912 = _T_1906 | _T_1860; // @[lsu_bus_buffer.scala 370:42]
  wire  _T_1913 = ~_T_1912; // @[lsu_bus_buffer.scala 369:78]
  wire  _T_1914 = _T_1853 & _T_1913; // @[lsu_bus_buffer.scala 369:76]
  wire  _T_1918 = WrPtr0_m == 2'h1; // @[lsu_bus_buffer.scala 370:33]
  wire  _T_1919 = io_lsu_busreq_m & _T_1918; // @[lsu_bus_buffer.scala 370:22]
  wire  _T_1920 = _T_1866 | _T_1919; // @[lsu_bus_buffer.scala 369:112]
  wire  _T_1926 = _T_1920 | _T_1871; // @[lsu_bus_buffer.scala 370:42]
  wire  _T_1927 = ~_T_1926; // @[lsu_bus_buffer.scala 369:78]
  wire  _T_1928 = _T_1864 & _T_1927; // @[lsu_bus_buffer.scala 369:76]
  wire  _T_1932 = WrPtr0_m == 2'h2; // @[lsu_bus_buffer.scala 370:33]
  wire  _T_1933 = io_lsu_busreq_m & _T_1932; // @[lsu_bus_buffer.scala 370:22]
  wire  _T_1934 = _T_1877 | _T_1933; // @[lsu_bus_buffer.scala 369:112]
  wire  _T_1940 = _T_1934 | _T_1882; // @[lsu_bus_buffer.scala 370:42]
  wire  _T_1941 = ~_T_1940; // @[lsu_bus_buffer.scala 369:78]
  wire  _T_1942 = _T_1875 & _T_1941; // @[lsu_bus_buffer.scala 369:76]
  reg [3:0] buf_rspageQ_0; // @[lsu_bus_buffer.scala 500:63]
  wire  _T_2746 = buf_state_3 == 3'h5; // @[lsu_bus_buffer.scala 413:102]
  wire  _T_2747 = buf_rspageQ_0[3] & _T_2746; // @[lsu_bus_buffer.scala 413:87]
  wire  _T_2743 = buf_state_2 == 3'h5; // @[lsu_bus_buffer.scala 413:102]
  wire  _T_2744 = buf_rspageQ_0[2] & _T_2743; // @[lsu_bus_buffer.scala 413:87]
  wire  _T_2740 = buf_state_1 == 3'h5; // @[lsu_bus_buffer.scala 413:102]
  wire  _T_2741 = buf_rspageQ_0[1] & _T_2740; // @[lsu_bus_buffer.scala 413:87]
  wire  _T_2737 = buf_state_0 == 3'h5; // @[lsu_bus_buffer.scala 413:102]
  wire  _T_2738 = buf_rspageQ_0[0] & _T_2737; // @[lsu_bus_buffer.scala 413:87]
  wire [3:0] buf_rsp_pickage_0 = {_T_2747,_T_2744,_T_2741,_T_2738}; // @[Cat.scala 29:58]
  wire  _T_2033 = |buf_rsp_pickage_0; // @[lsu_bus_buffer.scala 381:65]
  wire  _T_2034 = ~_T_2033; // @[lsu_bus_buffer.scala 381:44]
  wire  _T_2036 = _T_2034 & _T_2737; // @[lsu_bus_buffer.scala 381:70]
  reg [3:0] buf_rspageQ_1; // @[lsu_bus_buffer.scala 500:63]
  wire  _T_2762 = buf_rspageQ_1[3] & _T_2746; // @[lsu_bus_buffer.scala 413:87]
  wire  _T_2759 = buf_rspageQ_1[2] & _T_2743; // @[lsu_bus_buffer.scala 413:87]
  wire  _T_2756 = buf_rspageQ_1[1] & _T_2740; // @[lsu_bus_buffer.scala 413:87]
  wire  _T_2753 = buf_rspageQ_1[0] & _T_2737; // @[lsu_bus_buffer.scala 413:87]
  wire [3:0] buf_rsp_pickage_1 = {_T_2762,_T_2759,_T_2756,_T_2753}; // @[Cat.scala 29:58]
  wire  _T_2037 = |buf_rsp_pickage_1; // @[lsu_bus_buffer.scala 381:65]
  wire  _T_2038 = ~_T_2037; // @[lsu_bus_buffer.scala 381:44]
  wire  _T_2040 = _T_2038 & _T_2740; // @[lsu_bus_buffer.scala 381:70]
  reg [3:0] buf_rspageQ_2; // @[lsu_bus_buffer.scala 500:63]
  wire  _T_2777 = buf_rspageQ_2[3] & _T_2746; // @[lsu_bus_buffer.scala 413:87]
  wire  _T_2774 = buf_rspageQ_2[2] & _T_2743; // @[lsu_bus_buffer.scala 413:87]
  wire  _T_2771 = buf_rspageQ_2[1] & _T_2740; // @[lsu_bus_buffer.scala 413:87]
  wire  _T_2768 = buf_rspageQ_2[0] & _T_2737; // @[lsu_bus_buffer.scala 413:87]
  wire [3:0] buf_rsp_pickage_2 = {_T_2777,_T_2774,_T_2771,_T_2768}; // @[Cat.scala 29:58]
  wire  _T_2041 = |buf_rsp_pickage_2; // @[lsu_bus_buffer.scala 381:65]
  wire  _T_2042 = ~_T_2041; // @[lsu_bus_buffer.scala 381:44]
  wire  _T_2044 = _T_2042 & _T_2743; // @[lsu_bus_buffer.scala 381:70]
  reg [3:0] buf_rspageQ_3; // @[lsu_bus_buffer.scala 500:63]
  wire  _T_2792 = buf_rspageQ_3[3] & _T_2746; // @[lsu_bus_buffer.scala 413:87]
  wire  _T_2789 = buf_rspageQ_3[2] & _T_2743; // @[lsu_bus_buffer.scala 413:87]
  wire  _T_2786 = buf_rspageQ_3[1] & _T_2740; // @[lsu_bus_buffer.scala 413:87]
  wire  _T_2783 = buf_rspageQ_3[0] & _T_2737; // @[lsu_bus_buffer.scala 413:87]
  wire [3:0] buf_rsp_pickage_3 = {_T_2792,_T_2789,_T_2786,_T_2783}; // @[Cat.scala 29:58]
  wire  _T_2045 = |buf_rsp_pickage_3; // @[lsu_bus_buffer.scala 381:65]
  wire  _T_2046 = ~_T_2045; // @[lsu_bus_buffer.scala 381:44]
  wire  _T_2048 = _T_2046 & _T_2746; // @[lsu_bus_buffer.scala 381:70]
  wire [7:0] _T_2104 = {4'h0,_T_2048,_T_2044,_T_2040,_T_2036}; // @[Cat.scala 29:58]
  wire  _T_2107 = _T_2104[4] | _T_2104[5]; // @[lsu_bus_buffer.scala 385:42]
  wire  _T_2109 = _T_2107 | _T_2104[6]; // @[lsu_bus_buffer.scala 385:48]
  wire  _T_2111 = _T_2109 | _T_2104[7]; // @[lsu_bus_buffer.scala 385:54]
  wire  _T_2114 = _T_2104[2] | _T_2104[3]; // @[lsu_bus_buffer.scala 385:67]
  wire  _T_2116 = _T_2114 | _T_2104[6]; // @[lsu_bus_buffer.scala 385:73]
  wire  _T_2118 = _T_2116 | _T_2104[7]; // @[lsu_bus_buffer.scala 385:79]
  wire  _T_2121 = _T_2104[1] | _T_2104[3]; // @[lsu_bus_buffer.scala 385:92]
  wire  _T_2123 = _T_2121 | _T_2104[5]; // @[lsu_bus_buffer.scala 385:98]
  wire  _T_2125 = _T_2123 | _T_2104[7]; // @[lsu_bus_buffer.scala 385:104]
  wire [2:0] _T_2127 = {_T_2111,_T_2118,_T_2125}; // @[Cat.scala 29:58]
  wire  _T_3532 = ibuf_byp | io_ldst_dual_r; // @[lsu_bus_buffer.scala 443:77]
  wire  _T_3533 = ~ibuf_merge_en; // @[lsu_bus_buffer.scala 443:97]
  wire  _T_3534 = _T_3532 & _T_3533; // @[lsu_bus_buffer.scala 443:95]
  wire  _T_3535 = 2'h0 == WrPtr0_r; // @[lsu_bus_buffer.scala 443:117]
  wire  _T_3536 = _T_3534 & _T_3535; // @[lsu_bus_buffer.scala 443:112]
  wire  _T_3537 = ibuf_byp & io_ldst_dual_r; // @[lsu_bus_buffer.scala 443:144]
  wire  _T_3538 = 2'h0 == WrPtr1_r; // @[lsu_bus_buffer.scala 443:166]
  wire  _T_3539 = _T_3537 & _T_3538; // @[lsu_bus_buffer.scala 443:161]
  wire  _T_3540 = _T_3536 | _T_3539; // @[lsu_bus_buffer.scala 443:132]
  wire  _T_3541 = _T_853 & _T_3540; // @[lsu_bus_buffer.scala 443:63]
  wire  _T_3542 = 2'h0 == ibuf_tag; // @[lsu_bus_buffer.scala 443:206]
  wire  _T_3543 = ibuf_drain_vld & _T_3542; // @[lsu_bus_buffer.scala 443:201]
  wire  _T_3544 = _T_3541 | _T_3543; // @[lsu_bus_buffer.scala 443:183]
  wire  _T_3554 = io_lsu_bus_clk_en | io_dec_tlu_force_halt; // @[lsu_bus_buffer.scala 450:46]
  wire  _T_3589 = 3'h3 == buf_state_0; // @[Conditional.scala 37:30]
  reg  _T_4307; // @[Reg.scala 27:20]
  reg  _T_4305; // @[Reg.scala 27:20]
  reg  _T_4303; // @[Reg.scala 27:20]
  reg  _T_4301; // @[Reg.scala 27:20]
  wire [3:0] buf_ldfwd = {_T_4307,_T_4305,_T_4303,_T_4301}; // @[Cat.scala 29:58]
  wire  _T_3641 = buf_dual_0 & buf_dualhi_0; // @[lsu_bus_buffer.scala 471:26]
  wire  _T_3643 = ~buf_write[0]; // @[lsu_bus_buffer.scala 471:44]
  reg [1:0] buf_dualtag_0; // @[Reg.scala 27:20]
  wire  _T_3676 = 3'h4 == buf_state_0; // @[Conditional.scala 37:30]
  wire [3:0] _T_3686 = buf_ldfwd >> buf_dualtag_0; // @[lsu_bus_buffer.scala 483:21]
  wire  _GEN_53 = _T_3555 & buf_cmd_state_bus_en_0; // @[Conditional.scala 39:67]
  wire  _GEN_66 = _T_3551 ? 1'h0 : _GEN_53; // @[Conditional.scala 39:67]
  wire  buf_state_bus_en_0 = _T_3528 ? 1'h0 : _GEN_66; // @[Conditional.scala 40:58]
  wire  _T_3568 = buf_state_bus_en_0 & io_lsu_bus_clk_en; // @[lsu_bus_buffer.scala 456:49]
  wire  _T_3569 = _T_3568 | io_dec_tlu_force_halt; // @[lsu_bus_buffer.scala 456:70]
  wire  _T_3694 = 3'h5 == buf_state_0; // @[Conditional.scala 37:30]
  wire [1:0] RspPtr = _T_2127[1:0]; // @[lsu_bus_buffer.scala 393:10]
  wire  _T_3697 = RspPtr == 2'h0; // @[lsu_bus_buffer.scala 488:37]
  wire  _T_3698 = buf_dualtag_0 == RspPtr; // @[lsu_bus_buffer.scala 488:98]
  wire  _T_3699 = buf_dual_0 & _T_3698; // @[lsu_bus_buffer.scala 488:80]
  wire  _T_3700 = _T_3697 | _T_3699; // @[lsu_bus_buffer.scala 488:65]
  wire  _T_3701 = _T_3700 | io_dec_tlu_force_halt; // @[lsu_bus_buffer.scala 488:112]
  wire  _T_3702 = 3'h6 == buf_state_0; // @[Conditional.scala 37:30]
  wire  _GEN_31 = _T_3694 ? _T_3701 : _T_3702; // @[Conditional.scala 39:67]
  wire  _GEN_37 = _T_3676 ? _T_3569 : _GEN_31; // @[Conditional.scala 39:67]
  wire  _GEN_44 = _T_3589 ? _T_3569 : _GEN_37; // @[Conditional.scala 39:67]
  wire  _GEN_54 = _T_3555 ? _T_3569 : _GEN_44; // @[Conditional.scala 39:67]
  wire  _GEN_64 = _T_3551 ? _T_3554 : _GEN_54; // @[Conditional.scala 39:67]
  wire  buf_state_en_0 = _T_3528 ? _T_3544 : _GEN_64; // @[Conditional.scala 40:58]
  wire  _T_2129 = _T_1853 & buf_state_en_0; // @[lsu_bus_buffer.scala 405:94]
  wire  _T_2135 = ibuf_drain_vld & io_lsu_busreq_r; // @[lsu_bus_buffer.scala 407:23]
  wire  _T_2137 = _T_2135 & _T_3532; // @[lsu_bus_buffer.scala 407:41]
  wire  _T_2139 = _T_2137 & _T_1856; // @[lsu_bus_buffer.scala 407:71]
  wire  _T_2141 = _T_2139 & _T_1854; // @[lsu_bus_buffer.scala 407:92]
  wire  _T_2142 = _T_4471 | _T_2141; // @[lsu_bus_buffer.scala 406:86]
  wire  _T_2143 = ibuf_byp & io_lsu_busreq_r; // @[lsu_bus_buffer.scala 408:17]
  wire  _T_2144 = _T_2143 & io_ldst_dual_r; // @[lsu_bus_buffer.scala 408:35]
  wire  _T_2146 = _T_2144 & _T_1857; // @[lsu_bus_buffer.scala 408:52]
  wire  _T_2148 = _T_2146 & _T_1856; // @[lsu_bus_buffer.scala 408:73]
  wire  _T_2149 = _T_2142 | _T_2148; // @[lsu_bus_buffer.scala 407:114]
  wire  _T_2150 = _T_2129 & _T_2149; // @[lsu_bus_buffer.scala 405:113]
  wire  _T_2152 = _T_2150 | buf_age_0[0]; // @[lsu_bus_buffer.scala 408:97]
  wire  _T_2166 = _T_2139 & _T_1865; // @[lsu_bus_buffer.scala 407:92]
  wire  _T_2167 = _T_4476 | _T_2166; // @[lsu_bus_buffer.scala 406:86]
  wire  _T_2173 = _T_2146 & _T_1867; // @[lsu_bus_buffer.scala 408:73]
  wire  _T_2174 = _T_2167 | _T_2173; // @[lsu_bus_buffer.scala 407:114]
  wire  _T_2175 = _T_2129 & _T_2174; // @[lsu_bus_buffer.scala 405:113]
  wire  _T_2177 = _T_2175 | buf_age_0[1]; // @[lsu_bus_buffer.scala 408:97]
  wire  _T_2191 = _T_2139 & _T_1876; // @[lsu_bus_buffer.scala 407:92]
  wire  _T_2192 = _T_4481 | _T_2191; // @[lsu_bus_buffer.scala 406:86]
  wire  _T_2198 = _T_2146 & _T_1878; // @[lsu_bus_buffer.scala 408:73]
  wire  _T_2199 = _T_2192 | _T_2198; // @[lsu_bus_buffer.scala 407:114]
  wire  _T_2200 = _T_2129 & _T_2199; // @[lsu_bus_buffer.scala 405:113]
  wire  _T_2202 = _T_2200 | buf_age_0[2]; // @[lsu_bus_buffer.scala 408:97]
  wire  _T_2216 = _T_2139 & _T_1887; // @[lsu_bus_buffer.scala 407:92]
  wire  _T_2217 = _T_4486 | _T_2216; // @[lsu_bus_buffer.scala 406:86]
  wire  _T_2223 = _T_2146 & _T_1889; // @[lsu_bus_buffer.scala 408:73]
  wire  _T_2224 = _T_2217 | _T_2223; // @[lsu_bus_buffer.scala 407:114]
  wire  _T_2225 = _T_2129 & _T_2224; // @[lsu_bus_buffer.scala 405:113]
  wire  _T_2227 = _T_2225 | buf_age_0[3]; // @[lsu_bus_buffer.scala 408:97]
  wire [2:0] _T_2229 = {_T_2227,_T_2202,_T_2177}; // @[Cat.scala 29:58]
  wire  _T_3728 = 2'h1 == WrPtr0_r; // @[lsu_bus_buffer.scala 443:117]
  wire  _T_3729 = _T_3534 & _T_3728; // @[lsu_bus_buffer.scala 443:112]
  wire  _T_3731 = 2'h1 == WrPtr1_r; // @[lsu_bus_buffer.scala 443:166]
  wire  _T_3732 = _T_3537 & _T_3731; // @[lsu_bus_buffer.scala 443:161]
  wire  _T_3733 = _T_3729 | _T_3732; // @[lsu_bus_buffer.scala 443:132]
  wire  _T_3734 = _T_853 & _T_3733; // @[lsu_bus_buffer.scala 443:63]
  wire  _T_3735 = 2'h1 == ibuf_tag; // @[lsu_bus_buffer.scala 443:206]
  wire  _T_3736 = ibuf_drain_vld & _T_3735; // @[lsu_bus_buffer.scala 443:201]
  wire  _T_3737 = _T_3734 | _T_3736; // @[lsu_bus_buffer.scala 443:183]
  wire  _T_3782 = 3'h3 == buf_state_1; // @[Conditional.scala 37:30]
  wire  _T_3834 = buf_dual_1 & buf_dualhi_1; // @[lsu_bus_buffer.scala 471:26]
  wire  _T_3836 = ~buf_write[1]; // @[lsu_bus_buffer.scala 471:44]
  reg [1:0] buf_dualtag_1; // @[Reg.scala 27:20]
  wire  _T_3869 = 3'h4 == buf_state_1; // @[Conditional.scala 37:30]
  wire [3:0] _T_3879 = buf_ldfwd >> buf_dualtag_1; // @[lsu_bus_buffer.scala 483:21]
  wire  _GEN_129 = _T_3748 & buf_cmd_state_bus_en_1; // @[Conditional.scala 39:67]
  wire  _GEN_142 = _T_3744 ? 1'h0 : _GEN_129; // @[Conditional.scala 39:67]
  wire  buf_state_bus_en_1 = _T_3721 ? 1'h0 : _GEN_142; // @[Conditional.scala 40:58]
  wire  _T_3761 = buf_state_bus_en_1 & io_lsu_bus_clk_en; // @[lsu_bus_buffer.scala 456:49]
  wire  _T_3762 = _T_3761 | io_dec_tlu_force_halt; // @[lsu_bus_buffer.scala 456:70]
  wire  _T_3887 = 3'h5 == buf_state_1; // @[Conditional.scala 37:30]
  wire  _T_3890 = RspPtr == 2'h1; // @[lsu_bus_buffer.scala 488:37]
  wire  _T_3891 = buf_dualtag_1 == RspPtr; // @[lsu_bus_buffer.scala 488:98]
  wire  _T_3892 = buf_dual_1 & _T_3891; // @[lsu_bus_buffer.scala 488:80]
  wire  _T_3893 = _T_3890 | _T_3892; // @[lsu_bus_buffer.scala 488:65]
  wire  _T_3894 = _T_3893 | io_dec_tlu_force_halt; // @[lsu_bus_buffer.scala 488:112]
  wire  _T_3895 = 3'h6 == buf_state_1; // @[Conditional.scala 37:30]
  wire  _GEN_107 = _T_3887 ? _T_3894 : _T_3895; // @[Conditional.scala 39:67]
  wire  _GEN_113 = _T_3869 ? _T_3762 : _GEN_107; // @[Conditional.scala 39:67]
  wire  _GEN_120 = _T_3782 ? _T_3762 : _GEN_113; // @[Conditional.scala 39:67]
  wire  _GEN_130 = _T_3748 ? _T_3762 : _GEN_120; // @[Conditional.scala 39:67]
  wire  _GEN_140 = _T_3744 ? _T_3554 : _GEN_130; // @[Conditional.scala 39:67]
  wire  buf_state_en_1 = _T_3721 ? _T_3737 : _GEN_140; // @[Conditional.scala 40:58]
  wire  _T_2231 = _T_1864 & buf_state_en_1; // @[lsu_bus_buffer.scala 405:94]
  wire  _T_2241 = _T_2137 & _T_1867; // @[lsu_bus_buffer.scala 407:71]
  wire  _T_2243 = _T_2241 & _T_1854; // @[lsu_bus_buffer.scala 407:92]
  wire  _T_2244 = _T_4471 | _T_2243; // @[lsu_bus_buffer.scala 406:86]
  wire  _T_2248 = _T_2144 & _T_1868; // @[lsu_bus_buffer.scala 408:52]
  wire  _T_2250 = _T_2248 & _T_1856; // @[lsu_bus_buffer.scala 408:73]
  wire  _T_2251 = _T_2244 | _T_2250; // @[lsu_bus_buffer.scala 407:114]
  wire  _T_2252 = _T_2231 & _T_2251; // @[lsu_bus_buffer.scala 405:113]
  wire  _T_2254 = _T_2252 | buf_age_1[0]; // @[lsu_bus_buffer.scala 408:97]
  wire  _T_2268 = _T_2241 & _T_1865; // @[lsu_bus_buffer.scala 407:92]
  wire  _T_2269 = _T_4476 | _T_2268; // @[lsu_bus_buffer.scala 406:86]
  wire  _T_2275 = _T_2248 & _T_1867; // @[lsu_bus_buffer.scala 408:73]
  wire  _T_2276 = _T_2269 | _T_2275; // @[lsu_bus_buffer.scala 407:114]
  wire  _T_2277 = _T_2231 & _T_2276; // @[lsu_bus_buffer.scala 405:113]
  wire  _T_2279 = _T_2277 | buf_age_1[1]; // @[lsu_bus_buffer.scala 408:97]
  wire  _T_2293 = _T_2241 & _T_1876; // @[lsu_bus_buffer.scala 407:92]
  wire  _T_2294 = _T_4481 | _T_2293; // @[lsu_bus_buffer.scala 406:86]
  wire  _T_2300 = _T_2248 & _T_1878; // @[lsu_bus_buffer.scala 408:73]
  wire  _T_2301 = _T_2294 | _T_2300; // @[lsu_bus_buffer.scala 407:114]
  wire  _T_2302 = _T_2231 & _T_2301; // @[lsu_bus_buffer.scala 405:113]
  wire  _T_2304 = _T_2302 | buf_age_1[2]; // @[lsu_bus_buffer.scala 408:97]
  wire  _T_2318 = _T_2241 & _T_1887; // @[lsu_bus_buffer.scala 407:92]
  wire  _T_2319 = _T_4486 | _T_2318; // @[lsu_bus_buffer.scala 406:86]
  wire  _T_2325 = _T_2248 & _T_1889; // @[lsu_bus_buffer.scala 408:73]
  wire  _T_2326 = _T_2319 | _T_2325; // @[lsu_bus_buffer.scala 407:114]
  wire  _T_2327 = _T_2231 & _T_2326; // @[lsu_bus_buffer.scala 405:113]
  wire  _T_2329 = _T_2327 | buf_age_1[3]; // @[lsu_bus_buffer.scala 408:97]
  wire [2:0] _T_2331 = {_T_2329,_T_2304,_T_2279}; // @[Cat.scala 29:58]
  wire  _T_3921 = 2'h2 == WrPtr0_r; // @[lsu_bus_buffer.scala 443:117]
  wire  _T_3922 = _T_3534 & _T_3921; // @[lsu_bus_buffer.scala 443:112]
  wire  _T_3924 = 2'h2 == WrPtr1_r; // @[lsu_bus_buffer.scala 443:166]
  wire  _T_3925 = _T_3537 & _T_3924; // @[lsu_bus_buffer.scala 443:161]
  wire  _T_3926 = _T_3922 | _T_3925; // @[lsu_bus_buffer.scala 443:132]
  wire  _T_3927 = _T_853 & _T_3926; // @[lsu_bus_buffer.scala 443:63]
  wire  _T_3928 = 2'h2 == ibuf_tag; // @[lsu_bus_buffer.scala 443:206]
  wire  _T_3929 = ibuf_drain_vld & _T_3928; // @[lsu_bus_buffer.scala 443:201]
  wire  _T_3930 = _T_3927 | _T_3929; // @[lsu_bus_buffer.scala 443:183]
  wire  _T_3975 = 3'h3 == buf_state_2; // @[Conditional.scala 37:30]
  wire  _T_4027 = buf_dual_2 & buf_dualhi_2; // @[lsu_bus_buffer.scala 471:26]
  wire  _T_4029 = ~buf_write[2]; // @[lsu_bus_buffer.scala 471:44]
  reg [1:0] buf_dualtag_2; // @[Reg.scala 27:20]
  wire  _T_4062 = 3'h4 == buf_state_2; // @[Conditional.scala 37:30]
  wire [3:0] _T_4072 = buf_ldfwd >> buf_dualtag_2; // @[lsu_bus_buffer.scala 483:21]
  wire  _GEN_205 = _T_3941 & buf_cmd_state_bus_en_2; // @[Conditional.scala 39:67]
  wire  _GEN_218 = _T_3937 ? 1'h0 : _GEN_205; // @[Conditional.scala 39:67]
  wire  buf_state_bus_en_2 = _T_3914 ? 1'h0 : _GEN_218; // @[Conditional.scala 40:58]
  wire  _T_3954 = buf_state_bus_en_2 & io_lsu_bus_clk_en; // @[lsu_bus_buffer.scala 456:49]
  wire  _T_3955 = _T_3954 | io_dec_tlu_force_halt; // @[lsu_bus_buffer.scala 456:70]
  wire  _T_4080 = 3'h5 == buf_state_2; // @[Conditional.scala 37:30]
  wire  _T_4083 = RspPtr == 2'h2; // @[lsu_bus_buffer.scala 488:37]
  wire  _T_4084 = buf_dualtag_2 == RspPtr; // @[lsu_bus_buffer.scala 488:98]
  wire  _T_4085 = buf_dual_2 & _T_4084; // @[lsu_bus_buffer.scala 488:80]
  wire  _T_4086 = _T_4083 | _T_4085; // @[lsu_bus_buffer.scala 488:65]
  wire  _T_4087 = _T_4086 | io_dec_tlu_force_halt; // @[lsu_bus_buffer.scala 488:112]
  wire  _T_4088 = 3'h6 == buf_state_2; // @[Conditional.scala 37:30]
  wire  _GEN_183 = _T_4080 ? _T_4087 : _T_4088; // @[Conditional.scala 39:67]
  wire  _GEN_189 = _T_4062 ? _T_3955 : _GEN_183; // @[Conditional.scala 39:67]
  wire  _GEN_196 = _T_3975 ? _T_3955 : _GEN_189; // @[Conditional.scala 39:67]
  wire  _GEN_206 = _T_3941 ? _T_3955 : _GEN_196; // @[Conditional.scala 39:67]
  wire  _GEN_216 = _T_3937 ? _T_3554 : _GEN_206; // @[Conditional.scala 39:67]
  wire  buf_state_en_2 = _T_3914 ? _T_3930 : _GEN_216; // @[Conditional.scala 40:58]
  wire  _T_2333 = _T_1875 & buf_state_en_2; // @[lsu_bus_buffer.scala 405:94]
  wire  _T_2343 = _T_2137 & _T_1878; // @[lsu_bus_buffer.scala 407:71]
  wire  _T_2345 = _T_2343 & _T_1854; // @[lsu_bus_buffer.scala 407:92]
  wire  _T_2346 = _T_4471 | _T_2345; // @[lsu_bus_buffer.scala 406:86]
  wire  _T_2350 = _T_2144 & _T_1879; // @[lsu_bus_buffer.scala 408:52]
  wire  _T_2352 = _T_2350 & _T_1856; // @[lsu_bus_buffer.scala 408:73]
  wire  _T_2353 = _T_2346 | _T_2352; // @[lsu_bus_buffer.scala 407:114]
  wire  _T_2354 = _T_2333 & _T_2353; // @[lsu_bus_buffer.scala 405:113]
  wire  _T_2356 = _T_2354 | buf_age_2[0]; // @[lsu_bus_buffer.scala 408:97]
  wire  _T_2370 = _T_2343 & _T_1865; // @[lsu_bus_buffer.scala 407:92]
  wire  _T_2371 = _T_4476 | _T_2370; // @[lsu_bus_buffer.scala 406:86]
  wire  _T_2377 = _T_2350 & _T_1867; // @[lsu_bus_buffer.scala 408:73]
  wire  _T_2378 = _T_2371 | _T_2377; // @[lsu_bus_buffer.scala 407:114]
  wire  _T_2379 = _T_2333 & _T_2378; // @[lsu_bus_buffer.scala 405:113]
  wire  _T_2381 = _T_2379 | buf_age_2[1]; // @[lsu_bus_buffer.scala 408:97]
  wire  _T_2395 = _T_2343 & _T_1876; // @[lsu_bus_buffer.scala 407:92]
  wire  _T_2396 = _T_4481 | _T_2395; // @[lsu_bus_buffer.scala 406:86]
  wire  _T_2402 = _T_2350 & _T_1878; // @[lsu_bus_buffer.scala 408:73]
  wire  _T_2403 = _T_2396 | _T_2402; // @[lsu_bus_buffer.scala 407:114]
  wire  _T_2404 = _T_2333 & _T_2403; // @[lsu_bus_buffer.scala 405:113]
  wire  _T_2406 = _T_2404 | buf_age_2[2]; // @[lsu_bus_buffer.scala 408:97]
  wire  _T_2420 = _T_2343 & _T_1887; // @[lsu_bus_buffer.scala 407:92]
  wire  _T_2421 = _T_4486 | _T_2420; // @[lsu_bus_buffer.scala 406:86]
  wire  _T_2427 = _T_2350 & _T_1889; // @[lsu_bus_buffer.scala 408:73]
  wire  _T_2428 = _T_2421 | _T_2427; // @[lsu_bus_buffer.scala 407:114]
  wire  _T_2429 = _T_2333 & _T_2428; // @[lsu_bus_buffer.scala 405:113]
  wire  _T_2431 = _T_2429 | buf_age_2[3]; // @[lsu_bus_buffer.scala 408:97]
  wire [2:0] _T_2433 = {_T_2431,_T_2406,_T_2381}; // @[Cat.scala 29:58]
  wire  _T_4114 = 2'h3 == WrPtr0_r; // @[lsu_bus_buffer.scala 443:117]
  wire  _T_4115 = _T_3534 & _T_4114; // @[lsu_bus_buffer.scala 443:112]
  wire  _T_4117 = 2'h3 == WrPtr1_r; // @[lsu_bus_buffer.scala 443:166]
  wire  _T_4118 = _T_3537 & _T_4117; // @[lsu_bus_buffer.scala 443:161]
  wire  _T_4119 = _T_4115 | _T_4118; // @[lsu_bus_buffer.scala 443:132]
  wire  _T_4120 = _T_853 & _T_4119; // @[lsu_bus_buffer.scala 443:63]
  wire  _T_4121 = 2'h3 == ibuf_tag; // @[lsu_bus_buffer.scala 443:206]
  wire  _T_4122 = ibuf_drain_vld & _T_4121; // @[lsu_bus_buffer.scala 443:201]
  wire  _T_4123 = _T_4120 | _T_4122; // @[lsu_bus_buffer.scala 443:183]
  wire  _T_4168 = 3'h3 == buf_state_3; // @[Conditional.scala 37:30]
  wire  _T_4220 = buf_dual_3 & buf_dualhi_3; // @[lsu_bus_buffer.scala 471:26]
  wire  _T_4222 = ~buf_write[3]; // @[lsu_bus_buffer.scala 471:44]
  reg [1:0] buf_dualtag_3; // @[Reg.scala 27:20]
  wire  _T_4255 = 3'h4 == buf_state_3; // @[Conditional.scala 37:30]
  wire [3:0] _T_4265 = buf_ldfwd >> buf_dualtag_3; // @[lsu_bus_buffer.scala 483:21]
  wire  _GEN_281 = _T_4134 & buf_cmd_state_bus_en_3; // @[Conditional.scala 39:67]
  wire  _GEN_294 = _T_4130 ? 1'h0 : _GEN_281; // @[Conditional.scala 39:67]
  wire  buf_state_bus_en_3 = _T_4107 ? 1'h0 : _GEN_294; // @[Conditional.scala 40:58]
  wire  _T_4147 = buf_state_bus_en_3 & io_lsu_bus_clk_en; // @[lsu_bus_buffer.scala 456:49]
  wire  _T_4148 = _T_4147 | io_dec_tlu_force_halt; // @[lsu_bus_buffer.scala 456:70]
  wire  _T_4273 = 3'h5 == buf_state_3; // @[Conditional.scala 37:30]
  wire  _T_4276 = RspPtr == 2'h3; // @[lsu_bus_buffer.scala 488:37]
  wire  _T_4277 = buf_dualtag_3 == RspPtr; // @[lsu_bus_buffer.scala 488:98]
  wire  _T_4278 = buf_dual_3 & _T_4277; // @[lsu_bus_buffer.scala 488:80]
  wire  _T_4279 = _T_4276 | _T_4278; // @[lsu_bus_buffer.scala 488:65]
  wire  _T_4280 = _T_4279 | io_dec_tlu_force_halt; // @[lsu_bus_buffer.scala 488:112]
  wire  _T_4281 = 3'h6 == buf_state_3; // @[Conditional.scala 37:30]
  wire  _GEN_259 = _T_4273 ? _T_4280 : _T_4281; // @[Conditional.scala 39:67]
  wire  _GEN_265 = _T_4255 ? _T_4148 : _GEN_259; // @[Conditional.scala 39:67]
  wire  _GEN_272 = _T_4168 ? _T_4148 : _GEN_265; // @[Conditional.scala 39:67]
  wire  _GEN_282 = _T_4134 ? _T_4148 : _GEN_272; // @[Conditional.scala 39:67]
  wire  _GEN_292 = _T_4130 ? _T_3554 : _GEN_282; // @[Conditional.scala 39:67]
  wire  buf_state_en_3 = _T_4107 ? _T_4123 : _GEN_292; // @[Conditional.scala 40:58]
  wire  _T_2435 = _T_1886 & buf_state_en_3; // @[lsu_bus_buffer.scala 405:94]
  wire  _T_2445 = _T_2137 & _T_1889; // @[lsu_bus_buffer.scala 407:71]
  wire  _T_2447 = _T_2445 & _T_1854; // @[lsu_bus_buffer.scala 407:92]
  wire  _T_2448 = _T_4471 | _T_2447; // @[lsu_bus_buffer.scala 406:86]
  wire  _T_2452 = _T_2144 & _T_1890; // @[lsu_bus_buffer.scala 408:52]
  wire  _T_2454 = _T_2452 & _T_1856; // @[lsu_bus_buffer.scala 408:73]
  wire  _T_2455 = _T_2448 | _T_2454; // @[lsu_bus_buffer.scala 407:114]
  wire  _T_2456 = _T_2435 & _T_2455; // @[lsu_bus_buffer.scala 405:113]
  wire  _T_2458 = _T_2456 | buf_age_3[0]; // @[lsu_bus_buffer.scala 408:97]
  wire  _T_2472 = _T_2445 & _T_1865; // @[lsu_bus_buffer.scala 407:92]
  wire  _T_2473 = _T_4476 | _T_2472; // @[lsu_bus_buffer.scala 406:86]
  wire  _T_2479 = _T_2452 & _T_1867; // @[lsu_bus_buffer.scala 408:73]
  wire  _T_2480 = _T_2473 | _T_2479; // @[lsu_bus_buffer.scala 407:114]
  wire  _T_2481 = _T_2435 & _T_2480; // @[lsu_bus_buffer.scala 405:113]
  wire  _T_2483 = _T_2481 | buf_age_3[1]; // @[lsu_bus_buffer.scala 408:97]
  wire  _T_2497 = _T_2445 & _T_1876; // @[lsu_bus_buffer.scala 407:92]
  wire  _T_2498 = _T_4481 | _T_2497; // @[lsu_bus_buffer.scala 406:86]
  wire  _T_2504 = _T_2452 & _T_1878; // @[lsu_bus_buffer.scala 408:73]
  wire  _T_2505 = _T_2498 | _T_2504; // @[lsu_bus_buffer.scala 407:114]
  wire  _T_2506 = _T_2435 & _T_2505; // @[lsu_bus_buffer.scala 405:113]
  wire  _T_2508 = _T_2506 | buf_age_3[2]; // @[lsu_bus_buffer.scala 408:97]
  wire  _T_2522 = _T_2445 & _T_1887; // @[lsu_bus_buffer.scala 407:92]
  wire  _T_2523 = _T_4486 | _T_2522; // @[lsu_bus_buffer.scala 406:86]
  wire  _T_2529 = _T_2452 & _T_1889; // @[lsu_bus_buffer.scala 408:73]
  wire  _T_2530 = _T_2523 | _T_2529; // @[lsu_bus_buffer.scala 407:114]
  wire  _T_2531 = _T_2435 & _T_2530; // @[lsu_bus_buffer.scala 405:113]
  wire  _T_2533 = _T_2531 | buf_age_3[3]; // @[lsu_bus_buffer.scala 408:97]
  wire [2:0] _T_2535 = {_T_2533,_T_2508,_T_2483}; // @[Cat.scala 29:58]
  wire  _T_2799 = buf_state_0 == 3'h6; // @[lsu_bus_buffer.scala 416:47]
  wire  _T_2800 = _T_1853 | _T_2799; // @[lsu_bus_buffer.scala 416:32]
  wire  _T_2801 = ~_T_2800; // @[lsu_bus_buffer.scala 416:6]
  wire  _T_2809 = _T_2801 | _T_2141; // @[lsu_bus_buffer.scala 416:59]
  wire  _T_2816 = _T_2809 | _T_2148; // @[lsu_bus_buffer.scala 417:110]
  wire  _T_2817 = _T_2129 & _T_2816; // @[lsu_bus_buffer.scala 415:112]
  wire  _T_2821 = buf_state_1 == 3'h6; // @[lsu_bus_buffer.scala 416:47]
  wire  _T_2822 = _T_1864 | _T_2821; // @[lsu_bus_buffer.scala 416:32]
  wire  _T_2823 = ~_T_2822; // @[lsu_bus_buffer.scala 416:6]
  wire  _T_2831 = _T_2823 | _T_2166; // @[lsu_bus_buffer.scala 416:59]
  wire  _T_2838 = _T_2831 | _T_2173; // @[lsu_bus_buffer.scala 417:110]
  wire  _T_2839 = _T_2129 & _T_2838; // @[lsu_bus_buffer.scala 415:112]
  wire  _T_2843 = buf_state_2 == 3'h6; // @[lsu_bus_buffer.scala 416:47]
  wire  _T_2844 = _T_1875 | _T_2843; // @[lsu_bus_buffer.scala 416:32]
  wire  _T_2845 = ~_T_2844; // @[lsu_bus_buffer.scala 416:6]
  wire  _T_2853 = _T_2845 | _T_2191; // @[lsu_bus_buffer.scala 416:59]
  wire  _T_2860 = _T_2853 | _T_2198; // @[lsu_bus_buffer.scala 417:110]
  wire  _T_2861 = _T_2129 & _T_2860; // @[lsu_bus_buffer.scala 415:112]
  wire  _T_2865 = buf_state_3 == 3'h6; // @[lsu_bus_buffer.scala 416:47]
  wire  _T_2866 = _T_1886 | _T_2865; // @[lsu_bus_buffer.scala 416:32]
  wire  _T_2867 = ~_T_2866; // @[lsu_bus_buffer.scala 416:6]
  wire  _T_2875 = _T_2867 | _T_2216; // @[lsu_bus_buffer.scala 416:59]
  wire  _T_2882 = _T_2875 | _T_2223; // @[lsu_bus_buffer.scala 417:110]
  wire  _T_2883 = _T_2129 & _T_2882; // @[lsu_bus_buffer.scala 415:112]
  wire [3:0] buf_rspage_set_0 = {_T_2883,_T_2861,_T_2839,_T_2817}; // @[Cat.scala 29:58]
  wire  _T_2900 = _T_2801 | _T_2243; // @[lsu_bus_buffer.scala 416:59]
  wire  _T_2907 = _T_2900 | _T_2250; // @[lsu_bus_buffer.scala 417:110]
  wire  _T_2908 = _T_2231 & _T_2907; // @[lsu_bus_buffer.scala 415:112]
  wire  _T_2922 = _T_2823 | _T_2268; // @[lsu_bus_buffer.scala 416:59]
  wire  _T_2929 = _T_2922 | _T_2275; // @[lsu_bus_buffer.scala 417:110]
  wire  _T_2930 = _T_2231 & _T_2929; // @[lsu_bus_buffer.scala 415:112]
  wire  _T_2944 = _T_2845 | _T_2293; // @[lsu_bus_buffer.scala 416:59]
  wire  _T_2951 = _T_2944 | _T_2300; // @[lsu_bus_buffer.scala 417:110]
  wire  _T_2952 = _T_2231 & _T_2951; // @[lsu_bus_buffer.scala 415:112]
  wire  _T_2966 = _T_2867 | _T_2318; // @[lsu_bus_buffer.scala 416:59]
  wire  _T_2973 = _T_2966 | _T_2325; // @[lsu_bus_buffer.scala 417:110]
  wire  _T_2974 = _T_2231 & _T_2973; // @[lsu_bus_buffer.scala 415:112]
  wire [3:0] buf_rspage_set_1 = {_T_2974,_T_2952,_T_2930,_T_2908}; // @[Cat.scala 29:58]
  wire  _T_2991 = _T_2801 | _T_2345; // @[lsu_bus_buffer.scala 416:59]
  wire  _T_2998 = _T_2991 | _T_2352; // @[lsu_bus_buffer.scala 417:110]
  wire  _T_2999 = _T_2333 & _T_2998; // @[lsu_bus_buffer.scala 415:112]
  wire  _T_3013 = _T_2823 | _T_2370; // @[lsu_bus_buffer.scala 416:59]
  wire  _T_3020 = _T_3013 | _T_2377; // @[lsu_bus_buffer.scala 417:110]
  wire  _T_3021 = _T_2333 & _T_3020; // @[lsu_bus_buffer.scala 415:112]
  wire  _T_3035 = _T_2845 | _T_2395; // @[lsu_bus_buffer.scala 416:59]
  wire  _T_3042 = _T_3035 | _T_2402; // @[lsu_bus_buffer.scala 417:110]
  wire  _T_3043 = _T_2333 & _T_3042; // @[lsu_bus_buffer.scala 415:112]
  wire  _T_3057 = _T_2867 | _T_2420; // @[lsu_bus_buffer.scala 416:59]
  wire  _T_3064 = _T_3057 | _T_2427; // @[lsu_bus_buffer.scala 417:110]
  wire  _T_3065 = _T_2333 & _T_3064; // @[lsu_bus_buffer.scala 415:112]
  wire [3:0] buf_rspage_set_2 = {_T_3065,_T_3043,_T_3021,_T_2999}; // @[Cat.scala 29:58]
  wire  _T_3082 = _T_2801 | _T_2447; // @[lsu_bus_buffer.scala 416:59]
  wire  _T_3089 = _T_3082 | _T_2454; // @[lsu_bus_buffer.scala 417:110]
  wire  _T_3090 = _T_2435 & _T_3089; // @[lsu_bus_buffer.scala 415:112]
  wire  _T_3104 = _T_2823 | _T_2472; // @[lsu_bus_buffer.scala 416:59]
  wire  _T_3111 = _T_3104 | _T_2479; // @[lsu_bus_buffer.scala 417:110]
  wire  _T_3112 = _T_2435 & _T_3111; // @[lsu_bus_buffer.scala 415:112]
  wire  _T_3126 = _T_2845 | _T_2497; // @[lsu_bus_buffer.scala 416:59]
  wire  _T_3133 = _T_3126 | _T_2504; // @[lsu_bus_buffer.scala 417:110]
  wire  _T_3134 = _T_2435 & _T_3133; // @[lsu_bus_buffer.scala 415:112]
  wire  _T_3148 = _T_2867 | _T_2522; // @[lsu_bus_buffer.scala 416:59]
  wire  _T_3155 = _T_3148 | _T_2529; // @[lsu_bus_buffer.scala 417:110]
  wire  _T_3156 = _T_2435 & _T_3155; // @[lsu_bus_buffer.scala 415:112]
  wire [3:0] buf_rspage_set_3 = {_T_3156,_T_3134,_T_3112,_T_3090}; // @[Cat.scala 29:58]
  wire  _T_3241 = _T_2865 | _T_1886; // @[lsu_bus_buffer.scala 420:110]
  wire  _T_3242 = ~_T_3241; // @[lsu_bus_buffer.scala 420:84]
  wire  _T_3243 = buf_rspageQ_0[3] & _T_3242; // @[lsu_bus_buffer.scala 420:82]
  wire  _T_3235 = _T_2843 | _T_1875; // @[lsu_bus_buffer.scala 420:110]
  wire  _T_3236 = ~_T_3235; // @[lsu_bus_buffer.scala 420:84]
  wire  _T_3237 = buf_rspageQ_0[2] & _T_3236; // @[lsu_bus_buffer.scala 420:82]
  wire  _T_3229 = _T_2821 | _T_1864; // @[lsu_bus_buffer.scala 420:110]
  wire  _T_3230 = ~_T_3229; // @[lsu_bus_buffer.scala 420:84]
  wire  _T_3231 = buf_rspageQ_0[1] & _T_3230; // @[lsu_bus_buffer.scala 420:82]
  wire  _T_3223 = _T_2799 | _T_1853; // @[lsu_bus_buffer.scala 420:110]
  wire  _T_3224 = ~_T_3223; // @[lsu_bus_buffer.scala 420:84]
  wire  _T_3225 = buf_rspageQ_0[0] & _T_3224; // @[lsu_bus_buffer.scala 420:82]
  wire [3:0] buf_rspage_0 = {_T_3243,_T_3237,_T_3231,_T_3225}; // @[Cat.scala 29:58]
  wire  _T_3162 = buf_rspage_set_0[0] | buf_rspage_0[0]; // @[lsu_bus_buffer.scala 419:88]
  wire  _T_3165 = buf_rspage_set_0[1] | buf_rspage_0[1]; // @[lsu_bus_buffer.scala 419:88]
  wire  _T_3168 = buf_rspage_set_0[2] | buf_rspage_0[2]; // @[lsu_bus_buffer.scala 419:88]
  wire  _T_3171 = buf_rspage_set_0[3] | buf_rspage_0[3]; // @[lsu_bus_buffer.scala 419:88]
  wire [2:0] _T_3173 = {_T_3171,_T_3168,_T_3165}; // @[Cat.scala 29:58]
  wire  _T_3270 = buf_rspageQ_1[3] & _T_3242; // @[lsu_bus_buffer.scala 420:82]
  wire  _T_3264 = buf_rspageQ_1[2] & _T_3236; // @[lsu_bus_buffer.scala 420:82]
  wire  _T_3258 = buf_rspageQ_1[1] & _T_3230; // @[lsu_bus_buffer.scala 420:82]
  wire  _T_3252 = buf_rspageQ_1[0] & _T_3224; // @[lsu_bus_buffer.scala 420:82]
  wire [3:0] buf_rspage_1 = {_T_3270,_T_3264,_T_3258,_T_3252}; // @[Cat.scala 29:58]
  wire  _T_3177 = buf_rspage_set_1[0] | buf_rspage_1[0]; // @[lsu_bus_buffer.scala 419:88]
  wire  _T_3180 = buf_rspage_set_1[1] | buf_rspage_1[1]; // @[lsu_bus_buffer.scala 419:88]
  wire  _T_3183 = buf_rspage_set_1[2] | buf_rspage_1[2]; // @[lsu_bus_buffer.scala 419:88]
  wire  _T_3186 = buf_rspage_set_1[3] | buf_rspage_1[3]; // @[lsu_bus_buffer.scala 419:88]
  wire [2:0] _T_3188 = {_T_3186,_T_3183,_T_3180}; // @[Cat.scala 29:58]
  wire  _T_3297 = buf_rspageQ_2[3] & _T_3242; // @[lsu_bus_buffer.scala 420:82]
  wire  _T_3291 = buf_rspageQ_2[2] & _T_3236; // @[lsu_bus_buffer.scala 420:82]
  wire  _T_3285 = buf_rspageQ_2[1] & _T_3230; // @[lsu_bus_buffer.scala 420:82]
  wire  _T_3279 = buf_rspageQ_2[0] & _T_3224; // @[lsu_bus_buffer.scala 420:82]
  wire [3:0] buf_rspage_2 = {_T_3297,_T_3291,_T_3285,_T_3279}; // @[Cat.scala 29:58]
  wire  _T_3192 = buf_rspage_set_2[0] | buf_rspage_2[0]; // @[lsu_bus_buffer.scala 419:88]
  wire  _T_3195 = buf_rspage_set_2[1] | buf_rspage_2[1]; // @[lsu_bus_buffer.scala 419:88]
  wire  _T_3198 = buf_rspage_set_2[2] | buf_rspage_2[2]; // @[lsu_bus_buffer.scala 419:88]
  wire  _T_3201 = buf_rspage_set_2[3] | buf_rspage_2[3]; // @[lsu_bus_buffer.scala 419:88]
  wire [2:0] _T_3203 = {_T_3201,_T_3198,_T_3195}; // @[Cat.scala 29:58]
  wire  _T_3324 = buf_rspageQ_3[3] & _T_3242; // @[lsu_bus_buffer.scala 420:82]
  wire  _T_3318 = buf_rspageQ_3[2] & _T_3236; // @[lsu_bus_buffer.scala 420:82]
  wire  _T_3312 = buf_rspageQ_3[1] & _T_3230; // @[lsu_bus_buffer.scala 420:82]
  wire  _T_3306 = buf_rspageQ_3[0] & _T_3224; // @[lsu_bus_buffer.scala 420:82]
  wire [3:0] buf_rspage_3 = {_T_3324,_T_3318,_T_3312,_T_3306}; // @[Cat.scala 29:58]
  wire  _T_3207 = buf_rspage_set_3[0] | buf_rspage_3[0]; // @[lsu_bus_buffer.scala 419:88]
  wire  _T_3210 = buf_rspage_set_3[1] | buf_rspage_3[1]; // @[lsu_bus_buffer.scala 419:88]
  wire  _T_3213 = buf_rspage_set_3[2] | buf_rspage_3[2]; // @[lsu_bus_buffer.scala 419:88]
  wire  _T_3216 = buf_rspage_set_3[3] | buf_rspage_3[3]; // @[lsu_bus_buffer.scala 419:88]
  wire [2:0] _T_3218 = {_T_3216,_T_3213,_T_3210}; // @[Cat.scala 29:58]
  wire  _T_3329 = ibuf_drain_vld & _T_1854; // @[lsu_bus_buffer.scala 425:63]
  wire  _T_3331 = ibuf_drain_vld & _T_1865; // @[lsu_bus_buffer.scala 425:63]
  wire  _T_3333 = ibuf_drain_vld & _T_1876; // @[lsu_bus_buffer.scala 425:63]
  wire  _T_3335 = ibuf_drain_vld & _T_1887; // @[lsu_bus_buffer.scala 425:63]
  wire [3:0] ibuf_drainvec_vld = {_T_3335,_T_3333,_T_3331,_T_3329}; // @[Cat.scala 29:58]
  wire  _T_3343 = _T_3537 & _T_1857; // @[lsu_bus_buffer.scala 427:35]
  wire  _T_3352 = _T_3537 & _T_1868; // @[lsu_bus_buffer.scala 427:35]
  wire  _T_3361 = _T_3537 & _T_1879; // @[lsu_bus_buffer.scala 427:35]
  wire  _T_3370 = _T_3537 & _T_1890; // @[lsu_bus_buffer.scala 427:35]
  wire  _T_3400 = ibuf_drainvec_vld[0] ? ibuf_dual : io_ldst_dual_r; // @[lsu_bus_buffer.scala 429:45]
  wire  _T_3402 = ibuf_drainvec_vld[1] ? ibuf_dual : io_ldst_dual_r; // @[lsu_bus_buffer.scala 429:45]
  wire  _T_3404 = ibuf_drainvec_vld[2] ? ibuf_dual : io_ldst_dual_r; // @[lsu_bus_buffer.scala 429:45]
  wire  _T_3406 = ibuf_drainvec_vld[3] ? ibuf_dual : io_ldst_dual_r; // @[lsu_bus_buffer.scala 429:45]
  wire [3:0] buf_dual_in = {_T_3406,_T_3404,_T_3402,_T_3400}; // @[Cat.scala 29:58]
  wire  _T_3411 = ibuf_drainvec_vld[0] ? ibuf_samedw : ldst_samedw_r; // @[lsu_bus_buffer.scala 430:47]
  wire  _T_3413 = ibuf_drainvec_vld[1] ? ibuf_samedw : ldst_samedw_r; // @[lsu_bus_buffer.scala 430:47]
  wire  _T_3415 = ibuf_drainvec_vld[2] ? ibuf_samedw : ldst_samedw_r; // @[lsu_bus_buffer.scala 430:47]
  wire  _T_3417 = ibuf_drainvec_vld[3] ? ibuf_samedw : ldst_samedw_r; // @[lsu_bus_buffer.scala 430:47]
  wire [3:0] buf_samedw_in = {_T_3417,_T_3415,_T_3413,_T_3411}; // @[Cat.scala 29:58]
  wire  _T_3422 = ibuf_nomerge | ibuf_force_drain; // @[lsu_bus_buffer.scala 431:84]
  wire  _T_3423 = ibuf_drainvec_vld[0] ? _T_3422 : io_no_dword_merge_r; // @[lsu_bus_buffer.scala 431:48]
  wire  _T_3426 = ibuf_drainvec_vld[1] ? _T_3422 : io_no_dword_merge_r; // @[lsu_bus_buffer.scala 431:48]
  wire  _T_3429 = ibuf_drainvec_vld[2] ? _T_3422 : io_no_dword_merge_r; // @[lsu_bus_buffer.scala 431:48]
  wire  _T_3432 = ibuf_drainvec_vld[3] ? _T_3422 : io_no_dword_merge_r; // @[lsu_bus_buffer.scala 431:48]
  wire [3:0] buf_nomerge_in = {_T_3432,_T_3429,_T_3426,_T_3423}; // @[Cat.scala 29:58]
  wire  _T_3440 = ibuf_drainvec_vld[0] ? ibuf_dual : _T_3343; // @[lsu_bus_buffer.scala 432:47]
  wire  _T_3445 = ibuf_drainvec_vld[1] ? ibuf_dual : _T_3352; // @[lsu_bus_buffer.scala 432:47]
  wire  _T_3450 = ibuf_drainvec_vld[2] ? ibuf_dual : _T_3361; // @[lsu_bus_buffer.scala 432:47]
  wire  _T_3455 = ibuf_drainvec_vld[3] ? ibuf_dual : _T_3370; // @[lsu_bus_buffer.scala 432:47]
  wire [3:0] buf_dualhi_in = {_T_3455,_T_3450,_T_3445,_T_3440}; // @[Cat.scala 29:58]
  wire  _T_3484 = ibuf_drainvec_vld[0] ? ibuf_sideeffect : io_is_sideeffects_r; // @[lsu_bus_buffer.scala 434:51]
  wire  _T_3486 = ibuf_drainvec_vld[1] ? ibuf_sideeffect : io_is_sideeffects_r; // @[lsu_bus_buffer.scala 434:51]
  wire  _T_3488 = ibuf_drainvec_vld[2] ? ibuf_sideeffect : io_is_sideeffects_r; // @[lsu_bus_buffer.scala 434:51]
  wire  _T_3490 = ibuf_drainvec_vld[3] ? ibuf_sideeffect : io_is_sideeffects_r; // @[lsu_bus_buffer.scala 434:51]
  wire [3:0] buf_sideeffect_in = {_T_3490,_T_3488,_T_3486,_T_3484}; // @[Cat.scala 29:58]
  wire  _T_3495 = ibuf_drainvec_vld[0] ? ibuf_unsign : io_lsu_pkt_r_bits_unsign; // @[lsu_bus_buffer.scala 435:47]
  wire  _T_3497 = ibuf_drainvec_vld[1] ? ibuf_unsign : io_lsu_pkt_r_bits_unsign; // @[lsu_bus_buffer.scala 435:47]
  wire  _T_3499 = ibuf_drainvec_vld[2] ? ibuf_unsign : io_lsu_pkt_r_bits_unsign; // @[lsu_bus_buffer.scala 435:47]
  wire  _T_3501 = ibuf_drainvec_vld[3] ? ibuf_unsign : io_lsu_pkt_r_bits_unsign; // @[lsu_bus_buffer.scala 435:47]
  wire [3:0] buf_unsign_in = {_T_3501,_T_3499,_T_3497,_T_3495}; // @[Cat.scala 29:58]
  wire  _T_3518 = ibuf_drainvec_vld[0] ? ibuf_write : io_lsu_pkt_r_bits_store; // @[lsu_bus_buffer.scala 437:46]
  wire  _T_3520 = ibuf_drainvec_vld[1] ? ibuf_write : io_lsu_pkt_r_bits_store; // @[lsu_bus_buffer.scala 437:46]
  wire  _T_3522 = ibuf_drainvec_vld[2] ? ibuf_write : io_lsu_pkt_r_bits_store; // @[lsu_bus_buffer.scala 437:46]
  wire  _T_3524 = ibuf_drainvec_vld[3] ? ibuf_write : io_lsu_pkt_r_bits_store; // @[lsu_bus_buffer.scala 437:46]
  wire [3:0] buf_write_in = {_T_3524,_T_3522,_T_3520,_T_3518}; // @[Cat.scala 29:58]
  wire  _T_3572 = buf_state_en_0 & _T_3643; // @[lsu_bus_buffer.scala 458:44]
  wire  _T_3573 = _T_3572 & obuf_nosend; // @[lsu_bus_buffer.scala 458:60]
  wire  _T_3575 = _T_3573 & _T_1333; // @[lsu_bus_buffer.scala 458:74]
  wire  _T_3594 = io_dec_tlu_force_halt | buf_write[0]; // @[lsu_bus_buffer.scala 465:55]
  wire  _T_3596 = ~buf_samedw_0; // @[lsu_bus_buffer.scala 466:30]
  wire  _T_3597 = buf_dual_0 & _T_3596; // @[lsu_bus_buffer.scala 466:28]
  wire  _T_3600 = _T_3597 & _T_3643; // @[lsu_bus_buffer.scala 466:45]
  wire [2:0] _GEN_19 = 2'h1 == buf_dualtag_0 ? buf_state_1 : buf_state_0; // @[lsu_bus_buffer.scala 466:90]
  wire [2:0] _GEN_20 = 2'h2 == buf_dualtag_0 ? buf_state_2 : _GEN_19; // @[lsu_bus_buffer.scala 466:90]
  wire [2:0] _GEN_21 = 2'h3 == buf_dualtag_0 ? buf_state_3 : _GEN_20; // @[lsu_bus_buffer.scala 466:90]
  wire  _T_3601 = _GEN_21 != 3'h4; // @[lsu_bus_buffer.scala 466:90]
  wire  _T_3602 = _T_3600 & _T_3601; // @[lsu_bus_buffer.scala 466:61]
  wire  _T_4494 = _T_2746 | _T_2743; // @[lsu_bus_buffer.scala 524:93]
  wire  _T_4495 = _T_4494 | _T_2740; // @[lsu_bus_buffer.scala 524:93]
  wire  any_done_wait_state = _T_4495 | _T_2737; // @[lsu_bus_buffer.scala 524:93]
  wire  _T_3604 = buf_ldfwd[0] | any_done_wait_state; // @[lsu_bus_buffer.scala 467:31]
  wire  _T_3610 = buf_dualtag_0 == 2'h0; // @[lsu_bus_buffer.scala 56:118]
  wire  _T_3612 = buf_dualtag_0 == 2'h1; // @[lsu_bus_buffer.scala 56:118]
  wire  _T_3614 = buf_dualtag_0 == 2'h2; // @[lsu_bus_buffer.scala 56:118]
  wire  _T_3616 = buf_dualtag_0 == 2'h3; // @[lsu_bus_buffer.scala 56:118]
  wire  _T_3618 = _T_3610 & buf_ldfwd[0]; // @[Mux.scala 27:72]
  wire  _T_3619 = _T_3612 & buf_ldfwd[1]; // @[Mux.scala 27:72]
  wire  _T_3620 = _T_3614 & buf_ldfwd[2]; // @[Mux.scala 27:72]
  wire  _T_3621 = _T_3616 & buf_ldfwd[3]; // @[Mux.scala 27:72]
  wire  _T_3622 = _T_3618 | _T_3619; // @[Mux.scala 27:72]
  wire  _T_3623 = _T_3622 | _T_3620; // @[Mux.scala 27:72]
  wire  _T_3624 = _T_3623 | _T_3621; // @[Mux.scala 27:72]
  wire  _T_3626 = _T_3600 & _T_3624; // @[lsu_bus_buffer.scala 467:101]
  wire  _T_3627 = _GEN_21 == 3'h4; // @[lsu_bus_buffer.scala 467:167]
  wire  _T_3628 = _T_3626 & _T_3627; // @[lsu_bus_buffer.scala 467:138]
  wire  _T_3629 = _T_3628 & any_done_wait_state; // @[lsu_bus_buffer.scala 467:187]
  wire  _T_3630 = _T_3604 | _T_3629; // @[lsu_bus_buffer.scala 467:53]
  wire  _T_3681 = buf_ldfwd[0] | _T_3686[0]; // @[lsu_bus_buffer.scala 481:90]
  wire  _T_3682 = _T_3681 | any_done_wait_state; // @[lsu_bus_buffer.scala 481:118]
  wire  _GEN_29 = _T_3702 & buf_state_en_0; // @[Conditional.scala 39:67]
  wire  _GEN_32 = _T_3694 ? 1'h0 : _T_3702; // @[Conditional.scala 39:67]
  wire  _GEN_34 = _T_3694 ? 1'h0 : _GEN_29; // @[Conditional.scala 39:67]
  wire  _GEN_38 = _T_3676 ? 1'h0 : _GEN_32; // @[Conditional.scala 39:67]
  wire  _GEN_40 = _T_3676 ? 1'h0 : _GEN_34; // @[Conditional.scala 39:67]
  wire  _GEN_48 = _T_3589 ? 1'h0 : _GEN_38; // @[Conditional.scala 39:67]
  wire  _GEN_50 = _T_3589 ? 1'h0 : _GEN_40; // @[Conditional.scala 39:67]
  wire  _GEN_56 = _T_3555 ? _T_3575 : _GEN_50; // @[Conditional.scala 39:67]
  wire  _GEN_62 = _T_3555 ? 1'h0 : _GEN_48; // @[Conditional.scala 39:67]
  wire  _GEN_68 = _T_3551 ? 1'h0 : _GEN_56; // @[Conditional.scala 39:67]
  wire  _GEN_74 = _T_3551 ? 1'h0 : _GEN_62; // @[Conditional.scala 39:67]
  wire  buf_wr_en_0 = _T_3528 & buf_state_en_0; // @[Conditional.scala 40:58]
  wire  buf_ldfwd_en_0 = _T_3528 ? 1'h0 : _GEN_68; // @[Conditional.scala 40:58]
  wire  buf_rst_0 = _T_3528 ? 1'h0 : _GEN_74; // @[Conditional.scala 40:58]
  wire  _T_3765 = buf_state_en_1 & _T_3836; // @[lsu_bus_buffer.scala 458:44]
  wire  _T_3766 = _T_3765 & obuf_nosend; // @[lsu_bus_buffer.scala 458:60]
  wire  _T_3768 = _T_3766 & _T_1333; // @[lsu_bus_buffer.scala 458:74]
  wire  _T_3787 = io_dec_tlu_force_halt | buf_write[1]; // @[lsu_bus_buffer.scala 465:55]
  wire  _T_3789 = ~buf_samedw_1; // @[lsu_bus_buffer.scala 466:30]
  wire  _T_3790 = buf_dual_1 & _T_3789; // @[lsu_bus_buffer.scala 466:28]
  wire  _T_3793 = _T_3790 & _T_3836; // @[lsu_bus_buffer.scala 466:45]
  wire [2:0] _GEN_95 = 2'h1 == buf_dualtag_1 ? buf_state_1 : buf_state_0; // @[lsu_bus_buffer.scala 466:90]
  wire [2:0] _GEN_96 = 2'h2 == buf_dualtag_1 ? buf_state_2 : _GEN_95; // @[lsu_bus_buffer.scala 466:90]
  wire [2:0] _GEN_97 = 2'h3 == buf_dualtag_1 ? buf_state_3 : _GEN_96; // @[lsu_bus_buffer.scala 466:90]
  wire  _T_3794 = _GEN_97 != 3'h4; // @[lsu_bus_buffer.scala 466:90]
  wire  _T_3795 = _T_3793 & _T_3794; // @[lsu_bus_buffer.scala 466:61]
  wire  _T_3797 = buf_ldfwd[1] | any_done_wait_state; // @[lsu_bus_buffer.scala 467:31]
  wire  _T_3803 = buf_dualtag_1 == 2'h0; // @[lsu_bus_buffer.scala 56:118]
  wire  _T_3805 = buf_dualtag_1 == 2'h1; // @[lsu_bus_buffer.scala 56:118]
  wire  _T_3807 = buf_dualtag_1 == 2'h2; // @[lsu_bus_buffer.scala 56:118]
  wire  _T_3809 = buf_dualtag_1 == 2'h3; // @[lsu_bus_buffer.scala 56:118]
  wire  _T_3811 = _T_3803 & buf_ldfwd[0]; // @[Mux.scala 27:72]
  wire  _T_3812 = _T_3805 & buf_ldfwd[1]; // @[Mux.scala 27:72]
  wire  _T_3813 = _T_3807 & buf_ldfwd[2]; // @[Mux.scala 27:72]
  wire  _T_3814 = _T_3809 & buf_ldfwd[3]; // @[Mux.scala 27:72]
  wire  _T_3815 = _T_3811 | _T_3812; // @[Mux.scala 27:72]
  wire  _T_3816 = _T_3815 | _T_3813; // @[Mux.scala 27:72]
  wire  _T_3817 = _T_3816 | _T_3814; // @[Mux.scala 27:72]
  wire  _T_3819 = _T_3793 & _T_3817; // @[lsu_bus_buffer.scala 467:101]
  wire  _T_3820 = _GEN_97 == 3'h4; // @[lsu_bus_buffer.scala 467:167]
  wire  _T_3821 = _T_3819 & _T_3820; // @[lsu_bus_buffer.scala 467:138]
  wire  _T_3822 = _T_3821 & any_done_wait_state; // @[lsu_bus_buffer.scala 467:187]
  wire  _T_3823 = _T_3797 | _T_3822; // @[lsu_bus_buffer.scala 467:53]
  wire  _T_3874 = buf_ldfwd[1] | _T_3879[0]; // @[lsu_bus_buffer.scala 481:90]
  wire  _T_3875 = _T_3874 | any_done_wait_state; // @[lsu_bus_buffer.scala 481:118]
  wire  _GEN_105 = _T_3895 & buf_state_en_1; // @[Conditional.scala 39:67]
  wire  _GEN_108 = _T_3887 ? 1'h0 : _T_3895; // @[Conditional.scala 39:67]
  wire  _GEN_110 = _T_3887 ? 1'h0 : _GEN_105; // @[Conditional.scala 39:67]
  wire  _GEN_114 = _T_3869 ? 1'h0 : _GEN_108; // @[Conditional.scala 39:67]
  wire  _GEN_116 = _T_3869 ? 1'h0 : _GEN_110; // @[Conditional.scala 39:67]
  wire  _GEN_124 = _T_3782 ? 1'h0 : _GEN_114; // @[Conditional.scala 39:67]
  wire  _GEN_126 = _T_3782 ? 1'h0 : _GEN_116; // @[Conditional.scala 39:67]
  wire  _GEN_132 = _T_3748 ? _T_3768 : _GEN_126; // @[Conditional.scala 39:67]
  wire  _GEN_138 = _T_3748 ? 1'h0 : _GEN_124; // @[Conditional.scala 39:67]
  wire  _GEN_144 = _T_3744 ? 1'h0 : _GEN_132; // @[Conditional.scala 39:67]
  wire  _GEN_150 = _T_3744 ? 1'h0 : _GEN_138; // @[Conditional.scala 39:67]
  wire  buf_wr_en_1 = _T_3721 & buf_state_en_1; // @[Conditional.scala 40:58]
  wire  buf_ldfwd_en_1 = _T_3721 ? 1'h0 : _GEN_144; // @[Conditional.scala 40:58]
  wire  buf_rst_1 = _T_3721 ? 1'h0 : _GEN_150; // @[Conditional.scala 40:58]
  wire  _T_3958 = buf_state_en_2 & _T_4029; // @[lsu_bus_buffer.scala 458:44]
  wire  _T_3959 = _T_3958 & obuf_nosend; // @[lsu_bus_buffer.scala 458:60]
  wire  _T_3961 = _T_3959 & _T_1333; // @[lsu_bus_buffer.scala 458:74]
  wire  _T_3980 = io_dec_tlu_force_halt | buf_write[2]; // @[lsu_bus_buffer.scala 465:55]
  wire  _T_3982 = ~buf_samedw_2; // @[lsu_bus_buffer.scala 466:30]
  wire  _T_3983 = buf_dual_2 & _T_3982; // @[lsu_bus_buffer.scala 466:28]
  wire  _T_3986 = _T_3983 & _T_4029; // @[lsu_bus_buffer.scala 466:45]
  wire [2:0] _GEN_171 = 2'h1 == buf_dualtag_2 ? buf_state_1 : buf_state_0; // @[lsu_bus_buffer.scala 466:90]
  wire [2:0] _GEN_172 = 2'h2 == buf_dualtag_2 ? buf_state_2 : _GEN_171; // @[lsu_bus_buffer.scala 466:90]
  wire [2:0] _GEN_173 = 2'h3 == buf_dualtag_2 ? buf_state_3 : _GEN_172; // @[lsu_bus_buffer.scala 466:90]
  wire  _T_3987 = _GEN_173 != 3'h4; // @[lsu_bus_buffer.scala 466:90]
  wire  _T_3988 = _T_3986 & _T_3987; // @[lsu_bus_buffer.scala 466:61]
  wire  _T_3990 = buf_ldfwd[2] | any_done_wait_state; // @[lsu_bus_buffer.scala 467:31]
  wire  _T_3996 = buf_dualtag_2 == 2'h0; // @[lsu_bus_buffer.scala 56:118]
  wire  _T_3998 = buf_dualtag_2 == 2'h1; // @[lsu_bus_buffer.scala 56:118]
  wire  _T_4000 = buf_dualtag_2 == 2'h2; // @[lsu_bus_buffer.scala 56:118]
  wire  _T_4002 = buf_dualtag_2 == 2'h3; // @[lsu_bus_buffer.scala 56:118]
  wire  _T_4004 = _T_3996 & buf_ldfwd[0]; // @[Mux.scala 27:72]
  wire  _T_4005 = _T_3998 & buf_ldfwd[1]; // @[Mux.scala 27:72]
  wire  _T_4006 = _T_4000 & buf_ldfwd[2]; // @[Mux.scala 27:72]
  wire  _T_4007 = _T_4002 & buf_ldfwd[3]; // @[Mux.scala 27:72]
  wire  _T_4008 = _T_4004 | _T_4005; // @[Mux.scala 27:72]
  wire  _T_4009 = _T_4008 | _T_4006; // @[Mux.scala 27:72]
  wire  _T_4010 = _T_4009 | _T_4007; // @[Mux.scala 27:72]
  wire  _T_4012 = _T_3986 & _T_4010; // @[lsu_bus_buffer.scala 467:101]
  wire  _T_4013 = _GEN_173 == 3'h4; // @[lsu_bus_buffer.scala 467:167]
  wire  _T_4014 = _T_4012 & _T_4013; // @[lsu_bus_buffer.scala 467:138]
  wire  _T_4015 = _T_4014 & any_done_wait_state; // @[lsu_bus_buffer.scala 467:187]
  wire  _T_4016 = _T_3990 | _T_4015; // @[lsu_bus_buffer.scala 467:53]
  wire  _T_4067 = buf_ldfwd[2] | _T_4072[0]; // @[lsu_bus_buffer.scala 481:90]
  wire  _T_4068 = _T_4067 | any_done_wait_state; // @[lsu_bus_buffer.scala 481:118]
  wire  _GEN_181 = _T_4088 & buf_state_en_2; // @[Conditional.scala 39:67]
  wire  _GEN_184 = _T_4080 ? 1'h0 : _T_4088; // @[Conditional.scala 39:67]
  wire  _GEN_186 = _T_4080 ? 1'h0 : _GEN_181; // @[Conditional.scala 39:67]
  wire  _GEN_190 = _T_4062 ? 1'h0 : _GEN_184; // @[Conditional.scala 39:67]
  wire  _GEN_192 = _T_4062 ? 1'h0 : _GEN_186; // @[Conditional.scala 39:67]
  wire  _GEN_200 = _T_3975 ? 1'h0 : _GEN_190; // @[Conditional.scala 39:67]
  wire  _GEN_202 = _T_3975 ? 1'h0 : _GEN_192; // @[Conditional.scala 39:67]
  wire  _GEN_208 = _T_3941 ? _T_3961 : _GEN_202; // @[Conditional.scala 39:67]
  wire  _GEN_214 = _T_3941 ? 1'h0 : _GEN_200; // @[Conditional.scala 39:67]
  wire  _GEN_220 = _T_3937 ? 1'h0 : _GEN_208; // @[Conditional.scala 39:67]
  wire  _GEN_226 = _T_3937 ? 1'h0 : _GEN_214; // @[Conditional.scala 39:67]
  wire  buf_wr_en_2 = _T_3914 & buf_state_en_2; // @[Conditional.scala 40:58]
  wire  buf_ldfwd_en_2 = _T_3914 ? 1'h0 : _GEN_220; // @[Conditional.scala 40:58]
  wire  buf_rst_2 = _T_3914 ? 1'h0 : _GEN_226; // @[Conditional.scala 40:58]
  wire  _T_4151 = buf_state_en_3 & _T_4222; // @[lsu_bus_buffer.scala 458:44]
  wire  _T_4152 = _T_4151 & obuf_nosend; // @[lsu_bus_buffer.scala 458:60]
  wire  _T_4154 = _T_4152 & _T_1333; // @[lsu_bus_buffer.scala 458:74]
  wire  _T_4173 = io_dec_tlu_force_halt | buf_write[3]; // @[lsu_bus_buffer.scala 465:55]
  wire  _T_4175 = ~buf_samedw_3; // @[lsu_bus_buffer.scala 466:30]
  wire  _T_4176 = buf_dual_3 & _T_4175; // @[lsu_bus_buffer.scala 466:28]
  wire  _T_4179 = _T_4176 & _T_4222; // @[lsu_bus_buffer.scala 466:45]
  wire [2:0] _GEN_247 = 2'h1 == buf_dualtag_3 ? buf_state_1 : buf_state_0; // @[lsu_bus_buffer.scala 466:90]
  wire [2:0] _GEN_248 = 2'h2 == buf_dualtag_3 ? buf_state_2 : _GEN_247; // @[lsu_bus_buffer.scala 466:90]
  wire [2:0] _GEN_249 = 2'h3 == buf_dualtag_3 ? buf_state_3 : _GEN_248; // @[lsu_bus_buffer.scala 466:90]
  wire  _T_4180 = _GEN_249 != 3'h4; // @[lsu_bus_buffer.scala 466:90]
  wire  _T_4181 = _T_4179 & _T_4180; // @[lsu_bus_buffer.scala 466:61]
  wire  _T_4183 = buf_ldfwd[3] | any_done_wait_state; // @[lsu_bus_buffer.scala 467:31]
  wire  _T_4189 = buf_dualtag_3 == 2'h0; // @[lsu_bus_buffer.scala 56:118]
  wire  _T_4191 = buf_dualtag_3 == 2'h1; // @[lsu_bus_buffer.scala 56:118]
  wire  _T_4193 = buf_dualtag_3 == 2'h2; // @[lsu_bus_buffer.scala 56:118]
  wire  _T_4195 = buf_dualtag_3 == 2'h3; // @[lsu_bus_buffer.scala 56:118]
  wire  _T_4197 = _T_4189 & buf_ldfwd[0]; // @[Mux.scala 27:72]
  wire  _T_4198 = _T_4191 & buf_ldfwd[1]; // @[Mux.scala 27:72]
  wire  _T_4199 = _T_4193 & buf_ldfwd[2]; // @[Mux.scala 27:72]
  wire  _T_4200 = _T_4195 & buf_ldfwd[3]; // @[Mux.scala 27:72]
  wire  _T_4201 = _T_4197 | _T_4198; // @[Mux.scala 27:72]
  wire  _T_4202 = _T_4201 | _T_4199; // @[Mux.scala 27:72]
  wire  _T_4203 = _T_4202 | _T_4200; // @[Mux.scala 27:72]
  wire  _T_4205 = _T_4179 & _T_4203; // @[lsu_bus_buffer.scala 467:101]
  wire  _T_4206 = _GEN_249 == 3'h4; // @[lsu_bus_buffer.scala 467:167]
  wire  _T_4207 = _T_4205 & _T_4206; // @[lsu_bus_buffer.scala 467:138]
  wire  _T_4208 = _T_4207 & any_done_wait_state; // @[lsu_bus_buffer.scala 467:187]
  wire  _T_4209 = _T_4183 | _T_4208; // @[lsu_bus_buffer.scala 467:53]
  wire  _T_4260 = buf_ldfwd[3] | _T_4265[0]; // @[lsu_bus_buffer.scala 481:90]
  wire  _T_4261 = _T_4260 | any_done_wait_state; // @[lsu_bus_buffer.scala 481:118]
  wire  _GEN_257 = _T_4281 & buf_state_en_3; // @[Conditional.scala 39:67]
  wire  _GEN_260 = _T_4273 ? 1'h0 : _T_4281; // @[Conditional.scala 39:67]
  wire  _GEN_262 = _T_4273 ? 1'h0 : _GEN_257; // @[Conditional.scala 39:67]
  wire  _GEN_266 = _T_4255 ? 1'h0 : _GEN_260; // @[Conditional.scala 39:67]
  wire  _GEN_268 = _T_4255 ? 1'h0 : _GEN_262; // @[Conditional.scala 39:67]
  wire  _GEN_276 = _T_4168 ? 1'h0 : _GEN_266; // @[Conditional.scala 39:67]
  wire  _GEN_278 = _T_4168 ? 1'h0 : _GEN_268; // @[Conditional.scala 39:67]
  wire  _GEN_284 = _T_4134 ? _T_4154 : _GEN_278; // @[Conditional.scala 39:67]
  wire  _GEN_290 = _T_4134 ? 1'h0 : _GEN_276; // @[Conditional.scala 39:67]
  wire  _GEN_296 = _T_4130 ? 1'h0 : _GEN_284; // @[Conditional.scala 39:67]
  wire  _GEN_302 = _T_4130 ? 1'h0 : _GEN_290; // @[Conditional.scala 39:67]
  wire  buf_wr_en_3 = _T_4107 & buf_state_en_3; // @[Conditional.scala 40:58]
  wire  buf_ldfwd_en_3 = _T_4107 ? 1'h0 : _GEN_296; // @[Conditional.scala 40:58]
  wire  buf_rst_3 = _T_4107 ? 1'h0 : _GEN_302; // @[Conditional.scala 40:58]
  reg  _T_4336; // @[Reg.scala 27:20]
  reg  _T_4339; // @[Reg.scala 27:20]
  reg  _T_4342; // @[Reg.scala 27:20]
  reg  _T_4345; // @[Reg.scala 27:20]
  wire [3:0] buf_unsign = {_T_4345,_T_4342,_T_4339,_T_4336}; // @[Cat.scala 29:58]
  reg  _T_4411; // @[lsu_bus_buffer.scala 517:80]
  reg  _T_4406; // @[lsu_bus_buffer.scala 517:80]
  reg  _T_4401; // @[lsu_bus_buffer.scala 517:80]
  reg  _T_4396; // @[lsu_bus_buffer.scala 517:80]
  wire [3:0] buf_error = {_T_4411,_T_4406,_T_4401,_T_4396}; // @[Cat.scala 29:58]
  wire  _T_4394 = ~buf_rst_0; // @[lsu_bus_buffer.scala 517:126]
  wire  _T_4399 = ~buf_rst_1; // @[lsu_bus_buffer.scala 517:126]
  wire  _T_4404 = ~buf_rst_2; // @[lsu_bus_buffer.scala 517:126]
  wire  _T_4409 = ~buf_rst_3; // @[lsu_bus_buffer.scala 517:126]
  wire [1:0] _T_4415 = {io_lsu_busreq_m,1'h0}; // @[Cat.scala 29:58]
  wire [1:0] _T_4416 = io_ldst_dual_m ? _T_4415 : {{1'd0}, io_lsu_busreq_m}; // @[lsu_bus_buffer.scala 520:28]
  wire [1:0] _T_4417 = {io_lsu_busreq_r,1'h0}; // @[Cat.scala 29:58]
  wire [1:0] _T_4418 = io_ldst_dual_r ? _T_4417 : {{1'd0}, io_lsu_busreq_r}; // @[lsu_bus_buffer.scala 520:94]
  wire [2:0] _T_4419 = _T_4416 + _T_4418; // @[lsu_bus_buffer.scala 520:88]
  wire [2:0] _GEN_376 = {{2'd0}, ibuf_valid}; // @[lsu_bus_buffer.scala 520:154]
  wire [3:0] _T_4420 = _T_4419 + _GEN_376; // @[lsu_bus_buffer.scala 520:154]
  wire [1:0] _T_4425 = _T_5 + _T_12; // @[lsu_bus_buffer.scala 520:217]
  wire [1:0] _GEN_377 = {{1'd0}, _T_19}; // @[lsu_bus_buffer.scala 520:217]
  wire [2:0] _T_4426 = _T_4425 + _GEN_377; // @[lsu_bus_buffer.scala 520:217]
  wire [2:0] _GEN_378 = {{2'd0}, _T_26}; // @[lsu_bus_buffer.scala 520:217]
  wire [3:0] _T_4427 = _T_4426 + _GEN_378; // @[lsu_bus_buffer.scala 520:217]
  wire [3:0] buf_numvld_any = _T_4420 + _T_4427; // @[lsu_bus_buffer.scala 520:169]
  wire  _T_4498 = io_ldst_dual_d & io_dec_lsu_valid_raw_d; // @[lsu_bus_buffer.scala 526:52]
  wire  _T_4499 = buf_numvld_any >= 4'h3; // @[lsu_bus_buffer.scala 526:92]
  wire  _T_4500 = buf_numvld_any == 4'h4; // @[lsu_bus_buffer.scala 526:121]
  wire  _T_4502 = |buf_state_0; // @[lsu_bus_buffer.scala 527:52]
  wire  _T_4503 = |buf_state_1; // @[lsu_bus_buffer.scala 527:52]
  wire  _T_4504 = |buf_state_2; // @[lsu_bus_buffer.scala 527:52]
  wire  _T_4505 = |buf_state_3; // @[lsu_bus_buffer.scala 527:52]
  wire  _T_4506 = _T_4502 | _T_4503; // @[lsu_bus_buffer.scala 527:65]
  wire  _T_4507 = _T_4506 | _T_4504; // @[lsu_bus_buffer.scala 527:65]
  wire  _T_4508 = _T_4507 | _T_4505; // @[lsu_bus_buffer.scala 527:65]
  wire  _T_4509 = ~_T_4508; // @[lsu_bus_buffer.scala 527:34]
  wire  _T_4511 = _T_4509 & _T_852; // @[lsu_bus_buffer.scala 527:70]
  wire  _T_4514 = io_lsu_busreq_m & io_lsu_pkt_m_valid; // @[lsu_bus_buffer.scala 529:64]
  wire  _T_4515 = _T_4514 & io_lsu_pkt_m_bits_load; // @[lsu_bus_buffer.scala 529:85]
  wire  _T_4516 = ~io_flush_m_up; // @[lsu_bus_buffer.scala 529:112]
  wire  _T_4517 = _T_4515 & _T_4516; // @[lsu_bus_buffer.scala 529:110]
  wire  _T_4518 = ~io_ld_full_hit_m; // @[lsu_bus_buffer.scala 529:129]
  wire  _T_4520 = ~io_lsu_commit_r; // @[lsu_bus_buffer.scala 532:74]
  reg  lsu_nonblock_load_valid_r; // @[lsu_bus_buffer.scala 617:66]
  wire  _T_4538 = _T_2799 & _T_3643; // @[Mux.scala 27:72]
  wire  _T_4539 = _T_2821 & _T_3836; // @[Mux.scala 27:72]
  wire  _T_4540 = _T_2843 & _T_4029; // @[Mux.scala 27:72]
  wire  _T_4541 = _T_2865 & _T_4222; // @[Mux.scala 27:72]
  wire  _T_4542 = _T_4538 | _T_4539; // @[Mux.scala 27:72]
  wire  _T_4543 = _T_4542 | _T_4540; // @[Mux.scala 27:72]
  wire  lsu_nonblock_load_data_ready = _T_4543 | _T_4541; // @[Mux.scala 27:72]
  wire  _T_4549 = buf_error[0] & _T_3643; // @[lsu_bus_buffer.scala 535:121]
  wire  _T_4554 = buf_error[1] & _T_3836; // @[lsu_bus_buffer.scala 535:121]
  wire  _T_4559 = buf_error[2] & _T_4029; // @[lsu_bus_buffer.scala 535:121]
  wire  _T_4564 = buf_error[3] & _T_4222; // @[lsu_bus_buffer.scala 535:121]
  wire  _T_4565 = _T_2799 & _T_4549; // @[Mux.scala 27:72]
  wire  _T_4566 = _T_2821 & _T_4554; // @[Mux.scala 27:72]
  wire  _T_4567 = _T_2843 & _T_4559; // @[Mux.scala 27:72]
  wire  _T_4568 = _T_2865 & _T_4564; // @[Mux.scala 27:72]
  wire  _T_4569 = _T_4565 | _T_4566; // @[Mux.scala 27:72]
  wire  _T_4570 = _T_4569 | _T_4567; // @[Mux.scala 27:72]
  wire  _T_4577 = ~buf_dual_0; // @[lsu_bus_buffer.scala 536:122]
  wire  _T_4578 = ~buf_dualhi_0; // @[lsu_bus_buffer.scala 536:137]
  wire  _T_4579 = _T_4577 | _T_4578; // @[lsu_bus_buffer.scala 536:135]
  wire  _T_4580 = _T_4538 & _T_4579; // @[lsu_bus_buffer.scala 536:119]
  wire  _T_4585 = ~buf_dual_1; // @[lsu_bus_buffer.scala 536:122]
  wire  _T_4586 = ~buf_dualhi_1; // @[lsu_bus_buffer.scala 536:137]
  wire  _T_4587 = _T_4585 | _T_4586; // @[lsu_bus_buffer.scala 536:135]
  wire  _T_4588 = _T_4539 & _T_4587; // @[lsu_bus_buffer.scala 536:119]
  wire  _T_4593 = ~buf_dual_2; // @[lsu_bus_buffer.scala 536:122]
  wire  _T_4594 = ~buf_dualhi_2; // @[lsu_bus_buffer.scala 536:137]
  wire  _T_4595 = _T_4593 | _T_4594; // @[lsu_bus_buffer.scala 536:135]
  wire  _T_4596 = _T_4540 & _T_4595; // @[lsu_bus_buffer.scala 536:119]
  wire  _T_4601 = ~buf_dual_3; // @[lsu_bus_buffer.scala 536:122]
  wire  _T_4602 = ~buf_dualhi_3; // @[lsu_bus_buffer.scala 536:137]
  wire  _T_4603 = _T_4601 | _T_4602; // @[lsu_bus_buffer.scala 536:135]
  wire  _T_4604 = _T_4541 & _T_4603; // @[lsu_bus_buffer.scala 536:119]
  wire [1:0] _T_4607 = _T_4596 ? 2'h2 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_4608 = _T_4604 ? 2'h3 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _GEN_379 = {{1'd0}, _T_4588}; // @[Mux.scala 27:72]
  wire [1:0] _T_4610 = _GEN_379 | _T_4607; // @[Mux.scala 27:72]
  wire [31:0] _T_4645 = _T_4580 ? buf_data_0 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_4646 = _T_4588 ? buf_data_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_4647 = _T_4596 ? buf_data_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_4648 = _T_4604 ? buf_data_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_4649 = _T_4645 | _T_4646; // @[Mux.scala 27:72]
  wire [31:0] _T_4650 = _T_4649 | _T_4647; // @[Mux.scala 27:72]
  wire [31:0] lsu_nonblock_load_data_lo = _T_4650 | _T_4648; // @[Mux.scala 27:72]
  wire  _T_4657 = _T_4538 & _T_3641; // @[lsu_bus_buffer.scala 538:105]
  wire  _T_4663 = _T_4539 & _T_3834; // @[lsu_bus_buffer.scala 538:105]
  wire  _T_4669 = _T_4540 & _T_4027; // @[lsu_bus_buffer.scala 538:105]
  wire  _T_4675 = _T_4541 & _T_4220; // @[lsu_bus_buffer.scala 538:105]
  wire [31:0] _T_4676 = _T_4657 ? buf_data_0 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_4677 = _T_4663 ? buf_data_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_4678 = _T_4669 ? buf_data_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_4679 = _T_4675 ? buf_data_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_4680 = _T_4676 | _T_4677; // @[Mux.scala 27:72]
  wire [31:0] _T_4681 = _T_4680 | _T_4678; // @[Mux.scala 27:72]
  wire [31:0] lsu_nonblock_load_data_hi = _T_4681 | _T_4679; // @[Mux.scala 27:72]
  wire  _T_4683 = io_dctl_busbuff_lsu_nonblock_load_data_tag == 2'h0; // @[lsu_bus_buffer.scala 57:123]
  wire  _T_4684 = io_dctl_busbuff_lsu_nonblock_load_data_tag == 2'h1; // @[lsu_bus_buffer.scala 57:123]
  wire  _T_4685 = io_dctl_busbuff_lsu_nonblock_load_data_tag == 2'h2; // @[lsu_bus_buffer.scala 57:123]
  wire  _T_4686 = io_dctl_busbuff_lsu_nonblock_load_data_tag == 2'h3; // @[lsu_bus_buffer.scala 57:123]
  wire [31:0] _T_4687 = _T_4683 ? buf_addr_0 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_4688 = _T_4684 ? buf_addr_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_4689 = _T_4685 ? buf_addr_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_4690 = _T_4686 ? buf_addr_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_4691 = _T_4687 | _T_4688; // @[Mux.scala 27:72]
  wire [31:0] _T_4692 = _T_4691 | _T_4689; // @[Mux.scala 27:72]
  wire [31:0] _T_4693 = _T_4692 | _T_4690; // @[Mux.scala 27:72]
  wire [1:0] lsu_nonblock_addr_offset = _T_4693[1:0]; // @[lsu_bus_buffer.scala 539:96]
  wire [1:0] _T_4699 = _T_4683 ? buf_sz_0 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_4700 = _T_4684 ? buf_sz_1 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_4701 = _T_4685 ? buf_sz_2 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_4702 = _T_4686 ? buf_sz_3 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_4703 = _T_4699 | _T_4700; // @[Mux.scala 27:72]
  wire [1:0] _T_4704 = _T_4703 | _T_4701; // @[Mux.scala 27:72]
  wire [1:0] lsu_nonblock_sz = _T_4704 | _T_4702; // @[Mux.scala 27:72]
  wire  _T_4714 = _T_4683 & buf_unsign[0]; // @[Mux.scala 27:72]
  wire  _T_4715 = _T_4684 & buf_unsign[1]; // @[Mux.scala 27:72]
  wire  _T_4716 = _T_4685 & buf_unsign[2]; // @[Mux.scala 27:72]
  wire  _T_4717 = _T_4686 & buf_unsign[3]; // @[Mux.scala 27:72]
  wire  _T_4718 = _T_4714 | _T_4715; // @[Mux.scala 27:72]
  wire  _T_4719 = _T_4718 | _T_4716; // @[Mux.scala 27:72]
  wire  lsu_nonblock_unsign = _T_4719 | _T_4717; // @[Mux.scala 27:72]
  wire [63:0] _T_4739 = {lsu_nonblock_load_data_hi,lsu_nonblock_load_data_lo}; // @[Cat.scala 29:58]
  wire [3:0] _GEN_380 = {{2'd0}, lsu_nonblock_addr_offset}; // @[lsu_bus_buffer.scala 543:121]
  wire [5:0] _T_4740 = _GEN_380 * 4'h8; // @[lsu_bus_buffer.scala 543:121]
  wire [63:0] lsu_nonblock_data_unalgn = _T_4739 >> _T_4740; // @[lsu_bus_buffer.scala 543:92]
  wire  _T_4741 = ~io_dctl_busbuff_lsu_nonblock_load_data_error; // @[lsu_bus_buffer.scala 545:82]
  wire  _T_4743 = lsu_nonblock_sz == 2'h0; // @[lsu_bus_buffer.scala 546:94]
  wire  _T_4744 = lsu_nonblock_unsign & _T_4743; // @[lsu_bus_buffer.scala 546:76]
  wire [31:0] _T_4746 = {24'h0,lsu_nonblock_data_unalgn[7:0]}; // @[Cat.scala 29:58]
  wire  _T_4747 = lsu_nonblock_sz == 2'h1; // @[lsu_bus_buffer.scala 547:45]
  wire  _T_4748 = lsu_nonblock_unsign & _T_4747; // @[lsu_bus_buffer.scala 547:26]
  wire [31:0] _T_4750 = {16'h0,lsu_nonblock_data_unalgn[15:0]}; // @[Cat.scala 29:58]
  wire  _T_4751 = ~lsu_nonblock_unsign; // @[lsu_bus_buffer.scala 548:6]
  wire  _T_4753 = _T_4751 & _T_4743; // @[lsu_bus_buffer.scala 548:27]
  wire [23:0] _T_4756 = lsu_nonblock_data_unalgn[7] ? 24'hffffff : 24'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_4758 = {_T_4756,lsu_nonblock_data_unalgn[7:0]}; // @[Cat.scala 29:58]
  wire  _T_4761 = _T_4751 & _T_4747; // @[lsu_bus_buffer.scala 549:27]
  wire [15:0] _T_4764 = lsu_nonblock_data_unalgn[15] ? 16'hffff : 16'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_4766 = {_T_4764,lsu_nonblock_data_unalgn[15:0]}; // @[Cat.scala 29:58]
  wire  _T_4767 = lsu_nonblock_sz == 2'h2; // @[lsu_bus_buffer.scala 550:21]
  wire [31:0] _T_4768 = _T_4744 ? _T_4746 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_4769 = _T_4748 ? _T_4750 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_4770 = _T_4753 ? _T_4758 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_4771 = _T_4761 ? _T_4766 : 32'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_4772 = _T_4767 ? lsu_nonblock_data_unalgn : 64'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_4773 = _T_4768 | _T_4769; // @[Mux.scala 27:72]
  wire [31:0] _T_4774 = _T_4773 | _T_4770; // @[Mux.scala 27:72]
  wire [31:0] _T_4775 = _T_4774 | _T_4771; // @[Mux.scala 27:72]
  wire [63:0] _GEN_381 = {{32'd0}, _T_4775}; // @[Mux.scala 27:72]
  wire [63:0] _T_4776 = _GEN_381 | _T_4772; // @[Mux.scala 27:72]
  wire  _T_4874 = obuf_valid & obuf_write; // @[lsu_bus_buffer.scala 568:37]
  wire [31:0] _T_4880 = {obuf_addr[31:3],3'h0}; // @[Cat.scala 29:58]
  wire [2:0] _T_4882 = {1'h0,obuf_sz}; // @[Cat.scala 29:58]
  wire [7:0] _T_4892 = obuf_write ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire  _T_4895 = obuf_valid & _T_1343; // @[lsu_bus_buffer.scala 585:37]
  wire  _T_4897 = _T_4895 & _T_1349; // @[lsu_bus_buffer.scala 585:51]
  wire  _T_4909 = io_lsu_bus_clk_en_q & buf_error[0]; // @[lsu_bus_buffer.scala 598:126]
  wire  _T_4911 = _T_4909 & buf_write[0]; // @[lsu_bus_buffer.scala 598:141]
  wire  _T_4914 = io_lsu_bus_clk_en_q & buf_error[1]; // @[lsu_bus_buffer.scala 598:126]
  wire  _T_4916 = _T_4914 & buf_write[1]; // @[lsu_bus_buffer.scala 598:141]
  wire  _T_4919 = io_lsu_bus_clk_en_q & buf_error[2]; // @[lsu_bus_buffer.scala 598:126]
  wire  _T_4921 = _T_4919 & buf_write[2]; // @[lsu_bus_buffer.scala 598:141]
  wire  _T_4924 = io_lsu_bus_clk_en_q & buf_error[3]; // @[lsu_bus_buffer.scala 598:126]
  wire  _T_4926 = _T_4924 & buf_write[3]; // @[lsu_bus_buffer.scala 598:141]
  wire  _T_4927 = _T_2799 & _T_4911; // @[Mux.scala 27:72]
  wire  _T_4928 = _T_2821 & _T_4916; // @[Mux.scala 27:72]
  wire  _T_4929 = _T_2843 & _T_4921; // @[Mux.scala 27:72]
  wire  _T_4930 = _T_2865 & _T_4926; // @[Mux.scala 27:72]
  wire  _T_4931 = _T_4927 | _T_4928; // @[Mux.scala 27:72]
  wire  _T_4932 = _T_4931 | _T_4929; // @[Mux.scala 27:72]
  wire  _T_4942 = _T_2821 & buf_error[1]; // @[lsu_bus_buffer.scala 599:93]
  wire  _T_4944 = _T_4942 & buf_write[1]; // @[lsu_bus_buffer.scala 599:108]
  wire  _T_4947 = _T_2843 & buf_error[2]; // @[lsu_bus_buffer.scala 599:93]
  wire  _T_4949 = _T_4947 & buf_write[2]; // @[lsu_bus_buffer.scala 599:108]
  wire  _T_4952 = _T_2865 & buf_error[3]; // @[lsu_bus_buffer.scala 599:93]
  wire  _T_4954 = _T_4952 & buf_write[3]; // @[lsu_bus_buffer.scala 599:108]
  wire [1:0] _T_4957 = _T_4949 ? 2'h2 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_4958 = _T_4954 ? 2'h3 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _GEN_382 = {{1'd0}, _T_4944}; // @[Mux.scala 27:72]
  wire [1:0] _T_4960 = _GEN_382 | _T_4957; // @[Mux.scala 27:72]
  wire [1:0] lsu_imprecise_error_store_tag = _T_4960 | _T_4958; // @[Mux.scala 27:72]
  wire  _T_4962 = ~io_tlu_busbuff_lsu_imprecise_error_store_any; // @[lsu_bus_buffer.scala 601:97]
  wire [31:0] _GEN_351 = 2'h1 == lsu_imprecise_error_store_tag ? buf_addr_1 : buf_addr_0; // @[lsu_bus_buffer.scala 602:53]
  wire [31:0] _GEN_352 = 2'h2 == lsu_imprecise_error_store_tag ? buf_addr_2 : _GEN_351; // @[lsu_bus_buffer.scala 602:53]
  wire [31:0] _GEN_353 = 2'h3 == lsu_imprecise_error_store_tag ? buf_addr_3 : _GEN_352; // @[lsu_bus_buffer.scala 602:53]
  wire [31:0] _GEN_355 = 2'h1 == io_dctl_busbuff_lsu_nonblock_load_data_tag ? buf_addr_1 : buf_addr_0; // @[lsu_bus_buffer.scala 602:53]
  wire [31:0] _GEN_356 = 2'h2 == io_dctl_busbuff_lsu_nonblock_load_data_tag ? buf_addr_2 : _GEN_355; // @[lsu_bus_buffer.scala 602:53]
  wire [31:0] _GEN_357 = 2'h3 == io_dctl_busbuff_lsu_nonblock_load_data_tag ? buf_addr_3 : _GEN_356; // @[lsu_bus_buffer.scala 602:53]
  wire  _T_4970 = io_lsu_busreq_r & io_ldst_dual_r; // @[lsu_bus_buffer.scala 609:60]
  wire  _T_4977 = io_lsu_axi_aw_valid | io_lsu_axi_w_valid; // @[lsu_bus_buffer.scala 612:83]
  wire  _T_4983 = ~io_flush_r; // @[lsu_bus_buffer.scala 616:75]
  wire  _T_4984 = io_lsu_busreq_m & _T_4983; // @[lsu_bus_buffer.scala 616:73]
  reg  _T_4987; // @[lsu_bus_buffer.scala 616:56]
  rvclkhdr rvclkhdr ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_io_l1clk),
    .io_clk(rvclkhdr_io_clk),
    .io_en(rvclkhdr_io_en),
    .io_scan_mode(rvclkhdr_io_scan_mode)
  );
  rvclkhdr rvclkhdr_1 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_1_io_l1clk),
    .io_clk(rvclkhdr_1_io_clk),
    .io_en(rvclkhdr_1_io_en),
    .io_scan_mode(rvclkhdr_1_io_scan_mode)
  );
  rvclkhdr rvclkhdr_2 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_2_io_l1clk),
    .io_clk(rvclkhdr_2_io_clk),
    .io_en(rvclkhdr_2_io_en),
    .io_scan_mode(rvclkhdr_2_io_scan_mode)
  );
  rvclkhdr rvclkhdr_3 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_3_io_l1clk),
    .io_clk(rvclkhdr_3_io_clk),
    .io_en(rvclkhdr_3_io_en),
    .io_scan_mode(rvclkhdr_3_io_scan_mode)
  );
  rvclkhdr rvclkhdr_4 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_4_io_l1clk),
    .io_clk(rvclkhdr_4_io_clk),
    .io_en(rvclkhdr_4_io_en),
    .io_scan_mode(rvclkhdr_4_io_scan_mode)
  );
  rvclkhdr rvclkhdr_5 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_5_io_l1clk),
    .io_clk(rvclkhdr_5_io_clk),
    .io_en(rvclkhdr_5_io_en),
    .io_scan_mode(rvclkhdr_5_io_scan_mode)
  );
  rvclkhdr rvclkhdr_6 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_6_io_l1clk),
    .io_clk(rvclkhdr_6_io_clk),
    .io_en(rvclkhdr_6_io_en),
    .io_scan_mode(rvclkhdr_6_io_scan_mode)
  );
  rvclkhdr rvclkhdr_7 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_7_io_l1clk),
    .io_clk(rvclkhdr_7_io_clk),
    .io_en(rvclkhdr_7_io_en),
    .io_scan_mode(rvclkhdr_7_io_scan_mode)
  );
  rvclkhdr rvclkhdr_8 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_8_io_l1clk),
    .io_clk(rvclkhdr_8_io_clk),
    .io_en(rvclkhdr_8_io_en),
    .io_scan_mode(rvclkhdr_8_io_scan_mode)
  );
  rvclkhdr rvclkhdr_9 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_9_io_l1clk),
    .io_clk(rvclkhdr_9_io_clk),
    .io_en(rvclkhdr_9_io_en),
    .io_scan_mode(rvclkhdr_9_io_scan_mode)
  );
  rvclkhdr rvclkhdr_10 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_10_io_l1clk),
    .io_clk(rvclkhdr_10_io_clk),
    .io_en(rvclkhdr_10_io_en),
    .io_scan_mode(rvclkhdr_10_io_scan_mode)
  );
  rvclkhdr rvclkhdr_11 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_11_io_l1clk),
    .io_clk(rvclkhdr_11_io_clk),
    .io_en(rvclkhdr_11_io_en),
    .io_scan_mode(rvclkhdr_11_io_scan_mode)
  );
  assign io_tlu_busbuff_lsu_pmu_bus_misaligned = _T_4970 & io_lsu_commit_r; // @[lsu_bus_buffer.scala 609:41]
  assign io_tlu_busbuff_lsu_pmu_bus_error = io_tlu_busbuff_lsu_imprecise_error_load_any | io_tlu_busbuff_lsu_imprecise_error_store_any; // @[lsu_bus_buffer.scala 610:36]
  assign io_tlu_busbuff_lsu_pmu_bus_busy = _T_4977 | io_lsu_axi_ar_valid; // @[lsu_bus_buffer.scala 612:35]
  assign io_tlu_busbuff_lsu_imprecise_error_load_any = io_dctl_busbuff_lsu_nonblock_load_data_error & _T_4962; // @[lsu_bus_buffer.scala 601:47]
  assign io_tlu_busbuff_lsu_imprecise_error_store_any = _T_4932 | _T_4930; // @[lsu_bus_buffer.scala 598:48]
  assign io_tlu_busbuff_lsu_imprecise_error_addr_any = io_tlu_busbuff_lsu_imprecise_error_store_any ? _GEN_353 : _GEN_357; // @[lsu_bus_buffer.scala 602:47]
  assign io_dctl_busbuff_lsu_nonblock_load_valid_m = _T_4517 & _T_4518; // @[lsu_bus_buffer.scala 529:45]
  assign io_dctl_busbuff_lsu_nonblock_load_tag_m = _T_1863 ? 2'h0 : _T_1899; // @[lsu_bus_buffer.scala 530:43]
  assign io_dctl_busbuff_lsu_nonblock_load_inv_r = lsu_nonblock_load_valid_r & _T_4520; // @[lsu_bus_buffer.scala 532:43]
  assign io_dctl_busbuff_lsu_nonblock_load_inv_tag_r = WrPtr0_r; // @[lsu_bus_buffer.scala 533:47]
  assign io_dctl_busbuff_lsu_nonblock_load_data_valid = lsu_nonblock_load_data_ready & _T_4741; // @[lsu_bus_buffer.scala 545:48]
  assign io_dctl_busbuff_lsu_nonblock_load_data_error = _T_4570 | _T_4568; // @[lsu_bus_buffer.scala 535:48]
  assign io_dctl_busbuff_lsu_nonblock_load_data_tag = _T_4610 | _T_4608; // @[lsu_bus_buffer.scala 536:46]
  assign io_dctl_busbuff_lsu_nonblock_load_data = _T_4776[31:0]; // @[lsu_bus_buffer.scala 546:42]
  assign io_lsu_axi_aw_valid = _T_4874 & _T_1239; // @[lsu_bus_buffer.scala 568:23]
  assign io_lsu_axi_aw_bits_addr = obuf_sideeffect ? obuf_addr : _T_4880; // @[lsu_bus_buffer.scala 570:27]
  assign io_lsu_axi_aw_bits_size = obuf_sideeffect ? _T_4882 : 3'h3; // @[lsu_bus_buffer.scala 571:27]
  assign io_lsu_axi_w_valid = _T_4874 & _T_1239; // @[lsu_bus_buffer.scala 580:22]
  assign io_lsu_axi_w_bits_strb = obuf_byteen & _T_4892; // @[lsu_bus_buffer.scala 581:26]
  assign io_lsu_axi_ar_valid = _T_4897 & _T_1239; // @[lsu_bus_buffer.scala 585:23]
  assign io_lsu_axi_ar_bits_addr = obuf_sideeffect ? obuf_addr : _T_4880; // @[lsu_bus_buffer.scala 587:27]
  assign io_lsu_axi_ar_bits_size = obuf_sideeffect ? _T_4882 : 3'h3; // @[lsu_bus_buffer.scala 588:27]
  assign io_lsu_busreq_r = _T_4987; // @[lsu_bus_buffer.scala 616:19]
  assign io_lsu_bus_buffer_pend_any = |buf_numvld_pend_any; // @[lsu_bus_buffer.scala 525:30]
  assign io_lsu_bus_buffer_full_any = _T_4498 ? _T_4499 : _T_4500; // @[lsu_bus_buffer.scala 526:30]
  assign io_lsu_bus_buffer_empty_any = _T_4511 & _T_1231; // @[lsu_bus_buffer.scala 527:31]
  assign io_ld_byte_hit_buf_lo = {_T_69,_T_58}; // @[lsu_bus_buffer.scala 137:25]
  assign io_ld_byte_hit_buf_hi = {_T_84,_T_73}; // @[lsu_bus_buffer.scala 138:25]
  assign io_ld_fwddata_buf_lo = _T_650 | _T_651; // @[lsu_bus_buffer.scala 164:24]
  assign io_ld_fwddata_buf_hi = _T_747 | _T_748; // @[lsu_bus_buffer.scala 170:24]
  assign rvclkhdr_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_io_en = _T_853 & _T_854; // @[lib.scala 371:17]
  assign rvclkhdr_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_1_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_1_io_en = _T_853 & _T_854; // @[lib.scala 371:17]
  assign rvclkhdr_1_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_2_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_2_io_en = _T_1240 & io_lsu_bus_clk_en; // @[lib.scala 371:17]
  assign rvclkhdr_2_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_3_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_3_io_en = _T_1240 & io_lsu_bus_clk_en; // @[lib.scala 371:17]
  assign rvclkhdr_3_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_4_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_4_io_en = _T_3528 & buf_state_en_0; // @[lib.scala 371:17]
  assign rvclkhdr_4_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_5_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_5_io_en = _T_3721 & buf_state_en_1; // @[lib.scala 371:17]
  assign rvclkhdr_5_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_6_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_6_io_en = _T_3914 & buf_state_en_2; // @[lib.scala 371:17]
  assign rvclkhdr_6_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_7_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_7_io_en = _T_4107 & buf_state_en_3; // @[lib.scala 371:17]
  assign rvclkhdr_7_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_8_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_8_io_en = _T_3528 & buf_state_en_0; // @[lib.scala 371:17]
  assign rvclkhdr_8_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_9_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_9_io_en = _T_3721 & buf_state_en_1; // @[lib.scala 371:17]
  assign rvclkhdr_9_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_10_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_10_io_en = _T_3914 & buf_state_en_2; // @[lib.scala 371:17]
  assign rvclkhdr_10_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_11_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_11_io_en = _T_4107 & buf_state_en_3; // @[lib.scala 371:17]
  assign rvclkhdr_11_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  buf_addr_0 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  _T_4360 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  _T_4357 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  _T_4354 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  _T_4351 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  buf_state_0 = _RAND_5[2:0];
  _RAND_6 = {1{`RANDOM}};
  buf_addr_1 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  buf_state_1 = _RAND_7[2:0];
  _RAND_8 = {1{`RANDOM}};
  buf_addr_2 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  buf_state_2 = _RAND_9[2:0];
  _RAND_10 = {1{`RANDOM}};
  buf_addr_3 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  buf_state_3 = _RAND_11[2:0];
  _RAND_12 = {1{`RANDOM}};
  buf_byteen_3 = _RAND_12[3:0];
  _RAND_13 = {1{`RANDOM}};
  buf_byteen_2 = _RAND_13[3:0];
  _RAND_14 = {1{`RANDOM}};
  buf_byteen_1 = _RAND_14[3:0];
  _RAND_15 = {1{`RANDOM}};
  buf_byteen_0 = _RAND_15[3:0];
  _RAND_16 = {1{`RANDOM}};
  buf_ageQ_3 = _RAND_16[3:0];
  _RAND_17 = {1{`RANDOM}};
  _T_1848 = _RAND_17[1:0];
  _RAND_18 = {1{`RANDOM}};
  obuf_merge = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  obuf_tag1 = _RAND_19[1:0];
  _RAND_20 = {1{`RANDOM}};
  obuf_valid = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  obuf_wr_enQ = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  ibuf_addr = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  ibuf_write = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  ibuf_valid = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  ibuf_byteen = _RAND_25[3:0];
  _RAND_26 = {1{`RANDOM}};
  buf_ageQ_2 = _RAND_26[3:0];
  _RAND_27 = {1{`RANDOM}};
  buf_ageQ_1 = _RAND_27[3:0];
  _RAND_28 = {1{`RANDOM}};
  buf_ageQ_0 = _RAND_28[3:0];
  _RAND_29 = {1{`RANDOM}};
  buf_data_0 = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  buf_data_1 = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  buf_data_2 = _RAND_31[31:0];
  _RAND_32 = {1{`RANDOM}};
  buf_data_3 = _RAND_32[31:0];
  _RAND_33 = {1{`RANDOM}};
  ibuf_data = _RAND_33[31:0];
  _RAND_34 = {1{`RANDOM}};
  ibuf_timer = _RAND_34[2:0];
  _RAND_35 = {1{`RANDOM}};
  ibuf_sideeffect = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  WrPtr1_r = _RAND_36[1:0];
  _RAND_37 = {1{`RANDOM}};
  WrPtr0_r = _RAND_37[1:0];
  _RAND_38 = {1{`RANDOM}};
  ibuf_tag = _RAND_38[1:0];
  _RAND_39 = {1{`RANDOM}};
  ibuf_dualtag = _RAND_39[1:0];
  _RAND_40 = {1{`RANDOM}};
  ibuf_dual = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  ibuf_samedw = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  ibuf_nomerge = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  ibuf_unsign = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  ibuf_sz = _RAND_44[1:0];
  _RAND_45 = {1{`RANDOM}};
  obuf_wr_timer = _RAND_45[2:0];
  _RAND_46 = {1{`RANDOM}};
  buf_nomerge_0 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  buf_nomerge_1 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  buf_nomerge_2 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  buf_nomerge_3 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  _T_4330 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  _T_4327 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  _T_4324 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  _T_4321 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  obuf_sideeffect = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  buf_dual_3 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  buf_dual_2 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  buf_dual_1 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  buf_dual_0 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  buf_samedw_3 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  buf_samedw_2 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  buf_samedw_1 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  buf_samedw_0 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  obuf_write = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  obuf_nosend = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  obuf_addr = _RAND_65[31:0];
  _RAND_66 = {1{`RANDOM}};
  buf_sz_0 = _RAND_66[1:0];
  _RAND_67 = {1{`RANDOM}};
  buf_sz_1 = _RAND_67[1:0];
  _RAND_68 = {1{`RANDOM}};
  buf_sz_2 = _RAND_68[1:0];
  _RAND_69 = {1{`RANDOM}};
  buf_sz_3 = _RAND_69[1:0];
  _RAND_70 = {1{`RANDOM}};
  buf_dualhi_3 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  buf_dualhi_2 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  buf_dualhi_1 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  buf_dualhi_0 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  obuf_sz = _RAND_74[1:0];
  _RAND_75 = {1{`RANDOM}};
  obuf_byteen = _RAND_75[7:0];
  _RAND_76 = {1{`RANDOM}};
  buf_rspageQ_0 = _RAND_76[3:0];
  _RAND_77 = {1{`RANDOM}};
  buf_rspageQ_1 = _RAND_77[3:0];
  _RAND_78 = {1{`RANDOM}};
  buf_rspageQ_2 = _RAND_78[3:0];
  _RAND_79 = {1{`RANDOM}};
  buf_rspageQ_3 = _RAND_79[3:0];
  _RAND_80 = {1{`RANDOM}};
  _T_4307 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  _T_4305 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  _T_4303 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  _T_4301 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  buf_dualtag_0 = _RAND_84[1:0];
  _RAND_85 = {1{`RANDOM}};
  buf_dualtag_1 = _RAND_85[1:0];
  _RAND_86 = {1{`RANDOM}};
  buf_dualtag_2 = _RAND_86[1:0];
  _RAND_87 = {1{`RANDOM}};
  buf_dualtag_3 = _RAND_87[1:0];
  _RAND_88 = {1{`RANDOM}};
  _T_4336 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  _T_4339 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  _T_4342 = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  _T_4345 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  _T_4411 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  _T_4406 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  _T_4401 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  _T_4396 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  lsu_nonblock_load_valid_r = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  _T_4987 = _RAND_97[0:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    buf_addr_0 = 32'h0;
  end
  if (reset) begin
    _T_4360 = 1'h0;
  end
  if (reset) begin
    _T_4357 = 1'h0;
  end
  if (reset) begin
    _T_4354 = 1'h0;
  end
  if (reset) begin
    _T_4351 = 1'h0;
  end
  if (reset) begin
    buf_state_0 = 3'h0;
  end
  if (reset) begin
    buf_addr_1 = 32'h0;
  end
  if (reset) begin
    buf_state_1 = 3'h0;
  end
  if (reset) begin
    buf_addr_2 = 32'h0;
  end
  if (reset) begin
    buf_state_2 = 3'h0;
  end
  if (reset) begin
    buf_addr_3 = 32'h0;
  end
  if (reset) begin
    buf_state_3 = 3'h0;
  end
  if (reset) begin
    buf_byteen_3 = 4'h0;
  end
  if (reset) begin
    buf_byteen_2 = 4'h0;
  end
  if (reset) begin
    buf_byteen_1 = 4'h0;
  end
  if (reset) begin
    buf_byteen_0 = 4'h0;
  end
  if (reset) begin
    buf_ageQ_3 = 4'h0;
  end
  if (reset) begin
    _T_1848 = 2'h0;
  end
  if (reset) begin
    obuf_merge = 1'h0;
  end
  if (reset) begin
    obuf_tag1 = 2'h0;
  end
  if (reset) begin
    obuf_valid = 1'h0;
  end
  if (reset) begin
    obuf_wr_enQ = 1'h0;
  end
  if (reset) begin
    ibuf_addr = 32'h0;
  end
  if (reset) begin
    ibuf_write = 1'h0;
  end
  if (reset) begin
    ibuf_valid = 1'h0;
  end
  if (reset) begin
    ibuf_byteen = 4'h0;
  end
  if (reset) begin
    buf_ageQ_2 = 4'h0;
  end
  if (reset) begin
    buf_ageQ_1 = 4'h0;
  end
  if (reset) begin
    buf_ageQ_0 = 4'h0;
  end
  if (reset) begin
    buf_data_0 = 32'h0;
  end
  if (reset) begin
    buf_data_1 = 32'h0;
  end
  if (reset) begin
    buf_data_2 = 32'h0;
  end
  if (reset) begin
    buf_data_3 = 32'h0;
  end
  if (reset) begin
    ibuf_data = 32'h0;
  end
  if (reset) begin
    ibuf_timer = 3'h0;
  end
  if (reset) begin
    ibuf_sideeffect = 1'h0;
  end
  if (reset) begin
    WrPtr1_r = 2'h0;
  end
  if (reset) begin
    WrPtr0_r = 2'h0;
  end
  if (reset) begin
    ibuf_tag = 2'h0;
  end
  if (reset) begin
    ibuf_dualtag = 2'h0;
  end
  if (reset) begin
    ibuf_dual = 1'h0;
  end
  if (reset) begin
    ibuf_samedw = 1'h0;
  end
  if (reset) begin
    ibuf_nomerge = 1'h0;
  end
  if (reset) begin
    ibuf_unsign = 1'h0;
  end
  if (reset) begin
    ibuf_sz = 2'h0;
  end
  if (reset) begin
    obuf_wr_timer = 3'h0;
  end
  if (reset) begin
    buf_nomerge_0 = 1'h0;
  end
  if (reset) begin
    buf_nomerge_1 = 1'h0;
  end
  if (reset) begin
    buf_nomerge_2 = 1'h0;
  end
  if (reset) begin
    buf_nomerge_3 = 1'h0;
  end
  if (reset) begin
    _T_4330 = 1'h0;
  end
  if (reset) begin
    _T_4327 = 1'h0;
  end
  if (reset) begin
    _T_4324 = 1'h0;
  end
  if (reset) begin
    _T_4321 = 1'h0;
  end
  if (reset) begin
    obuf_sideeffect = 1'h0;
  end
  if (reset) begin
    buf_dual_3 = 1'h0;
  end
  if (reset) begin
    buf_dual_2 = 1'h0;
  end
  if (reset) begin
    buf_dual_1 = 1'h0;
  end
  if (reset) begin
    buf_dual_0 = 1'h0;
  end
  if (reset) begin
    buf_samedw_3 = 1'h0;
  end
  if (reset) begin
    buf_samedw_2 = 1'h0;
  end
  if (reset) begin
    buf_samedw_1 = 1'h0;
  end
  if (reset) begin
    buf_samedw_0 = 1'h0;
  end
  if (reset) begin
    obuf_write = 1'h0;
  end
  if (reset) begin
    obuf_nosend = 1'h0;
  end
  if (reset) begin
    obuf_addr = 32'h0;
  end
  if (reset) begin
    buf_sz_0 = 2'h0;
  end
  if (reset) begin
    buf_sz_1 = 2'h0;
  end
  if (reset) begin
    buf_sz_2 = 2'h0;
  end
  if (reset) begin
    buf_sz_3 = 2'h0;
  end
  if (reset) begin
    buf_dualhi_3 = 1'h0;
  end
  if (reset) begin
    buf_dualhi_2 = 1'h0;
  end
  if (reset) begin
    buf_dualhi_1 = 1'h0;
  end
  if (reset) begin
    buf_dualhi_0 = 1'h0;
  end
  if (reset) begin
    obuf_sz = 2'h0;
  end
  if (reset) begin
    obuf_byteen = 8'h0;
  end
  if (reset) begin
    buf_rspageQ_0 = 4'h0;
  end
  if (reset) begin
    buf_rspageQ_1 = 4'h0;
  end
  if (reset) begin
    buf_rspageQ_2 = 4'h0;
  end
  if (reset) begin
    buf_rspageQ_3 = 4'h0;
  end
  if (reset) begin
    _T_4307 = 1'h0;
  end
  if (reset) begin
    _T_4305 = 1'h0;
  end
  if (reset) begin
    _T_4303 = 1'h0;
  end
  if (reset) begin
    _T_4301 = 1'h0;
  end
  if (reset) begin
    buf_dualtag_0 = 2'h0;
  end
  if (reset) begin
    buf_dualtag_1 = 2'h0;
  end
  if (reset) begin
    buf_dualtag_2 = 2'h0;
  end
  if (reset) begin
    buf_dualtag_3 = 2'h0;
  end
  if (reset) begin
    _T_4336 = 1'h0;
  end
  if (reset) begin
    _T_4339 = 1'h0;
  end
  if (reset) begin
    _T_4342 = 1'h0;
  end
  if (reset) begin
    _T_4345 = 1'h0;
  end
  if (reset) begin
    _T_4411 = 1'h0;
  end
  if (reset) begin
    _T_4406 = 1'h0;
  end
  if (reset) begin
    _T_4401 = 1'h0;
  end
  if (reset) begin
    _T_4396 = 1'h0;
  end
  if (reset) begin
    lsu_nonblock_load_valid_r = 1'h0;
  end
  if (reset) begin
    _T_4987 = 1'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge rvclkhdr_4_io_l1clk or posedge reset) begin
    if (reset) begin
      buf_addr_0 <= 32'h0;
    end else if (ibuf_drainvec_vld[0]) begin
      buf_addr_0 <= ibuf_addr;
    end else if (_T_3343) begin
      buf_addr_0 <= io_end_addr_r;
    end else begin
      buf_addr_0 <= io_lsu_addr_r;
    end
  end
  always @(posedge io_lsu_bus_buf_c1_clk or posedge reset) begin
    if (reset) begin
      _T_4360 <= 1'h0;
    end else if (buf_wr_en_3) begin
      _T_4360 <= buf_write_in[3];
    end
  end
  always @(posedge io_lsu_bus_buf_c1_clk or posedge reset) begin
    if (reset) begin
      _T_4357 <= 1'h0;
    end else if (buf_wr_en_2) begin
      _T_4357 <= buf_write_in[2];
    end
  end
  always @(posedge io_lsu_bus_buf_c1_clk or posedge reset) begin
    if (reset) begin
      _T_4354 <= 1'h0;
    end else if (buf_wr_en_1) begin
      _T_4354 <= buf_write_in[1];
    end
  end
  always @(posedge io_lsu_bus_buf_c1_clk or posedge reset) begin
    if (reset) begin
      _T_4351 <= 1'h0;
    end else if (buf_wr_en_0) begin
      _T_4351 <= buf_write_in[0];
    end
  end
  always @(posedge io_lsu_bus_buf_c1_clk or posedge reset) begin
    if (reset) begin
      buf_state_0 <= 3'h0;
    end else if (buf_state_en_0) begin
      if (_T_3528) begin
        if (io_lsu_bus_clk_en) begin
          buf_state_0 <= 3'h2;
        end else begin
          buf_state_0 <= 3'h1;
        end
      end else if (_T_3551) begin
        if (io_dec_tlu_force_halt) begin
          buf_state_0 <= 3'h0;
        end else begin
          buf_state_0 <= 3'h2;
        end
      end else if (_T_3555) begin
        if (io_dec_tlu_force_halt) begin
          buf_state_0 <= 3'h0;
        end else begin
          buf_state_0 <= 3'h3;
        end
      end else if (_T_3589) begin
        if (_T_3594) begin
          buf_state_0 <= 3'h0;
        end else if (_T_3602) begin
          buf_state_0 <= 3'h4;
        end else if (_T_3630) begin
          buf_state_0 <= 3'h5;
        end else begin
          buf_state_0 <= 3'h6;
        end
      end else if (_T_3676) begin
        if (io_dec_tlu_force_halt) begin
          buf_state_0 <= 3'h0;
        end else if (_T_3682) begin
          buf_state_0 <= 3'h5;
        end else begin
          buf_state_0 <= 3'h6;
        end
      end else if (_T_3694) begin
        if (io_dec_tlu_force_halt) begin
          buf_state_0 <= 3'h0;
        end else begin
          buf_state_0 <= 3'h6;
        end
      end else begin
        buf_state_0 <= 3'h0;
      end
    end
  end
  always @(posedge rvclkhdr_5_io_l1clk or posedge reset) begin
    if (reset) begin
      buf_addr_1 <= 32'h0;
    end else if (ibuf_drainvec_vld[1]) begin
      buf_addr_1 <= ibuf_addr;
    end else if (_T_3352) begin
      buf_addr_1 <= io_end_addr_r;
    end else begin
      buf_addr_1 <= io_lsu_addr_r;
    end
  end
  always @(posedge io_lsu_bus_buf_c1_clk or posedge reset) begin
    if (reset) begin
      buf_state_1 <= 3'h0;
    end else if (buf_state_en_1) begin
      if (_T_3721) begin
        if (io_lsu_bus_clk_en) begin
          buf_state_1 <= 3'h2;
        end else begin
          buf_state_1 <= 3'h1;
        end
      end else if (_T_3744) begin
        if (io_dec_tlu_force_halt) begin
          buf_state_1 <= 3'h0;
        end else begin
          buf_state_1 <= 3'h2;
        end
      end else if (_T_3748) begin
        if (io_dec_tlu_force_halt) begin
          buf_state_1 <= 3'h0;
        end else begin
          buf_state_1 <= 3'h3;
        end
      end else if (_T_3782) begin
        if (_T_3787) begin
          buf_state_1 <= 3'h0;
        end else if (_T_3795) begin
          buf_state_1 <= 3'h4;
        end else if (_T_3823) begin
          buf_state_1 <= 3'h5;
        end else begin
          buf_state_1 <= 3'h6;
        end
      end else if (_T_3869) begin
        if (io_dec_tlu_force_halt) begin
          buf_state_1 <= 3'h0;
        end else if (_T_3875) begin
          buf_state_1 <= 3'h5;
        end else begin
          buf_state_1 <= 3'h6;
        end
      end else if (_T_3887) begin
        if (io_dec_tlu_force_halt) begin
          buf_state_1 <= 3'h0;
        end else begin
          buf_state_1 <= 3'h6;
        end
      end else begin
        buf_state_1 <= 3'h0;
      end
    end
  end
  always @(posedge rvclkhdr_6_io_l1clk or posedge reset) begin
    if (reset) begin
      buf_addr_2 <= 32'h0;
    end else if (ibuf_drainvec_vld[2]) begin
      buf_addr_2 <= ibuf_addr;
    end else if (_T_3361) begin
      buf_addr_2 <= io_end_addr_r;
    end else begin
      buf_addr_2 <= io_lsu_addr_r;
    end
  end
  always @(posedge io_lsu_bus_buf_c1_clk or posedge reset) begin
    if (reset) begin
      buf_state_2 <= 3'h0;
    end else if (buf_state_en_2) begin
      if (_T_3914) begin
        if (io_lsu_bus_clk_en) begin
          buf_state_2 <= 3'h2;
        end else begin
          buf_state_2 <= 3'h1;
        end
      end else if (_T_3937) begin
        if (io_dec_tlu_force_halt) begin
          buf_state_2 <= 3'h0;
        end else begin
          buf_state_2 <= 3'h2;
        end
      end else if (_T_3941) begin
        if (io_dec_tlu_force_halt) begin
          buf_state_2 <= 3'h0;
        end else begin
          buf_state_2 <= 3'h3;
        end
      end else if (_T_3975) begin
        if (_T_3980) begin
          buf_state_2 <= 3'h0;
        end else if (_T_3988) begin
          buf_state_2 <= 3'h4;
        end else if (_T_4016) begin
          buf_state_2 <= 3'h5;
        end else begin
          buf_state_2 <= 3'h6;
        end
      end else if (_T_4062) begin
        if (io_dec_tlu_force_halt) begin
          buf_state_2 <= 3'h0;
        end else if (_T_4068) begin
          buf_state_2 <= 3'h5;
        end else begin
          buf_state_2 <= 3'h6;
        end
      end else if (_T_4080) begin
        if (io_dec_tlu_force_halt) begin
          buf_state_2 <= 3'h0;
        end else begin
          buf_state_2 <= 3'h6;
        end
      end else begin
        buf_state_2 <= 3'h0;
      end
    end
  end
  always @(posedge rvclkhdr_7_io_l1clk or posedge reset) begin
    if (reset) begin
      buf_addr_3 <= 32'h0;
    end else if (ibuf_drainvec_vld[3]) begin
      buf_addr_3 <= ibuf_addr;
    end else if (_T_3370) begin
      buf_addr_3 <= io_end_addr_r;
    end else begin
      buf_addr_3 <= io_lsu_addr_r;
    end
  end
  always @(posedge io_lsu_bus_buf_c1_clk or posedge reset) begin
    if (reset) begin
      buf_state_3 <= 3'h0;
    end else if (buf_state_en_3) begin
      if (_T_4107) begin
        if (io_lsu_bus_clk_en) begin
          buf_state_3 <= 3'h2;
        end else begin
          buf_state_3 <= 3'h1;
        end
      end else if (_T_4130) begin
        if (io_dec_tlu_force_halt) begin
          buf_state_3 <= 3'h0;
        end else begin
          buf_state_3 <= 3'h2;
        end
      end else if (_T_4134) begin
        if (io_dec_tlu_force_halt) begin
          buf_state_3 <= 3'h0;
        end else begin
          buf_state_3 <= 3'h3;
        end
      end else if (_T_4168) begin
        if (_T_4173) begin
          buf_state_3 <= 3'h0;
        end else if (_T_4181) begin
          buf_state_3 <= 3'h4;
        end else if (_T_4209) begin
          buf_state_3 <= 3'h5;
        end else begin
          buf_state_3 <= 3'h6;
        end
      end else if (_T_4255) begin
        if (io_dec_tlu_force_halt) begin
          buf_state_3 <= 3'h0;
        end else if (_T_4261) begin
          buf_state_3 <= 3'h5;
        end else begin
          buf_state_3 <= 3'h6;
        end
      end else if (_T_4273) begin
        if (io_dec_tlu_force_halt) begin
          buf_state_3 <= 3'h0;
        end else begin
          buf_state_3 <= 3'h6;
        end
      end else begin
        buf_state_3 <= 3'h0;
      end
    end
  end
  always @(posedge io_lsu_bus_buf_c1_clk or posedge reset) begin
    if (reset) begin
      buf_byteen_3 <= 4'h0;
    end else if (buf_wr_en_3) begin
      if (ibuf_drainvec_vld[3]) begin
        buf_byteen_3 <= ibuf_byteen_out;
      end else if (_T_3370) begin
        buf_byteen_3 <= ldst_byteen_hi_r;
      end else begin
        buf_byteen_3 <= ldst_byteen_lo_r;
      end
    end
  end
  always @(posedge io_lsu_bus_buf_c1_clk or posedge reset) begin
    if (reset) begin
      buf_byteen_2 <= 4'h0;
    end else if (buf_wr_en_2) begin
      if (ibuf_drainvec_vld[2]) begin
        buf_byteen_2 <= ibuf_byteen_out;
      end else if (_T_3361) begin
        buf_byteen_2 <= ldst_byteen_hi_r;
      end else begin
        buf_byteen_2 <= ldst_byteen_lo_r;
      end
    end
  end
  always @(posedge io_lsu_bus_buf_c1_clk or posedge reset) begin
    if (reset) begin
      buf_byteen_1 <= 4'h0;
    end else if (buf_wr_en_1) begin
      if (ibuf_drainvec_vld[1]) begin
        buf_byteen_1 <= ibuf_byteen_out;
      end else if (_T_3352) begin
        buf_byteen_1 <= ldst_byteen_hi_r;
      end else begin
        buf_byteen_1 <= ldst_byteen_lo_r;
      end
    end
  end
  always @(posedge io_lsu_bus_buf_c1_clk or posedge reset) begin
    if (reset) begin
      buf_byteen_0 <= 4'h0;
    end else if (buf_wr_en_0) begin
      if (ibuf_drainvec_vld[0]) begin
        buf_byteen_0 <= ibuf_byteen_out;
      end else if (_T_3343) begin
        buf_byteen_0 <= ldst_byteen_hi_r;
      end else begin
        buf_byteen_0 <= ldst_byteen_lo_r;
      end
    end
  end
  always @(posedge io_lsu_bus_buf_c1_clk or posedge reset) begin
    if (reset) begin
      buf_ageQ_3 <= 4'h0;
    end else begin
      buf_ageQ_3 <= {_T_2535,_T_2458};
    end
  end
  always @(posedge io_lsu_bus_obuf_c1_clk or posedge reset) begin
    if (reset) begin
      _T_1848 <= 2'h0;
    end else if (obuf_wr_en) begin
      if (ibuf_buf_byp) begin
        _T_1848 <= WrPtr0_r;
      end else begin
        _T_1848 <= CmdPtr0;
      end
    end
  end
  always @(posedge io_lsu_bus_obuf_c1_clk or posedge reset) begin
    if (reset) begin
      obuf_merge <= 1'h0;
    end else if (obuf_wr_en) begin
      obuf_merge <= obuf_merge_en;
    end
  end
  always @(posedge io_lsu_bus_obuf_c1_clk or posedge reset) begin
    if (reset) begin
      obuf_tag1 <= 2'h0;
    end else if (obuf_wr_en) begin
      if (ibuf_buf_byp) begin
        obuf_tag1 <= WrPtr1_r;
      end else begin
        obuf_tag1 <= CmdPtr1;
      end
    end
  end
  always @(posedge io_lsu_free_c2_clk or posedge reset) begin
    if (reset) begin
      obuf_valid <= 1'h0;
    end else begin
      obuf_valid <= _T_1839 & _T_1840;
    end
  end
  always @(posedge io_lsu_busm_clk or posedge reset) begin
    if (reset) begin
      obuf_wr_enQ <= 1'h0;
    end else begin
      obuf_wr_enQ <= _T_1240 & io_lsu_bus_clk_en;
    end
  end
  always @(posedge rvclkhdr_io_l1clk or posedge reset) begin
    if (reset) begin
      ibuf_addr <= 32'h0;
    end else if (io_ldst_dual_r) begin
      ibuf_addr <= io_end_addr_r;
    end else begin
      ibuf_addr <= io_lsu_addr_r;
    end
  end
  always @(posedge io_lsu_bus_ibuf_c1_clk or posedge reset) begin
    if (reset) begin
      ibuf_write <= 1'h0;
    end else if (ibuf_wr_en) begin
      ibuf_write <= io_lsu_pkt_r_bits_store;
    end
  end
  always @(posedge io_lsu_free_c2_clk or posedge reset) begin
    if (reset) begin
      ibuf_valid <= 1'h0;
    end else begin
      ibuf_valid <= _T_1005 & _T_1006;
    end
  end
  always @(posedge io_lsu_bus_ibuf_c1_clk or posedge reset) begin
    if (reset) begin
      ibuf_byteen <= 4'h0;
    end else if (ibuf_wr_en) begin
      if (_T_866) begin
        ibuf_byteen <= _T_881;
      end else if (io_ldst_dual_r) begin
        ibuf_byteen <= ldst_byteen_hi_r;
      end else begin
        ibuf_byteen <= ldst_byteen_lo_r;
      end
    end
  end
  always @(posedge io_lsu_bus_buf_c1_clk or posedge reset) begin
    if (reset) begin
      buf_ageQ_2 <= 4'h0;
    end else begin
      buf_ageQ_2 <= {_T_2433,_T_2356};
    end
  end
  always @(posedge io_lsu_bus_buf_c1_clk or posedge reset) begin
    if (reset) begin
      buf_ageQ_1 <= 4'h0;
    end else begin
      buf_ageQ_1 <= {_T_2331,_T_2254};
    end
  end
  always @(posedge io_lsu_bus_buf_c1_clk or posedge reset) begin
    if (reset) begin
      buf_ageQ_0 <= 4'h0;
    end else begin
      buf_ageQ_0 <= {_T_2229,_T_2152};
    end
  end
  always @(posedge rvclkhdr_8_io_l1clk or posedge reset) begin
    if (reset) begin
      buf_data_0 <= 32'h0;
    end else if (_T_3528) begin
      if (_T_3543) begin
        buf_data_0 <= ibuf_data_out;
      end else begin
        buf_data_0 <= store_data_lo_r;
      end
    end else begin
      buf_data_0 <= 32'h0;
    end
  end
  always @(posedge rvclkhdr_9_io_l1clk or posedge reset) begin
    if (reset) begin
      buf_data_1 <= 32'h0;
    end else if (_T_3721) begin
      if (_T_3736) begin
        buf_data_1 <= ibuf_data_out;
      end else begin
        buf_data_1 <= store_data_lo_r;
      end
    end else begin
      buf_data_1 <= 32'h0;
    end
  end
  always @(posedge rvclkhdr_10_io_l1clk or posedge reset) begin
    if (reset) begin
      buf_data_2 <= 32'h0;
    end else if (_T_3914) begin
      if (_T_3929) begin
        buf_data_2 <= ibuf_data_out;
      end else begin
        buf_data_2 <= store_data_lo_r;
      end
    end else begin
      buf_data_2 <= 32'h0;
    end
  end
  always @(posedge rvclkhdr_11_io_l1clk or posedge reset) begin
    if (reset) begin
      buf_data_3 <= 32'h0;
    end else if (_T_4107) begin
      if (_T_4122) begin
        buf_data_3 <= ibuf_data_out;
      end else begin
        buf_data_3 <= store_data_lo_r;
      end
    end else begin
      buf_data_3 <= 32'h0;
    end
  end
  always @(posedge rvclkhdr_1_io_l1clk or posedge reset) begin
    if (reset) begin
      ibuf_data <= 32'h0;
    end else begin
      ibuf_data <= {_T_922,_T_893};
    end
  end
  always @(posedge io_lsu_free_c2_clk or posedge reset) begin
    if (reset) begin
      ibuf_timer <= 3'h0;
    end else if (ibuf_wr_en) begin
      ibuf_timer <= 3'h0;
    end else if (_T_923) begin
      ibuf_timer <= _T_926;
    end
  end
  always @(posedge io_lsu_bus_ibuf_c1_clk or posedge reset) begin
    if (reset) begin
      ibuf_sideeffect <= 1'h0;
    end else if (ibuf_wr_en) begin
      ibuf_sideeffect <= io_is_sideeffects_r;
    end
  end
  always @(posedge io_lsu_c2_r_clk or posedge reset) begin
    if (reset) begin
      WrPtr1_r <= 2'h0;
    end else if (_T_1914) begin
      WrPtr1_r <= 2'h0;
    end else if (_T_1928) begin
      WrPtr1_r <= 2'h1;
    end else if (_T_1942) begin
      WrPtr1_r <= 2'h2;
    end else begin
      WrPtr1_r <= 2'h3;
    end
  end
  always @(posedge io_lsu_c2_r_clk or posedge reset) begin
    if (reset) begin
      WrPtr0_r <= 2'h0;
    end else if (_T_1863) begin
      WrPtr0_r <= 2'h0;
    end else if (_T_1874) begin
      WrPtr0_r <= 2'h1;
    end else if (_T_1885) begin
      WrPtr0_r <= 2'h2;
    end else begin
      WrPtr0_r <= 2'h3;
    end
  end
  always @(posedge io_lsu_bus_ibuf_c1_clk or posedge reset) begin
    if (reset) begin
      ibuf_tag <= 2'h0;
    end else if (ibuf_wr_en) begin
      if (!(_T_866)) begin
        if (io_ldst_dual_r) begin
          ibuf_tag <= WrPtr1_r;
        end else begin
          ibuf_tag <= WrPtr0_r;
        end
      end
    end
  end
  always @(posedge io_lsu_bus_ibuf_c1_clk or posedge reset) begin
    if (reset) begin
      ibuf_dualtag <= 2'h0;
    end else if (ibuf_wr_en) begin
      ibuf_dualtag <= WrPtr0_r;
    end
  end
  always @(posedge io_lsu_bus_ibuf_c1_clk or posedge reset) begin
    if (reset) begin
      ibuf_dual <= 1'h0;
    end else if (ibuf_wr_en) begin
      ibuf_dual <= io_ldst_dual_r;
    end
  end
  always @(posedge io_lsu_bus_ibuf_c1_clk or posedge reset) begin
    if (reset) begin
      ibuf_samedw <= 1'h0;
    end else if (ibuf_wr_en) begin
      ibuf_samedw <= ldst_samedw_r;
    end
  end
  always @(posedge io_lsu_bus_ibuf_c1_clk or posedge reset) begin
    if (reset) begin
      ibuf_nomerge <= 1'h0;
    end else if (ibuf_wr_en) begin
      ibuf_nomerge <= io_no_dword_merge_r;
    end
  end
  always @(posedge io_lsu_bus_ibuf_c1_clk or posedge reset) begin
    if (reset) begin
      ibuf_unsign <= 1'h0;
    end else if (ibuf_wr_en) begin
      ibuf_unsign <= io_lsu_pkt_r_bits_unsign;
    end
  end
  always @(posedge io_lsu_bus_ibuf_c1_clk or posedge reset) begin
    if (reset) begin
      ibuf_sz <= 2'h0;
    end else if (ibuf_wr_en) begin
      ibuf_sz <= ibuf_sz_in;
    end
  end
  always @(posedge io_lsu_busm_clk or posedge reset) begin
    if (reset) begin
      obuf_wr_timer <= 3'h0;
    end else if (obuf_wr_en) begin
      obuf_wr_timer <= 3'h0;
    end else if (_T_1058) begin
      obuf_wr_timer <= _T_1060;
    end
  end
  always @(posedge io_lsu_bus_buf_c1_clk or posedge reset) begin
    if (reset) begin
      buf_nomerge_0 <= 1'h0;
    end else if (buf_wr_en_0) begin
      buf_nomerge_0 <= buf_nomerge_in[0];
    end
  end
  always @(posedge io_lsu_bus_buf_c1_clk or posedge reset) begin
    if (reset) begin
      buf_nomerge_1 <= 1'h0;
    end else if (buf_wr_en_1) begin
      buf_nomerge_1 <= buf_nomerge_in[1];
    end
  end
  always @(posedge io_lsu_bus_buf_c1_clk or posedge reset) begin
    if (reset) begin
      buf_nomerge_2 <= 1'h0;
    end else if (buf_wr_en_2) begin
      buf_nomerge_2 <= buf_nomerge_in[2];
    end
  end
  always @(posedge io_lsu_bus_buf_c1_clk or posedge reset) begin
    if (reset) begin
      buf_nomerge_3 <= 1'h0;
    end else if (buf_wr_en_3) begin
      buf_nomerge_3 <= buf_nomerge_in[3];
    end
  end
  always @(posedge io_lsu_bus_buf_c1_clk or posedge reset) begin
    if (reset) begin
      _T_4330 <= 1'h0;
    end else if (buf_wr_en_3) begin
      _T_4330 <= buf_sideeffect_in[3];
    end
  end
  always @(posedge io_lsu_bus_buf_c1_clk or posedge reset) begin
    if (reset) begin
      _T_4327 <= 1'h0;
    end else if (buf_wr_en_2) begin
      _T_4327 <= buf_sideeffect_in[2];
    end
  end
  always @(posedge io_lsu_bus_buf_c1_clk or posedge reset) begin
    if (reset) begin
      _T_4324 <= 1'h0;
    end else if (buf_wr_en_1) begin
      _T_4324 <= buf_sideeffect_in[1];
    end
  end
  always @(posedge io_lsu_bus_buf_c1_clk or posedge reset) begin
    if (reset) begin
      _T_4321 <= 1'h0;
    end else if (buf_wr_en_0) begin
      _T_4321 <= buf_sideeffect_in[0];
    end
  end
  always @(posedge io_lsu_bus_obuf_c1_clk or posedge reset) begin
    if (reset) begin
      obuf_sideeffect <= 1'h0;
    end else if (obuf_wr_en) begin
      if (ibuf_buf_byp) begin
        obuf_sideeffect <= io_is_sideeffects_r;
      end else begin
        obuf_sideeffect <= _T_1051;
      end
    end
  end
  always @(posedge io_lsu_bus_buf_c1_clk or posedge reset) begin
    if (reset) begin
      buf_dual_3 <= 1'h0;
    end else if (buf_wr_en_3) begin
      buf_dual_3 <= buf_dual_in[3];
    end
  end
  always @(posedge io_lsu_bus_buf_c1_clk or posedge reset) begin
    if (reset) begin
      buf_dual_2 <= 1'h0;
    end else if (buf_wr_en_2) begin
      buf_dual_2 <= buf_dual_in[2];
    end
  end
  always @(posedge io_lsu_bus_buf_c1_clk or posedge reset) begin
    if (reset) begin
      buf_dual_1 <= 1'h0;
    end else if (buf_wr_en_1) begin
      buf_dual_1 <= buf_dual_in[1];
    end
  end
  always @(posedge io_lsu_bus_buf_c1_clk or posedge reset) begin
    if (reset) begin
      buf_dual_0 <= 1'h0;
    end else if (buf_wr_en_0) begin
      buf_dual_0 <= buf_dual_in[0];
    end
  end
  always @(posedge io_lsu_bus_buf_c1_clk or posedge reset) begin
    if (reset) begin
      buf_samedw_3 <= 1'h0;
    end else if (buf_wr_en_3) begin
      buf_samedw_3 <= buf_samedw_in[3];
    end
  end
  always @(posedge io_lsu_bus_buf_c1_clk or posedge reset) begin
    if (reset) begin
      buf_samedw_2 <= 1'h0;
    end else if (buf_wr_en_2) begin
      buf_samedw_2 <= buf_samedw_in[2];
    end
  end
  always @(posedge io_lsu_bus_buf_c1_clk or posedge reset) begin
    if (reset) begin
      buf_samedw_1 <= 1'h0;
    end else if (buf_wr_en_1) begin
      buf_samedw_1 <= buf_samedw_in[1];
    end
  end
  always @(posedge io_lsu_bus_buf_c1_clk or posedge reset) begin
    if (reset) begin
      buf_samedw_0 <= 1'h0;
    end else if (buf_wr_en_0) begin
      buf_samedw_0 <= buf_samedw_in[0];
    end
  end
  always @(posedge io_lsu_bus_obuf_c1_clk or posedge reset) begin
    if (reset) begin
      obuf_write <= 1'h0;
    end else if (obuf_wr_en) begin
      if (ibuf_buf_byp) begin
        obuf_write <= io_lsu_pkt_r_bits_store;
      end else begin
        obuf_write <= _T_1202;
      end
    end
  end
  always @(posedge io_lsu_free_c2_clk or posedge reset) begin
    if (reset) begin
      obuf_nosend <= 1'h0;
    end else if (obuf_wr_en) begin
      obuf_nosend <= obuf_nosend_in;
    end
  end
  always @(posedge rvclkhdr_2_io_l1clk or posedge reset) begin
    if (reset) begin
      obuf_addr <= 32'h0;
    end else if (ibuf_buf_byp) begin
      obuf_addr <= io_lsu_addr_r;
    end else begin
      obuf_addr <= _T_1289;
    end
  end
  always @(posedge io_lsu_bus_buf_c1_clk or posedge reset) begin
    if (reset) begin
      buf_sz_0 <= 2'h0;
    end else if (buf_wr_en_0) begin
      if (ibuf_drainvec_vld[0]) begin
        buf_sz_0 <= ibuf_sz;
      end else begin
        buf_sz_0 <= ibuf_sz_in;
      end
    end
  end
  always @(posedge io_lsu_bus_buf_c1_clk or posedge reset) begin
    if (reset) begin
      buf_sz_1 <= 2'h0;
    end else if (buf_wr_en_1) begin
      if (ibuf_drainvec_vld[1]) begin
        buf_sz_1 <= ibuf_sz;
      end else begin
        buf_sz_1 <= ibuf_sz_in;
      end
    end
  end
  always @(posedge io_lsu_bus_buf_c1_clk or posedge reset) begin
    if (reset) begin
      buf_sz_2 <= 2'h0;
    end else if (buf_wr_en_2) begin
      if (ibuf_drainvec_vld[2]) begin
        buf_sz_2 <= ibuf_sz;
      end else begin
        buf_sz_2 <= ibuf_sz_in;
      end
    end
  end
  always @(posedge io_lsu_bus_buf_c1_clk or posedge reset) begin
    if (reset) begin
      buf_sz_3 <= 2'h0;
    end else if (buf_wr_en_3) begin
      if (ibuf_drainvec_vld[3]) begin
        buf_sz_3 <= ibuf_sz;
      end else begin
        buf_sz_3 <= ibuf_sz_in;
      end
    end
  end
  always @(posedge io_lsu_bus_buf_c1_clk or posedge reset) begin
    if (reset) begin
      buf_dualhi_3 <= 1'h0;
    end else if (buf_wr_en_3) begin
      buf_dualhi_3 <= buf_dualhi_in[3];
    end
  end
  always @(posedge io_lsu_bus_buf_c1_clk or posedge reset) begin
    if (reset) begin
      buf_dualhi_2 <= 1'h0;
    end else if (buf_wr_en_2) begin
      buf_dualhi_2 <= buf_dualhi_in[2];
    end
  end
  always @(posedge io_lsu_bus_buf_c1_clk or posedge reset) begin
    if (reset) begin
      buf_dualhi_1 <= 1'h0;
    end else if (buf_wr_en_1) begin
      buf_dualhi_1 <= buf_dualhi_in[1];
    end
  end
  always @(posedge io_lsu_bus_buf_c1_clk or posedge reset) begin
    if (reset) begin
      buf_dualhi_0 <= 1'h0;
    end else if (buf_wr_en_0) begin
      buf_dualhi_0 <= buf_dualhi_in[0];
    end
  end
  always @(posedge io_lsu_bus_obuf_c1_clk or posedge reset) begin
    if (reset) begin
      obuf_sz <= 2'h0;
    end else if (obuf_wr_en) begin
      if (ibuf_buf_byp) begin
        obuf_sz <= ibuf_sz_in;
      end else begin
        obuf_sz <= _T_1302;
      end
    end
  end
  always @(posedge io_lsu_bus_obuf_c1_clk or posedge reset) begin
    if (reset) begin
      obuf_byteen <= 8'h0;
    end else if (obuf_wr_en) begin
      obuf_byteen <= obuf_byteen_in;
    end
  end
  always @(posedge io_lsu_bus_buf_c1_clk or posedge reset) begin
    if (reset) begin
      buf_rspageQ_0 <= 4'h0;
    end else begin
      buf_rspageQ_0 <= {_T_3173,_T_3162};
    end
  end
  always @(posedge io_lsu_bus_buf_c1_clk or posedge reset) begin
    if (reset) begin
      buf_rspageQ_1 <= 4'h0;
    end else begin
      buf_rspageQ_1 <= {_T_3188,_T_3177};
    end
  end
  always @(posedge io_lsu_bus_buf_c1_clk or posedge reset) begin
    if (reset) begin
      buf_rspageQ_2 <= 4'h0;
    end else begin
      buf_rspageQ_2 <= {_T_3203,_T_3192};
    end
  end
  always @(posedge io_lsu_bus_buf_c1_clk or posedge reset) begin
    if (reset) begin
      buf_rspageQ_3 <= 4'h0;
    end else begin
      buf_rspageQ_3 <= {_T_3218,_T_3207};
    end
  end
  always @(posedge io_lsu_bus_buf_c1_clk or posedge reset) begin
    if (reset) begin
      _T_4307 <= 1'h0;
    end else if (buf_ldfwd_en_3) begin
      if (_T_4107) begin
        _T_4307 <= 1'h0;
      end else if (_T_4130) begin
        _T_4307 <= 1'h0;
      end else begin
        _T_4307 <= _T_4134;
      end
    end
  end
  always @(posedge io_lsu_bus_buf_c1_clk or posedge reset) begin
    if (reset) begin
      _T_4305 <= 1'h0;
    end else if (buf_ldfwd_en_2) begin
      if (_T_3914) begin
        _T_4305 <= 1'h0;
      end else if (_T_3937) begin
        _T_4305 <= 1'h0;
      end else begin
        _T_4305 <= _T_3941;
      end
    end
  end
  always @(posedge io_lsu_bus_buf_c1_clk or posedge reset) begin
    if (reset) begin
      _T_4303 <= 1'h0;
    end else if (buf_ldfwd_en_1) begin
      if (_T_3721) begin
        _T_4303 <= 1'h0;
      end else if (_T_3744) begin
        _T_4303 <= 1'h0;
      end else begin
        _T_4303 <= _T_3748;
      end
    end
  end
  always @(posedge io_lsu_bus_buf_c1_clk or posedge reset) begin
    if (reset) begin
      _T_4301 <= 1'h0;
    end else if (buf_ldfwd_en_0) begin
      if (_T_3528) begin
        _T_4301 <= 1'h0;
      end else if (_T_3551) begin
        _T_4301 <= 1'h0;
      end else begin
        _T_4301 <= _T_3555;
      end
    end
  end
  always @(posedge io_lsu_bus_buf_c1_clk or posedge reset) begin
    if (reset) begin
      buf_dualtag_0 <= 2'h0;
    end else if (buf_wr_en_0) begin
      if (ibuf_drainvec_vld[0]) begin
        buf_dualtag_0 <= ibuf_dualtag;
      end else if (_T_3343) begin
        buf_dualtag_0 <= WrPtr0_r;
      end else begin
        buf_dualtag_0 <= WrPtr1_r;
      end
    end
  end
  always @(posedge io_lsu_bus_buf_c1_clk or posedge reset) begin
    if (reset) begin
      buf_dualtag_1 <= 2'h0;
    end else if (buf_wr_en_1) begin
      if (ibuf_drainvec_vld[1]) begin
        buf_dualtag_1 <= ibuf_dualtag;
      end else if (_T_3352) begin
        buf_dualtag_1 <= WrPtr0_r;
      end else begin
        buf_dualtag_1 <= WrPtr1_r;
      end
    end
  end
  always @(posedge io_lsu_bus_buf_c1_clk or posedge reset) begin
    if (reset) begin
      buf_dualtag_2 <= 2'h0;
    end else if (buf_wr_en_2) begin
      if (ibuf_drainvec_vld[2]) begin
        buf_dualtag_2 <= ibuf_dualtag;
      end else if (_T_3361) begin
        buf_dualtag_2 <= WrPtr0_r;
      end else begin
        buf_dualtag_2 <= WrPtr1_r;
      end
    end
  end
  always @(posedge io_lsu_bus_buf_c1_clk or posedge reset) begin
    if (reset) begin
      buf_dualtag_3 <= 2'h0;
    end else if (buf_wr_en_3) begin
      if (ibuf_drainvec_vld[3]) begin
        buf_dualtag_3 <= ibuf_dualtag;
      end else if (_T_3370) begin
        buf_dualtag_3 <= WrPtr0_r;
      end else begin
        buf_dualtag_3 <= WrPtr1_r;
      end
    end
  end
  always @(posedge io_lsu_bus_buf_c1_clk or posedge reset) begin
    if (reset) begin
      _T_4336 <= 1'h0;
    end else if (buf_wr_en_0) begin
      _T_4336 <= buf_unsign_in[0];
    end
  end
  always @(posedge io_lsu_bus_buf_c1_clk or posedge reset) begin
    if (reset) begin
      _T_4339 <= 1'h0;
    end else if (buf_wr_en_1) begin
      _T_4339 <= buf_unsign_in[1];
    end
  end
  always @(posedge io_lsu_bus_buf_c1_clk or posedge reset) begin
    if (reset) begin
      _T_4342 <= 1'h0;
    end else if (buf_wr_en_2) begin
      _T_4342 <= buf_unsign_in[2];
    end
  end
  always @(posedge io_lsu_bus_buf_c1_clk or posedge reset) begin
    if (reset) begin
      _T_4345 <= 1'h0;
    end else if (buf_wr_en_3) begin
      _T_4345 <= buf_unsign_in[3];
    end
  end
  always @(posedge io_lsu_bus_buf_c1_clk or posedge reset) begin
    if (reset) begin
      _T_4411 <= 1'h0;
    end else begin
      _T_4411 <= buf_error[3] & _T_4409;
    end
  end
  always @(posedge io_lsu_bus_buf_c1_clk or posedge reset) begin
    if (reset) begin
      _T_4406 <= 1'h0;
    end else begin
      _T_4406 <= buf_error[2] & _T_4404;
    end
  end
  always @(posedge io_lsu_bus_buf_c1_clk or posedge reset) begin
    if (reset) begin
      _T_4401 <= 1'h0;
    end else begin
      _T_4401 <= buf_error[1] & _T_4399;
    end
  end
  always @(posedge io_lsu_bus_buf_c1_clk or posedge reset) begin
    if (reset) begin
      _T_4396 <= 1'h0;
    end else begin
      _T_4396 <= buf_error[0] & _T_4394;
    end
  end
  always @(posedge io_lsu_c2_r_clk or posedge reset) begin
    if (reset) begin
      lsu_nonblock_load_valid_r <= 1'h0;
    end else begin
      lsu_nonblock_load_valid_r <= io_dctl_busbuff_lsu_nonblock_load_valid_m;
    end
  end
  always @(posedge io_lsu_c2_r_clk or posedge reset) begin
    if (reset) begin
      _T_4987 <= 1'h0;
    end else begin
      _T_4987 <= _T_4984 & _T_4518;
    end
  end
endmodule
module lsu_bus_intf(
  input         clock,
  input         reset,
  input         io_scan_mode,
  output        io_tlu_busbuff_lsu_pmu_bus_misaligned,
  output        io_tlu_busbuff_lsu_pmu_bus_error,
  output        io_tlu_busbuff_lsu_pmu_bus_busy,
  input         io_tlu_busbuff_dec_tlu_external_ldfwd_disable,
  input         io_tlu_busbuff_dec_tlu_wb_coalescing_disable,
  input         io_tlu_busbuff_dec_tlu_sideeffect_posted_disable,
  output        io_tlu_busbuff_lsu_imprecise_error_load_any,
  output        io_tlu_busbuff_lsu_imprecise_error_store_any,
  output [31:0] io_tlu_busbuff_lsu_imprecise_error_addr_any,
  input         io_lsu_c1_m_clk,
  input         io_lsu_c1_r_clk,
  input         io_lsu_c2_r_clk,
  input         io_lsu_bus_ibuf_c1_clk,
  input         io_lsu_bus_obuf_c1_clk,
  input         io_lsu_bus_buf_c1_clk,
  input         io_lsu_free_c2_clk,
  input         io_free_clk,
  input         io_lsu_busm_clk,
  output        io_axi_aw_valid,
  output [31:0] io_axi_aw_bits_addr,
  output [2:0]  io_axi_aw_bits_size,
  output        io_axi_w_valid,
  output [7:0]  io_axi_w_bits_strb,
  output        io_axi_ar_valid,
  output [31:0] io_axi_ar_bits_addr,
  output [2:0]  io_axi_ar_bits_size,
  input         io_dec_lsu_valid_raw_d,
  input         io_lsu_busreq_m,
  input         io_lsu_pkt_m_valid,
  input         io_lsu_pkt_m_bits_by,
  input         io_lsu_pkt_m_bits_half,
  input         io_lsu_pkt_m_bits_word,
  input         io_lsu_pkt_m_bits_load,
  input         io_lsu_pkt_r_valid,
  input         io_lsu_pkt_r_bits_by,
  input         io_lsu_pkt_r_bits_half,
  input         io_lsu_pkt_r_bits_word,
  input         io_lsu_pkt_r_bits_load,
  input         io_lsu_pkt_r_bits_store,
  input         io_lsu_pkt_r_bits_unsign,
  input  [31:0] io_lsu_addr_d,
  input  [31:0] io_lsu_addr_m,
  input  [31:0] io_lsu_addr_r,
  input  [31:0] io_end_addr_d,
  input  [31:0] io_end_addr_m,
  input  [31:0] io_end_addr_r,
  input  [31:0] io_store_data_r,
  input         io_dec_tlu_force_halt,
  input         io_lsu_commit_r,
  input         io_is_sideeffects_m,
  input         io_flush_m_up,
  input         io_flush_r,
  output        io_lsu_busreq_r,
  output        io_lsu_bus_buffer_pend_any,
  output        io_lsu_bus_buffer_full_any,
  output        io_lsu_bus_buffer_empty_any,
  output [31:0] io_bus_read_data_m,
  output        io_dctl_busbuff_lsu_nonblock_load_valid_m,
  output [1:0]  io_dctl_busbuff_lsu_nonblock_load_tag_m,
  output        io_dctl_busbuff_lsu_nonblock_load_inv_r,
  output [1:0]  io_dctl_busbuff_lsu_nonblock_load_inv_tag_r,
  output        io_dctl_busbuff_lsu_nonblock_load_data_valid,
  output        io_dctl_busbuff_lsu_nonblock_load_data_error,
  output [1:0]  io_dctl_busbuff_lsu_nonblock_load_data_tag,
  output [31:0] io_dctl_busbuff_lsu_nonblock_load_data,
  input         io_lsu_bus_clk_en
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  wire  bus_buffer_clock; // @[lsu_bus_intf.scala 101:39]
  wire  bus_buffer_reset; // @[lsu_bus_intf.scala 101:39]
  wire  bus_buffer_io_scan_mode; // @[lsu_bus_intf.scala 101:39]
  wire  bus_buffer_io_tlu_busbuff_lsu_pmu_bus_misaligned; // @[lsu_bus_intf.scala 101:39]
  wire  bus_buffer_io_tlu_busbuff_lsu_pmu_bus_error; // @[lsu_bus_intf.scala 101:39]
  wire  bus_buffer_io_tlu_busbuff_lsu_pmu_bus_busy; // @[lsu_bus_intf.scala 101:39]
  wire  bus_buffer_io_tlu_busbuff_dec_tlu_external_ldfwd_disable; // @[lsu_bus_intf.scala 101:39]
  wire  bus_buffer_io_tlu_busbuff_dec_tlu_wb_coalescing_disable; // @[lsu_bus_intf.scala 101:39]
  wire  bus_buffer_io_tlu_busbuff_dec_tlu_sideeffect_posted_disable; // @[lsu_bus_intf.scala 101:39]
  wire  bus_buffer_io_tlu_busbuff_lsu_imprecise_error_load_any; // @[lsu_bus_intf.scala 101:39]
  wire  bus_buffer_io_tlu_busbuff_lsu_imprecise_error_store_any; // @[lsu_bus_intf.scala 101:39]
  wire [31:0] bus_buffer_io_tlu_busbuff_lsu_imprecise_error_addr_any; // @[lsu_bus_intf.scala 101:39]
  wire  bus_buffer_io_dctl_busbuff_lsu_nonblock_load_valid_m; // @[lsu_bus_intf.scala 101:39]
  wire [1:0] bus_buffer_io_dctl_busbuff_lsu_nonblock_load_tag_m; // @[lsu_bus_intf.scala 101:39]
  wire  bus_buffer_io_dctl_busbuff_lsu_nonblock_load_inv_r; // @[lsu_bus_intf.scala 101:39]
  wire [1:0] bus_buffer_io_dctl_busbuff_lsu_nonblock_load_inv_tag_r; // @[lsu_bus_intf.scala 101:39]
  wire  bus_buffer_io_dctl_busbuff_lsu_nonblock_load_data_valid; // @[lsu_bus_intf.scala 101:39]
  wire  bus_buffer_io_dctl_busbuff_lsu_nonblock_load_data_error; // @[lsu_bus_intf.scala 101:39]
  wire [1:0] bus_buffer_io_dctl_busbuff_lsu_nonblock_load_data_tag; // @[lsu_bus_intf.scala 101:39]
  wire [31:0] bus_buffer_io_dctl_busbuff_lsu_nonblock_load_data; // @[lsu_bus_intf.scala 101:39]
  wire  bus_buffer_io_dec_tlu_force_halt; // @[lsu_bus_intf.scala 101:39]
  wire  bus_buffer_io_lsu_c2_r_clk; // @[lsu_bus_intf.scala 101:39]
  wire  bus_buffer_io_lsu_bus_ibuf_c1_clk; // @[lsu_bus_intf.scala 101:39]
  wire  bus_buffer_io_lsu_bus_obuf_c1_clk; // @[lsu_bus_intf.scala 101:39]
  wire  bus_buffer_io_lsu_bus_buf_c1_clk; // @[lsu_bus_intf.scala 101:39]
  wire  bus_buffer_io_lsu_free_c2_clk; // @[lsu_bus_intf.scala 101:39]
  wire  bus_buffer_io_lsu_busm_clk; // @[lsu_bus_intf.scala 101:39]
  wire  bus_buffer_io_dec_lsu_valid_raw_d; // @[lsu_bus_intf.scala 101:39]
  wire  bus_buffer_io_lsu_pkt_m_valid; // @[lsu_bus_intf.scala 101:39]
  wire  bus_buffer_io_lsu_pkt_m_bits_load; // @[lsu_bus_intf.scala 101:39]
  wire  bus_buffer_io_lsu_pkt_r_bits_by; // @[lsu_bus_intf.scala 101:39]
  wire  bus_buffer_io_lsu_pkt_r_bits_half; // @[lsu_bus_intf.scala 101:39]
  wire  bus_buffer_io_lsu_pkt_r_bits_word; // @[lsu_bus_intf.scala 101:39]
  wire  bus_buffer_io_lsu_pkt_r_bits_load; // @[lsu_bus_intf.scala 101:39]
  wire  bus_buffer_io_lsu_pkt_r_bits_store; // @[lsu_bus_intf.scala 101:39]
  wire  bus_buffer_io_lsu_pkt_r_bits_unsign; // @[lsu_bus_intf.scala 101:39]
  wire [31:0] bus_buffer_io_lsu_addr_m; // @[lsu_bus_intf.scala 101:39]
  wire [31:0] bus_buffer_io_end_addr_m; // @[lsu_bus_intf.scala 101:39]
  wire [31:0] bus_buffer_io_lsu_addr_r; // @[lsu_bus_intf.scala 101:39]
  wire [31:0] bus_buffer_io_end_addr_r; // @[lsu_bus_intf.scala 101:39]
  wire [31:0] bus_buffer_io_store_data_r; // @[lsu_bus_intf.scala 101:39]
  wire  bus_buffer_io_no_word_merge_r; // @[lsu_bus_intf.scala 101:39]
  wire  bus_buffer_io_no_dword_merge_r; // @[lsu_bus_intf.scala 101:39]
  wire  bus_buffer_io_lsu_busreq_m; // @[lsu_bus_intf.scala 101:39]
  wire  bus_buffer_io_ld_full_hit_m; // @[lsu_bus_intf.scala 101:39]
  wire  bus_buffer_io_flush_m_up; // @[lsu_bus_intf.scala 101:39]
  wire  bus_buffer_io_flush_r; // @[lsu_bus_intf.scala 101:39]
  wire  bus_buffer_io_lsu_commit_r; // @[lsu_bus_intf.scala 101:39]
  wire  bus_buffer_io_is_sideeffects_r; // @[lsu_bus_intf.scala 101:39]
  wire  bus_buffer_io_ldst_dual_d; // @[lsu_bus_intf.scala 101:39]
  wire  bus_buffer_io_ldst_dual_m; // @[lsu_bus_intf.scala 101:39]
  wire  bus_buffer_io_ldst_dual_r; // @[lsu_bus_intf.scala 101:39]
  wire [7:0] bus_buffer_io_ldst_byteen_ext_m; // @[lsu_bus_intf.scala 101:39]
  wire  bus_buffer_io_lsu_axi_aw_valid; // @[lsu_bus_intf.scala 101:39]
  wire [31:0] bus_buffer_io_lsu_axi_aw_bits_addr; // @[lsu_bus_intf.scala 101:39]
  wire [2:0] bus_buffer_io_lsu_axi_aw_bits_size; // @[lsu_bus_intf.scala 101:39]
  wire  bus_buffer_io_lsu_axi_w_valid; // @[lsu_bus_intf.scala 101:39]
  wire [7:0] bus_buffer_io_lsu_axi_w_bits_strb; // @[lsu_bus_intf.scala 101:39]
  wire  bus_buffer_io_lsu_axi_ar_valid; // @[lsu_bus_intf.scala 101:39]
  wire [31:0] bus_buffer_io_lsu_axi_ar_bits_addr; // @[lsu_bus_intf.scala 101:39]
  wire [2:0] bus_buffer_io_lsu_axi_ar_bits_size; // @[lsu_bus_intf.scala 101:39]
  wire  bus_buffer_io_lsu_bus_clk_en; // @[lsu_bus_intf.scala 101:39]
  wire  bus_buffer_io_lsu_bus_clk_en_q; // @[lsu_bus_intf.scala 101:39]
  wire  bus_buffer_io_lsu_busreq_r; // @[lsu_bus_intf.scala 101:39]
  wire  bus_buffer_io_lsu_bus_buffer_pend_any; // @[lsu_bus_intf.scala 101:39]
  wire  bus_buffer_io_lsu_bus_buffer_full_any; // @[lsu_bus_intf.scala 101:39]
  wire  bus_buffer_io_lsu_bus_buffer_empty_any; // @[lsu_bus_intf.scala 101:39]
  wire [3:0] bus_buffer_io_ld_byte_hit_buf_lo; // @[lsu_bus_intf.scala 101:39]
  wire [3:0] bus_buffer_io_ld_byte_hit_buf_hi; // @[lsu_bus_intf.scala 101:39]
  wire [31:0] bus_buffer_io_ld_fwddata_buf_lo; // @[lsu_bus_intf.scala 101:39]
  wire [31:0] bus_buffer_io_ld_fwddata_buf_hi; // @[lsu_bus_intf.scala 101:39]
  wire [3:0] _T_3 = io_lsu_pkt_m_bits_word ? 4'hf : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_4 = io_lsu_pkt_m_bits_half ? 4'h3 : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_5 = io_lsu_pkt_m_bits_by ? 4'h1 : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_6 = _T_3 | _T_4; // @[Mux.scala 27:72]
  wire [3:0] ldst_byteen_m = _T_6 | _T_5; // @[Mux.scala 27:72]
  wire  addr_match_dw_lo_r_m = io_lsu_addr_r[31:3] == io_lsu_addr_m[31:3]; // @[lsu_bus_intf.scala 155:51]
  wire  _T_17 = io_lsu_addr_r[2] ^ io_lsu_addr_m[2]; // @[lsu_bus_intf.scala 156:71]
  wire  _T_18 = ~_T_17; // @[lsu_bus_intf.scala 156:53]
  wire  addr_match_word_lo_r_m = addr_match_dw_lo_r_m & _T_18; // @[lsu_bus_intf.scala 156:51]
  reg  ldst_dual_r; // @[lsu_bus_intf.scala 201:33]
  wire  _T_20 = ~ldst_dual_r; // @[lsu_bus_intf.scala 157:48]
  wire  _T_21 = io_lsu_busreq_r & _T_20; // @[lsu_bus_intf.scala 157:46]
  wire  _T_22 = _T_21 & io_lsu_busreq_m; // @[lsu_bus_intf.scala 157:61]
  wire  _T_23 = ~addr_match_word_lo_r_m; // @[lsu_bus_intf.scala 157:107]
  wire  _T_24 = io_lsu_pkt_m_bits_load | _T_23; // @[lsu_bus_intf.scala 157:105]
  wire  _T_29 = ~addr_match_dw_lo_r_m; // @[lsu_bus_intf.scala 158:107]
  wire  _T_30 = io_lsu_pkt_m_bits_load | _T_29; // @[lsu_bus_intf.scala 158:105]
  wire [6:0] _GEN_0 = {{3'd0}, ldst_byteen_m}; // @[lsu_bus_intf.scala 160:49]
  wire [6:0] _T_34 = _GEN_0 << io_lsu_addr_m[1:0]; // @[lsu_bus_intf.scala 160:49]
  reg [3:0] ldst_byteen_r; // @[lsu_bus_intf.scala 203:33]
  wire [6:0] _GEN_1 = {{3'd0}, ldst_byteen_r}; // @[lsu_bus_intf.scala 161:49]
  wire [6:0] _T_37 = _GEN_1 << io_lsu_addr_r[1:0]; // @[lsu_bus_intf.scala 161:49]
  wire [4:0] _T_40 = {io_lsu_addr_r[1:0],3'h0}; // @[Cat.scala 29:58]
  wire [62:0] _GEN_2 = {{31'd0}, io_store_data_r}; // @[lsu_bus_intf.scala 162:52]
  wire [62:0] _T_41 = _GEN_2 << _T_40; // @[lsu_bus_intf.scala 162:52]
  wire [7:0] ldst_byteen_ext_m = {{1'd0}, _T_34}; // @[lsu_bus_intf.scala 160:27]
  wire [3:0] ldst_byteen_hi_m = ldst_byteen_ext_m[7:4]; // @[lsu_bus_intf.scala 163:47]
  wire [3:0] ldst_byteen_lo_m = ldst_byteen_ext_m[3:0]; // @[lsu_bus_intf.scala 164:47]
  wire [7:0] ldst_byteen_ext_r = {{1'd0}, _T_37}; // @[lsu_bus_intf.scala 161:27]
  wire [3:0] ldst_byteen_hi_r = ldst_byteen_ext_r[7:4]; // @[lsu_bus_intf.scala 165:47]
  wire [3:0] ldst_byteen_lo_r = ldst_byteen_ext_r[3:0]; // @[lsu_bus_intf.scala 166:47]
  wire [63:0] store_data_ext_r = {{1'd0}, _T_41}; // @[lsu_bus_intf.scala 162:27]
  wire [31:0] store_data_hi_r = store_data_ext_r[63:32]; // @[lsu_bus_intf.scala 168:46]
  wire [31:0] store_data_lo_r = store_data_ext_r[31:0]; // @[lsu_bus_intf.scala 169:46]
  wire  _T_50 = io_lsu_addr_m[31:2] == io_lsu_addr_r[31:2]; // @[lsu_bus_intf.scala 170:51]
  wire  _T_51 = _T_50 & io_lsu_pkt_r_valid; // @[lsu_bus_intf.scala 170:76]
  wire  _T_52 = _T_51 & io_lsu_pkt_r_bits_store; // @[lsu_bus_intf.scala 170:97]
  wire  ld_addr_rhit_lo_lo = _T_52 & io_lsu_busreq_m; // @[lsu_bus_intf.scala 170:123]
  wire  _T_56 = io_end_addr_m[31:2] == io_lsu_addr_r[31:2]; // @[lsu_bus_intf.scala 171:51]
  wire  _T_57 = _T_56 & io_lsu_pkt_r_valid; // @[lsu_bus_intf.scala 171:76]
  wire  _T_58 = _T_57 & io_lsu_pkt_r_bits_store; // @[lsu_bus_intf.scala 171:97]
  wire  ld_addr_rhit_lo_hi = _T_58 & io_lsu_busreq_m; // @[lsu_bus_intf.scala 171:123]
  wire  _T_62 = io_lsu_addr_m[31:2] == io_end_addr_r[31:2]; // @[lsu_bus_intf.scala 172:51]
  wire  _T_63 = _T_62 & io_lsu_pkt_r_valid; // @[lsu_bus_intf.scala 172:76]
  wire  _T_64 = _T_63 & io_lsu_pkt_r_bits_store; // @[lsu_bus_intf.scala 172:97]
  wire  ld_addr_rhit_hi_lo = _T_64 & io_lsu_busreq_m; // @[lsu_bus_intf.scala 172:123]
  wire  _T_68 = io_end_addr_m[31:2] == io_end_addr_r[31:2]; // @[lsu_bus_intf.scala 173:51]
  wire  _T_69 = _T_68 & io_lsu_pkt_r_valid; // @[lsu_bus_intf.scala 173:76]
  wire  _T_70 = _T_69 & io_lsu_pkt_r_bits_store; // @[lsu_bus_intf.scala 173:97]
  wire  ld_addr_rhit_hi_hi = _T_70 & io_lsu_busreq_m; // @[lsu_bus_intf.scala 173:123]
  wire  _T_73 = ld_addr_rhit_lo_lo & ldst_byteen_lo_r[0]; // @[lsu_bus_intf.scala 175:70]
  wire  _T_75 = _T_73 & ldst_byteen_lo_m[0]; // @[lsu_bus_intf.scala 175:92]
  wire  _T_77 = ld_addr_rhit_lo_lo & ldst_byteen_lo_r[1]; // @[lsu_bus_intf.scala 175:70]
  wire  _T_79 = _T_77 & ldst_byteen_lo_m[1]; // @[lsu_bus_intf.scala 175:92]
  wire  _T_81 = ld_addr_rhit_lo_lo & ldst_byteen_lo_r[2]; // @[lsu_bus_intf.scala 175:70]
  wire  _T_83 = _T_81 & ldst_byteen_lo_m[2]; // @[lsu_bus_intf.scala 175:92]
  wire  _T_85 = ld_addr_rhit_lo_lo & ldst_byteen_lo_r[3]; // @[lsu_bus_intf.scala 175:70]
  wire  _T_87 = _T_85 & ldst_byteen_lo_m[3]; // @[lsu_bus_intf.scala 175:92]
  wire [3:0] ld_byte_rhit_lo_lo = {_T_87,_T_83,_T_79,_T_75}; // @[Cat.scala 29:58]
  wire  _T_92 = ld_addr_rhit_lo_hi & ldst_byteen_lo_r[0]; // @[lsu_bus_intf.scala 176:70]
  wire  _T_94 = _T_92 & ldst_byteen_hi_m[0]; // @[lsu_bus_intf.scala 176:92]
  wire  _T_96 = ld_addr_rhit_lo_hi & ldst_byteen_lo_r[1]; // @[lsu_bus_intf.scala 176:70]
  wire  _T_98 = _T_96 & ldst_byteen_hi_m[1]; // @[lsu_bus_intf.scala 176:92]
  wire  _T_100 = ld_addr_rhit_lo_hi & ldst_byteen_lo_r[2]; // @[lsu_bus_intf.scala 176:70]
  wire  _T_102 = _T_100 & ldst_byteen_hi_m[2]; // @[lsu_bus_intf.scala 176:92]
  wire  _T_104 = ld_addr_rhit_lo_hi & ldst_byteen_lo_r[3]; // @[lsu_bus_intf.scala 176:70]
  wire  _T_106 = _T_104 & ldst_byteen_hi_m[3]; // @[lsu_bus_intf.scala 176:92]
  wire [3:0] ld_byte_rhit_lo_hi = {_T_106,_T_102,_T_98,_T_94}; // @[Cat.scala 29:58]
  wire  _T_111 = ld_addr_rhit_hi_lo & ldst_byteen_hi_r[0]; // @[lsu_bus_intf.scala 177:70]
  wire  _T_113 = _T_111 & ldst_byteen_lo_m[0]; // @[lsu_bus_intf.scala 177:92]
  wire  _T_115 = ld_addr_rhit_hi_lo & ldst_byteen_hi_r[1]; // @[lsu_bus_intf.scala 177:70]
  wire  _T_117 = _T_115 & ldst_byteen_lo_m[1]; // @[lsu_bus_intf.scala 177:92]
  wire  _T_119 = ld_addr_rhit_hi_lo & ldst_byteen_hi_r[2]; // @[lsu_bus_intf.scala 177:70]
  wire  _T_121 = _T_119 & ldst_byteen_lo_m[2]; // @[lsu_bus_intf.scala 177:92]
  wire  _T_123 = ld_addr_rhit_hi_lo & ldst_byteen_hi_r[3]; // @[lsu_bus_intf.scala 177:70]
  wire  _T_125 = _T_123 & ldst_byteen_lo_m[3]; // @[lsu_bus_intf.scala 177:92]
  wire [3:0] ld_byte_rhit_hi_lo = {_T_125,_T_121,_T_117,_T_113}; // @[Cat.scala 29:58]
  wire  _T_130 = ld_addr_rhit_hi_hi & ldst_byteen_hi_r[0]; // @[lsu_bus_intf.scala 178:70]
  wire  _T_132 = _T_130 & ldst_byteen_hi_m[0]; // @[lsu_bus_intf.scala 178:92]
  wire  _T_134 = ld_addr_rhit_hi_hi & ldst_byteen_hi_r[1]; // @[lsu_bus_intf.scala 178:70]
  wire  _T_136 = _T_134 & ldst_byteen_hi_m[1]; // @[lsu_bus_intf.scala 178:92]
  wire  _T_138 = ld_addr_rhit_hi_hi & ldst_byteen_hi_r[2]; // @[lsu_bus_intf.scala 178:70]
  wire  _T_140 = _T_138 & ldst_byteen_hi_m[2]; // @[lsu_bus_intf.scala 178:92]
  wire  _T_142 = ld_addr_rhit_hi_hi & ldst_byteen_hi_r[3]; // @[lsu_bus_intf.scala 178:70]
  wire  _T_144 = _T_142 & ldst_byteen_hi_m[3]; // @[lsu_bus_intf.scala 178:92]
  wire [3:0] ld_byte_rhit_hi_hi = {_T_144,_T_140,_T_136,_T_132}; // @[Cat.scala 29:58]
  wire  _T_150 = ld_byte_rhit_lo_lo[0] | ld_byte_rhit_hi_lo[0]; // @[lsu_bus_intf.scala 180:73]
  wire [3:0] ld_byte_hit_buf_lo = bus_buffer_io_ld_byte_hit_buf_lo; // @[lsu_bus_intf.scala 138:38]
  wire  _T_152 = _T_150 | ld_byte_hit_buf_lo[0]; // @[lsu_bus_intf.scala 180:97]
  wire  _T_155 = ld_byte_rhit_lo_lo[1] | ld_byte_rhit_hi_lo[1]; // @[lsu_bus_intf.scala 180:73]
  wire  _T_157 = _T_155 | ld_byte_hit_buf_lo[1]; // @[lsu_bus_intf.scala 180:97]
  wire  _T_160 = ld_byte_rhit_lo_lo[2] | ld_byte_rhit_hi_lo[2]; // @[lsu_bus_intf.scala 180:73]
  wire  _T_162 = _T_160 | ld_byte_hit_buf_lo[2]; // @[lsu_bus_intf.scala 180:97]
  wire  _T_165 = ld_byte_rhit_lo_lo[3] | ld_byte_rhit_hi_lo[3]; // @[lsu_bus_intf.scala 180:73]
  wire  _T_167 = _T_165 | ld_byte_hit_buf_lo[3]; // @[lsu_bus_intf.scala 180:97]
  wire [3:0] ld_byte_hit_lo = {_T_167,_T_162,_T_157,_T_152}; // @[Cat.scala 29:58]
  wire  _T_173 = ld_byte_rhit_lo_hi[0] | ld_byte_rhit_hi_hi[0]; // @[lsu_bus_intf.scala 181:73]
  wire [3:0] ld_byte_hit_buf_hi = bus_buffer_io_ld_byte_hit_buf_hi; // @[lsu_bus_intf.scala 139:38]
  wire  _T_175 = _T_173 | ld_byte_hit_buf_hi[0]; // @[lsu_bus_intf.scala 181:97]
  wire  _T_178 = ld_byte_rhit_lo_hi[1] | ld_byte_rhit_hi_hi[1]; // @[lsu_bus_intf.scala 181:73]
  wire  _T_180 = _T_178 | ld_byte_hit_buf_hi[1]; // @[lsu_bus_intf.scala 181:97]
  wire  _T_183 = ld_byte_rhit_lo_hi[2] | ld_byte_rhit_hi_hi[2]; // @[lsu_bus_intf.scala 181:73]
  wire  _T_185 = _T_183 | ld_byte_hit_buf_hi[2]; // @[lsu_bus_intf.scala 181:97]
  wire  _T_188 = ld_byte_rhit_lo_hi[3] | ld_byte_rhit_hi_hi[3]; // @[lsu_bus_intf.scala 181:73]
  wire  _T_190 = _T_188 | ld_byte_hit_buf_hi[3]; // @[lsu_bus_intf.scala 181:97]
  wire [3:0] ld_byte_hit_hi = {_T_190,_T_185,_T_180,_T_175}; // @[Cat.scala 29:58]
  wire [3:0] ld_byte_rhit_lo = {_T_165,_T_160,_T_155,_T_150}; // @[Cat.scala 29:58]
  wire [3:0] ld_byte_rhit_hi = {_T_188,_T_183,_T_178,_T_173}; // @[Cat.scala 29:58]
  wire [7:0] _T_228 = ld_byte_rhit_lo_lo[0] ? store_data_lo_r[7:0] : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_229 = ld_byte_rhit_hi_lo[0] ? store_data_hi_r[7:0] : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_230 = _T_228 | _T_229; // @[Mux.scala 27:72]
  wire [7:0] _T_236 = ld_byte_rhit_lo_lo[1] ? store_data_lo_r[15:8] : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_237 = ld_byte_rhit_hi_lo[1] ? store_data_hi_r[15:8] : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_238 = _T_236 | _T_237; // @[Mux.scala 27:72]
  wire [7:0] _T_244 = ld_byte_rhit_lo_lo[2] ? store_data_lo_r[23:16] : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_245 = ld_byte_rhit_hi_lo[2] ? store_data_hi_r[23:16] : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_246 = _T_244 | _T_245; // @[Mux.scala 27:72]
  wire [7:0] _T_252 = ld_byte_rhit_lo_lo[3] ? store_data_lo_r[31:24] : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_253 = ld_byte_rhit_hi_lo[3] ? store_data_hi_r[31:24] : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_254 = _T_252 | _T_253; // @[Mux.scala 27:72]
  wire [31:0] ld_fwddata_rpipe_lo = {_T_254,_T_246,_T_238,_T_230}; // @[Cat.scala 29:58]
  wire [7:0] _T_263 = ld_byte_rhit_lo_hi[0] ? store_data_lo_r[7:0] : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_264 = ld_byte_rhit_hi_hi[0] ? store_data_hi_r[7:0] : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_265 = _T_263 | _T_264; // @[Mux.scala 27:72]
  wire [7:0] _T_271 = ld_byte_rhit_lo_hi[1] ? store_data_lo_r[15:8] : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_272 = ld_byte_rhit_hi_hi[1] ? store_data_hi_r[15:8] : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_273 = _T_271 | _T_272; // @[Mux.scala 27:72]
  wire [7:0] _T_279 = ld_byte_rhit_lo_hi[2] ? store_data_lo_r[23:16] : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_280 = ld_byte_rhit_hi_hi[2] ? store_data_hi_r[23:16] : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_281 = _T_279 | _T_280; // @[Mux.scala 27:72]
  wire [7:0] _T_287 = ld_byte_rhit_lo_hi[3] ? store_data_lo_r[31:24] : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_288 = ld_byte_rhit_hi_hi[3] ? store_data_hi_r[31:24] : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_289 = _T_287 | _T_288; // @[Mux.scala 27:72]
  wire [31:0] ld_fwddata_rpipe_hi = {_T_289,_T_281,_T_273,_T_265}; // @[Cat.scala 29:58]
  wire [31:0] ld_fwddata_buf_lo = bus_buffer_io_ld_fwddata_buf_lo; // @[lsu_bus_intf.scala 140:38]
  wire [7:0] _T_297 = ld_byte_rhit_lo[0] ? ld_fwddata_rpipe_lo[7:0] : ld_fwddata_buf_lo[7:0]; // @[lsu_bus_intf.scala 186:54]
  wire [7:0] _T_301 = ld_byte_rhit_lo[1] ? ld_fwddata_rpipe_lo[15:8] : ld_fwddata_buf_lo[15:8]; // @[lsu_bus_intf.scala 186:54]
  wire [7:0] _T_305 = ld_byte_rhit_lo[2] ? ld_fwddata_rpipe_lo[23:16] : ld_fwddata_buf_lo[23:16]; // @[lsu_bus_intf.scala 186:54]
  wire [7:0] _T_309 = ld_byte_rhit_lo[3] ? ld_fwddata_rpipe_lo[31:24] : ld_fwddata_buf_lo[31:24]; // @[lsu_bus_intf.scala 186:54]
  wire [31:0] _T_312 = {_T_309,_T_305,_T_301,_T_297}; // @[Cat.scala 29:58]
  wire [31:0] ld_fwddata_buf_hi = bus_buffer_io_ld_fwddata_buf_hi; // @[lsu_bus_intf.scala 141:38]
  wire [7:0] _T_316 = ld_byte_rhit_hi[0] ? ld_fwddata_rpipe_hi[7:0] : ld_fwddata_buf_hi[7:0]; // @[lsu_bus_intf.scala 187:54]
  wire [7:0] _T_320 = ld_byte_rhit_hi[1] ? ld_fwddata_rpipe_hi[15:8] : ld_fwddata_buf_hi[15:8]; // @[lsu_bus_intf.scala 187:54]
  wire [7:0] _T_324 = ld_byte_rhit_hi[2] ? ld_fwddata_rpipe_hi[23:16] : ld_fwddata_buf_hi[23:16]; // @[lsu_bus_intf.scala 187:54]
  wire [7:0] _T_328 = ld_byte_rhit_hi[3] ? ld_fwddata_rpipe_hi[31:24] : ld_fwddata_buf_hi[31:24]; // @[lsu_bus_intf.scala 187:54]
  wire [31:0] _T_331 = {_T_328,_T_324,_T_320,_T_316}; // @[Cat.scala 29:58]
  wire  _T_334 = ~ldst_byteen_lo_m[0]; // @[lsu_bus_intf.scala 188:72]
  wire  _T_335 = ld_byte_hit_lo[0] | _T_334; // @[lsu_bus_intf.scala 188:70]
  wire  _T_338 = ~ldst_byteen_lo_m[1]; // @[lsu_bus_intf.scala 188:72]
  wire  _T_339 = ld_byte_hit_lo[1] | _T_338; // @[lsu_bus_intf.scala 188:70]
  wire  _T_342 = ~ldst_byteen_lo_m[2]; // @[lsu_bus_intf.scala 188:72]
  wire  _T_343 = ld_byte_hit_lo[2] | _T_342; // @[lsu_bus_intf.scala 188:70]
  wire  _T_346 = ~ldst_byteen_lo_m[3]; // @[lsu_bus_intf.scala 188:72]
  wire  _T_347 = ld_byte_hit_lo[3] | _T_346; // @[lsu_bus_intf.scala 188:70]
  wire  _T_348 = _T_335 & _T_339; // @[lsu_bus_intf.scala 188:111]
  wire  _T_349 = _T_348 & _T_343; // @[lsu_bus_intf.scala 188:111]
  wire  ld_full_hit_lo_m = _T_349 & _T_347; // @[lsu_bus_intf.scala 188:111]
  wire  _T_353 = ~ldst_byteen_hi_m[0]; // @[lsu_bus_intf.scala 189:72]
  wire  _T_354 = ld_byte_hit_hi[0] | _T_353; // @[lsu_bus_intf.scala 189:70]
  wire  _T_357 = ~ldst_byteen_hi_m[1]; // @[lsu_bus_intf.scala 189:72]
  wire  _T_358 = ld_byte_hit_hi[1] | _T_357; // @[lsu_bus_intf.scala 189:70]
  wire  _T_361 = ~ldst_byteen_hi_m[2]; // @[lsu_bus_intf.scala 189:72]
  wire  _T_362 = ld_byte_hit_hi[2] | _T_361; // @[lsu_bus_intf.scala 189:70]
  wire  _T_365 = ~ldst_byteen_hi_m[3]; // @[lsu_bus_intf.scala 189:72]
  wire  _T_366 = ld_byte_hit_hi[3] | _T_365; // @[lsu_bus_intf.scala 189:70]
  wire  _T_367 = _T_354 & _T_358; // @[lsu_bus_intf.scala 189:111]
  wire  _T_368 = _T_367 & _T_362; // @[lsu_bus_intf.scala 189:111]
  wire  ld_full_hit_hi_m = _T_368 & _T_366; // @[lsu_bus_intf.scala 189:111]
  wire  _T_370 = ld_full_hit_lo_m & ld_full_hit_hi_m; // @[lsu_bus_intf.scala 190:47]
  wire  _T_371 = _T_370 & io_lsu_busreq_m; // @[lsu_bus_intf.scala 190:66]
  wire  _T_372 = _T_371 & io_lsu_pkt_m_bits_load; // @[lsu_bus_intf.scala 190:84]
  wire  _T_373 = ~io_is_sideeffects_m; // @[lsu_bus_intf.scala 190:111]
  wire [63:0] ld_fwddata_hi = {{32'd0}, _T_331}; // @[lsu_bus_intf.scala 187:27]
  wire [63:0] ld_fwddata_lo = {{32'd0}, _T_312}; // @[lsu_bus_intf.scala 186:27]
  wire [63:0] _T_377 = {ld_fwddata_hi[31:0],ld_fwddata_lo[31:0]}; // @[Cat.scala 29:58]
  wire [3:0] _GEN_3 = {{2'd0}, io_lsu_addr_m[1:0]}; // @[lsu_bus_intf.scala 191:83]
  wire [5:0] _T_379 = 4'h8 * _GEN_3; // @[lsu_bus_intf.scala 191:83]
  wire [63:0] ld_fwddata_m = _T_377 >> _T_379; // @[lsu_bus_intf.scala 191:76]
  reg  lsu_bus_clk_en_q; // @[lsu_bus_intf.scala 195:32]
  reg  ldst_dual_m; // @[lsu_bus_intf.scala 198:27]
  reg  is_sideeffects_r; // @[lsu_bus_intf.scala 202:33]
  lsu_bus_buffer bus_buffer ( // @[lsu_bus_intf.scala 101:39]
    .clock(bus_buffer_clock),
    .reset(bus_buffer_reset),
    .io_scan_mode(bus_buffer_io_scan_mode),
    .io_tlu_busbuff_lsu_pmu_bus_misaligned(bus_buffer_io_tlu_busbuff_lsu_pmu_bus_misaligned),
    .io_tlu_busbuff_lsu_pmu_bus_error(bus_buffer_io_tlu_busbuff_lsu_pmu_bus_error),
    .io_tlu_busbuff_lsu_pmu_bus_busy(bus_buffer_io_tlu_busbuff_lsu_pmu_bus_busy),
    .io_tlu_busbuff_dec_tlu_external_ldfwd_disable(bus_buffer_io_tlu_busbuff_dec_tlu_external_ldfwd_disable),
    .io_tlu_busbuff_dec_tlu_wb_coalescing_disable(bus_buffer_io_tlu_busbuff_dec_tlu_wb_coalescing_disable),
    .io_tlu_busbuff_dec_tlu_sideeffect_posted_disable(bus_buffer_io_tlu_busbuff_dec_tlu_sideeffect_posted_disable),
    .io_tlu_busbuff_lsu_imprecise_error_load_any(bus_buffer_io_tlu_busbuff_lsu_imprecise_error_load_any),
    .io_tlu_busbuff_lsu_imprecise_error_store_any(bus_buffer_io_tlu_busbuff_lsu_imprecise_error_store_any),
    .io_tlu_busbuff_lsu_imprecise_error_addr_any(bus_buffer_io_tlu_busbuff_lsu_imprecise_error_addr_any),
    .io_dctl_busbuff_lsu_nonblock_load_valid_m(bus_buffer_io_dctl_busbuff_lsu_nonblock_load_valid_m),
    .io_dctl_busbuff_lsu_nonblock_load_tag_m(bus_buffer_io_dctl_busbuff_lsu_nonblock_load_tag_m),
    .io_dctl_busbuff_lsu_nonblock_load_inv_r(bus_buffer_io_dctl_busbuff_lsu_nonblock_load_inv_r),
    .io_dctl_busbuff_lsu_nonblock_load_inv_tag_r(bus_buffer_io_dctl_busbuff_lsu_nonblock_load_inv_tag_r),
    .io_dctl_busbuff_lsu_nonblock_load_data_valid(bus_buffer_io_dctl_busbuff_lsu_nonblock_load_data_valid),
    .io_dctl_busbuff_lsu_nonblock_load_data_error(bus_buffer_io_dctl_busbuff_lsu_nonblock_load_data_error),
    .io_dctl_busbuff_lsu_nonblock_load_data_tag(bus_buffer_io_dctl_busbuff_lsu_nonblock_load_data_tag),
    .io_dctl_busbuff_lsu_nonblock_load_data(bus_buffer_io_dctl_busbuff_lsu_nonblock_load_data),
    .io_dec_tlu_force_halt(bus_buffer_io_dec_tlu_force_halt),
    .io_lsu_c2_r_clk(bus_buffer_io_lsu_c2_r_clk),
    .io_lsu_bus_ibuf_c1_clk(bus_buffer_io_lsu_bus_ibuf_c1_clk),
    .io_lsu_bus_obuf_c1_clk(bus_buffer_io_lsu_bus_obuf_c1_clk),
    .io_lsu_bus_buf_c1_clk(bus_buffer_io_lsu_bus_buf_c1_clk),
    .io_lsu_free_c2_clk(bus_buffer_io_lsu_free_c2_clk),
    .io_lsu_busm_clk(bus_buffer_io_lsu_busm_clk),
    .io_dec_lsu_valid_raw_d(bus_buffer_io_dec_lsu_valid_raw_d),
    .io_lsu_pkt_m_valid(bus_buffer_io_lsu_pkt_m_valid),
    .io_lsu_pkt_m_bits_load(bus_buffer_io_lsu_pkt_m_bits_load),
    .io_lsu_pkt_r_bits_by(bus_buffer_io_lsu_pkt_r_bits_by),
    .io_lsu_pkt_r_bits_half(bus_buffer_io_lsu_pkt_r_bits_half),
    .io_lsu_pkt_r_bits_word(bus_buffer_io_lsu_pkt_r_bits_word),
    .io_lsu_pkt_r_bits_load(bus_buffer_io_lsu_pkt_r_bits_load),
    .io_lsu_pkt_r_bits_store(bus_buffer_io_lsu_pkt_r_bits_store),
    .io_lsu_pkt_r_bits_unsign(bus_buffer_io_lsu_pkt_r_bits_unsign),
    .io_lsu_addr_m(bus_buffer_io_lsu_addr_m),
    .io_end_addr_m(bus_buffer_io_end_addr_m),
    .io_lsu_addr_r(bus_buffer_io_lsu_addr_r),
    .io_end_addr_r(bus_buffer_io_end_addr_r),
    .io_store_data_r(bus_buffer_io_store_data_r),
    .io_no_word_merge_r(bus_buffer_io_no_word_merge_r),
    .io_no_dword_merge_r(bus_buffer_io_no_dword_merge_r),
    .io_lsu_busreq_m(bus_buffer_io_lsu_busreq_m),
    .io_ld_full_hit_m(bus_buffer_io_ld_full_hit_m),
    .io_flush_m_up(bus_buffer_io_flush_m_up),
    .io_flush_r(bus_buffer_io_flush_r),
    .io_lsu_commit_r(bus_buffer_io_lsu_commit_r),
    .io_is_sideeffects_r(bus_buffer_io_is_sideeffects_r),
    .io_ldst_dual_d(bus_buffer_io_ldst_dual_d),
    .io_ldst_dual_m(bus_buffer_io_ldst_dual_m),
    .io_ldst_dual_r(bus_buffer_io_ldst_dual_r),
    .io_ldst_byteen_ext_m(bus_buffer_io_ldst_byteen_ext_m),
    .io_lsu_axi_aw_valid(bus_buffer_io_lsu_axi_aw_valid),
    .io_lsu_axi_aw_bits_addr(bus_buffer_io_lsu_axi_aw_bits_addr),
    .io_lsu_axi_aw_bits_size(bus_buffer_io_lsu_axi_aw_bits_size),
    .io_lsu_axi_w_valid(bus_buffer_io_lsu_axi_w_valid),
    .io_lsu_axi_w_bits_strb(bus_buffer_io_lsu_axi_w_bits_strb),
    .io_lsu_axi_ar_valid(bus_buffer_io_lsu_axi_ar_valid),
    .io_lsu_axi_ar_bits_addr(bus_buffer_io_lsu_axi_ar_bits_addr),
    .io_lsu_axi_ar_bits_size(bus_buffer_io_lsu_axi_ar_bits_size),
    .io_lsu_bus_clk_en(bus_buffer_io_lsu_bus_clk_en),
    .io_lsu_bus_clk_en_q(bus_buffer_io_lsu_bus_clk_en_q),
    .io_lsu_busreq_r(bus_buffer_io_lsu_busreq_r),
    .io_lsu_bus_buffer_pend_any(bus_buffer_io_lsu_bus_buffer_pend_any),
    .io_lsu_bus_buffer_full_any(bus_buffer_io_lsu_bus_buffer_full_any),
    .io_lsu_bus_buffer_empty_any(bus_buffer_io_lsu_bus_buffer_empty_any),
    .io_ld_byte_hit_buf_lo(bus_buffer_io_ld_byte_hit_buf_lo),
    .io_ld_byte_hit_buf_hi(bus_buffer_io_ld_byte_hit_buf_hi),
    .io_ld_fwddata_buf_lo(bus_buffer_io_ld_fwddata_buf_lo),
    .io_ld_fwddata_buf_hi(bus_buffer_io_ld_fwddata_buf_hi)
  );
  assign io_tlu_busbuff_lsu_pmu_bus_misaligned = bus_buffer_io_tlu_busbuff_lsu_pmu_bus_misaligned; // @[lsu_bus_intf.scala 104:18]
  assign io_tlu_busbuff_lsu_pmu_bus_error = bus_buffer_io_tlu_busbuff_lsu_pmu_bus_error; // @[lsu_bus_intf.scala 104:18]
  assign io_tlu_busbuff_lsu_pmu_bus_busy = bus_buffer_io_tlu_busbuff_lsu_pmu_bus_busy; // @[lsu_bus_intf.scala 104:18]
  assign io_tlu_busbuff_lsu_imprecise_error_load_any = bus_buffer_io_tlu_busbuff_lsu_imprecise_error_load_any; // @[lsu_bus_intf.scala 104:18]
  assign io_tlu_busbuff_lsu_imprecise_error_store_any = bus_buffer_io_tlu_busbuff_lsu_imprecise_error_store_any; // @[lsu_bus_intf.scala 104:18]
  assign io_tlu_busbuff_lsu_imprecise_error_addr_any = bus_buffer_io_tlu_busbuff_lsu_imprecise_error_addr_any; // @[lsu_bus_intf.scala 104:18]
  assign io_axi_aw_valid = bus_buffer_io_lsu_axi_aw_valid; // @[lsu_bus_intf.scala 130:43]
  assign io_axi_aw_bits_addr = bus_buffer_io_lsu_axi_aw_bits_addr; // @[lsu_bus_intf.scala 130:43]
  assign io_axi_aw_bits_size = bus_buffer_io_lsu_axi_aw_bits_size; // @[lsu_bus_intf.scala 130:43]
  assign io_axi_w_valid = bus_buffer_io_lsu_axi_w_valid; // @[lsu_bus_intf.scala 130:43]
  assign io_axi_w_bits_strb = bus_buffer_io_lsu_axi_w_bits_strb; // @[lsu_bus_intf.scala 130:43]
  assign io_axi_ar_valid = bus_buffer_io_lsu_axi_ar_valid; // @[lsu_bus_intf.scala 130:43]
  assign io_axi_ar_bits_addr = bus_buffer_io_lsu_axi_ar_bits_addr; // @[lsu_bus_intf.scala 130:43]
  assign io_axi_ar_bits_size = bus_buffer_io_lsu_axi_ar_bits_size; // @[lsu_bus_intf.scala 130:43]
  assign io_lsu_busreq_r = bus_buffer_io_lsu_busreq_r; // @[lsu_bus_intf.scala 133:38]
  assign io_lsu_bus_buffer_pend_any = bus_buffer_io_lsu_bus_buffer_pend_any; // @[lsu_bus_intf.scala 134:38]
  assign io_lsu_bus_buffer_full_any = bus_buffer_io_lsu_bus_buffer_full_any; // @[lsu_bus_intf.scala 135:38]
  assign io_lsu_bus_buffer_empty_any = bus_buffer_io_lsu_bus_buffer_empty_any; // @[lsu_bus_intf.scala 136:38]
  assign io_bus_read_data_m = ld_fwddata_m[31:0]; // @[lsu_bus_intf.scala 192:27]
  assign io_dctl_busbuff_lsu_nonblock_load_valid_m = bus_buffer_io_dctl_busbuff_lsu_nonblock_load_valid_m; // @[lsu_bus_intf.scala 142:19]
  assign io_dctl_busbuff_lsu_nonblock_load_tag_m = bus_buffer_io_dctl_busbuff_lsu_nonblock_load_tag_m; // @[lsu_bus_intf.scala 142:19]
  assign io_dctl_busbuff_lsu_nonblock_load_inv_r = bus_buffer_io_dctl_busbuff_lsu_nonblock_load_inv_r; // @[lsu_bus_intf.scala 142:19]
  assign io_dctl_busbuff_lsu_nonblock_load_inv_tag_r = bus_buffer_io_dctl_busbuff_lsu_nonblock_load_inv_tag_r; // @[lsu_bus_intf.scala 142:19]
  assign io_dctl_busbuff_lsu_nonblock_load_data_valid = bus_buffer_io_dctl_busbuff_lsu_nonblock_load_data_valid; // @[lsu_bus_intf.scala 142:19]
  assign io_dctl_busbuff_lsu_nonblock_load_data_error = bus_buffer_io_dctl_busbuff_lsu_nonblock_load_data_error; // @[lsu_bus_intf.scala 142:19]
  assign io_dctl_busbuff_lsu_nonblock_load_data_tag = bus_buffer_io_dctl_busbuff_lsu_nonblock_load_data_tag; // @[lsu_bus_intf.scala 142:19]
  assign io_dctl_busbuff_lsu_nonblock_load_data = bus_buffer_io_dctl_busbuff_lsu_nonblock_load_data; // @[lsu_bus_intf.scala 142:19]
  assign bus_buffer_clock = clock;
  assign bus_buffer_reset = reset;
  assign bus_buffer_io_scan_mode = io_scan_mode; // @[lsu_bus_intf.scala 103:29]
  assign bus_buffer_io_tlu_busbuff_dec_tlu_external_ldfwd_disable = io_tlu_busbuff_dec_tlu_external_ldfwd_disable; // @[lsu_bus_intf.scala 104:18]
  assign bus_buffer_io_tlu_busbuff_dec_tlu_wb_coalescing_disable = io_tlu_busbuff_dec_tlu_wb_coalescing_disable; // @[lsu_bus_intf.scala 104:18]
  assign bus_buffer_io_tlu_busbuff_dec_tlu_sideeffect_posted_disable = io_tlu_busbuff_dec_tlu_sideeffect_posted_disable; // @[lsu_bus_intf.scala 104:18]
  assign bus_buffer_io_dec_tlu_force_halt = io_dec_tlu_force_halt; // @[lsu_bus_intf.scala 106:51]
  assign bus_buffer_io_lsu_c2_r_clk = io_lsu_c2_r_clk; // @[lsu_bus_intf.scala 107:51]
  assign bus_buffer_io_lsu_bus_ibuf_c1_clk = io_lsu_bus_ibuf_c1_clk; // @[lsu_bus_intf.scala 108:51]
  assign bus_buffer_io_lsu_bus_obuf_c1_clk = io_lsu_bus_obuf_c1_clk; // @[lsu_bus_intf.scala 109:51]
  assign bus_buffer_io_lsu_bus_buf_c1_clk = io_lsu_bus_buf_c1_clk; // @[lsu_bus_intf.scala 110:51]
  assign bus_buffer_io_lsu_free_c2_clk = io_lsu_free_c2_clk; // @[lsu_bus_intf.scala 111:51]
  assign bus_buffer_io_lsu_busm_clk = io_lsu_busm_clk; // @[lsu_bus_intf.scala 112:51]
  assign bus_buffer_io_dec_lsu_valid_raw_d = io_dec_lsu_valid_raw_d; // @[lsu_bus_intf.scala 113:51]
  assign bus_buffer_io_lsu_pkt_m_valid = io_lsu_pkt_m_valid; // @[lsu_bus_intf.scala 116:27]
  assign bus_buffer_io_lsu_pkt_m_bits_load = io_lsu_pkt_m_bits_load; // @[lsu_bus_intf.scala 116:27]
  assign bus_buffer_io_lsu_pkt_r_bits_by = io_lsu_pkt_r_bits_by; // @[lsu_bus_intf.scala 117:27]
  assign bus_buffer_io_lsu_pkt_r_bits_half = io_lsu_pkt_r_bits_half; // @[lsu_bus_intf.scala 117:27]
  assign bus_buffer_io_lsu_pkt_r_bits_word = io_lsu_pkt_r_bits_word; // @[lsu_bus_intf.scala 117:27]
  assign bus_buffer_io_lsu_pkt_r_bits_load = io_lsu_pkt_r_bits_load; // @[lsu_bus_intf.scala 117:27]
  assign bus_buffer_io_lsu_pkt_r_bits_store = io_lsu_pkt_r_bits_store; // @[lsu_bus_intf.scala 117:27]
  assign bus_buffer_io_lsu_pkt_r_bits_unsign = io_lsu_pkt_r_bits_unsign; // @[lsu_bus_intf.scala 117:27]
  assign bus_buffer_io_lsu_addr_m = io_lsu_addr_m; // @[lsu_bus_intf.scala 120:51]
  assign bus_buffer_io_end_addr_m = io_end_addr_m; // @[lsu_bus_intf.scala 121:51]
  assign bus_buffer_io_lsu_addr_r = io_lsu_addr_r; // @[lsu_bus_intf.scala 122:51]
  assign bus_buffer_io_end_addr_r = io_end_addr_r; // @[lsu_bus_intf.scala 123:51]
  assign bus_buffer_io_store_data_r = io_store_data_r; // @[lsu_bus_intf.scala 124:51]
  assign bus_buffer_io_no_word_merge_r = _T_22 & _T_24; // @[lsu_bus_intf.scala 143:51]
  assign bus_buffer_io_no_dword_merge_r = _T_22 & _T_30; // @[lsu_bus_intf.scala 144:51]
  assign bus_buffer_io_lsu_busreq_m = io_lsu_busreq_m; // @[lsu_bus_intf.scala 126:51]
  assign bus_buffer_io_ld_full_hit_m = _T_372 & _T_373; // @[lsu_bus_intf.scala 150:51]
  assign bus_buffer_io_flush_m_up = io_flush_m_up; // @[lsu_bus_intf.scala 127:51]
  assign bus_buffer_io_flush_r = io_flush_r; // @[lsu_bus_intf.scala 128:51]
  assign bus_buffer_io_lsu_commit_r = io_lsu_commit_r; // @[lsu_bus_intf.scala 129:51]
  assign bus_buffer_io_is_sideeffects_r = is_sideeffects_r; // @[lsu_bus_intf.scala 145:51]
  assign bus_buffer_io_ldst_dual_d = io_lsu_addr_d[2] != io_end_addr_d[2]; // @[lsu_bus_intf.scala 146:51]
  assign bus_buffer_io_ldst_dual_m = ldst_dual_m; // @[lsu_bus_intf.scala 147:51]
  assign bus_buffer_io_ldst_dual_r = ldst_dual_r; // @[lsu_bus_intf.scala 148:51]
  assign bus_buffer_io_ldst_byteen_ext_m = {{1'd0}, _T_34}; // @[lsu_bus_intf.scala 149:51]
  assign bus_buffer_io_lsu_bus_clk_en = io_lsu_bus_clk_en; // @[lsu_bus_intf.scala 131:51]
  assign bus_buffer_io_lsu_bus_clk_en_q = lsu_bus_clk_en_q; // @[lsu_bus_intf.scala 151:51]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ldst_dual_r = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  ldst_byteen_r = _RAND_1[3:0];
  _RAND_2 = {1{`RANDOM}};
  lsu_bus_clk_en_q = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  ldst_dual_m = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  is_sideeffects_r = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    ldst_dual_r = 1'h0;
  end
  if (reset) begin
    ldst_byteen_r = 4'h0;
  end
  if (reset) begin
    lsu_bus_clk_en_q = 1'h0;
  end
  if (reset) begin
    ldst_dual_m = 1'h0;
  end
  if (reset) begin
    is_sideeffects_r = 1'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge io_lsu_c1_r_clk or posedge reset) begin
    if (reset) begin
      ldst_dual_r <= 1'h0;
    end else begin
      ldst_dual_r <= ldst_dual_m;
    end
  end
  always @(posedge io_lsu_c1_r_clk or posedge reset) begin
    if (reset) begin
      ldst_byteen_r <= 4'h0;
    end else begin
      ldst_byteen_r <= _T_6 | _T_5;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      lsu_bus_clk_en_q <= 1'h0;
    end else begin
      lsu_bus_clk_en_q <= io_lsu_bus_clk_en;
    end
  end
  always @(posedge io_lsu_c1_m_clk or posedge reset) begin
    if (reset) begin
      ldst_dual_m <= 1'h0;
    end else begin
      ldst_dual_m <= io_lsu_addr_d[2] != io_end_addr_d[2];
    end
  end
  always @(posedge io_lsu_c1_r_clk or posedge reset) begin
    if (reset) begin
      is_sideeffects_r <= 1'h0;
    end else begin
      is_sideeffects_r <= io_is_sideeffects_m;
    end
  end
endmodule
module lsu(
  input         clock,
  input         reset,
  input         io_clk_override,
  input         io_lsu_dma_dma_lsc_ctl_dma_dccm_req,
  input  [31:0] io_lsu_dma_dma_lsc_ctl_dma_mem_addr,
  input  [2:0]  io_lsu_dma_dma_lsc_ctl_dma_mem_sz,
  input         io_lsu_dma_dma_lsc_ctl_dma_mem_write,
  input  [63:0] io_lsu_dma_dma_lsc_ctl_dma_mem_wdata,
  input  [31:0] io_lsu_dma_dma_dccm_ctl_dma_mem_addr,
  input  [63:0] io_lsu_dma_dma_dccm_ctl_dma_mem_wdata,
  output        io_lsu_dma_dma_dccm_ctl_dccm_dma_rvalid,
  output        io_lsu_dma_dma_dccm_ctl_dccm_dma_ecc_error,
  output [2:0]  io_lsu_dma_dma_dccm_ctl_dccm_dma_rtag,
  output [63:0] io_lsu_dma_dma_dccm_ctl_dccm_dma_rdata,
  output        io_lsu_dma_dccm_ready,
  input  [2:0]  io_lsu_dma_dma_mem_tag,
  output        io_lsu_pic_picm_wren,
  output        io_lsu_pic_picm_rden,
  output        io_lsu_pic_picm_mken,
  output [31:0] io_lsu_pic_picm_rdaddr,
  output [31:0] io_lsu_pic_picm_wraddr,
  output [31:0] io_lsu_pic_picm_wr_data,
  input  [31:0] io_lsu_pic_picm_rd_data,
  input  [31:0] io_lsu_exu_exu_lsu_rs1_d,
  input  [31:0] io_lsu_exu_exu_lsu_rs2_d,
  output        io_lsu_dec_tlu_busbuff_lsu_pmu_bus_misaligned,
  output        io_lsu_dec_tlu_busbuff_lsu_pmu_bus_error,
  output        io_lsu_dec_tlu_busbuff_lsu_pmu_bus_busy,
  input         io_lsu_dec_tlu_busbuff_dec_tlu_external_ldfwd_disable,
  input         io_lsu_dec_tlu_busbuff_dec_tlu_wb_coalescing_disable,
  input         io_lsu_dec_tlu_busbuff_dec_tlu_sideeffect_posted_disable,
  output        io_lsu_dec_tlu_busbuff_lsu_imprecise_error_load_any,
  output        io_lsu_dec_tlu_busbuff_lsu_imprecise_error_store_any,
  output [31:0] io_lsu_dec_tlu_busbuff_lsu_imprecise_error_addr_any,
  output        io_lsu_dec_dctl_busbuff_lsu_nonblock_load_valid_m,
  output [1:0]  io_lsu_dec_dctl_busbuff_lsu_nonblock_load_tag_m,
  output        io_lsu_dec_dctl_busbuff_lsu_nonblock_load_inv_r,
  output [1:0]  io_lsu_dec_dctl_busbuff_lsu_nonblock_load_inv_tag_r,
  output        io_lsu_dec_dctl_busbuff_lsu_nonblock_load_data_valid,
  output        io_lsu_dec_dctl_busbuff_lsu_nonblock_load_data_error,
  output [1:0]  io_lsu_dec_dctl_busbuff_lsu_nonblock_load_data_tag,
  output [31:0] io_lsu_dec_dctl_busbuff_lsu_nonblock_load_data,
  output        io_dccm_wren,
  output        io_dccm_rden,
  output [15:0] io_dccm_wr_addr_lo,
  output [15:0] io_dccm_wr_addr_hi,
  output [15:0] io_dccm_rd_addr_lo,
  output [15:0] io_dccm_rd_addr_hi,
  output [38:0] io_dccm_wr_data_lo,
  output [38:0] io_dccm_wr_data_hi,
  input  [38:0] io_dccm_rd_data_lo,
  input  [38:0] io_dccm_rd_data_hi,
  output        io_lsu_tlu_lsu_pmu_load_external_m,
  output        io_lsu_tlu_lsu_pmu_store_external_m,
  output        io_axi_aw_valid,
  output [31:0] io_axi_aw_bits_addr,
  output [2:0]  io_axi_aw_bits_size,
  output        io_axi_w_valid,
  output [7:0]  io_axi_w_bits_strb,
  output        io_axi_ar_valid,
  output [31:0] io_axi_ar_bits_addr,
  output [2:0]  io_axi_ar_bits_size,
  input         io_dec_tlu_flush_lower_r,
  input         io_dec_tlu_i0_kill_writeb_r,
  input         io_dec_tlu_force_halt,
  input         io_dec_tlu_core_ecc_disable,
  input  [11:0] io_dec_lsu_offset_d,
  input         io_lsu_p_valid,
  input         io_lsu_p_bits_fast_int,
  input         io_lsu_p_bits_by,
  input         io_lsu_p_bits_half,
  input         io_lsu_p_bits_word,
  input         io_lsu_p_bits_load,
  input         io_lsu_p_bits_store,
  input         io_lsu_p_bits_unsign,
  input         io_lsu_p_bits_store_data_bypass_d,
  input         io_lsu_p_bits_load_ldst_bypass_d,
  input         io_trigger_pkt_any_0_select,
  input         io_trigger_pkt_any_0_match_pkt,
  input         io_trigger_pkt_any_0_store,
  input         io_trigger_pkt_any_0_load,
  input  [31:0] io_trigger_pkt_any_0_tdata2,
  input         io_trigger_pkt_any_1_select,
  input         io_trigger_pkt_any_1_match_pkt,
  input         io_trigger_pkt_any_1_store,
  input         io_trigger_pkt_any_1_load,
  input  [31:0] io_trigger_pkt_any_1_tdata2,
  input         io_trigger_pkt_any_2_select,
  input         io_trigger_pkt_any_2_match_pkt,
  input         io_trigger_pkt_any_2_store,
  input         io_trigger_pkt_any_2_load,
  input  [31:0] io_trigger_pkt_any_2_tdata2,
  input         io_trigger_pkt_any_3_select,
  input         io_trigger_pkt_any_3_match_pkt,
  input         io_trigger_pkt_any_3_store,
  input         io_trigger_pkt_any_3_load,
  input  [31:0] io_trigger_pkt_any_3_tdata2,
  input         io_dec_lsu_valid_raw_d,
  input  [31:0] io_dec_tlu_mrac_ff,
  output [31:0] io_lsu_result_m,
  output [31:0] io_lsu_result_corr_r,
  output        io_lsu_load_stall_any,
  output        io_lsu_store_stall_any,
  output        io_lsu_fastint_stall_any,
  output        io_lsu_idle_any,
  output [30:0] io_lsu_fir_addr,
  output [1:0]  io_lsu_fir_error,
  output        io_lsu_single_ecc_error_incr,
  output        io_lsu_error_pkt_r_valid,
  output        io_lsu_error_pkt_r_bits_single_ecc_error,
  output        io_lsu_error_pkt_r_bits_inst_type,
  output        io_lsu_error_pkt_r_bits_exc_type,
  output [3:0]  io_lsu_error_pkt_r_bits_mscause,
  output [31:0] io_lsu_error_pkt_r_bits_addr,
  output        io_lsu_pmu_misaligned_m,
  output [3:0]  io_lsu_trigger_match_m,
  input         io_lsu_bus_clk_en,
  input         io_scan_mode,
  input         io_free_clk
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire  lsu_lsc_ctl_reset; // @[lsu.scala 60:30]
  wire  lsu_lsc_ctl_io_lsu_c1_m_clk; // @[lsu.scala 60:30]
  wire  lsu_lsc_ctl_io_lsu_c1_r_clk; // @[lsu.scala 60:30]
  wire  lsu_lsc_ctl_io_lsu_c2_m_clk; // @[lsu.scala 60:30]
  wire  lsu_lsc_ctl_io_lsu_c2_r_clk; // @[lsu.scala 60:30]
  wire  lsu_lsc_ctl_io_lsu_store_c1_m_clk; // @[lsu.scala 60:30]
  wire [31:0] lsu_lsc_ctl_io_lsu_ld_data_corr_r; // @[lsu.scala 60:30]
  wire  lsu_lsc_ctl_io_lsu_single_ecc_error_r; // @[lsu.scala 60:30]
  wire  lsu_lsc_ctl_io_lsu_double_ecc_error_r; // @[lsu.scala 60:30]
  wire [31:0] lsu_lsc_ctl_io_lsu_ld_data_m; // @[lsu.scala 60:30]
  wire  lsu_lsc_ctl_io_lsu_single_ecc_error_m; // @[lsu.scala 60:30]
  wire  lsu_lsc_ctl_io_lsu_double_ecc_error_m; // @[lsu.scala 60:30]
  wire  lsu_lsc_ctl_io_flush_m_up; // @[lsu.scala 60:30]
  wire  lsu_lsc_ctl_io_flush_r; // @[lsu.scala 60:30]
  wire [31:0] lsu_lsc_ctl_io_lsu_exu_exu_lsu_rs1_d; // @[lsu.scala 60:30]
  wire [31:0] lsu_lsc_ctl_io_lsu_exu_exu_lsu_rs2_d; // @[lsu.scala 60:30]
  wire  lsu_lsc_ctl_io_lsu_p_valid; // @[lsu.scala 60:30]
  wire  lsu_lsc_ctl_io_lsu_p_bits_fast_int; // @[lsu.scala 60:30]
  wire  lsu_lsc_ctl_io_lsu_p_bits_by; // @[lsu.scala 60:30]
  wire  lsu_lsc_ctl_io_lsu_p_bits_half; // @[lsu.scala 60:30]
  wire  lsu_lsc_ctl_io_lsu_p_bits_word; // @[lsu.scala 60:30]
  wire  lsu_lsc_ctl_io_lsu_p_bits_load; // @[lsu.scala 60:30]
  wire  lsu_lsc_ctl_io_lsu_p_bits_store; // @[lsu.scala 60:30]
  wire  lsu_lsc_ctl_io_lsu_p_bits_unsign; // @[lsu.scala 60:30]
  wire  lsu_lsc_ctl_io_lsu_p_bits_store_data_bypass_d; // @[lsu.scala 60:30]
  wire  lsu_lsc_ctl_io_lsu_p_bits_load_ldst_bypass_d; // @[lsu.scala 60:30]
  wire  lsu_lsc_ctl_io_dec_lsu_valid_raw_d; // @[lsu.scala 60:30]
  wire [11:0] lsu_lsc_ctl_io_dec_lsu_offset_d; // @[lsu.scala 60:30]
  wire [31:0] lsu_lsc_ctl_io_picm_mask_data_m; // @[lsu.scala 60:30]
  wire [31:0] lsu_lsc_ctl_io_bus_read_data_m; // @[lsu.scala 60:30]
  wire [31:0] lsu_lsc_ctl_io_lsu_result_m; // @[lsu.scala 60:30]
  wire [31:0] lsu_lsc_ctl_io_lsu_result_corr_r; // @[lsu.scala 60:30]
  wire [31:0] lsu_lsc_ctl_io_lsu_addr_d; // @[lsu.scala 60:30]
  wire [31:0] lsu_lsc_ctl_io_lsu_addr_m; // @[lsu.scala 60:30]
  wire [31:0] lsu_lsc_ctl_io_lsu_addr_r; // @[lsu.scala 60:30]
  wire [31:0] lsu_lsc_ctl_io_end_addr_d; // @[lsu.scala 60:30]
  wire [31:0] lsu_lsc_ctl_io_end_addr_m; // @[lsu.scala 60:30]
  wire [31:0] lsu_lsc_ctl_io_end_addr_r; // @[lsu.scala 60:30]
  wire [31:0] lsu_lsc_ctl_io_store_data_m; // @[lsu.scala 60:30]
  wire [31:0] lsu_lsc_ctl_io_dec_tlu_mrac_ff; // @[lsu.scala 60:30]
  wire  lsu_lsc_ctl_io_lsu_exc_m; // @[lsu.scala 60:30]
  wire  lsu_lsc_ctl_io_is_sideeffects_m; // @[lsu.scala 60:30]
  wire  lsu_lsc_ctl_io_lsu_commit_r; // @[lsu.scala 60:30]
  wire  lsu_lsc_ctl_io_lsu_single_ecc_error_incr; // @[lsu.scala 60:30]
  wire  lsu_lsc_ctl_io_lsu_error_pkt_r_valid; // @[lsu.scala 60:30]
  wire  lsu_lsc_ctl_io_lsu_error_pkt_r_bits_single_ecc_error; // @[lsu.scala 60:30]
  wire  lsu_lsc_ctl_io_lsu_error_pkt_r_bits_inst_type; // @[lsu.scala 60:30]
  wire  lsu_lsc_ctl_io_lsu_error_pkt_r_bits_exc_type; // @[lsu.scala 60:30]
  wire [3:0] lsu_lsc_ctl_io_lsu_error_pkt_r_bits_mscause; // @[lsu.scala 60:30]
  wire [31:0] lsu_lsc_ctl_io_lsu_error_pkt_r_bits_addr; // @[lsu.scala 60:30]
  wire [30:0] lsu_lsc_ctl_io_lsu_fir_addr; // @[lsu.scala 60:30]
  wire [1:0] lsu_lsc_ctl_io_lsu_fir_error; // @[lsu.scala 60:30]
  wire  lsu_lsc_ctl_io_addr_in_dccm_d; // @[lsu.scala 60:30]
  wire  lsu_lsc_ctl_io_addr_in_dccm_m; // @[lsu.scala 60:30]
  wire  lsu_lsc_ctl_io_addr_in_dccm_r; // @[lsu.scala 60:30]
  wire  lsu_lsc_ctl_io_addr_in_pic_d; // @[lsu.scala 60:30]
  wire  lsu_lsc_ctl_io_addr_in_pic_m; // @[lsu.scala 60:30]
  wire  lsu_lsc_ctl_io_addr_in_pic_r; // @[lsu.scala 60:30]
  wire  lsu_lsc_ctl_io_addr_external_m; // @[lsu.scala 60:30]
  wire  lsu_lsc_ctl_io_dma_lsc_ctl_dma_dccm_req; // @[lsu.scala 60:30]
  wire [31:0] lsu_lsc_ctl_io_dma_lsc_ctl_dma_mem_addr; // @[lsu.scala 60:30]
  wire [2:0] lsu_lsc_ctl_io_dma_lsc_ctl_dma_mem_sz; // @[lsu.scala 60:30]
  wire  lsu_lsc_ctl_io_dma_lsc_ctl_dma_mem_write; // @[lsu.scala 60:30]
  wire [63:0] lsu_lsc_ctl_io_dma_lsc_ctl_dma_mem_wdata; // @[lsu.scala 60:30]
  wire  lsu_lsc_ctl_io_lsu_pkt_d_valid; // @[lsu.scala 60:30]
  wire  lsu_lsc_ctl_io_lsu_pkt_d_bits_fast_int; // @[lsu.scala 60:30]
  wire  lsu_lsc_ctl_io_lsu_pkt_d_bits_by; // @[lsu.scala 60:30]
  wire  lsu_lsc_ctl_io_lsu_pkt_d_bits_half; // @[lsu.scala 60:30]
  wire  lsu_lsc_ctl_io_lsu_pkt_d_bits_word; // @[lsu.scala 60:30]
  wire  lsu_lsc_ctl_io_lsu_pkt_d_bits_dword; // @[lsu.scala 60:30]
  wire  lsu_lsc_ctl_io_lsu_pkt_d_bits_load; // @[lsu.scala 60:30]
  wire  lsu_lsc_ctl_io_lsu_pkt_d_bits_store; // @[lsu.scala 60:30]
  wire  lsu_lsc_ctl_io_lsu_pkt_d_bits_unsign; // @[lsu.scala 60:30]
  wire  lsu_lsc_ctl_io_lsu_pkt_d_bits_dma; // @[lsu.scala 60:30]
  wire  lsu_lsc_ctl_io_lsu_pkt_d_bits_store_data_bypass_d; // @[lsu.scala 60:30]
  wire  lsu_lsc_ctl_io_lsu_pkt_d_bits_load_ldst_bypass_d; // @[lsu.scala 60:30]
  wire  lsu_lsc_ctl_io_lsu_pkt_d_bits_store_data_bypass_m; // @[lsu.scala 60:30]
  wire  lsu_lsc_ctl_io_lsu_pkt_m_valid; // @[lsu.scala 60:30]
  wire  lsu_lsc_ctl_io_lsu_pkt_m_bits_fast_int; // @[lsu.scala 60:30]
  wire  lsu_lsc_ctl_io_lsu_pkt_m_bits_by; // @[lsu.scala 60:30]
  wire  lsu_lsc_ctl_io_lsu_pkt_m_bits_half; // @[lsu.scala 60:30]
  wire  lsu_lsc_ctl_io_lsu_pkt_m_bits_word; // @[lsu.scala 60:30]
  wire  lsu_lsc_ctl_io_lsu_pkt_m_bits_dword; // @[lsu.scala 60:30]
  wire  lsu_lsc_ctl_io_lsu_pkt_m_bits_load; // @[lsu.scala 60:30]
  wire  lsu_lsc_ctl_io_lsu_pkt_m_bits_store; // @[lsu.scala 60:30]
  wire  lsu_lsc_ctl_io_lsu_pkt_m_bits_unsign; // @[lsu.scala 60:30]
  wire  lsu_lsc_ctl_io_lsu_pkt_m_bits_dma; // @[lsu.scala 60:30]
  wire  lsu_lsc_ctl_io_lsu_pkt_m_bits_store_data_bypass_m; // @[lsu.scala 60:30]
  wire  lsu_lsc_ctl_io_lsu_pkt_r_valid; // @[lsu.scala 60:30]
  wire  lsu_lsc_ctl_io_lsu_pkt_r_bits_by; // @[lsu.scala 60:30]
  wire  lsu_lsc_ctl_io_lsu_pkt_r_bits_half; // @[lsu.scala 60:30]
  wire  lsu_lsc_ctl_io_lsu_pkt_r_bits_word; // @[lsu.scala 60:30]
  wire  lsu_lsc_ctl_io_lsu_pkt_r_bits_dword; // @[lsu.scala 60:30]
  wire  lsu_lsc_ctl_io_lsu_pkt_r_bits_load; // @[lsu.scala 60:30]
  wire  lsu_lsc_ctl_io_lsu_pkt_r_bits_store; // @[lsu.scala 60:30]
  wire  lsu_lsc_ctl_io_lsu_pkt_r_bits_unsign; // @[lsu.scala 60:30]
  wire  lsu_lsc_ctl_io_lsu_pkt_r_bits_dma; // @[lsu.scala 60:30]
  wire  dccm_ctl_clock; // @[lsu.scala 63:30]
  wire  dccm_ctl_reset; // @[lsu.scala 63:30]
  wire  dccm_ctl_io_lsu_c2_m_clk; // @[lsu.scala 63:30]
  wire  dccm_ctl_io_lsu_c2_r_clk; // @[lsu.scala 63:30]
  wire  dccm_ctl_io_lsu_free_c2_clk; // @[lsu.scala 63:30]
  wire  dccm_ctl_io_lsu_store_c1_r_clk; // @[lsu.scala 63:30]
  wire  dccm_ctl_io_lsu_pkt_d_valid; // @[lsu.scala 63:30]
  wire  dccm_ctl_io_lsu_pkt_d_bits_word; // @[lsu.scala 63:30]
  wire  dccm_ctl_io_lsu_pkt_d_bits_dword; // @[lsu.scala 63:30]
  wire  dccm_ctl_io_lsu_pkt_d_bits_load; // @[lsu.scala 63:30]
  wire  dccm_ctl_io_lsu_pkt_d_bits_store; // @[lsu.scala 63:30]
  wire  dccm_ctl_io_lsu_pkt_d_bits_dma; // @[lsu.scala 63:30]
  wire  dccm_ctl_io_lsu_pkt_m_valid; // @[lsu.scala 63:30]
  wire  dccm_ctl_io_lsu_pkt_m_bits_by; // @[lsu.scala 63:30]
  wire  dccm_ctl_io_lsu_pkt_m_bits_half; // @[lsu.scala 63:30]
  wire  dccm_ctl_io_lsu_pkt_m_bits_word; // @[lsu.scala 63:30]
  wire  dccm_ctl_io_lsu_pkt_m_bits_load; // @[lsu.scala 63:30]
  wire  dccm_ctl_io_lsu_pkt_m_bits_store; // @[lsu.scala 63:30]
  wire  dccm_ctl_io_lsu_pkt_m_bits_dma; // @[lsu.scala 63:30]
  wire  dccm_ctl_io_lsu_pkt_r_valid; // @[lsu.scala 63:30]
  wire  dccm_ctl_io_lsu_pkt_r_bits_by; // @[lsu.scala 63:30]
  wire  dccm_ctl_io_lsu_pkt_r_bits_half; // @[lsu.scala 63:30]
  wire  dccm_ctl_io_lsu_pkt_r_bits_word; // @[lsu.scala 63:30]
  wire  dccm_ctl_io_lsu_pkt_r_bits_load; // @[lsu.scala 63:30]
  wire  dccm_ctl_io_lsu_pkt_r_bits_store; // @[lsu.scala 63:30]
  wire  dccm_ctl_io_lsu_pkt_r_bits_dma; // @[lsu.scala 63:30]
  wire  dccm_ctl_io_addr_in_dccm_d; // @[lsu.scala 63:30]
  wire  dccm_ctl_io_addr_in_dccm_m; // @[lsu.scala 63:30]
  wire  dccm_ctl_io_addr_in_dccm_r; // @[lsu.scala 63:30]
  wire  dccm_ctl_io_addr_in_pic_d; // @[lsu.scala 63:30]
  wire  dccm_ctl_io_addr_in_pic_m; // @[lsu.scala 63:30]
  wire  dccm_ctl_io_addr_in_pic_r; // @[lsu.scala 63:30]
  wire  dccm_ctl_io_lsu_raw_fwd_lo_r; // @[lsu.scala 63:30]
  wire  dccm_ctl_io_lsu_raw_fwd_hi_r; // @[lsu.scala 63:30]
  wire  dccm_ctl_io_lsu_commit_r; // @[lsu.scala 63:30]
  wire [31:0] dccm_ctl_io_lsu_addr_d; // @[lsu.scala 63:30]
  wire [15:0] dccm_ctl_io_lsu_addr_m; // @[lsu.scala 63:30]
  wire [31:0] dccm_ctl_io_lsu_addr_r; // @[lsu.scala 63:30]
  wire [15:0] dccm_ctl_io_end_addr_d; // @[lsu.scala 63:30]
  wire [15:0] dccm_ctl_io_end_addr_m; // @[lsu.scala 63:30]
  wire [15:0] dccm_ctl_io_end_addr_r; // @[lsu.scala 63:30]
  wire  dccm_ctl_io_stbuf_reqvld_any; // @[lsu.scala 63:30]
  wire [15:0] dccm_ctl_io_stbuf_addr_any; // @[lsu.scala 63:30]
  wire [31:0] dccm_ctl_io_stbuf_data_any; // @[lsu.scala 63:30]
  wire [6:0] dccm_ctl_io_stbuf_ecc_any; // @[lsu.scala 63:30]
  wire [31:0] dccm_ctl_io_stbuf_fwddata_hi_m; // @[lsu.scala 63:30]
  wire [31:0] dccm_ctl_io_stbuf_fwddata_lo_m; // @[lsu.scala 63:30]
  wire [3:0] dccm_ctl_io_stbuf_fwdbyteen_lo_m; // @[lsu.scala 63:30]
  wire [3:0] dccm_ctl_io_stbuf_fwdbyteen_hi_m; // @[lsu.scala 63:30]
  wire [31:0] dccm_ctl_io_lsu_ld_data_corr_r; // @[lsu.scala 63:30]
  wire  dccm_ctl_io_lsu_double_ecc_error_r; // @[lsu.scala 63:30]
  wire  dccm_ctl_io_single_ecc_error_hi_r; // @[lsu.scala 63:30]
  wire  dccm_ctl_io_single_ecc_error_lo_r; // @[lsu.scala 63:30]
  wire [31:0] dccm_ctl_io_sec_data_hi_r_ff; // @[lsu.scala 63:30]
  wire [31:0] dccm_ctl_io_sec_data_lo_r_ff; // @[lsu.scala 63:30]
  wire [6:0] dccm_ctl_io_sec_data_ecc_hi_r_ff; // @[lsu.scala 63:30]
  wire [6:0] dccm_ctl_io_sec_data_ecc_lo_r_ff; // @[lsu.scala 63:30]
  wire [31:0] dccm_ctl_io_dccm_rdata_hi_m; // @[lsu.scala 63:30]
  wire [31:0] dccm_ctl_io_dccm_rdata_lo_m; // @[lsu.scala 63:30]
  wire [6:0] dccm_ctl_io_dccm_data_ecc_hi_m; // @[lsu.scala 63:30]
  wire [6:0] dccm_ctl_io_dccm_data_ecc_lo_m; // @[lsu.scala 63:30]
  wire [31:0] dccm_ctl_io_lsu_ld_data_m; // @[lsu.scala 63:30]
  wire  dccm_ctl_io_lsu_double_ecc_error_m; // @[lsu.scala 63:30]
  wire [31:0] dccm_ctl_io_sec_data_hi_m; // @[lsu.scala 63:30]
  wire [31:0] dccm_ctl_io_sec_data_lo_m; // @[lsu.scala 63:30]
  wire [31:0] dccm_ctl_io_store_data_m; // @[lsu.scala 63:30]
  wire  dccm_ctl_io_dma_dccm_wen; // @[lsu.scala 63:30]
  wire  dccm_ctl_io_dma_pic_wen; // @[lsu.scala 63:30]
  wire [2:0] dccm_ctl_io_dma_mem_tag_m; // @[lsu.scala 63:30]
  wire [31:0] dccm_ctl_io_dma_dccm_wdata_lo; // @[lsu.scala 63:30]
  wire [31:0] dccm_ctl_io_dma_dccm_wdata_hi; // @[lsu.scala 63:30]
  wire [6:0] dccm_ctl_io_dma_dccm_wdata_ecc_hi; // @[lsu.scala 63:30]
  wire [6:0] dccm_ctl_io_dma_dccm_wdata_ecc_lo; // @[lsu.scala 63:30]
  wire [31:0] dccm_ctl_io_store_data_hi_r; // @[lsu.scala 63:30]
  wire [31:0] dccm_ctl_io_store_data_lo_r; // @[lsu.scala 63:30]
  wire [31:0] dccm_ctl_io_store_datafn_hi_r; // @[lsu.scala 63:30]
  wire [31:0] dccm_ctl_io_store_datafn_lo_r; // @[lsu.scala 63:30]
  wire [31:0] dccm_ctl_io_store_data_r; // @[lsu.scala 63:30]
  wire  dccm_ctl_io_ld_single_ecc_error_r; // @[lsu.scala 63:30]
  wire  dccm_ctl_io_ld_single_ecc_error_r_ff; // @[lsu.scala 63:30]
  wire [31:0] dccm_ctl_io_picm_mask_data_m; // @[lsu.scala 63:30]
  wire  dccm_ctl_io_lsu_stbuf_commit_any; // @[lsu.scala 63:30]
  wire  dccm_ctl_io_lsu_dccm_rden_m; // @[lsu.scala 63:30]
  wire [31:0] dccm_ctl_io_dma_dccm_ctl_dma_mem_addr; // @[lsu.scala 63:30]
  wire [63:0] dccm_ctl_io_dma_dccm_ctl_dma_mem_wdata; // @[lsu.scala 63:30]
  wire  dccm_ctl_io_dma_dccm_ctl_dccm_dma_rvalid; // @[lsu.scala 63:30]
  wire  dccm_ctl_io_dma_dccm_ctl_dccm_dma_ecc_error; // @[lsu.scala 63:30]
  wire [2:0] dccm_ctl_io_dma_dccm_ctl_dccm_dma_rtag; // @[lsu.scala 63:30]
  wire [63:0] dccm_ctl_io_dma_dccm_ctl_dccm_dma_rdata; // @[lsu.scala 63:30]
  wire  dccm_ctl_io_dccm_wren; // @[lsu.scala 63:30]
  wire  dccm_ctl_io_dccm_rden; // @[lsu.scala 63:30]
  wire [15:0] dccm_ctl_io_dccm_wr_addr_lo; // @[lsu.scala 63:30]
  wire [15:0] dccm_ctl_io_dccm_wr_addr_hi; // @[lsu.scala 63:30]
  wire [15:0] dccm_ctl_io_dccm_rd_addr_lo; // @[lsu.scala 63:30]
  wire [15:0] dccm_ctl_io_dccm_rd_addr_hi; // @[lsu.scala 63:30]
  wire [38:0] dccm_ctl_io_dccm_wr_data_lo; // @[lsu.scala 63:30]
  wire [38:0] dccm_ctl_io_dccm_wr_data_hi; // @[lsu.scala 63:30]
  wire [38:0] dccm_ctl_io_dccm_rd_data_lo; // @[lsu.scala 63:30]
  wire [38:0] dccm_ctl_io_dccm_rd_data_hi; // @[lsu.scala 63:30]
  wire  dccm_ctl_io_lsu_pic_picm_wren; // @[lsu.scala 63:30]
  wire  dccm_ctl_io_lsu_pic_picm_rden; // @[lsu.scala 63:30]
  wire  dccm_ctl_io_lsu_pic_picm_mken; // @[lsu.scala 63:30]
  wire [31:0] dccm_ctl_io_lsu_pic_picm_rdaddr; // @[lsu.scala 63:30]
  wire [31:0] dccm_ctl_io_lsu_pic_picm_wraddr; // @[lsu.scala 63:30]
  wire [31:0] dccm_ctl_io_lsu_pic_picm_wr_data; // @[lsu.scala 63:30]
  wire [31:0] dccm_ctl_io_lsu_pic_picm_rd_data; // @[lsu.scala 63:30]
  wire  dccm_ctl_io_scan_mode; // @[lsu.scala 63:30]
  wire  stbuf_clock; // @[lsu.scala 64:30]
  wire  stbuf_reset; // @[lsu.scala 64:30]
  wire  stbuf_io_lsu_c1_m_clk; // @[lsu.scala 64:30]
  wire  stbuf_io_lsu_c1_r_clk; // @[lsu.scala 64:30]
  wire  stbuf_io_lsu_stbuf_c1_clk; // @[lsu.scala 64:30]
  wire  stbuf_io_lsu_free_c2_clk; // @[lsu.scala 64:30]
  wire  stbuf_io_lsu_pkt_m_valid; // @[lsu.scala 64:30]
  wire  stbuf_io_lsu_pkt_m_bits_store; // @[lsu.scala 64:30]
  wire  stbuf_io_lsu_pkt_m_bits_dma; // @[lsu.scala 64:30]
  wire  stbuf_io_lsu_pkt_r_valid; // @[lsu.scala 64:30]
  wire  stbuf_io_lsu_pkt_r_bits_by; // @[lsu.scala 64:30]
  wire  stbuf_io_lsu_pkt_r_bits_half; // @[lsu.scala 64:30]
  wire  stbuf_io_lsu_pkt_r_bits_word; // @[lsu.scala 64:30]
  wire  stbuf_io_lsu_pkt_r_bits_dword; // @[lsu.scala 64:30]
  wire  stbuf_io_lsu_pkt_r_bits_store; // @[lsu.scala 64:30]
  wire  stbuf_io_lsu_pkt_r_bits_dma; // @[lsu.scala 64:30]
  wire  stbuf_io_store_stbuf_reqvld_r; // @[lsu.scala 64:30]
  wire  stbuf_io_lsu_commit_r; // @[lsu.scala 64:30]
  wire  stbuf_io_dec_lsu_valid_raw_d; // @[lsu.scala 64:30]
  wire [31:0] stbuf_io_store_data_hi_r; // @[lsu.scala 64:30]
  wire [31:0] stbuf_io_store_data_lo_r; // @[lsu.scala 64:30]
  wire [31:0] stbuf_io_store_datafn_hi_r; // @[lsu.scala 64:30]
  wire [31:0] stbuf_io_store_datafn_lo_r; // @[lsu.scala 64:30]
  wire  stbuf_io_lsu_stbuf_commit_any; // @[lsu.scala 64:30]
  wire [15:0] stbuf_io_lsu_addr_d; // @[lsu.scala 64:30]
  wire [31:0] stbuf_io_lsu_addr_m; // @[lsu.scala 64:30]
  wire [31:0] stbuf_io_lsu_addr_r; // @[lsu.scala 64:30]
  wire [15:0] stbuf_io_end_addr_d; // @[lsu.scala 64:30]
  wire [31:0] stbuf_io_end_addr_m; // @[lsu.scala 64:30]
  wire [31:0] stbuf_io_end_addr_r; // @[lsu.scala 64:30]
  wire  stbuf_io_addr_in_dccm_m; // @[lsu.scala 64:30]
  wire  stbuf_io_addr_in_dccm_r; // @[lsu.scala 64:30]
  wire  stbuf_io_scan_mode; // @[lsu.scala 64:30]
  wire  stbuf_io_stbuf_reqvld_any; // @[lsu.scala 64:30]
  wire  stbuf_io_stbuf_reqvld_flushed_any; // @[lsu.scala 64:30]
  wire [15:0] stbuf_io_stbuf_addr_any; // @[lsu.scala 64:30]
  wire [31:0] stbuf_io_stbuf_data_any; // @[lsu.scala 64:30]
  wire  stbuf_io_lsu_stbuf_full_any; // @[lsu.scala 64:30]
  wire  stbuf_io_lsu_stbuf_empty_any; // @[lsu.scala 64:30]
  wire  stbuf_io_ldst_stbuf_reqvld_r; // @[lsu.scala 64:30]
  wire [31:0] stbuf_io_stbuf_fwddata_hi_m; // @[lsu.scala 64:30]
  wire [31:0] stbuf_io_stbuf_fwddata_lo_m; // @[lsu.scala 64:30]
  wire [3:0] stbuf_io_stbuf_fwdbyteen_hi_m; // @[lsu.scala 64:30]
  wire [3:0] stbuf_io_stbuf_fwdbyteen_lo_m; // @[lsu.scala 64:30]
  wire  ecc_clock; // @[lsu.scala 65:30]
  wire  ecc_reset; // @[lsu.scala 65:30]
  wire  ecc_io_lsu_c2_r_clk; // @[lsu.scala 65:30]
  wire  ecc_io_lsu_pkt_m_valid; // @[lsu.scala 65:30]
  wire  ecc_io_lsu_pkt_m_bits_load; // @[lsu.scala 65:30]
  wire  ecc_io_lsu_pkt_m_bits_store; // @[lsu.scala 65:30]
  wire  ecc_io_lsu_pkt_m_bits_dma; // @[lsu.scala 65:30]
  wire [31:0] ecc_io_stbuf_data_any; // @[lsu.scala 65:30]
  wire  ecc_io_dec_tlu_core_ecc_disable; // @[lsu.scala 65:30]
  wire [15:0] ecc_io_lsu_addr_m; // @[lsu.scala 65:30]
  wire [15:0] ecc_io_end_addr_m; // @[lsu.scala 65:30]
  wire [31:0] ecc_io_dccm_rdata_hi_m; // @[lsu.scala 65:30]
  wire [31:0] ecc_io_dccm_rdata_lo_m; // @[lsu.scala 65:30]
  wire [6:0] ecc_io_dccm_data_ecc_hi_m; // @[lsu.scala 65:30]
  wire [6:0] ecc_io_dccm_data_ecc_lo_m; // @[lsu.scala 65:30]
  wire  ecc_io_ld_single_ecc_error_r; // @[lsu.scala 65:30]
  wire  ecc_io_ld_single_ecc_error_r_ff; // @[lsu.scala 65:30]
  wire  ecc_io_lsu_dccm_rden_m; // @[lsu.scala 65:30]
  wire  ecc_io_addr_in_dccm_m; // @[lsu.scala 65:30]
  wire  ecc_io_dma_dccm_wen; // @[lsu.scala 65:30]
  wire [31:0] ecc_io_dma_dccm_wdata_lo; // @[lsu.scala 65:30]
  wire [31:0] ecc_io_dma_dccm_wdata_hi; // @[lsu.scala 65:30]
  wire  ecc_io_scan_mode; // @[lsu.scala 65:30]
  wire [31:0] ecc_io_sec_data_hi_r; // @[lsu.scala 65:30]
  wire [31:0] ecc_io_sec_data_lo_r; // @[lsu.scala 65:30]
  wire [31:0] ecc_io_sec_data_hi_m; // @[lsu.scala 65:30]
  wire [31:0] ecc_io_sec_data_lo_m; // @[lsu.scala 65:30]
  wire [31:0] ecc_io_sec_data_hi_r_ff; // @[lsu.scala 65:30]
  wire [31:0] ecc_io_sec_data_lo_r_ff; // @[lsu.scala 65:30]
  wire [6:0] ecc_io_dma_dccm_wdata_ecc_hi; // @[lsu.scala 65:30]
  wire [6:0] ecc_io_dma_dccm_wdata_ecc_lo; // @[lsu.scala 65:30]
  wire [6:0] ecc_io_stbuf_ecc_any; // @[lsu.scala 65:30]
  wire [6:0] ecc_io_sec_data_ecc_hi_r_ff; // @[lsu.scala 65:30]
  wire [6:0] ecc_io_sec_data_ecc_lo_r_ff; // @[lsu.scala 65:30]
  wire  ecc_io_single_ecc_error_hi_r; // @[lsu.scala 65:30]
  wire  ecc_io_single_ecc_error_lo_r; // @[lsu.scala 65:30]
  wire  ecc_io_lsu_single_ecc_error_r; // @[lsu.scala 65:30]
  wire  ecc_io_lsu_double_ecc_error_r; // @[lsu.scala 65:30]
  wire  ecc_io_lsu_single_ecc_error_m; // @[lsu.scala 65:30]
  wire  ecc_io_lsu_double_ecc_error_m; // @[lsu.scala 65:30]
  wire  trigger_io_trigger_pkt_any_0_select; // @[lsu.scala 66:30]
  wire  trigger_io_trigger_pkt_any_0_match_pkt; // @[lsu.scala 66:30]
  wire  trigger_io_trigger_pkt_any_0_store; // @[lsu.scala 66:30]
  wire  trigger_io_trigger_pkt_any_0_load; // @[lsu.scala 66:30]
  wire [31:0] trigger_io_trigger_pkt_any_0_tdata2; // @[lsu.scala 66:30]
  wire  trigger_io_trigger_pkt_any_1_select; // @[lsu.scala 66:30]
  wire  trigger_io_trigger_pkt_any_1_match_pkt; // @[lsu.scala 66:30]
  wire  trigger_io_trigger_pkt_any_1_store; // @[lsu.scala 66:30]
  wire  trigger_io_trigger_pkt_any_1_load; // @[lsu.scala 66:30]
  wire [31:0] trigger_io_trigger_pkt_any_1_tdata2; // @[lsu.scala 66:30]
  wire  trigger_io_trigger_pkt_any_2_select; // @[lsu.scala 66:30]
  wire  trigger_io_trigger_pkt_any_2_match_pkt; // @[lsu.scala 66:30]
  wire  trigger_io_trigger_pkt_any_2_store; // @[lsu.scala 66:30]
  wire  trigger_io_trigger_pkt_any_2_load; // @[lsu.scala 66:30]
  wire [31:0] trigger_io_trigger_pkt_any_2_tdata2; // @[lsu.scala 66:30]
  wire  trigger_io_trigger_pkt_any_3_select; // @[lsu.scala 66:30]
  wire  trigger_io_trigger_pkt_any_3_match_pkt; // @[lsu.scala 66:30]
  wire  trigger_io_trigger_pkt_any_3_store; // @[lsu.scala 66:30]
  wire  trigger_io_trigger_pkt_any_3_load; // @[lsu.scala 66:30]
  wire [31:0] trigger_io_trigger_pkt_any_3_tdata2; // @[lsu.scala 66:30]
  wire  trigger_io_lsu_pkt_m_valid; // @[lsu.scala 66:30]
  wire  trigger_io_lsu_pkt_m_bits_half; // @[lsu.scala 66:30]
  wire  trigger_io_lsu_pkt_m_bits_word; // @[lsu.scala 66:30]
  wire  trigger_io_lsu_pkt_m_bits_load; // @[lsu.scala 66:30]
  wire  trigger_io_lsu_pkt_m_bits_store; // @[lsu.scala 66:30]
  wire  trigger_io_lsu_pkt_m_bits_dma; // @[lsu.scala 66:30]
  wire [31:0] trigger_io_lsu_addr_m; // @[lsu.scala 66:30]
  wire [31:0] trigger_io_store_data_m; // @[lsu.scala 66:30]
  wire [3:0] trigger_io_lsu_trigger_match_m; // @[lsu.scala 66:30]
  wire  clkdomain_clock; // @[lsu.scala 67:30]
  wire  clkdomain_reset; // @[lsu.scala 67:30]
  wire  clkdomain_io_free_clk; // @[lsu.scala 67:30]
  wire  clkdomain_io_clk_override; // @[lsu.scala 67:30]
  wire  clkdomain_io_dma_dccm_req; // @[lsu.scala 67:30]
  wire  clkdomain_io_ldst_stbuf_reqvld_r; // @[lsu.scala 67:30]
  wire  clkdomain_io_stbuf_reqvld_any; // @[lsu.scala 67:30]
  wire  clkdomain_io_stbuf_reqvld_flushed_any; // @[lsu.scala 67:30]
  wire  clkdomain_io_lsu_busreq_r; // @[lsu.scala 67:30]
  wire  clkdomain_io_lsu_bus_buffer_pend_any; // @[lsu.scala 67:30]
  wire  clkdomain_io_lsu_bus_buffer_empty_any; // @[lsu.scala 67:30]
  wire  clkdomain_io_lsu_stbuf_empty_any; // @[lsu.scala 67:30]
  wire  clkdomain_io_lsu_bus_clk_en; // @[lsu.scala 67:30]
  wire  clkdomain_io_lsu_p_valid; // @[lsu.scala 67:30]
  wire  clkdomain_io_lsu_pkt_d_valid; // @[lsu.scala 67:30]
  wire  clkdomain_io_lsu_pkt_d_bits_store; // @[lsu.scala 67:30]
  wire  clkdomain_io_lsu_pkt_m_valid; // @[lsu.scala 67:30]
  wire  clkdomain_io_lsu_pkt_m_bits_store; // @[lsu.scala 67:30]
  wire  clkdomain_io_lsu_pkt_r_valid; // @[lsu.scala 67:30]
  wire  clkdomain_io_lsu_c1_m_clk; // @[lsu.scala 67:30]
  wire  clkdomain_io_lsu_c1_r_clk; // @[lsu.scala 67:30]
  wire  clkdomain_io_lsu_c2_m_clk; // @[lsu.scala 67:30]
  wire  clkdomain_io_lsu_c2_r_clk; // @[lsu.scala 67:30]
  wire  clkdomain_io_lsu_store_c1_m_clk; // @[lsu.scala 67:30]
  wire  clkdomain_io_lsu_store_c1_r_clk; // @[lsu.scala 67:30]
  wire  clkdomain_io_lsu_stbuf_c1_clk; // @[lsu.scala 67:30]
  wire  clkdomain_io_lsu_bus_obuf_c1_clk; // @[lsu.scala 67:30]
  wire  clkdomain_io_lsu_bus_ibuf_c1_clk; // @[lsu.scala 67:30]
  wire  clkdomain_io_lsu_bus_buf_c1_clk; // @[lsu.scala 67:30]
  wire  clkdomain_io_lsu_busm_clk; // @[lsu.scala 67:30]
  wire  clkdomain_io_lsu_free_c2_clk; // @[lsu.scala 67:30]
  wire  clkdomain_io_scan_mode; // @[lsu.scala 67:30]
  wire  bus_intf_clock; // @[lsu.scala 68:30]
  wire  bus_intf_reset; // @[lsu.scala 68:30]
  wire  bus_intf_io_scan_mode; // @[lsu.scala 68:30]
  wire  bus_intf_io_tlu_busbuff_lsu_pmu_bus_misaligned; // @[lsu.scala 68:30]
  wire  bus_intf_io_tlu_busbuff_lsu_pmu_bus_error; // @[lsu.scala 68:30]
  wire  bus_intf_io_tlu_busbuff_lsu_pmu_bus_busy; // @[lsu.scala 68:30]
  wire  bus_intf_io_tlu_busbuff_dec_tlu_external_ldfwd_disable; // @[lsu.scala 68:30]
  wire  bus_intf_io_tlu_busbuff_dec_tlu_wb_coalescing_disable; // @[lsu.scala 68:30]
  wire  bus_intf_io_tlu_busbuff_dec_tlu_sideeffect_posted_disable; // @[lsu.scala 68:30]
  wire  bus_intf_io_tlu_busbuff_lsu_imprecise_error_load_any; // @[lsu.scala 68:30]
  wire  bus_intf_io_tlu_busbuff_lsu_imprecise_error_store_any; // @[lsu.scala 68:30]
  wire [31:0] bus_intf_io_tlu_busbuff_lsu_imprecise_error_addr_any; // @[lsu.scala 68:30]
  wire  bus_intf_io_lsu_c1_m_clk; // @[lsu.scala 68:30]
  wire  bus_intf_io_lsu_c1_r_clk; // @[lsu.scala 68:30]
  wire  bus_intf_io_lsu_c2_r_clk; // @[lsu.scala 68:30]
  wire  bus_intf_io_lsu_bus_ibuf_c1_clk; // @[lsu.scala 68:30]
  wire  bus_intf_io_lsu_bus_obuf_c1_clk; // @[lsu.scala 68:30]
  wire  bus_intf_io_lsu_bus_buf_c1_clk; // @[lsu.scala 68:30]
  wire  bus_intf_io_lsu_free_c2_clk; // @[lsu.scala 68:30]
  wire  bus_intf_io_free_clk; // @[lsu.scala 68:30]
  wire  bus_intf_io_lsu_busm_clk; // @[lsu.scala 68:30]
  wire  bus_intf_io_axi_aw_valid; // @[lsu.scala 68:30]
  wire [31:0] bus_intf_io_axi_aw_bits_addr; // @[lsu.scala 68:30]
  wire [2:0] bus_intf_io_axi_aw_bits_size; // @[lsu.scala 68:30]
  wire  bus_intf_io_axi_w_valid; // @[lsu.scala 68:30]
  wire [7:0] bus_intf_io_axi_w_bits_strb; // @[lsu.scala 68:30]
  wire  bus_intf_io_axi_ar_valid; // @[lsu.scala 68:30]
  wire [31:0] bus_intf_io_axi_ar_bits_addr; // @[lsu.scala 68:30]
  wire [2:0] bus_intf_io_axi_ar_bits_size; // @[lsu.scala 68:30]
  wire  bus_intf_io_dec_lsu_valid_raw_d; // @[lsu.scala 68:30]
  wire  bus_intf_io_lsu_busreq_m; // @[lsu.scala 68:30]
  wire  bus_intf_io_lsu_pkt_m_valid; // @[lsu.scala 68:30]
  wire  bus_intf_io_lsu_pkt_m_bits_by; // @[lsu.scala 68:30]
  wire  bus_intf_io_lsu_pkt_m_bits_half; // @[lsu.scala 68:30]
  wire  bus_intf_io_lsu_pkt_m_bits_word; // @[lsu.scala 68:30]
  wire  bus_intf_io_lsu_pkt_m_bits_load; // @[lsu.scala 68:30]
  wire  bus_intf_io_lsu_pkt_r_valid; // @[lsu.scala 68:30]
  wire  bus_intf_io_lsu_pkt_r_bits_by; // @[lsu.scala 68:30]
  wire  bus_intf_io_lsu_pkt_r_bits_half; // @[lsu.scala 68:30]
  wire  bus_intf_io_lsu_pkt_r_bits_word; // @[lsu.scala 68:30]
  wire  bus_intf_io_lsu_pkt_r_bits_load; // @[lsu.scala 68:30]
  wire  bus_intf_io_lsu_pkt_r_bits_store; // @[lsu.scala 68:30]
  wire  bus_intf_io_lsu_pkt_r_bits_unsign; // @[lsu.scala 68:30]
  wire [31:0] bus_intf_io_lsu_addr_d; // @[lsu.scala 68:30]
  wire [31:0] bus_intf_io_lsu_addr_m; // @[lsu.scala 68:30]
  wire [31:0] bus_intf_io_lsu_addr_r; // @[lsu.scala 68:30]
  wire [31:0] bus_intf_io_end_addr_d; // @[lsu.scala 68:30]
  wire [31:0] bus_intf_io_end_addr_m; // @[lsu.scala 68:30]
  wire [31:0] bus_intf_io_end_addr_r; // @[lsu.scala 68:30]
  wire [31:0] bus_intf_io_store_data_r; // @[lsu.scala 68:30]
  wire  bus_intf_io_dec_tlu_force_halt; // @[lsu.scala 68:30]
  wire  bus_intf_io_lsu_commit_r; // @[lsu.scala 68:30]
  wire  bus_intf_io_is_sideeffects_m; // @[lsu.scala 68:30]
  wire  bus_intf_io_flush_m_up; // @[lsu.scala 68:30]
  wire  bus_intf_io_flush_r; // @[lsu.scala 68:30]
  wire  bus_intf_io_lsu_busreq_r; // @[lsu.scala 68:30]
  wire  bus_intf_io_lsu_bus_buffer_pend_any; // @[lsu.scala 68:30]
  wire  bus_intf_io_lsu_bus_buffer_full_any; // @[lsu.scala 68:30]
  wire  bus_intf_io_lsu_bus_buffer_empty_any; // @[lsu.scala 68:30]
  wire [31:0] bus_intf_io_bus_read_data_m; // @[lsu.scala 68:30]
  wire  bus_intf_io_dctl_busbuff_lsu_nonblock_load_valid_m; // @[lsu.scala 68:30]
  wire [1:0] bus_intf_io_dctl_busbuff_lsu_nonblock_load_tag_m; // @[lsu.scala 68:30]
  wire  bus_intf_io_dctl_busbuff_lsu_nonblock_load_inv_r; // @[lsu.scala 68:30]
  wire [1:0] bus_intf_io_dctl_busbuff_lsu_nonblock_load_inv_tag_r; // @[lsu.scala 68:30]
  wire  bus_intf_io_dctl_busbuff_lsu_nonblock_load_data_valid; // @[lsu.scala 68:30]
  wire  bus_intf_io_dctl_busbuff_lsu_nonblock_load_data_error; // @[lsu.scala 68:30]
  wire [1:0] bus_intf_io_dctl_busbuff_lsu_nonblock_load_data_tag; // @[lsu.scala 68:30]
  wire [31:0] bus_intf_io_dctl_busbuff_lsu_nonblock_load_data; // @[lsu.scala 68:30]
  wire  bus_intf_io_lsu_bus_clk_en; // @[lsu.scala 68:30]
  wire  _T = stbuf_io_lsu_stbuf_full_any | bus_intf_io_lsu_bus_buffer_full_any; // @[lsu.scala 74:57]
  wire  _T_3 = ~lsu_lsc_ctl_io_lsu_pkt_m_bits_dma; // @[lsu.scala 81:58]
  wire  _T_4 = lsu_lsc_ctl_io_lsu_pkt_m_valid & _T_3; // @[lsu.scala 81:56]
  wire  _T_5 = lsu_lsc_ctl_io_addr_in_dccm_m | lsu_lsc_ctl_io_addr_in_pic_m; // @[lsu.scala 81:126]
  wire  _T_6 = _T_4 & _T_5; // @[lsu.scala 81:93]
  wire  ldst_nodma_mtor = _T_6 & lsu_lsc_ctl_io_lsu_pkt_m_bits_store; // @[lsu.scala 81:158]
  wire  _T_7 = io_dec_lsu_valid_raw_d | ldst_nodma_mtor; // @[lsu.scala 82:53]
  wire  _T_8 = _T_7 | dccm_ctl_io_ld_single_ecc_error_r_ff; // @[lsu.scala 82:71]
  wire  _T_10 = io_lsu_dma_dma_lsc_ctl_dma_dccm_req & io_lsu_dma_dma_lsc_ctl_dma_mem_write; // @[lsu.scala 83:58]
  wire [5:0] _T_13 = {io_lsu_dma_dma_lsc_ctl_dma_mem_addr[2:0],3'h0}; // @[Cat.scala 29:58]
  wire [63:0] dma_dccm_wdata = io_lsu_dma_dma_lsc_ctl_dma_mem_wdata >> _T_13; // @[lsu.scala 85:58]
  wire  _T_19 = ~lsu_lsc_ctl_io_lsu_pkt_r_bits_dma; // @[lsu.scala 96:130]
  wire  _T_20 = lsu_lsc_ctl_io_lsu_pkt_r_valid & _T_19; // @[lsu.scala 96:128]
  wire  _T_21 = _T_4 | _T_20; // @[lsu.scala 96:94]
  wire  _T_22 = ~_T_21; // @[lsu.scala 96:22]
  wire  _T_25 = lsu_lsc_ctl_io_lsu_pkt_r_valid & lsu_lsc_ctl_io_lsu_pkt_r_bits_store; // @[lsu.scala 98:61]
  wire  _T_26 = _T_25 & lsu_lsc_ctl_io_addr_in_dccm_r; // @[lsu.scala 98:99]
  wire  _T_27 = ~io_dec_tlu_i0_kill_writeb_r; // @[lsu.scala 98:133]
  wire  _T_28 = _T_26 & _T_27; // @[lsu.scala 98:131]
  wire  _T_30 = lsu_lsc_ctl_io_lsu_pkt_m_bits_load | lsu_lsc_ctl_io_lsu_pkt_m_bits_store; // @[lsu.scala 100:90]
  wire  _T_34 = _T_30 & lsu_lsc_ctl_io_addr_external_m; // @[lsu.scala 102:131]
  wire  _T_35 = lsu_lsc_ctl_io_lsu_pkt_m_valid & _T_34; // @[lsu.scala 102:53]
  wire  _T_36 = ~io_dec_tlu_flush_lower_r; // @[lsu.scala 102:167]
  wire  _T_37 = _T_35 & _T_36; // @[lsu.scala 102:165]
  wire  _T_38 = ~lsu_lsc_ctl_io_lsu_exc_m; // @[lsu.scala 102:181]
  wire  _T_39 = _T_37 & _T_38; // @[lsu.scala 102:179]
  wire  _T_40 = ~lsu_lsc_ctl_io_lsu_pkt_m_bits_fast_int; // @[lsu.scala 102:209]
  wire  _T_42 = lsu_lsc_ctl_io_lsu_pkt_m_bits_half & lsu_lsc_ctl_io_lsu_addr_m[0]; // @[lsu.scala 104:100]
  wire  _T_44 = |lsu_lsc_ctl_io_lsu_addr_m[1:0]; // @[lsu.scala 104:203]
  wire  _T_45 = lsu_lsc_ctl_io_lsu_pkt_m_bits_word & _T_44; // @[lsu.scala 104:170]
  wire  _T_46 = _T_42 | _T_45; // @[lsu.scala 104:132]
  wire  _T_48 = lsu_lsc_ctl_io_lsu_pkt_m_valid & lsu_lsc_ctl_io_lsu_pkt_m_bits_load; // @[lsu.scala 105:73]
  wire  _T_50 = lsu_lsc_ctl_io_lsu_pkt_m_valid & lsu_lsc_ctl_io_lsu_pkt_m_bits_store; // @[lsu.scala 106:73]
  reg [2:0] dma_mem_tag_m; // @[lsu.scala 317:67]
  reg  lsu_raw_fwd_hi_r; // @[lsu.scala 318:67]
  reg  lsu_raw_fwd_lo_r; // @[lsu.scala 319:67]
  lsu_lsc_ctl lsu_lsc_ctl ( // @[lsu.scala 60:30]
    .reset(lsu_lsc_ctl_reset),
    .io_lsu_c1_m_clk(lsu_lsc_ctl_io_lsu_c1_m_clk),
    .io_lsu_c1_r_clk(lsu_lsc_ctl_io_lsu_c1_r_clk),
    .io_lsu_c2_m_clk(lsu_lsc_ctl_io_lsu_c2_m_clk),
    .io_lsu_c2_r_clk(lsu_lsc_ctl_io_lsu_c2_r_clk),
    .io_lsu_store_c1_m_clk(lsu_lsc_ctl_io_lsu_store_c1_m_clk),
    .io_lsu_ld_data_corr_r(lsu_lsc_ctl_io_lsu_ld_data_corr_r),
    .io_lsu_single_ecc_error_r(lsu_lsc_ctl_io_lsu_single_ecc_error_r),
    .io_lsu_double_ecc_error_r(lsu_lsc_ctl_io_lsu_double_ecc_error_r),
    .io_lsu_ld_data_m(lsu_lsc_ctl_io_lsu_ld_data_m),
    .io_lsu_single_ecc_error_m(lsu_lsc_ctl_io_lsu_single_ecc_error_m),
    .io_lsu_double_ecc_error_m(lsu_lsc_ctl_io_lsu_double_ecc_error_m),
    .io_flush_m_up(lsu_lsc_ctl_io_flush_m_up),
    .io_flush_r(lsu_lsc_ctl_io_flush_r),
    .io_lsu_exu_exu_lsu_rs1_d(lsu_lsc_ctl_io_lsu_exu_exu_lsu_rs1_d),
    .io_lsu_exu_exu_lsu_rs2_d(lsu_lsc_ctl_io_lsu_exu_exu_lsu_rs2_d),
    .io_lsu_p_valid(lsu_lsc_ctl_io_lsu_p_valid),
    .io_lsu_p_bits_fast_int(lsu_lsc_ctl_io_lsu_p_bits_fast_int),
    .io_lsu_p_bits_by(lsu_lsc_ctl_io_lsu_p_bits_by),
    .io_lsu_p_bits_half(lsu_lsc_ctl_io_lsu_p_bits_half),
    .io_lsu_p_bits_word(lsu_lsc_ctl_io_lsu_p_bits_word),
    .io_lsu_p_bits_load(lsu_lsc_ctl_io_lsu_p_bits_load),
    .io_lsu_p_bits_store(lsu_lsc_ctl_io_lsu_p_bits_store),
    .io_lsu_p_bits_unsign(lsu_lsc_ctl_io_lsu_p_bits_unsign),
    .io_lsu_p_bits_store_data_bypass_d(lsu_lsc_ctl_io_lsu_p_bits_store_data_bypass_d),
    .io_lsu_p_bits_load_ldst_bypass_d(lsu_lsc_ctl_io_lsu_p_bits_load_ldst_bypass_d),
    .io_dec_lsu_valid_raw_d(lsu_lsc_ctl_io_dec_lsu_valid_raw_d),
    .io_dec_lsu_offset_d(lsu_lsc_ctl_io_dec_lsu_offset_d),
    .io_picm_mask_data_m(lsu_lsc_ctl_io_picm_mask_data_m),
    .io_bus_read_data_m(lsu_lsc_ctl_io_bus_read_data_m),
    .io_lsu_result_m(lsu_lsc_ctl_io_lsu_result_m),
    .io_lsu_result_corr_r(lsu_lsc_ctl_io_lsu_result_corr_r),
    .io_lsu_addr_d(lsu_lsc_ctl_io_lsu_addr_d),
    .io_lsu_addr_m(lsu_lsc_ctl_io_lsu_addr_m),
    .io_lsu_addr_r(lsu_lsc_ctl_io_lsu_addr_r),
    .io_end_addr_d(lsu_lsc_ctl_io_end_addr_d),
    .io_end_addr_m(lsu_lsc_ctl_io_end_addr_m),
    .io_end_addr_r(lsu_lsc_ctl_io_end_addr_r),
    .io_store_data_m(lsu_lsc_ctl_io_store_data_m),
    .io_dec_tlu_mrac_ff(lsu_lsc_ctl_io_dec_tlu_mrac_ff),
    .io_lsu_exc_m(lsu_lsc_ctl_io_lsu_exc_m),
    .io_is_sideeffects_m(lsu_lsc_ctl_io_is_sideeffects_m),
    .io_lsu_commit_r(lsu_lsc_ctl_io_lsu_commit_r),
    .io_lsu_single_ecc_error_incr(lsu_lsc_ctl_io_lsu_single_ecc_error_incr),
    .io_lsu_error_pkt_r_valid(lsu_lsc_ctl_io_lsu_error_pkt_r_valid),
    .io_lsu_error_pkt_r_bits_single_ecc_error(lsu_lsc_ctl_io_lsu_error_pkt_r_bits_single_ecc_error),
    .io_lsu_error_pkt_r_bits_inst_type(lsu_lsc_ctl_io_lsu_error_pkt_r_bits_inst_type),
    .io_lsu_error_pkt_r_bits_exc_type(lsu_lsc_ctl_io_lsu_error_pkt_r_bits_exc_type),
    .io_lsu_error_pkt_r_bits_mscause(lsu_lsc_ctl_io_lsu_error_pkt_r_bits_mscause),
    .io_lsu_error_pkt_r_bits_addr(lsu_lsc_ctl_io_lsu_error_pkt_r_bits_addr),
    .io_lsu_fir_addr(lsu_lsc_ctl_io_lsu_fir_addr),
    .io_lsu_fir_error(lsu_lsc_ctl_io_lsu_fir_error),
    .io_addr_in_dccm_d(lsu_lsc_ctl_io_addr_in_dccm_d),
    .io_addr_in_dccm_m(lsu_lsc_ctl_io_addr_in_dccm_m),
    .io_addr_in_dccm_r(lsu_lsc_ctl_io_addr_in_dccm_r),
    .io_addr_in_pic_d(lsu_lsc_ctl_io_addr_in_pic_d),
    .io_addr_in_pic_m(lsu_lsc_ctl_io_addr_in_pic_m),
    .io_addr_in_pic_r(lsu_lsc_ctl_io_addr_in_pic_r),
    .io_addr_external_m(lsu_lsc_ctl_io_addr_external_m),
    .io_dma_lsc_ctl_dma_dccm_req(lsu_lsc_ctl_io_dma_lsc_ctl_dma_dccm_req),
    .io_dma_lsc_ctl_dma_mem_addr(lsu_lsc_ctl_io_dma_lsc_ctl_dma_mem_addr),
    .io_dma_lsc_ctl_dma_mem_sz(lsu_lsc_ctl_io_dma_lsc_ctl_dma_mem_sz),
    .io_dma_lsc_ctl_dma_mem_write(lsu_lsc_ctl_io_dma_lsc_ctl_dma_mem_write),
    .io_dma_lsc_ctl_dma_mem_wdata(lsu_lsc_ctl_io_dma_lsc_ctl_dma_mem_wdata),
    .io_lsu_pkt_d_valid(lsu_lsc_ctl_io_lsu_pkt_d_valid),
    .io_lsu_pkt_d_bits_fast_int(lsu_lsc_ctl_io_lsu_pkt_d_bits_fast_int),
    .io_lsu_pkt_d_bits_by(lsu_lsc_ctl_io_lsu_pkt_d_bits_by),
    .io_lsu_pkt_d_bits_half(lsu_lsc_ctl_io_lsu_pkt_d_bits_half),
    .io_lsu_pkt_d_bits_word(lsu_lsc_ctl_io_lsu_pkt_d_bits_word),
    .io_lsu_pkt_d_bits_dword(lsu_lsc_ctl_io_lsu_pkt_d_bits_dword),
    .io_lsu_pkt_d_bits_load(lsu_lsc_ctl_io_lsu_pkt_d_bits_load),
    .io_lsu_pkt_d_bits_store(lsu_lsc_ctl_io_lsu_pkt_d_bits_store),
    .io_lsu_pkt_d_bits_unsign(lsu_lsc_ctl_io_lsu_pkt_d_bits_unsign),
    .io_lsu_pkt_d_bits_dma(lsu_lsc_ctl_io_lsu_pkt_d_bits_dma),
    .io_lsu_pkt_d_bits_store_data_bypass_d(lsu_lsc_ctl_io_lsu_pkt_d_bits_store_data_bypass_d),
    .io_lsu_pkt_d_bits_load_ldst_bypass_d(lsu_lsc_ctl_io_lsu_pkt_d_bits_load_ldst_bypass_d),
    .io_lsu_pkt_d_bits_store_data_bypass_m(lsu_lsc_ctl_io_lsu_pkt_d_bits_store_data_bypass_m),
    .io_lsu_pkt_m_valid(lsu_lsc_ctl_io_lsu_pkt_m_valid),
    .io_lsu_pkt_m_bits_fast_int(lsu_lsc_ctl_io_lsu_pkt_m_bits_fast_int),
    .io_lsu_pkt_m_bits_by(lsu_lsc_ctl_io_lsu_pkt_m_bits_by),
    .io_lsu_pkt_m_bits_half(lsu_lsc_ctl_io_lsu_pkt_m_bits_half),
    .io_lsu_pkt_m_bits_word(lsu_lsc_ctl_io_lsu_pkt_m_bits_word),
    .io_lsu_pkt_m_bits_dword(lsu_lsc_ctl_io_lsu_pkt_m_bits_dword),
    .io_lsu_pkt_m_bits_load(lsu_lsc_ctl_io_lsu_pkt_m_bits_load),
    .io_lsu_pkt_m_bits_store(lsu_lsc_ctl_io_lsu_pkt_m_bits_store),
    .io_lsu_pkt_m_bits_unsign(lsu_lsc_ctl_io_lsu_pkt_m_bits_unsign),
    .io_lsu_pkt_m_bits_dma(lsu_lsc_ctl_io_lsu_pkt_m_bits_dma),
    .io_lsu_pkt_m_bits_store_data_bypass_m(lsu_lsc_ctl_io_lsu_pkt_m_bits_store_data_bypass_m),
    .io_lsu_pkt_r_valid(lsu_lsc_ctl_io_lsu_pkt_r_valid),
    .io_lsu_pkt_r_bits_by(lsu_lsc_ctl_io_lsu_pkt_r_bits_by),
    .io_lsu_pkt_r_bits_half(lsu_lsc_ctl_io_lsu_pkt_r_bits_half),
    .io_lsu_pkt_r_bits_word(lsu_lsc_ctl_io_lsu_pkt_r_bits_word),
    .io_lsu_pkt_r_bits_dword(lsu_lsc_ctl_io_lsu_pkt_r_bits_dword),
    .io_lsu_pkt_r_bits_load(lsu_lsc_ctl_io_lsu_pkt_r_bits_load),
    .io_lsu_pkt_r_bits_store(lsu_lsc_ctl_io_lsu_pkt_r_bits_store),
    .io_lsu_pkt_r_bits_unsign(lsu_lsc_ctl_io_lsu_pkt_r_bits_unsign),
    .io_lsu_pkt_r_bits_dma(lsu_lsc_ctl_io_lsu_pkt_r_bits_dma)
  );
  lsu_dccm_ctl dccm_ctl ( // @[lsu.scala 63:30]
    .clock(dccm_ctl_clock),
    .reset(dccm_ctl_reset),
    .io_lsu_c2_m_clk(dccm_ctl_io_lsu_c2_m_clk),
    .io_lsu_c2_r_clk(dccm_ctl_io_lsu_c2_r_clk),
    .io_lsu_free_c2_clk(dccm_ctl_io_lsu_free_c2_clk),
    .io_lsu_store_c1_r_clk(dccm_ctl_io_lsu_store_c1_r_clk),
    .io_lsu_pkt_d_valid(dccm_ctl_io_lsu_pkt_d_valid),
    .io_lsu_pkt_d_bits_word(dccm_ctl_io_lsu_pkt_d_bits_word),
    .io_lsu_pkt_d_bits_dword(dccm_ctl_io_lsu_pkt_d_bits_dword),
    .io_lsu_pkt_d_bits_load(dccm_ctl_io_lsu_pkt_d_bits_load),
    .io_lsu_pkt_d_bits_store(dccm_ctl_io_lsu_pkt_d_bits_store),
    .io_lsu_pkt_d_bits_dma(dccm_ctl_io_lsu_pkt_d_bits_dma),
    .io_lsu_pkt_m_valid(dccm_ctl_io_lsu_pkt_m_valid),
    .io_lsu_pkt_m_bits_by(dccm_ctl_io_lsu_pkt_m_bits_by),
    .io_lsu_pkt_m_bits_half(dccm_ctl_io_lsu_pkt_m_bits_half),
    .io_lsu_pkt_m_bits_word(dccm_ctl_io_lsu_pkt_m_bits_word),
    .io_lsu_pkt_m_bits_load(dccm_ctl_io_lsu_pkt_m_bits_load),
    .io_lsu_pkt_m_bits_store(dccm_ctl_io_lsu_pkt_m_bits_store),
    .io_lsu_pkt_m_bits_dma(dccm_ctl_io_lsu_pkt_m_bits_dma),
    .io_lsu_pkt_r_valid(dccm_ctl_io_lsu_pkt_r_valid),
    .io_lsu_pkt_r_bits_by(dccm_ctl_io_lsu_pkt_r_bits_by),
    .io_lsu_pkt_r_bits_half(dccm_ctl_io_lsu_pkt_r_bits_half),
    .io_lsu_pkt_r_bits_word(dccm_ctl_io_lsu_pkt_r_bits_word),
    .io_lsu_pkt_r_bits_load(dccm_ctl_io_lsu_pkt_r_bits_load),
    .io_lsu_pkt_r_bits_store(dccm_ctl_io_lsu_pkt_r_bits_store),
    .io_lsu_pkt_r_bits_dma(dccm_ctl_io_lsu_pkt_r_bits_dma),
    .io_addr_in_dccm_d(dccm_ctl_io_addr_in_dccm_d),
    .io_addr_in_dccm_m(dccm_ctl_io_addr_in_dccm_m),
    .io_addr_in_dccm_r(dccm_ctl_io_addr_in_dccm_r),
    .io_addr_in_pic_d(dccm_ctl_io_addr_in_pic_d),
    .io_addr_in_pic_m(dccm_ctl_io_addr_in_pic_m),
    .io_addr_in_pic_r(dccm_ctl_io_addr_in_pic_r),
    .io_lsu_raw_fwd_lo_r(dccm_ctl_io_lsu_raw_fwd_lo_r),
    .io_lsu_raw_fwd_hi_r(dccm_ctl_io_lsu_raw_fwd_hi_r),
    .io_lsu_commit_r(dccm_ctl_io_lsu_commit_r),
    .io_lsu_addr_d(dccm_ctl_io_lsu_addr_d),
    .io_lsu_addr_m(dccm_ctl_io_lsu_addr_m),
    .io_lsu_addr_r(dccm_ctl_io_lsu_addr_r),
    .io_end_addr_d(dccm_ctl_io_end_addr_d),
    .io_end_addr_m(dccm_ctl_io_end_addr_m),
    .io_end_addr_r(dccm_ctl_io_end_addr_r),
    .io_stbuf_reqvld_any(dccm_ctl_io_stbuf_reqvld_any),
    .io_stbuf_addr_any(dccm_ctl_io_stbuf_addr_any),
    .io_stbuf_data_any(dccm_ctl_io_stbuf_data_any),
    .io_stbuf_ecc_any(dccm_ctl_io_stbuf_ecc_any),
    .io_stbuf_fwddata_hi_m(dccm_ctl_io_stbuf_fwddata_hi_m),
    .io_stbuf_fwddata_lo_m(dccm_ctl_io_stbuf_fwddata_lo_m),
    .io_stbuf_fwdbyteen_lo_m(dccm_ctl_io_stbuf_fwdbyteen_lo_m),
    .io_stbuf_fwdbyteen_hi_m(dccm_ctl_io_stbuf_fwdbyteen_hi_m),
    .io_lsu_ld_data_corr_r(dccm_ctl_io_lsu_ld_data_corr_r),
    .io_lsu_double_ecc_error_r(dccm_ctl_io_lsu_double_ecc_error_r),
    .io_single_ecc_error_hi_r(dccm_ctl_io_single_ecc_error_hi_r),
    .io_single_ecc_error_lo_r(dccm_ctl_io_single_ecc_error_lo_r),
    .io_sec_data_hi_r_ff(dccm_ctl_io_sec_data_hi_r_ff),
    .io_sec_data_lo_r_ff(dccm_ctl_io_sec_data_lo_r_ff),
    .io_sec_data_ecc_hi_r_ff(dccm_ctl_io_sec_data_ecc_hi_r_ff),
    .io_sec_data_ecc_lo_r_ff(dccm_ctl_io_sec_data_ecc_lo_r_ff),
    .io_dccm_rdata_hi_m(dccm_ctl_io_dccm_rdata_hi_m),
    .io_dccm_rdata_lo_m(dccm_ctl_io_dccm_rdata_lo_m),
    .io_dccm_data_ecc_hi_m(dccm_ctl_io_dccm_data_ecc_hi_m),
    .io_dccm_data_ecc_lo_m(dccm_ctl_io_dccm_data_ecc_lo_m),
    .io_lsu_ld_data_m(dccm_ctl_io_lsu_ld_data_m),
    .io_lsu_double_ecc_error_m(dccm_ctl_io_lsu_double_ecc_error_m),
    .io_sec_data_hi_m(dccm_ctl_io_sec_data_hi_m),
    .io_sec_data_lo_m(dccm_ctl_io_sec_data_lo_m),
    .io_store_data_m(dccm_ctl_io_store_data_m),
    .io_dma_dccm_wen(dccm_ctl_io_dma_dccm_wen),
    .io_dma_pic_wen(dccm_ctl_io_dma_pic_wen),
    .io_dma_mem_tag_m(dccm_ctl_io_dma_mem_tag_m),
    .io_dma_dccm_wdata_lo(dccm_ctl_io_dma_dccm_wdata_lo),
    .io_dma_dccm_wdata_hi(dccm_ctl_io_dma_dccm_wdata_hi),
    .io_dma_dccm_wdata_ecc_hi(dccm_ctl_io_dma_dccm_wdata_ecc_hi),
    .io_dma_dccm_wdata_ecc_lo(dccm_ctl_io_dma_dccm_wdata_ecc_lo),
    .io_store_data_hi_r(dccm_ctl_io_store_data_hi_r),
    .io_store_data_lo_r(dccm_ctl_io_store_data_lo_r),
    .io_store_datafn_hi_r(dccm_ctl_io_store_datafn_hi_r),
    .io_store_datafn_lo_r(dccm_ctl_io_store_datafn_lo_r),
    .io_store_data_r(dccm_ctl_io_store_data_r),
    .io_ld_single_ecc_error_r(dccm_ctl_io_ld_single_ecc_error_r),
    .io_ld_single_ecc_error_r_ff(dccm_ctl_io_ld_single_ecc_error_r_ff),
    .io_picm_mask_data_m(dccm_ctl_io_picm_mask_data_m),
    .io_lsu_stbuf_commit_any(dccm_ctl_io_lsu_stbuf_commit_any),
    .io_lsu_dccm_rden_m(dccm_ctl_io_lsu_dccm_rden_m),
    .io_dma_dccm_ctl_dma_mem_addr(dccm_ctl_io_dma_dccm_ctl_dma_mem_addr),
    .io_dma_dccm_ctl_dma_mem_wdata(dccm_ctl_io_dma_dccm_ctl_dma_mem_wdata),
    .io_dma_dccm_ctl_dccm_dma_rvalid(dccm_ctl_io_dma_dccm_ctl_dccm_dma_rvalid),
    .io_dma_dccm_ctl_dccm_dma_ecc_error(dccm_ctl_io_dma_dccm_ctl_dccm_dma_ecc_error),
    .io_dma_dccm_ctl_dccm_dma_rtag(dccm_ctl_io_dma_dccm_ctl_dccm_dma_rtag),
    .io_dma_dccm_ctl_dccm_dma_rdata(dccm_ctl_io_dma_dccm_ctl_dccm_dma_rdata),
    .io_dccm_wren(dccm_ctl_io_dccm_wren),
    .io_dccm_rden(dccm_ctl_io_dccm_rden),
    .io_dccm_wr_addr_lo(dccm_ctl_io_dccm_wr_addr_lo),
    .io_dccm_wr_addr_hi(dccm_ctl_io_dccm_wr_addr_hi),
    .io_dccm_rd_addr_lo(dccm_ctl_io_dccm_rd_addr_lo),
    .io_dccm_rd_addr_hi(dccm_ctl_io_dccm_rd_addr_hi),
    .io_dccm_wr_data_lo(dccm_ctl_io_dccm_wr_data_lo),
    .io_dccm_wr_data_hi(dccm_ctl_io_dccm_wr_data_hi),
    .io_dccm_rd_data_lo(dccm_ctl_io_dccm_rd_data_lo),
    .io_dccm_rd_data_hi(dccm_ctl_io_dccm_rd_data_hi),
    .io_lsu_pic_picm_wren(dccm_ctl_io_lsu_pic_picm_wren),
    .io_lsu_pic_picm_rden(dccm_ctl_io_lsu_pic_picm_rden),
    .io_lsu_pic_picm_mken(dccm_ctl_io_lsu_pic_picm_mken),
    .io_lsu_pic_picm_rdaddr(dccm_ctl_io_lsu_pic_picm_rdaddr),
    .io_lsu_pic_picm_wraddr(dccm_ctl_io_lsu_pic_picm_wraddr),
    .io_lsu_pic_picm_wr_data(dccm_ctl_io_lsu_pic_picm_wr_data),
    .io_lsu_pic_picm_rd_data(dccm_ctl_io_lsu_pic_picm_rd_data),
    .io_scan_mode(dccm_ctl_io_scan_mode)
  );
  lsu_stbuf stbuf ( // @[lsu.scala 64:30]
    .clock(stbuf_clock),
    .reset(stbuf_reset),
    .io_lsu_c1_m_clk(stbuf_io_lsu_c1_m_clk),
    .io_lsu_c1_r_clk(stbuf_io_lsu_c1_r_clk),
    .io_lsu_stbuf_c1_clk(stbuf_io_lsu_stbuf_c1_clk),
    .io_lsu_free_c2_clk(stbuf_io_lsu_free_c2_clk),
    .io_lsu_pkt_m_valid(stbuf_io_lsu_pkt_m_valid),
    .io_lsu_pkt_m_bits_store(stbuf_io_lsu_pkt_m_bits_store),
    .io_lsu_pkt_m_bits_dma(stbuf_io_lsu_pkt_m_bits_dma),
    .io_lsu_pkt_r_valid(stbuf_io_lsu_pkt_r_valid),
    .io_lsu_pkt_r_bits_by(stbuf_io_lsu_pkt_r_bits_by),
    .io_lsu_pkt_r_bits_half(stbuf_io_lsu_pkt_r_bits_half),
    .io_lsu_pkt_r_bits_word(stbuf_io_lsu_pkt_r_bits_word),
    .io_lsu_pkt_r_bits_dword(stbuf_io_lsu_pkt_r_bits_dword),
    .io_lsu_pkt_r_bits_store(stbuf_io_lsu_pkt_r_bits_store),
    .io_lsu_pkt_r_bits_dma(stbuf_io_lsu_pkt_r_bits_dma),
    .io_store_stbuf_reqvld_r(stbuf_io_store_stbuf_reqvld_r),
    .io_lsu_commit_r(stbuf_io_lsu_commit_r),
    .io_dec_lsu_valid_raw_d(stbuf_io_dec_lsu_valid_raw_d),
    .io_store_data_hi_r(stbuf_io_store_data_hi_r),
    .io_store_data_lo_r(stbuf_io_store_data_lo_r),
    .io_store_datafn_hi_r(stbuf_io_store_datafn_hi_r),
    .io_store_datafn_lo_r(stbuf_io_store_datafn_lo_r),
    .io_lsu_stbuf_commit_any(stbuf_io_lsu_stbuf_commit_any),
    .io_lsu_addr_d(stbuf_io_lsu_addr_d),
    .io_lsu_addr_m(stbuf_io_lsu_addr_m),
    .io_lsu_addr_r(stbuf_io_lsu_addr_r),
    .io_end_addr_d(stbuf_io_end_addr_d),
    .io_end_addr_m(stbuf_io_end_addr_m),
    .io_end_addr_r(stbuf_io_end_addr_r),
    .io_addr_in_dccm_m(stbuf_io_addr_in_dccm_m),
    .io_addr_in_dccm_r(stbuf_io_addr_in_dccm_r),
    .io_scan_mode(stbuf_io_scan_mode),
    .io_stbuf_reqvld_any(stbuf_io_stbuf_reqvld_any),
    .io_stbuf_reqvld_flushed_any(stbuf_io_stbuf_reqvld_flushed_any),
    .io_stbuf_addr_any(stbuf_io_stbuf_addr_any),
    .io_stbuf_data_any(stbuf_io_stbuf_data_any),
    .io_lsu_stbuf_full_any(stbuf_io_lsu_stbuf_full_any),
    .io_lsu_stbuf_empty_any(stbuf_io_lsu_stbuf_empty_any),
    .io_ldst_stbuf_reqvld_r(stbuf_io_ldst_stbuf_reqvld_r),
    .io_stbuf_fwddata_hi_m(stbuf_io_stbuf_fwddata_hi_m),
    .io_stbuf_fwddata_lo_m(stbuf_io_stbuf_fwddata_lo_m),
    .io_stbuf_fwdbyteen_hi_m(stbuf_io_stbuf_fwdbyteen_hi_m),
    .io_stbuf_fwdbyteen_lo_m(stbuf_io_stbuf_fwdbyteen_lo_m)
  );
  lsu_ecc ecc ( // @[lsu.scala 65:30]
    .clock(ecc_clock),
    .reset(ecc_reset),
    .io_lsu_c2_r_clk(ecc_io_lsu_c2_r_clk),
    .io_lsu_pkt_m_valid(ecc_io_lsu_pkt_m_valid),
    .io_lsu_pkt_m_bits_load(ecc_io_lsu_pkt_m_bits_load),
    .io_lsu_pkt_m_bits_store(ecc_io_lsu_pkt_m_bits_store),
    .io_lsu_pkt_m_bits_dma(ecc_io_lsu_pkt_m_bits_dma),
    .io_stbuf_data_any(ecc_io_stbuf_data_any),
    .io_dec_tlu_core_ecc_disable(ecc_io_dec_tlu_core_ecc_disable),
    .io_lsu_addr_m(ecc_io_lsu_addr_m),
    .io_end_addr_m(ecc_io_end_addr_m),
    .io_dccm_rdata_hi_m(ecc_io_dccm_rdata_hi_m),
    .io_dccm_rdata_lo_m(ecc_io_dccm_rdata_lo_m),
    .io_dccm_data_ecc_hi_m(ecc_io_dccm_data_ecc_hi_m),
    .io_dccm_data_ecc_lo_m(ecc_io_dccm_data_ecc_lo_m),
    .io_ld_single_ecc_error_r(ecc_io_ld_single_ecc_error_r),
    .io_ld_single_ecc_error_r_ff(ecc_io_ld_single_ecc_error_r_ff),
    .io_lsu_dccm_rden_m(ecc_io_lsu_dccm_rden_m),
    .io_addr_in_dccm_m(ecc_io_addr_in_dccm_m),
    .io_dma_dccm_wen(ecc_io_dma_dccm_wen),
    .io_dma_dccm_wdata_lo(ecc_io_dma_dccm_wdata_lo),
    .io_dma_dccm_wdata_hi(ecc_io_dma_dccm_wdata_hi),
    .io_scan_mode(ecc_io_scan_mode),
    .io_sec_data_hi_r(ecc_io_sec_data_hi_r),
    .io_sec_data_lo_r(ecc_io_sec_data_lo_r),
    .io_sec_data_hi_m(ecc_io_sec_data_hi_m),
    .io_sec_data_lo_m(ecc_io_sec_data_lo_m),
    .io_sec_data_hi_r_ff(ecc_io_sec_data_hi_r_ff),
    .io_sec_data_lo_r_ff(ecc_io_sec_data_lo_r_ff),
    .io_dma_dccm_wdata_ecc_hi(ecc_io_dma_dccm_wdata_ecc_hi),
    .io_dma_dccm_wdata_ecc_lo(ecc_io_dma_dccm_wdata_ecc_lo),
    .io_stbuf_ecc_any(ecc_io_stbuf_ecc_any),
    .io_sec_data_ecc_hi_r_ff(ecc_io_sec_data_ecc_hi_r_ff),
    .io_sec_data_ecc_lo_r_ff(ecc_io_sec_data_ecc_lo_r_ff),
    .io_single_ecc_error_hi_r(ecc_io_single_ecc_error_hi_r),
    .io_single_ecc_error_lo_r(ecc_io_single_ecc_error_lo_r),
    .io_lsu_single_ecc_error_r(ecc_io_lsu_single_ecc_error_r),
    .io_lsu_double_ecc_error_r(ecc_io_lsu_double_ecc_error_r),
    .io_lsu_single_ecc_error_m(ecc_io_lsu_single_ecc_error_m),
    .io_lsu_double_ecc_error_m(ecc_io_lsu_double_ecc_error_m)
  );
  lsu_trigger trigger ( // @[lsu.scala 66:30]
    .io_trigger_pkt_any_0_select(trigger_io_trigger_pkt_any_0_select),
    .io_trigger_pkt_any_0_match_pkt(trigger_io_trigger_pkt_any_0_match_pkt),
    .io_trigger_pkt_any_0_store(trigger_io_trigger_pkt_any_0_store),
    .io_trigger_pkt_any_0_load(trigger_io_trigger_pkt_any_0_load),
    .io_trigger_pkt_any_0_tdata2(trigger_io_trigger_pkt_any_0_tdata2),
    .io_trigger_pkt_any_1_select(trigger_io_trigger_pkt_any_1_select),
    .io_trigger_pkt_any_1_match_pkt(trigger_io_trigger_pkt_any_1_match_pkt),
    .io_trigger_pkt_any_1_store(trigger_io_trigger_pkt_any_1_store),
    .io_trigger_pkt_any_1_load(trigger_io_trigger_pkt_any_1_load),
    .io_trigger_pkt_any_1_tdata2(trigger_io_trigger_pkt_any_1_tdata2),
    .io_trigger_pkt_any_2_select(trigger_io_trigger_pkt_any_2_select),
    .io_trigger_pkt_any_2_match_pkt(trigger_io_trigger_pkt_any_2_match_pkt),
    .io_trigger_pkt_any_2_store(trigger_io_trigger_pkt_any_2_store),
    .io_trigger_pkt_any_2_load(trigger_io_trigger_pkt_any_2_load),
    .io_trigger_pkt_any_2_tdata2(trigger_io_trigger_pkt_any_2_tdata2),
    .io_trigger_pkt_any_3_select(trigger_io_trigger_pkt_any_3_select),
    .io_trigger_pkt_any_3_match_pkt(trigger_io_trigger_pkt_any_3_match_pkt),
    .io_trigger_pkt_any_3_store(trigger_io_trigger_pkt_any_3_store),
    .io_trigger_pkt_any_3_load(trigger_io_trigger_pkt_any_3_load),
    .io_trigger_pkt_any_3_tdata2(trigger_io_trigger_pkt_any_3_tdata2),
    .io_lsu_pkt_m_valid(trigger_io_lsu_pkt_m_valid),
    .io_lsu_pkt_m_bits_half(trigger_io_lsu_pkt_m_bits_half),
    .io_lsu_pkt_m_bits_word(trigger_io_lsu_pkt_m_bits_word),
    .io_lsu_pkt_m_bits_load(trigger_io_lsu_pkt_m_bits_load),
    .io_lsu_pkt_m_bits_store(trigger_io_lsu_pkt_m_bits_store),
    .io_lsu_pkt_m_bits_dma(trigger_io_lsu_pkt_m_bits_dma),
    .io_lsu_addr_m(trigger_io_lsu_addr_m),
    .io_store_data_m(trigger_io_store_data_m),
    .io_lsu_trigger_match_m(trigger_io_lsu_trigger_match_m)
  );
  lsu_clkdomain clkdomain ( // @[lsu.scala 67:30]
    .clock(clkdomain_clock),
    .reset(clkdomain_reset),
    .io_free_clk(clkdomain_io_free_clk),
    .io_clk_override(clkdomain_io_clk_override),
    .io_dma_dccm_req(clkdomain_io_dma_dccm_req),
    .io_ldst_stbuf_reqvld_r(clkdomain_io_ldst_stbuf_reqvld_r),
    .io_stbuf_reqvld_any(clkdomain_io_stbuf_reqvld_any),
    .io_stbuf_reqvld_flushed_any(clkdomain_io_stbuf_reqvld_flushed_any),
    .io_lsu_busreq_r(clkdomain_io_lsu_busreq_r),
    .io_lsu_bus_buffer_pend_any(clkdomain_io_lsu_bus_buffer_pend_any),
    .io_lsu_bus_buffer_empty_any(clkdomain_io_lsu_bus_buffer_empty_any),
    .io_lsu_stbuf_empty_any(clkdomain_io_lsu_stbuf_empty_any),
    .io_lsu_bus_clk_en(clkdomain_io_lsu_bus_clk_en),
    .io_lsu_p_valid(clkdomain_io_lsu_p_valid),
    .io_lsu_pkt_d_valid(clkdomain_io_lsu_pkt_d_valid),
    .io_lsu_pkt_d_bits_store(clkdomain_io_lsu_pkt_d_bits_store),
    .io_lsu_pkt_m_valid(clkdomain_io_lsu_pkt_m_valid),
    .io_lsu_pkt_m_bits_store(clkdomain_io_lsu_pkt_m_bits_store),
    .io_lsu_pkt_r_valid(clkdomain_io_lsu_pkt_r_valid),
    .io_lsu_c1_m_clk(clkdomain_io_lsu_c1_m_clk),
    .io_lsu_c1_r_clk(clkdomain_io_lsu_c1_r_clk),
    .io_lsu_c2_m_clk(clkdomain_io_lsu_c2_m_clk),
    .io_lsu_c2_r_clk(clkdomain_io_lsu_c2_r_clk),
    .io_lsu_store_c1_m_clk(clkdomain_io_lsu_store_c1_m_clk),
    .io_lsu_store_c1_r_clk(clkdomain_io_lsu_store_c1_r_clk),
    .io_lsu_stbuf_c1_clk(clkdomain_io_lsu_stbuf_c1_clk),
    .io_lsu_bus_obuf_c1_clk(clkdomain_io_lsu_bus_obuf_c1_clk),
    .io_lsu_bus_ibuf_c1_clk(clkdomain_io_lsu_bus_ibuf_c1_clk),
    .io_lsu_bus_buf_c1_clk(clkdomain_io_lsu_bus_buf_c1_clk),
    .io_lsu_busm_clk(clkdomain_io_lsu_busm_clk),
    .io_lsu_free_c2_clk(clkdomain_io_lsu_free_c2_clk),
    .io_scan_mode(clkdomain_io_scan_mode)
  );
  lsu_bus_intf bus_intf ( // @[lsu.scala 68:30]
    .clock(bus_intf_clock),
    .reset(bus_intf_reset),
    .io_scan_mode(bus_intf_io_scan_mode),
    .io_tlu_busbuff_lsu_pmu_bus_misaligned(bus_intf_io_tlu_busbuff_lsu_pmu_bus_misaligned),
    .io_tlu_busbuff_lsu_pmu_bus_error(bus_intf_io_tlu_busbuff_lsu_pmu_bus_error),
    .io_tlu_busbuff_lsu_pmu_bus_busy(bus_intf_io_tlu_busbuff_lsu_pmu_bus_busy),
    .io_tlu_busbuff_dec_tlu_external_ldfwd_disable(bus_intf_io_tlu_busbuff_dec_tlu_external_ldfwd_disable),
    .io_tlu_busbuff_dec_tlu_wb_coalescing_disable(bus_intf_io_tlu_busbuff_dec_tlu_wb_coalescing_disable),
    .io_tlu_busbuff_dec_tlu_sideeffect_posted_disable(bus_intf_io_tlu_busbuff_dec_tlu_sideeffect_posted_disable),
    .io_tlu_busbuff_lsu_imprecise_error_load_any(bus_intf_io_tlu_busbuff_lsu_imprecise_error_load_any),
    .io_tlu_busbuff_lsu_imprecise_error_store_any(bus_intf_io_tlu_busbuff_lsu_imprecise_error_store_any),
    .io_tlu_busbuff_lsu_imprecise_error_addr_any(bus_intf_io_tlu_busbuff_lsu_imprecise_error_addr_any),
    .io_lsu_c1_m_clk(bus_intf_io_lsu_c1_m_clk),
    .io_lsu_c1_r_clk(bus_intf_io_lsu_c1_r_clk),
    .io_lsu_c2_r_clk(bus_intf_io_lsu_c2_r_clk),
    .io_lsu_bus_ibuf_c1_clk(bus_intf_io_lsu_bus_ibuf_c1_clk),
    .io_lsu_bus_obuf_c1_clk(bus_intf_io_lsu_bus_obuf_c1_clk),
    .io_lsu_bus_buf_c1_clk(bus_intf_io_lsu_bus_buf_c1_clk),
    .io_lsu_free_c2_clk(bus_intf_io_lsu_free_c2_clk),
    .io_free_clk(bus_intf_io_free_clk),
    .io_lsu_busm_clk(bus_intf_io_lsu_busm_clk),
    .io_axi_aw_valid(bus_intf_io_axi_aw_valid),
    .io_axi_aw_bits_addr(bus_intf_io_axi_aw_bits_addr),
    .io_axi_aw_bits_size(bus_intf_io_axi_aw_bits_size),
    .io_axi_w_valid(bus_intf_io_axi_w_valid),
    .io_axi_w_bits_strb(bus_intf_io_axi_w_bits_strb),
    .io_axi_ar_valid(bus_intf_io_axi_ar_valid),
    .io_axi_ar_bits_addr(bus_intf_io_axi_ar_bits_addr),
    .io_axi_ar_bits_size(bus_intf_io_axi_ar_bits_size),
    .io_dec_lsu_valid_raw_d(bus_intf_io_dec_lsu_valid_raw_d),
    .io_lsu_busreq_m(bus_intf_io_lsu_busreq_m),
    .io_lsu_pkt_m_valid(bus_intf_io_lsu_pkt_m_valid),
    .io_lsu_pkt_m_bits_by(bus_intf_io_lsu_pkt_m_bits_by),
    .io_lsu_pkt_m_bits_half(bus_intf_io_lsu_pkt_m_bits_half),
    .io_lsu_pkt_m_bits_word(bus_intf_io_lsu_pkt_m_bits_word),
    .io_lsu_pkt_m_bits_load(bus_intf_io_lsu_pkt_m_bits_load),
    .io_lsu_pkt_r_valid(bus_intf_io_lsu_pkt_r_valid),
    .io_lsu_pkt_r_bits_by(bus_intf_io_lsu_pkt_r_bits_by),
    .io_lsu_pkt_r_bits_half(bus_intf_io_lsu_pkt_r_bits_half),
    .io_lsu_pkt_r_bits_word(bus_intf_io_lsu_pkt_r_bits_word),
    .io_lsu_pkt_r_bits_load(bus_intf_io_lsu_pkt_r_bits_load),
    .io_lsu_pkt_r_bits_store(bus_intf_io_lsu_pkt_r_bits_store),
    .io_lsu_pkt_r_bits_unsign(bus_intf_io_lsu_pkt_r_bits_unsign),
    .io_lsu_addr_d(bus_intf_io_lsu_addr_d),
    .io_lsu_addr_m(bus_intf_io_lsu_addr_m),
    .io_lsu_addr_r(bus_intf_io_lsu_addr_r),
    .io_end_addr_d(bus_intf_io_end_addr_d),
    .io_end_addr_m(bus_intf_io_end_addr_m),
    .io_end_addr_r(bus_intf_io_end_addr_r),
    .io_store_data_r(bus_intf_io_store_data_r),
    .io_dec_tlu_force_halt(bus_intf_io_dec_tlu_force_halt),
    .io_lsu_commit_r(bus_intf_io_lsu_commit_r),
    .io_is_sideeffects_m(bus_intf_io_is_sideeffects_m),
    .io_flush_m_up(bus_intf_io_flush_m_up),
    .io_flush_r(bus_intf_io_flush_r),
    .io_lsu_busreq_r(bus_intf_io_lsu_busreq_r),
    .io_lsu_bus_buffer_pend_any(bus_intf_io_lsu_bus_buffer_pend_any),
    .io_lsu_bus_buffer_full_any(bus_intf_io_lsu_bus_buffer_full_any),
    .io_lsu_bus_buffer_empty_any(bus_intf_io_lsu_bus_buffer_empty_any),
    .io_bus_read_data_m(bus_intf_io_bus_read_data_m),
    .io_dctl_busbuff_lsu_nonblock_load_valid_m(bus_intf_io_dctl_busbuff_lsu_nonblock_load_valid_m),
    .io_dctl_busbuff_lsu_nonblock_load_tag_m(bus_intf_io_dctl_busbuff_lsu_nonblock_load_tag_m),
    .io_dctl_busbuff_lsu_nonblock_load_inv_r(bus_intf_io_dctl_busbuff_lsu_nonblock_load_inv_r),
    .io_dctl_busbuff_lsu_nonblock_load_inv_tag_r(bus_intf_io_dctl_busbuff_lsu_nonblock_load_inv_tag_r),
    .io_dctl_busbuff_lsu_nonblock_load_data_valid(bus_intf_io_dctl_busbuff_lsu_nonblock_load_data_valid),
    .io_dctl_busbuff_lsu_nonblock_load_data_error(bus_intf_io_dctl_busbuff_lsu_nonblock_load_data_error),
    .io_dctl_busbuff_lsu_nonblock_load_data_tag(bus_intf_io_dctl_busbuff_lsu_nonblock_load_data_tag),
    .io_dctl_busbuff_lsu_nonblock_load_data(bus_intf_io_dctl_busbuff_lsu_nonblock_load_data),
    .io_lsu_bus_clk_en(bus_intf_io_lsu_bus_clk_en)
  );
  assign io_lsu_dma_dma_dccm_ctl_dccm_dma_rvalid = dccm_ctl_io_dma_dccm_ctl_dccm_dma_rvalid; // @[lsu.scala 194:27]
  assign io_lsu_dma_dma_dccm_ctl_dccm_dma_ecc_error = dccm_ctl_io_dma_dccm_ctl_dccm_dma_ecc_error; // @[lsu.scala 194:27]
  assign io_lsu_dma_dma_dccm_ctl_dccm_dma_rtag = dccm_ctl_io_dma_dccm_ctl_dccm_dma_rtag; // @[lsu.scala 194:27]
  assign io_lsu_dma_dma_dccm_ctl_dccm_dma_rdata = dccm_ctl_io_dma_dccm_ctl_dccm_dma_rdata; // @[lsu.scala 194:27]
  assign io_lsu_dma_dccm_ready = ~_T_8; // @[lsu.scala 82:25]
  assign io_lsu_pic_picm_wren = dccm_ctl_io_lsu_pic_picm_wren; // @[lsu.scala 196:14]
  assign io_lsu_pic_picm_rden = dccm_ctl_io_lsu_pic_picm_rden; // @[lsu.scala 196:14]
  assign io_lsu_pic_picm_mken = dccm_ctl_io_lsu_pic_picm_mken; // @[lsu.scala 196:14]
  assign io_lsu_pic_picm_rdaddr = dccm_ctl_io_lsu_pic_picm_rdaddr; // @[lsu.scala 196:14]
  assign io_lsu_pic_picm_wraddr = dccm_ctl_io_lsu_pic_picm_wraddr; // @[lsu.scala 196:14]
  assign io_lsu_pic_picm_wr_data = dccm_ctl_io_lsu_pic_picm_wr_data; // @[lsu.scala 196:14]
  assign io_lsu_dec_tlu_busbuff_lsu_pmu_bus_misaligned = bus_intf_io_tlu_busbuff_lsu_pmu_bus_misaligned; // @[lsu.scala 286:26]
  assign io_lsu_dec_tlu_busbuff_lsu_pmu_bus_error = bus_intf_io_tlu_busbuff_lsu_pmu_bus_error; // @[lsu.scala 286:26]
  assign io_lsu_dec_tlu_busbuff_lsu_pmu_bus_busy = bus_intf_io_tlu_busbuff_lsu_pmu_bus_busy; // @[lsu.scala 286:26]
  assign io_lsu_dec_tlu_busbuff_lsu_imprecise_error_load_any = bus_intf_io_tlu_busbuff_lsu_imprecise_error_load_any; // @[lsu.scala 286:26]
  assign io_lsu_dec_tlu_busbuff_lsu_imprecise_error_store_any = bus_intf_io_tlu_busbuff_lsu_imprecise_error_store_any; // @[lsu.scala 286:26]
  assign io_lsu_dec_tlu_busbuff_lsu_imprecise_error_addr_any = bus_intf_io_tlu_busbuff_lsu_imprecise_error_addr_any; // @[lsu.scala 286:26]
  assign io_lsu_dec_dctl_busbuff_lsu_nonblock_load_valid_m = bus_intf_io_dctl_busbuff_lsu_nonblock_load_valid_m; // @[lsu.scala 313:27]
  assign io_lsu_dec_dctl_busbuff_lsu_nonblock_load_tag_m = bus_intf_io_dctl_busbuff_lsu_nonblock_load_tag_m; // @[lsu.scala 313:27]
  assign io_lsu_dec_dctl_busbuff_lsu_nonblock_load_inv_r = bus_intf_io_dctl_busbuff_lsu_nonblock_load_inv_r; // @[lsu.scala 313:27]
  assign io_lsu_dec_dctl_busbuff_lsu_nonblock_load_inv_tag_r = bus_intf_io_dctl_busbuff_lsu_nonblock_load_inv_tag_r; // @[lsu.scala 313:27]
  assign io_lsu_dec_dctl_busbuff_lsu_nonblock_load_data_valid = bus_intf_io_dctl_busbuff_lsu_nonblock_load_data_valid; // @[lsu.scala 313:27]
  assign io_lsu_dec_dctl_busbuff_lsu_nonblock_load_data_error = bus_intf_io_dctl_busbuff_lsu_nonblock_load_data_error; // @[lsu.scala 313:27]
  assign io_lsu_dec_dctl_busbuff_lsu_nonblock_load_data_tag = bus_intf_io_dctl_busbuff_lsu_nonblock_load_data_tag; // @[lsu.scala 313:27]
  assign io_lsu_dec_dctl_busbuff_lsu_nonblock_load_data = bus_intf_io_dctl_busbuff_lsu_nonblock_load_data; // @[lsu.scala 313:27]
  assign io_dccm_wren = dccm_ctl_io_dccm_wren; // @[lsu.scala 195:11]
  assign io_dccm_rden = dccm_ctl_io_dccm_rden; // @[lsu.scala 195:11]
  assign io_dccm_wr_addr_lo = dccm_ctl_io_dccm_wr_addr_lo; // @[lsu.scala 195:11]
  assign io_dccm_wr_addr_hi = dccm_ctl_io_dccm_wr_addr_hi; // @[lsu.scala 195:11]
  assign io_dccm_rd_addr_lo = dccm_ctl_io_dccm_rd_addr_lo; // @[lsu.scala 195:11]
  assign io_dccm_rd_addr_hi = dccm_ctl_io_dccm_rd_addr_hi; // @[lsu.scala 195:11]
  assign io_dccm_wr_data_lo = dccm_ctl_io_dccm_wr_data_lo; // @[lsu.scala 195:11]
  assign io_dccm_wr_data_hi = dccm_ctl_io_dccm_wr_data_hi; // @[lsu.scala 195:11]
  assign io_lsu_tlu_lsu_pmu_load_external_m = _T_48 & lsu_lsc_ctl_io_addr_external_m; // @[lsu.scala 105:39]
  assign io_lsu_tlu_lsu_pmu_store_external_m = _T_50 & lsu_lsc_ctl_io_addr_external_m; // @[lsu.scala 106:39]
  assign io_axi_aw_valid = bus_intf_io_axi_aw_valid; // @[lsu.scala 314:49]
  assign io_axi_aw_bits_addr = bus_intf_io_axi_aw_bits_addr; // @[lsu.scala 314:49]
  assign io_axi_aw_bits_size = bus_intf_io_axi_aw_bits_size; // @[lsu.scala 314:49]
  assign io_axi_w_valid = bus_intf_io_axi_w_valid; // @[lsu.scala 314:49]
  assign io_axi_w_bits_strb = bus_intf_io_axi_w_bits_strb; // @[lsu.scala 314:49]
  assign io_axi_ar_valid = bus_intf_io_axi_ar_valid; // @[lsu.scala 314:49]
  assign io_axi_ar_bits_addr = bus_intf_io_axi_ar_bits_addr; // @[lsu.scala 314:49]
  assign io_axi_ar_bits_size = bus_intf_io_axi_ar_bits_size; // @[lsu.scala 314:49]
  assign io_lsu_result_m = lsu_lsc_ctl_io_lsu_result_m; // @[lsu.scala 61:19]
  assign io_lsu_result_corr_r = lsu_lsc_ctl_io_lsu_result_corr_r; // @[lsu.scala 62:24]
  assign io_lsu_load_stall_any = bus_intf_io_lsu_bus_buffer_full_any | dccm_ctl_io_ld_single_ecc_error_r_ff; // @[lsu.scala 75:25]
  assign io_lsu_store_stall_any = _T | dccm_ctl_io_ld_single_ecc_error_r_ff; // @[lsu.scala 74:26]
  assign io_lsu_fastint_stall_any = dccm_ctl_io_ld_single_ecc_error_r; // @[lsu.scala 76:28]
  assign io_lsu_idle_any = _T_22 & bus_intf_io_lsu_bus_buffer_empty_any; // @[lsu.scala 96:19]
  assign io_lsu_fir_addr = lsu_lsc_ctl_io_lsu_fir_addr; // @[lsu.scala 137:49]
  assign io_lsu_fir_error = lsu_lsc_ctl_io_lsu_fir_error; // @[lsu.scala 138:49]
  assign io_lsu_single_ecc_error_incr = lsu_lsc_ctl_io_lsu_single_ecc_error_incr; // @[lsu.scala 135:49]
  assign io_lsu_error_pkt_r_valid = lsu_lsc_ctl_io_lsu_error_pkt_r_valid; // @[lsu.scala 136:49]
  assign io_lsu_error_pkt_r_bits_single_ecc_error = lsu_lsc_ctl_io_lsu_error_pkt_r_bits_single_ecc_error; // @[lsu.scala 136:49]
  assign io_lsu_error_pkt_r_bits_inst_type = lsu_lsc_ctl_io_lsu_error_pkt_r_bits_inst_type; // @[lsu.scala 136:49]
  assign io_lsu_error_pkt_r_bits_exc_type = lsu_lsc_ctl_io_lsu_error_pkt_r_bits_exc_type; // @[lsu.scala 136:49]
  assign io_lsu_error_pkt_r_bits_mscause = lsu_lsc_ctl_io_lsu_error_pkt_r_bits_mscause; // @[lsu.scala 136:49]
  assign io_lsu_error_pkt_r_bits_addr = lsu_lsc_ctl_io_lsu_error_pkt_r_bits_addr; // @[lsu.scala 136:49]
  assign io_lsu_pmu_misaligned_m = lsu_lsc_ctl_io_lsu_pkt_m_valid & _T_46; // @[lsu.scala 104:27]
  assign io_lsu_trigger_match_m = trigger_io_lsu_trigger_match_m; // @[lsu.scala 261:50]
  assign lsu_lsc_ctl_reset = reset;
  assign lsu_lsc_ctl_io_lsu_c1_m_clk = clkdomain_io_lsu_c1_m_clk; // @[lsu.scala 110:46]
  assign lsu_lsc_ctl_io_lsu_c1_r_clk = clkdomain_io_lsu_c1_r_clk; // @[lsu.scala 111:46]
  assign lsu_lsc_ctl_io_lsu_c2_m_clk = clkdomain_io_lsu_c2_m_clk; // @[lsu.scala 112:46]
  assign lsu_lsc_ctl_io_lsu_c2_r_clk = clkdomain_io_lsu_c2_r_clk; // @[lsu.scala 113:46]
  assign lsu_lsc_ctl_io_lsu_store_c1_m_clk = clkdomain_io_lsu_store_c1_m_clk; // @[lsu.scala 114:46]
  assign lsu_lsc_ctl_io_lsu_ld_data_corr_r = dccm_ctl_io_lsu_ld_data_corr_r; // @[lsu.scala 116:46]
  assign lsu_lsc_ctl_io_lsu_single_ecc_error_r = ecc_io_lsu_single_ecc_error_r; // @[lsu.scala 117:46]
  assign lsu_lsc_ctl_io_lsu_double_ecc_error_r = ecc_io_lsu_double_ecc_error_r; // @[lsu.scala 118:46]
  assign lsu_lsc_ctl_io_lsu_ld_data_m = dccm_ctl_io_lsu_ld_data_m; // @[lsu.scala 119:46]
  assign lsu_lsc_ctl_io_lsu_single_ecc_error_m = ecc_io_lsu_single_ecc_error_m; // @[lsu.scala 120:46]
  assign lsu_lsc_ctl_io_lsu_double_ecc_error_m = ecc_io_lsu_double_ecc_error_m; // @[lsu.scala 121:46]
  assign lsu_lsc_ctl_io_flush_m_up = io_dec_tlu_flush_lower_r; // @[lsu.scala 122:46]
  assign lsu_lsc_ctl_io_flush_r = io_dec_tlu_i0_kill_writeb_r; // @[lsu.scala 123:46]
  assign lsu_lsc_ctl_io_lsu_exu_exu_lsu_rs1_d = io_lsu_exu_exu_lsu_rs1_d; // @[lsu.scala 124:46]
  assign lsu_lsc_ctl_io_lsu_exu_exu_lsu_rs2_d = io_lsu_exu_exu_lsu_rs2_d; // @[lsu.scala 124:46]
  assign lsu_lsc_ctl_io_lsu_p_valid = io_lsu_p_valid; // @[lsu.scala 125:46]
  assign lsu_lsc_ctl_io_lsu_p_bits_fast_int = io_lsu_p_bits_fast_int; // @[lsu.scala 125:46]
  assign lsu_lsc_ctl_io_lsu_p_bits_by = io_lsu_p_bits_by; // @[lsu.scala 125:46]
  assign lsu_lsc_ctl_io_lsu_p_bits_half = io_lsu_p_bits_half; // @[lsu.scala 125:46]
  assign lsu_lsc_ctl_io_lsu_p_bits_word = io_lsu_p_bits_word; // @[lsu.scala 125:46]
  assign lsu_lsc_ctl_io_lsu_p_bits_load = io_lsu_p_bits_load; // @[lsu.scala 125:46]
  assign lsu_lsc_ctl_io_lsu_p_bits_store = io_lsu_p_bits_store; // @[lsu.scala 125:46]
  assign lsu_lsc_ctl_io_lsu_p_bits_unsign = io_lsu_p_bits_unsign; // @[lsu.scala 125:46]
  assign lsu_lsc_ctl_io_lsu_p_bits_store_data_bypass_d = io_lsu_p_bits_store_data_bypass_d; // @[lsu.scala 125:46]
  assign lsu_lsc_ctl_io_lsu_p_bits_load_ldst_bypass_d = io_lsu_p_bits_load_ldst_bypass_d; // @[lsu.scala 125:46]
  assign lsu_lsc_ctl_io_dec_lsu_valid_raw_d = io_dec_lsu_valid_raw_d; // @[lsu.scala 126:46]
  assign lsu_lsc_ctl_io_dec_lsu_offset_d = io_dec_lsu_offset_d; // @[lsu.scala 127:46]
  assign lsu_lsc_ctl_io_picm_mask_data_m = dccm_ctl_io_picm_mask_data_m; // @[lsu.scala 128:46]
  assign lsu_lsc_ctl_io_bus_read_data_m = bus_intf_io_bus_read_data_m; // @[lsu.scala 129:46]
  assign lsu_lsc_ctl_io_dec_tlu_mrac_ff = io_dec_tlu_mrac_ff; // @[lsu.scala 131:46]
  assign lsu_lsc_ctl_io_dma_lsc_ctl_dma_dccm_req = io_lsu_dma_dma_lsc_ctl_dma_dccm_req; // @[lsu.scala 130:38]
  assign lsu_lsc_ctl_io_dma_lsc_ctl_dma_mem_addr = io_lsu_dma_dma_lsc_ctl_dma_mem_addr; // @[lsu.scala 130:38]
  assign lsu_lsc_ctl_io_dma_lsc_ctl_dma_mem_sz = io_lsu_dma_dma_lsc_ctl_dma_mem_sz; // @[lsu.scala 130:38]
  assign lsu_lsc_ctl_io_dma_lsc_ctl_dma_mem_write = io_lsu_dma_dma_lsc_ctl_dma_mem_write; // @[lsu.scala 130:38]
  assign lsu_lsc_ctl_io_dma_lsc_ctl_dma_mem_wdata = io_lsu_dma_dma_lsc_ctl_dma_mem_wdata; // @[lsu.scala 130:38]
  assign dccm_ctl_clock = clock;
  assign dccm_ctl_reset = reset;
  assign dccm_ctl_io_lsu_c2_m_clk = clkdomain_io_lsu_c2_m_clk; // @[lsu.scala 141:46]
  assign dccm_ctl_io_lsu_c2_r_clk = clkdomain_io_lsu_c2_r_clk; // @[lsu.scala 142:46]
  assign dccm_ctl_io_lsu_free_c2_clk = clkdomain_io_lsu_free_c2_clk; // @[lsu.scala 143:46]
  assign dccm_ctl_io_lsu_store_c1_r_clk = clkdomain_io_lsu_store_c1_r_clk; // @[lsu.scala 145:46]
  assign dccm_ctl_io_lsu_pkt_d_valid = lsu_lsc_ctl_io_lsu_pkt_d_valid; // @[lsu.scala 146:46]
  assign dccm_ctl_io_lsu_pkt_d_bits_word = lsu_lsc_ctl_io_lsu_pkt_d_bits_word; // @[lsu.scala 146:46]
  assign dccm_ctl_io_lsu_pkt_d_bits_dword = lsu_lsc_ctl_io_lsu_pkt_d_bits_dword; // @[lsu.scala 146:46]
  assign dccm_ctl_io_lsu_pkt_d_bits_load = lsu_lsc_ctl_io_lsu_pkt_d_bits_load; // @[lsu.scala 146:46]
  assign dccm_ctl_io_lsu_pkt_d_bits_store = lsu_lsc_ctl_io_lsu_pkt_d_bits_store; // @[lsu.scala 146:46]
  assign dccm_ctl_io_lsu_pkt_d_bits_dma = lsu_lsc_ctl_io_lsu_pkt_d_bits_dma; // @[lsu.scala 146:46]
  assign dccm_ctl_io_lsu_pkt_m_valid = lsu_lsc_ctl_io_lsu_pkt_m_valid; // @[lsu.scala 147:46]
  assign dccm_ctl_io_lsu_pkt_m_bits_by = lsu_lsc_ctl_io_lsu_pkt_m_bits_by; // @[lsu.scala 147:46]
  assign dccm_ctl_io_lsu_pkt_m_bits_half = lsu_lsc_ctl_io_lsu_pkt_m_bits_half; // @[lsu.scala 147:46]
  assign dccm_ctl_io_lsu_pkt_m_bits_word = lsu_lsc_ctl_io_lsu_pkt_m_bits_word; // @[lsu.scala 147:46]
  assign dccm_ctl_io_lsu_pkt_m_bits_load = lsu_lsc_ctl_io_lsu_pkt_m_bits_load; // @[lsu.scala 147:46]
  assign dccm_ctl_io_lsu_pkt_m_bits_store = lsu_lsc_ctl_io_lsu_pkt_m_bits_store; // @[lsu.scala 147:46]
  assign dccm_ctl_io_lsu_pkt_m_bits_dma = lsu_lsc_ctl_io_lsu_pkt_m_bits_dma; // @[lsu.scala 147:46]
  assign dccm_ctl_io_lsu_pkt_r_valid = lsu_lsc_ctl_io_lsu_pkt_r_valid; // @[lsu.scala 148:46]
  assign dccm_ctl_io_lsu_pkt_r_bits_by = lsu_lsc_ctl_io_lsu_pkt_r_bits_by; // @[lsu.scala 148:46]
  assign dccm_ctl_io_lsu_pkt_r_bits_half = lsu_lsc_ctl_io_lsu_pkt_r_bits_half; // @[lsu.scala 148:46]
  assign dccm_ctl_io_lsu_pkt_r_bits_word = lsu_lsc_ctl_io_lsu_pkt_r_bits_word; // @[lsu.scala 148:46]
  assign dccm_ctl_io_lsu_pkt_r_bits_load = lsu_lsc_ctl_io_lsu_pkt_r_bits_load; // @[lsu.scala 148:46]
  assign dccm_ctl_io_lsu_pkt_r_bits_store = lsu_lsc_ctl_io_lsu_pkt_r_bits_store; // @[lsu.scala 148:46]
  assign dccm_ctl_io_lsu_pkt_r_bits_dma = lsu_lsc_ctl_io_lsu_pkt_r_bits_dma; // @[lsu.scala 148:46]
  assign dccm_ctl_io_addr_in_dccm_d = lsu_lsc_ctl_io_addr_in_dccm_d; // @[lsu.scala 149:46]
  assign dccm_ctl_io_addr_in_dccm_m = lsu_lsc_ctl_io_addr_in_dccm_m; // @[lsu.scala 150:46]
  assign dccm_ctl_io_addr_in_dccm_r = lsu_lsc_ctl_io_addr_in_dccm_r; // @[lsu.scala 151:46]
  assign dccm_ctl_io_addr_in_pic_d = lsu_lsc_ctl_io_addr_in_pic_d; // @[lsu.scala 152:46]
  assign dccm_ctl_io_addr_in_pic_m = lsu_lsc_ctl_io_addr_in_pic_m; // @[lsu.scala 153:46]
  assign dccm_ctl_io_addr_in_pic_r = lsu_lsc_ctl_io_addr_in_pic_r; // @[lsu.scala 154:46]
  assign dccm_ctl_io_lsu_raw_fwd_lo_r = lsu_raw_fwd_lo_r; // @[lsu.scala 155:46]
  assign dccm_ctl_io_lsu_raw_fwd_hi_r = lsu_raw_fwd_hi_r; // @[lsu.scala 156:46]
  assign dccm_ctl_io_lsu_commit_r = lsu_lsc_ctl_io_lsu_commit_r; // @[lsu.scala 157:46]
  assign dccm_ctl_io_lsu_addr_d = lsu_lsc_ctl_io_lsu_addr_d; // @[lsu.scala 158:46]
  assign dccm_ctl_io_lsu_addr_m = lsu_lsc_ctl_io_lsu_addr_m[15:0]; // @[lsu.scala 159:46]
  assign dccm_ctl_io_lsu_addr_r = lsu_lsc_ctl_io_lsu_addr_r; // @[lsu.scala 160:46]
  assign dccm_ctl_io_end_addr_d = lsu_lsc_ctl_io_end_addr_d[15:0]; // @[lsu.scala 161:46]
  assign dccm_ctl_io_end_addr_m = lsu_lsc_ctl_io_end_addr_m[15:0]; // @[lsu.scala 162:46]
  assign dccm_ctl_io_end_addr_r = lsu_lsc_ctl_io_end_addr_r[15:0]; // @[lsu.scala 163:46]
  assign dccm_ctl_io_stbuf_reqvld_any = stbuf_io_stbuf_reqvld_any; // @[lsu.scala 164:46]
  assign dccm_ctl_io_stbuf_addr_any = stbuf_io_stbuf_addr_any; // @[lsu.scala 165:46]
  assign dccm_ctl_io_stbuf_data_any = stbuf_io_stbuf_data_any; // @[lsu.scala 166:46]
  assign dccm_ctl_io_stbuf_ecc_any = ecc_io_stbuf_ecc_any; // @[lsu.scala 167:46]
  assign dccm_ctl_io_stbuf_fwddata_hi_m = stbuf_io_stbuf_fwddata_hi_m; // @[lsu.scala 168:46]
  assign dccm_ctl_io_stbuf_fwddata_lo_m = stbuf_io_stbuf_fwddata_lo_m; // @[lsu.scala 169:46]
  assign dccm_ctl_io_stbuf_fwdbyteen_lo_m = stbuf_io_stbuf_fwdbyteen_lo_m; // @[lsu.scala 170:46]
  assign dccm_ctl_io_stbuf_fwdbyteen_hi_m = stbuf_io_stbuf_fwdbyteen_hi_m; // @[lsu.scala 171:46]
  assign dccm_ctl_io_lsu_double_ecc_error_r = ecc_io_lsu_double_ecc_error_r; // @[lsu.scala 172:46]
  assign dccm_ctl_io_single_ecc_error_hi_r = ecc_io_single_ecc_error_hi_r; // @[lsu.scala 173:46]
  assign dccm_ctl_io_single_ecc_error_lo_r = ecc_io_single_ecc_error_lo_r; // @[lsu.scala 174:46]
  assign dccm_ctl_io_sec_data_hi_r_ff = ecc_io_sec_data_hi_r_ff; // @[lsu.scala 177:46]
  assign dccm_ctl_io_sec_data_lo_r_ff = ecc_io_sec_data_lo_r_ff; // @[lsu.scala 178:46]
  assign dccm_ctl_io_sec_data_ecc_hi_r_ff = ecc_io_sec_data_ecc_hi_r_ff; // @[lsu.scala 179:46]
  assign dccm_ctl_io_sec_data_ecc_lo_r_ff = ecc_io_sec_data_ecc_lo_r_ff; // @[lsu.scala 180:46]
  assign dccm_ctl_io_lsu_double_ecc_error_m = ecc_io_lsu_double_ecc_error_m; // @[lsu.scala 181:46]
  assign dccm_ctl_io_sec_data_hi_m = ecc_io_sec_data_hi_m; // @[lsu.scala 182:46]
  assign dccm_ctl_io_sec_data_lo_m = ecc_io_sec_data_lo_m; // @[lsu.scala 183:46]
  assign dccm_ctl_io_store_data_m = lsu_lsc_ctl_io_store_data_m; // @[lsu.scala 184:46]
  assign dccm_ctl_io_dma_dccm_wen = _T_10 & lsu_lsc_ctl_io_addr_in_dccm_d; // @[lsu.scala 185:46]
  assign dccm_ctl_io_dma_pic_wen = _T_10 & lsu_lsc_ctl_io_addr_in_pic_d; // @[lsu.scala 186:46]
  assign dccm_ctl_io_dma_mem_tag_m = dma_mem_tag_m; // @[lsu.scala 187:46]
  assign dccm_ctl_io_dma_dccm_wdata_lo = dma_dccm_wdata[31:0]; // @[lsu.scala 188:46]
  assign dccm_ctl_io_dma_dccm_wdata_hi = dma_dccm_wdata[63:32]; // @[lsu.scala 189:46]
  assign dccm_ctl_io_dma_dccm_wdata_ecc_hi = ecc_io_dma_dccm_wdata_ecc_hi; // @[lsu.scala 190:46]
  assign dccm_ctl_io_dma_dccm_wdata_ecc_lo = ecc_io_dma_dccm_wdata_ecc_lo; // @[lsu.scala 191:46]
  assign dccm_ctl_io_dma_dccm_ctl_dma_mem_addr = io_lsu_dma_dma_dccm_ctl_dma_mem_addr; // @[lsu.scala 194:27]
  assign dccm_ctl_io_dma_dccm_ctl_dma_mem_wdata = io_lsu_dma_dma_dccm_ctl_dma_mem_wdata; // @[lsu.scala 194:27]
  assign dccm_ctl_io_dccm_rd_data_lo = io_dccm_rd_data_lo; // @[lsu.scala 195:11]
  assign dccm_ctl_io_dccm_rd_data_hi = io_dccm_rd_data_hi; // @[lsu.scala 195:11]
  assign dccm_ctl_io_lsu_pic_picm_rd_data = io_lsu_pic_picm_rd_data; // @[lsu.scala 196:14]
  assign dccm_ctl_io_scan_mode = io_scan_mode; // @[lsu.scala 192:46]
  assign stbuf_clock = clock;
  assign stbuf_reset = reset;
  assign stbuf_io_lsu_c1_m_clk = clkdomain_io_lsu_c1_m_clk; // @[lsu.scala 199:49]
  assign stbuf_io_lsu_c1_r_clk = clkdomain_io_lsu_c1_r_clk; // @[lsu.scala 200:48]
  assign stbuf_io_lsu_stbuf_c1_clk = clkdomain_io_lsu_stbuf_c1_clk; // @[lsu.scala 201:54]
  assign stbuf_io_lsu_free_c2_clk = clkdomain_io_lsu_free_c2_clk; // @[lsu.scala 202:54]
  assign stbuf_io_lsu_pkt_m_valid = lsu_lsc_ctl_io_lsu_pkt_m_valid; // @[lsu.scala 203:48]
  assign stbuf_io_lsu_pkt_m_bits_store = lsu_lsc_ctl_io_lsu_pkt_m_bits_store; // @[lsu.scala 203:48]
  assign stbuf_io_lsu_pkt_m_bits_dma = lsu_lsc_ctl_io_lsu_pkt_m_bits_dma; // @[lsu.scala 203:48]
  assign stbuf_io_lsu_pkt_r_valid = lsu_lsc_ctl_io_lsu_pkt_r_valid; // @[lsu.scala 204:48]
  assign stbuf_io_lsu_pkt_r_bits_by = lsu_lsc_ctl_io_lsu_pkt_r_bits_by; // @[lsu.scala 204:48]
  assign stbuf_io_lsu_pkt_r_bits_half = lsu_lsc_ctl_io_lsu_pkt_r_bits_half; // @[lsu.scala 204:48]
  assign stbuf_io_lsu_pkt_r_bits_word = lsu_lsc_ctl_io_lsu_pkt_r_bits_word; // @[lsu.scala 204:48]
  assign stbuf_io_lsu_pkt_r_bits_dword = lsu_lsc_ctl_io_lsu_pkt_r_bits_dword; // @[lsu.scala 204:48]
  assign stbuf_io_lsu_pkt_r_bits_store = lsu_lsc_ctl_io_lsu_pkt_r_bits_store; // @[lsu.scala 204:48]
  assign stbuf_io_lsu_pkt_r_bits_dma = lsu_lsc_ctl_io_lsu_pkt_r_bits_dma; // @[lsu.scala 204:48]
  assign stbuf_io_store_stbuf_reqvld_r = _T_28 & _T_19; // @[lsu.scala 205:48]
  assign stbuf_io_lsu_commit_r = lsu_lsc_ctl_io_lsu_commit_r; // @[lsu.scala 206:49]
  assign stbuf_io_dec_lsu_valid_raw_d = io_dec_lsu_valid_raw_d; // @[lsu.scala 207:49]
  assign stbuf_io_store_data_hi_r = dccm_ctl_io_store_data_hi_r; // @[lsu.scala 208:62]
  assign stbuf_io_store_data_lo_r = dccm_ctl_io_store_data_lo_r; // @[lsu.scala 209:62]
  assign stbuf_io_store_datafn_hi_r = dccm_ctl_io_store_datafn_hi_r; // @[lsu.scala 210:49]
  assign stbuf_io_store_datafn_lo_r = dccm_ctl_io_store_datafn_lo_r; // @[lsu.scala 211:56]
  assign stbuf_io_lsu_stbuf_commit_any = dccm_ctl_io_lsu_stbuf_commit_any; // @[lsu.scala 212:52]
  assign stbuf_io_lsu_addr_d = lsu_lsc_ctl_io_lsu_addr_d[15:0]; // @[lsu.scala 213:64]
  assign stbuf_io_lsu_addr_m = lsu_lsc_ctl_io_lsu_addr_m; // @[lsu.scala 214:64]
  assign stbuf_io_lsu_addr_r = lsu_lsc_ctl_io_lsu_addr_r; // @[lsu.scala 215:64]
  assign stbuf_io_end_addr_d = lsu_lsc_ctl_io_end_addr_d[15:0]; // @[lsu.scala 216:64]
  assign stbuf_io_end_addr_m = lsu_lsc_ctl_io_end_addr_m; // @[lsu.scala 217:64]
  assign stbuf_io_end_addr_r = lsu_lsc_ctl_io_end_addr_r; // @[lsu.scala 218:64]
  assign stbuf_io_addr_in_dccm_m = lsu_lsc_ctl_io_addr_in_dccm_m; // @[lsu.scala 219:49]
  assign stbuf_io_addr_in_dccm_r = lsu_lsc_ctl_io_addr_in_dccm_r; // @[lsu.scala 220:56]
  assign stbuf_io_scan_mode = io_scan_mode; // @[lsu.scala 222:49]
  assign ecc_clock = clock;
  assign ecc_reset = reset;
  assign ecc_io_lsu_c2_r_clk = clkdomain_io_lsu_c2_r_clk; // @[lsu.scala 226:52]
  assign ecc_io_lsu_pkt_m_valid = lsu_lsc_ctl_io_lsu_pkt_m_valid; // @[lsu.scala 227:52]
  assign ecc_io_lsu_pkt_m_bits_load = lsu_lsc_ctl_io_lsu_pkt_m_bits_load; // @[lsu.scala 227:52]
  assign ecc_io_lsu_pkt_m_bits_store = lsu_lsc_ctl_io_lsu_pkt_m_bits_store; // @[lsu.scala 227:52]
  assign ecc_io_lsu_pkt_m_bits_dma = lsu_lsc_ctl_io_lsu_pkt_m_bits_dma; // @[lsu.scala 227:52]
  assign ecc_io_stbuf_data_any = stbuf_io_stbuf_data_any; // @[lsu.scala 229:54]
  assign ecc_io_dec_tlu_core_ecc_disable = io_dec_tlu_core_ecc_disable; // @[lsu.scala 230:50]
  assign ecc_io_lsu_addr_m = lsu_lsc_ctl_io_lsu_addr_m[15:0]; // @[lsu.scala 235:58]
  assign ecc_io_end_addr_m = lsu_lsc_ctl_io_end_addr_m[15:0]; // @[lsu.scala 236:58]
  assign ecc_io_dccm_rdata_hi_m = dccm_ctl_io_dccm_rdata_hi_m; // @[lsu.scala 239:54]
  assign ecc_io_dccm_rdata_lo_m = dccm_ctl_io_dccm_rdata_lo_m; // @[lsu.scala 240:54]
  assign ecc_io_dccm_data_ecc_hi_m = dccm_ctl_io_dccm_data_ecc_hi_m; // @[lsu.scala 243:50]
  assign ecc_io_dccm_data_ecc_lo_m = dccm_ctl_io_dccm_data_ecc_lo_m; // @[lsu.scala 244:50]
  assign ecc_io_ld_single_ecc_error_r = dccm_ctl_io_ld_single_ecc_error_r; // @[lsu.scala 245:50]
  assign ecc_io_ld_single_ecc_error_r_ff = dccm_ctl_io_ld_single_ecc_error_r_ff; // @[lsu.scala 246:50]
  assign ecc_io_lsu_dccm_rden_m = dccm_ctl_io_lsu_dccm_rden_m; // @[lsu.scala 247:50]
  assign ecc_io_addr_in_dccm_m = lsu_lsc_ctl_io_addr_in_dccm_m; // @[lsu.scala 248:50]
  assign ecc_io_dma_dccm_wen = _T_10 & lsu_lsc_ctl_io_addr_in_dccm_d; // @[lsu.scala 249:50]
  assign ecc_io_dma_dccm_wdata_lo = dma_dccm_wdata[31:0]; // @[lsu.scala 250:50]
  assign ecc_io_dma_dccm_wdata_hi = dma_dccm_wdata[63:32]; // @[lsu.scala 251:50]
  assign ecc_io_scan_mode = io_scan_mode; // @[lsu.scala 252:50]
  assign trigger_io_trigger_pkt_any_0_select = io_trigger_pkt_any_0_select; // @[lsu.scala 256:50]
  assign trigger_io_trigger_pkt_any_0_match_pkt = io_trigger_pkt_any_0_match_pkt; // @[lsu.scala 256:50]
  assign trigger_io_trigger_pkt_any_0_store = io_trigger_pkt_any_0_store; // @[lsu.scala 256:50]
  assign trigger_io_trigger_pkt_any_0_load = io_trigger_pkt_any_0_load; // @[lsu.scala 256:50]
  assign trigger_io_trigger_pkt_any_0_tdata2 = io_trigger_pkt_any_0_tdata2; // @[lsu.scala 256:50]
  assign trigger_io_trigger_pkt_any_1_select = io_trigger_pkt_any_1_select; // @[lsu.scala 256:50]
  assign trigger_io_trigger_pkt_any_1_match_pkt = io_trigger_pkt_any_1_match_pkt; // @[lsu.scala 256:50]
  assign trigger_io_trigger_pkt_any_1_store = io_trigger_pkt_any_1_store; // @[lsu.scala 256:50]
  assign trigger_io_trigger_pkt_any_1_load = io_trigger_pkt_any_1_load; // @[lsu.scala 256:50]
  assign trigger_io_trigger_pkt_any_1_tdata2 = io_trigger_pkt_any_1_tdata2; // @[lsu.scala 256:50]
  assign trigger_io_trigger_pkt_any_2_select = io_trigger_pkt_any_2_select; // @[lsu.scala 256:50]
  assign trigger_io_trigger_pkt_any_2_match_pkt = io_trigger_pkt_any_2_match_pkt; // @[lsu.scala 256:50]
  assign trigger_io_trigger_pkt_any_2_store = io_trigger_pkt_any_2_store; // @[lsu.scala 256:50]
  assign trigger_io_trigger_pkt_any_2_load = io_trigger_pkt_any_2_load; // @[lsu.scala 256:50]
  assign trigger_io_trigger_pkt_any_2_tdata2 = io_trigger_pkt_any_2_tdata2; // @[lsu.scala 256:50]
  assign trigger_io_trigger_pkt_any_3_select = io_trigger_pkt_any_3_select; // @[lsu.scala 256:50]
  assign trigger_io_trigger_pkt_any_3_match_pkt = io_trigger_pkt_any_3_match_pkt; // @[lsu.scala 256:50]
  assign trigger_io_trigger_pkt_any_3_store = io_trigger_pkt_any_3_store; // @[lsu.scala 256:50]
  assign trigger_io_trigger_pkt_any_3_load = io_trigger_pkt_any_3_load; // @[lsu.scala 256:50]
  assign trigger_io_trigger_pkt_any_3_tdata2 = io_trigger_pkt_any_3_tdata2; // @[lsu.scala 256:50]
  assign trigger_io_lsu_pkt_m_valid = lsu_lsc_ctl_io_lsu_pkt_m_valid; // @[lsu.scala 257:50]
  assign trigger_io_lsu_pkt_m_bits_half = lsu_lsc_ctl_io_lsu_pkt_m_bits_half; // @[lsu.scala 257:50]
  assign trigger_io_lsu_pkt_m_bits_word = lsu_lsc_ctl_io_lsu_pkt_m_bits_word; // @[lsu.scala 257:50]
  assign trigger_io_lsu_pkt_m_bits_load = lsu_lsc_ctl_io_lsu_pkt_m_bits_load; // @[lsu.scala 257:50]
  assign trigger_io_lsu_pkt_m_bits_store = lsu_lsc_ctl_io_lsu_pkt_m_bits_store; // @[lsu.scala 257:50]
  assign trigger_io_lsu_pkt_m_bits_dma = lsu_lsc_ctl_io_lsu_pkt_m_bits_dma; // @[lsu.scala 257:50]
  assign trigger_io_lsu_addr_m = lsu_lsc_ctl_io_lsu_addr_m; // @[lsu.scala 258:50]
  assign trigger_io_store_data_m = lsu_lsc_ctl_io_store_data_m; // @[lsu.scala 259:50]
  assign clkdomain_clock = clock;
  assign clkdomain_reset = reset;
  assign clkdomain_io_free_clk = io_free_clk; // @[lsu.scala 265:50]
  assign clkdomain_io_clk_override = io_clk_override; // @[lsu.scala 266:50]
  assign clkdomain_io_dma_dccm_req = io_lsu_dma_dma_lsc_ctl_dma_dccm_req; // @[lsu.scala 268:50]
  assign clkdomain_io_ldst_stbuf_reqvld_r = stbuf_io_ldst_stbuf_reqvld_r; // @[lsu.scala 269:50]
  assign clkdomain_io_stbuf_reqvld_any = stbuf_io_stbuf_reqvld_any; // @[lsu.scala 270:50]
  assign clkdomain_io_stbuf_reqvld_flushed_any = stbuf_io_stbuf_reqvld_flushed_any; // @[lsu.scala 271:50]
  assign clkdomain_io_lsu_busreq_r = bus_intf_io_lsu_busreq_r; // @[lsu.scala 272:50]
  assign clkdomain_io_lsu_bus_buffer_pend_any = bus_intf_io_lsu_bus_buffer_pend_any; // @[lsu.scala 273:50]
  assign clkdomain_io_lsu_bus_buffer_empty_any = bus_intf_io_lsu_bus_buffer_empty_any; // @[lsu.scala 274:50]
  assign clkdomain_io_lsu_stbuf_empty_any = stbuf_io_lsu_stbuf_empty_any; // @[lsu.scala 275:50]
  assign clkdomain_io_lsu_bus_clk_en = io_lsu_bus_clk_en; // @[lsu.scala 276:50]
  assign clkdomain_io_lsu_p_valid = io_lsu_p_valid; // @[lsu.scala 277:50]
  assign clkdomain_io_lsu_pkt_d_valid = lsu_lsc_ctl_io_lsu_pkt_d_valid; // @[lsu.scala 278:50]
  assign clkdomain_io_lsu_pkt_d_bits_store = lsu_lsc_ctl_io_lsu_pkt_d_bits_store; // @[lsu.scala 278:50]
  assign clkdomain_io_lsu_pkt_m_valid = lsu_lsc_ctl_io_lsu_pkt_m_valid; // @[lsu.scala 279:50]
  assign clkdomain_io_lsu_pkt_m_bits_store = lsu_lsc_ctl_io_lsu_pkt_m_bits_store; // @[lsu.scala 279:50]
  assign clkdomain_io_lsu_pkt_r_valid = lsu_lsc_ctl_io_lsu_pkt_r_valid; // @[lsu.scala 280:50]
  assign clkdomain_io_scan_mode = io_scan_mode; // @[lsu.scala 281:50]
  assign bus_intf_clock = clock;
  assign bus_intf_reset = reset;
  assign bus_intf_io_scan_mode = io_scan_mode; // @[lsu.scala 285:49]
  assign bus_intf_io_tlu_busbuff_dec_tlu_external_ldfwd_disable = io_lsu_dec_tlu_busbuff_dec_tlu_external_ldfwd_disable; // @[lsu.scala 286:26]
  assign bus_intf_io_tlu_busbuff_dec_tlu_wb_coalescing_disable = io_lsu_dec_tlu_busbuff_dec_tlu_wb_coalescing_disable; // @[lsu.scala 286:26]
  assign bus_intf_io_tlu_busbuff_dec_tlu_sideeffect_posted_disable = io_lsu_dec_tlu_busbuff_dec_tlu_sideeffect_posted_disable; // @[lsu.scala 286:26]
  assign bus_intf_io_lsu_c1_m_clk = clkdomain_io_lsu_c1_m_clk; // @[lsu.scala 287:49]
  assign bus_intf_io_lsu_c1_r_clk = clkdomain_io_lsu_c1_r_clk; // @[lsu.scala 288:49]
  assign bus_intf_io_lsu_c2_r_clk = clkdomain_io_lsu_c2_r_clk; // @[lsu.scala 289:49]
  assign bus_intf_io_lsu_bus_ibuf_c1_clk = clkdomain_io_lsu_bus_ibuf_c1_clk; // @[lsu.scala 290:49]
  assign bus_intf_io_lsu_bus_obuf_c1_clk = clkdomain_io_lsu_bus_obuf_c1_clk; // @[lsu.scala 291:49]
  assign bus_intf_io_lsu_bus_buf_c1_clk = clkdomain_io_lsu_bus_buf_c1_clk; // @[lsu.scala 292:49]
  assign bus_intf_io_lsu_free_c2_clk = clkdomain_io_lsu_free_c2_clk; // @[lsu.scala 293:49]
  assign bus_intf_io_free_clk = io_free_clk; // @[lsu.scala 294:49]
  assign bus_intf_io_lsu_busm_clk = clkdomain_io_lsu_busm_clk; // @[lsu.scala 295:49]
  assign bus_intf_io_dec_lsu_valid_raw_d = io_dec_lsu_valid_raw_d; // @[lsu.scala 296:49]
  assign bus_intf_io_lsu_busreq_m = _T_39 & _T_40; // @[lsu.scala 297:49]
  assign bus_intf_io_lsu_pkt_m_valid = lsu_lsc_ctl_io_lsu_pkt_m_valid; // @[lsu.scala 305:49]
  assign bus_intf_io_lsu_pkt_m_bits_by = lsu_lsc_ctl_io_lsu_pkt_m_bits_by; // @[lsu.scala 305:49]
  assign bus_intf_io_lsu_pkt_m_bits_half = lsu_lsc_ctl_io_lsu_pkt_m_bits_half; // @[lsu.scala 305:49]
  assign bus_intf_io_lsu_pkt_m_bits_word = lsu_lsc_ctl_io_lsu_pkt_m_bits_word; // @[lsu.scala 305:49]
  assign bus_intf_io_lsu_pkt_m_bits_load = lsu_lsc_ctl_io_lsu_pkt_m_bits_load; // @[lsu.scala 305:49]
  assign bus_intf_io_lsu_pkt_r_valid = lsu_lsc_ctl_io_lsu_pkt_r_valid; // @[lsu.scala 306:49]
  assign bus_intf_io_lsu_pkt_r_bits_by = lsu_lsc_ctl_io_lsu_pkt_r_bits_by; // @[lsu.scala 306:49]
  assign bus_intf_io_lsu_pkt_r_bits_half = lsu_lsc_ctl_io_lsu_pkt_r_bits_half; // @[lsu.scala 306:49]
  assign bus_intf_io_lsu_pkt_r_bits_word = lsu_lsc_ctl_io_lsu_pkt_r_bits_word; // @[lsu.scala 306:49]
  assign bus_intf_io_lsu_pkt_r_bits_load = lsu_lsc_ctl_io_lsu_pkt_r_bits_load; // @[lsu.scala 306:49]
  assign bus_intf_io_lsu_pkt_r_bits_store = lsu_lsc_ctl_io_lsu_pkt_r_bits_store; // @[lsu.scala 306:49]
  assign bus_intf_io_lsu_pkt_r_bits_unsign = lsu_lsc_ctl_io_lsu_pkt_r_bits_unsign; // @[lsu.scala 306:49]
  assign bus_intf_io_lsu_addr_d = lsu_lsc_ctl_io_lsu_addr_d; // @[lsu.scala 298:49]
  assign bus_intf_io_lsu_addr_m = lsu_lsc_ctl_io_lsu_addr_m; // @[lsu.scala 299:49]
  assign bus_intf_io_lsu_addr_r = lsu_lsc_ctl_io_lsu_addr_r; // @[lsu.scala 300:49]
  assign bus_intf_io_end_addr_d = lsu_lsc_ctl_io_end_addr_d; // @[lsu.scala 301:49]
  assign bus_intf_io_end_addr_m = lsu_lsc_ctl_io_end_addr_m; // @[lsu.scala 302:49]
  assign bus_intf_io_end_addr_r = lsu_lsc_ctl_io_end_addr_r; // @[lsu.scala 303:49]
  assign bus_intf_io_store_data_r = dccm_ctl_io_store_data_r; // @[lsu.scala 304:49]
  assign bus_intf_io_dec_tlu_force_halt = io_dec_tlu_force_halt; // @[lsu.scala 307:49]
  assign bus_intf_io_lsu_commit_r = lsu_lsc_ctl_io_lsu_commit_r; // @[lsu.scala 308:49]
  assign bus_intf_io_is_sideeffects_m = lsu_lsc_ctl_io_is_sideeffects_m; // @[lsu.scala 309:49]
  assign bus_intf_io_flush_m_up = io_dec_tlu_flush_lower_r; // @[lsu.scala 310:49]
  assign bus_intf_io_flush_r = io_dec_tlu_i0_kill_writeb_r; // @[lsu.scala 311:49]
  assign bus_intf_io_lsu_bus_clk_en = io_lsu_bus_clk_en; // @[lsu.scala 315:49]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  dma_mem_tag_m = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  lsu_raw_fwd_hi_r = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  lsu_raw_fwd_lo_r = _RAND_2[0:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    dma_mem_tag_m = 3'h0;
  end
  if (reset) begin
    lsu_raw_fwd_hi_r = 1'h0;
  end
  if (reset) begin
    lsu_raw_fwd_lo_r = 1'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clkdomain_io_lsu_c1_m_clk or posedge reset) begin
    if (reset) begin
      dma_mem_tag_m <= 3'h0;
    end else begin
      dma_mem_tag_m <= io_lsu_dma_dma_mem_tag;
    end
  end
  always @(posedge clkdomain_io_lsu_c2_r_clk or posedge reset) begin
    if (reset) begin
      lsu_raw_fwd_hi_r <= 1'h0;
    end else begin
      lsu_raw_fwd_hi_r <= |stbuf_io_stbuf_fwdbyteen_hi_m;
    end
  end
  always @(posedge clkdomain_io_lsu_c2_r_clk or posedge reset) begin
    if (reset) begin
      lsu_raw_fwd_lo_r <= 1'h0;
    end else begin
      lsu_raw_fwd_lo_r <= |stbuf_io_stbuf_fwdbyteen_lo_m;
    end
  end
endmodule
module pic_ctrl(
  input         clock,
  input         reset,
  input         io_scan_mode,
  input         io_free_clk,
  input         io_active_clk,
  input         io_clk_override,
  input  [31:0] io_extintsrc_req,
  input         io_lsu_pic_picm_wren,
  input         io_lsu_pic_picm_rden,
  input         io_lsu_pic_picm_mken,
  input  [31:0] io_lsu_pic_picm_rdaddr,
  input  [31:0] io_lsu_pic_picm_wraddr,
  input  [31:0] io_lsu_pic_picm_wr_data,
  output [31:0] io_lsu_pic_picm_rd_data,
  output [7:0]  io_dec_pic_pic_claimid,
  output [3:0]  io_dec_pic_pic_pl,
  output        io_dec_pic_mhwakeup,
  input  [3:0]  io_dec_pic_dec_tlu_meicurpl,
  input  [3:0]  io_dec_pic_dec_tlu_meipt,
  output        io_dec_pic_mexintpend
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
`endif // RANDOMIZE_REG_INIT
  wire  rvclkhdr_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_1_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_1_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_1_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_1_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_2_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_2_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_2_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_2_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_3_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_3_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_3_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_3_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_4_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_4_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_4_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_4_io_scan_mode; // @[lib.scala 343:22]
  wire  pic_raddr_c1_clk = rvclkhdr_io_l1clk; // @[pic_ctrl.scala 95:42 pic_ctrl.scala 132:21]
  reg [31:0] picm_raddr_ff; // @[pic_ctrl.scala 101:56]
  wire  pic_data_c1_clk = rvclkhdr_1_io_l1clk; // @[pic_ctrl.scala 96:42 pic_ctrl.scala 133:21]
  reg [31:0] picm_waddr_ff; // @[pic_ctrl.scala 102:57]
  reg  picm_wren_ff; // @[pic_ctrl.scala 103:55]
  reg  picm_rden_ff; // @[pic_ctrl.scala 104:55]
  reg  picm_mken_ff; // @[pic_ctrl.scala 105:55]
  reg [31:0] picm_wr_data_ff; // @[pic_ctrl.scala 106:58]
  wire [31:0] _T_6 = picm_raddr_ff ^ 32'hf00c2000; // @[pic_ctrl.scala 108:59]
  wire [31:0] temp_raddr_intenable_base_match = ~_T_6; // @[pic_ctrl.scala 108:43]
  wire  raddr_intenable_base_match = &temp_raddr_intenable_base_match[31:7]; // @[pic_ctrl.scala 109:89]
  wire  raddr_intpriority_base_match = picm_raddr_ff[31:7] == 25'h1e01800; // @[pic_ctrl.scala 111:71]
  wire  raddr_config_gw_base_match = picm_raddr_ff[31:7] == 25'h1e01880; // @[pic_ctrl.scala 112:71]
  wire  raddr_config_pic_match = picm_raddr_ff == 32'hf00c3000; // @[pic_ctrl.scala 113:71]
  wire  addr_intpend_base_match = picm_raddr_ff[31:6] == 26'h3c03040; // @[pic_ctrl.scala 114:71]
  wire  waddr_config_pic_match = picm_waddr_ff == 32'hf00c3000; // @[pic_ctrl.scala 116:71]
  wire  addr_clear_gw_base_match = picm_waddr_ff[31:7] == 25'h1e018a0; // @[pic_ctrl.scala 117:71]
  wire  waddr_intpriority_base_match = picm_waddr_ff[31:7] == 25'h1e01800; // @[pic_ctrl.scala 118:71]
  wire  waddr_intenable_base_match = picm_waddr_ff[31:7] == 25'h1e01840; // @[pic_ctrl.scala 119:71]
  wire  waddr_config_gw_base_match = picm_waddr_ff[31:7] == 25'h1e01880; // @[pic_ctrl.scala 120:71]
  wire  _T_17 = picm_rden_ff & picm_wren_ff; // @[pic_ctrl.scala 121:53]
  wire  _T_18 = picm_raddr_ff == picm_waddr_ff; // @[pic_ctrl.scala 121:86]
  wire  picm_bypass_ff = _T_17 & _T_18; // @[pic_ctrl.scala 121:68]
  wire  _T_19 = io_lsu_pic_picm_mken | io_lsu_pic_picm_rden; // @[pic_ctrl.scala 125:50]
  wire  _T_20 = waddr_intpriority_base_match & picm_wren_ff; // @[pic_ctrl.scala 127:59]
  wire  _T_21 = raddr_intpriority_base_match & picm_rden_ff; // @[pic_ctrl.scala 127:108]
  wire  _T_22 = _T_20 | _T_21; // @[pic_ctrl.scala 127:76]
  wire  _T_23 = waddr_intenable_base_match & picm_wren_ff; // @[pic_ctrl.scala 128:57]
  wire  _T_24 = raddr_intenable_base_match & picm_rden_ff; // @[pic_ctrl.scala 128:104]
  wire  _T_25 = _T_23 | _T_24; // @[pic_ctrl.scala 128:74]
  wire  _T_26 = waddr_config_gw_base_match & picm_wren_ff; // @[pic_ctrl.scala 129:59]
  wire  _T_27 = raddr_config_gw_base_match & picm_rden_ff; // @[pic_ctrl.scala 129:108]
  wire  _T_28 = _T_26 | _T_27; // @[pic_ctrl.scala 129:76]
  reg [30:0] _T_33; // @[lib.scala 37:81]
  reg [30:0] _T_34; // @[lib.scala 37:58]
  wire [31:0] extintsrc_req_sync = {_T_34,io_extintsrc_req[0]}; // @[Cat.scala 29:58]
  wire  _T_37 = picm_waddr_ff[6:2] == 5'h1; // @[pic_ctrl.scala 141:139]
  wire  _T_38 = waddr_intpriority_base_match & _T_37; // @[pic_ctrl.scala 141:106]
  wire  intpriority_reg_we_1 = _T_38 & picm_wren_ff; // @[pic_ctrl.scala 141:153]
  wire  _T_40 = picm_waddr_ff[6:2] == 5'h2; // @[pic_ctrl.scala 141:139]
  wire  _T_41 = waddr_intpriority_base_match & _T_40; // @[pic_ctrl.scala 141:106]
  wire  intpriority_reg_we_2 = _T_41 & picm_wren_ff; // @[pic_ctrl.scala 141:153]
  wire  _T_43 = picm_waddr_ff[6:2] == 5'h3; // @[pic_ctrl.scala 141:139]
  wire  _T_44 = waddr_intpriority_base_match & _T_43; // @[pic_ctrl.scala 141:106]
  wire  intpriority_reg_we_3 = _T_44 & picm_wren_ff; // @[pic_ctrl.scala 141:153]
  wire  _T_46 = picm_waddr_ff[6:2] == 5'h4; // @[pic_ctrl.scala 141:139]
  wire  _T_47 = waddr_intpriority_base_match & _T_46; // @[pic_ctrl.scala 141:106]
  wire  intpriority_reg_we_4 = _T_47 & picm_wren_ff; // @[pic_ctrl.scala 141:153]
  wire  _T_49 = picm_waddr_ff[6:2] == 5'h5; // @[pic_ctrl.scala 141:139]
  wire  _T_50 = waddr_intpriority_base_match & _T_49; // @[pic_ctrl.scala 141:106]
  wire  intpriority_reg_we_5 = _T_50 & picm_wren_ff; // @[pic_ctrl.scala 141:153]
  wire  _T_52 = picm_waddr_ff[6:2] == 5'h6; // @[pic_ctrl.scala 141:139]
  wire  _T_53 = waddr_intpriority_base_match & _T_52; // @[pic_ctrl.scala 141:106]
  wire  intpriority_reg_we_6 = _T_53 & picm_wren_ff; // @[pic_ctrl.scala 141:153]
  wire  _T_55 = picm_waddr_ff[6:2] == 5'h7; // @[pic_ctrl.scala 141:139]
  wire  _T_56 = waddr_intpriority_base_match & _T_55; // @[pic_ctrl.scala 141:106]
  wire  intpriority_reg_we_7 = _T_56 & picm_wren_ff; // @[pic_ctrl.scala 141:153]
  wire  _T_58 = picm_waddr_ff[6:2] == 5'h8; // @[pic_ctrl.scala 141:139]
  wire  _T_59 = waddr_intpriority_base_match & _T_58; // @[pic_ctrl.scala 141:106]
  wire  intpriority_reg_we_8 = _T_59 & picm_wren_ff; // @[pic_ctrl.scala 141:153]
  wire  _T_61 = picm_waddr_ff[6:2] == 5'h9; // @[pic_ctrl.scala 141:139]
  wire  _T_62 = waddr_intpriority_base_match & _T_61; // @[pic_ctrl.scala 141:106]
  wire  intpriority_reg_we_9 = _T_62 & picm_wren_ff; // @[pic_ctrl.scala 141:153]
  wire  _T_64 = picm_waddr_ff[6:2] == 5'ha; // @[pic_ctrl.scala 141:139]
  wire  _T_65 = waddr_intpriority_base_match & _T_64; // @[pic_ctrl.scala 141:106]
  wire  intpriority_reg_we_10 = _T_65 & picm_wren_ff; // @[pic_ctrl.scala 141:153]
  wire  _T_67 = picm_waddr_ff[6:2] == 5'hb; // @[pic_ctrl.scala 141:139]
  wire  _T_68 = waddr_intpriority_base_match & _T_67; // @[pic_ctrl.scala 141:106]
  wire  intpriority_reg_we_11 = _T_68 & picm_wren_ff; // @[pic_ctrl.scala 141:153]
  wire  _T_70 = picm_waddr_ff[6:2] == 5'hc; // @[pic_ctrl.scala 141:139]
  wire  _T_71 = waddr_intpriority_base_match & _T_70; // @[pic_ctrl.scala 141:106]
  wire  intpriority_reg_we_12 = _T_71 & picm_wren_ff; // @[pic_ctrl.scala 141:153]
  wire  _T_73 = picm_waddr_ff[6:2] == 5'hd; // @[pic_ctrl.scala 141:139]
  wire  _T_74 = waddr_intpriority_base_match & _T_73; // @[pic_ctrl.scala 141:106]
  wire  intpriority_reg_we_13 = _T_74 & picm_wren_ff; // @[pic_ctrl.scala 141:153]
  wire  _T_76 = picm_waddr_ff[6:2] == 5'he; // @[pic_ctrl.scala 141:139]
  wire  _T_77 = waddr_intpriority_base_match & _T_76; // @[pic_ctrl.scala 141:106]
  wire  intpriority_reg_we_14 = _T_77 & picm_wren_ff; // @[pic_ctrl.scala 141:153]
  wire  _T_79 = picm_waddr_ff[6:2] == 5'hf; // @[pic_ctrl.scala 141:139]
  wire  _T_80 = waddr_intpriority_base_match & _T_79; // @[pic_ctrl.scala 141:106]
  wire  intpriority_reg_we_15 = _T_80 & picm_wren_ff; // @[pic_ctrl.scala 141:153]
  wire  _T_82 = picm_waddr_ff[6:2] == 5'h10; // @[pic_ctrl.scala 141:139]
  wire  _T_83 = waddr_intpriority_base_match & _T_82; // @[pic_ctrl.scala 141:106]
  wire  intpriority_reg_we_16 = _T_83 & picm_wren_ff; // @[pic_ctrl.scala 141:153]
  wire  _T_85 = picm_waddr_ff[6:2] == 5'h11; // @[pic_ctrl.scala 141:139]
  wire  _T_86 = waddr_intpriority_base_match & _T_85; // @[pic_ctrl.scala 141:106]
  wire  intpriority_reg_we_17 = _T_86 & picm_wren_ff; // @[pic_ctrl.scala 141:153]
  wire  _T_88 = picm_waddr_ff[6:2] == 5'h12; // @[pic_ctrl.scala 141:139]
  wire  _T_89 = waddr_intpriority_base_match & _T_88; // @[pic_ctrl.scala 141:106]
  wire  intpriority_reg_we_18 = _T_89 & picm_wren_ff; // @[pic_ctrl.scala 141:153]
  wire  _T_91 = picm_waddr_ff[6:2] == 5'h13; // @[pic_ctrl.scala 141:139]
  wire  _T_92 = waddr_intpriority_base_match & _T_91; // @[pic_ctrl.scala 141:106]
  wire  intpriority_reg_we_19 = _T_92 & picm_wren_ff; // @[pic_ctrl.scala 141:153]
  wire  _T_94 = picm_waddr_ff[6:2] == 5'h14; // @[pic_ctrl.scala 141:139]
  wire  _T_95 = waddr_intpriority_base_match & _T_94; // @[pic_ctrl.scala 141:106]
  wire  intpriority_reg_we_20 = _T_95 & picm_wren_ff; // @[pic_ctrl.scala 141:153]
  wire  _T_97 = picm_waddr_ff[6:2] == 5'h15; // @[pic_ctrl.scala 141:139]
  wire  _T_98 = waddr_intpriority_base_match & _T_97; // @[pic_ctrl.scala 141:106]
  wire  intpriority_reg_we_21 = _T_98 & picm_wren_ff; // @[pic_ctrl.scala 141:153]
  wire  _T_100 = picm_waddr_ff[6:2] == 5'h16; // @[pic_ctrl.scala 141:139]
  wire  _T_101 = waddr_intpriority_base_match & _T_100; // @[pic_ctrl.scala 141:106]
  wire  intpriority_reg_we_22 = _T_101 & picm_wren_ff; // @[pic_ctrl.scala 141:153]
  wire  _T_103 = picm_waddr_ff[6:2] == 5'h17; // @[pic_ctrl.scala 141:139]
  wire  _T_104 = waddr_intpriority_base_match & _T_103; // @[pic_ctrl.scala 141:106]
  wire  intpriority_reg_we_23 = _T_104 & picm_wren_ff; // @[pic_ctrl.scala 141:153]
  wire  _T_106 = picm_waddr_ff[6:2] == 5'h18; // @[pic_ctrl.scala 141:139]
  wire  _T_107 = waddr_intpriority_base_match & _T_106; // @[pic_ctrl.scala 141:106]
  wire  intpriority_reg_we_24 = _T_107 & picm_wren_ff; // @[pic_ctrl.scala 141:153]
  wire  _T_109 = picm_waddr_ff[6:2] == 5'h19; // @[pic_ctrl.scala 141:139]
  wire  _T_110 = waddr_intpriority_base_match & _T_109; // @[pic_ctrl.scala 141:106]
  wire  intpriority_reg_we_25 = _T_110 & picm_wren_ff; // @[pic_ctrl.scala 141:153]
  wire  _T_112 = picm_waddr_ff[6:2] == 5'h1a; // @[pic_ctrl.scala 141:139]
  wire  _T_113 = waddr_intpriority_base_match & _T_112; // @[pic_ctrl.scala 141:106]
  wire  intpriority_reg_we_26 = _T_113 & picm_wren_ff; // @[pic_ctrl.scala 141:153]
  wire  _T_115 = picm_waddr_ff[6:2] == 5'h1b; // @[pic_ctrl.scala 141:139]
  wire  _T_116 = waddr_intpriority_base_match & _T_115; // @[pic_ctrl.scala 141:106]
  wire  intpriority_reg_we_27 = _T_116 & picm_wren_ff; // @[pic_ctrl.scala 141:153]
  wire  _T_118 = picm_waddr_ff[6:2] == 5'h1c; // @[pic_ctrl.scala 141:139]
  wire  _T_119 = waddr_intpriority_base_match & _T_118; // @[pic_ctrl.scala 141:106]
  wire  intpriority_reg_we_28 = _T_119 & picm_wren_ff; // @[pic_ctrl.scala 141:153]
  wire  _T_121 = picm_waddr_ff[6:2] == 5'h1d; // @[pic_ctrl.scala 141:139]
  wire  _T_122 = waddr_intpriority_base_match & _T_121; // @[pic_ctrl.scala 141:106]
  wire  intpriority_reg_we_29 = _T_122 & picm_wren_ff; // @[pic_ctrl.scala 141:153]
  wire  _T_124 = picm_waddr_ff[6:2] == 5'h1e; // @[pic_ctrl.scala 141:139]
  wire  _T_125 = waddr_intpriority_base_match & _T_124; // @[pic_ctrl.scala 141:106]
  wire  intpriority_reg_we_30 = _T_125 & picm_wren_ff; // @[pic_ctrl.scala 141:153]
  wire  _T_127 = picm_waddr_ff[6:2] == 5'h1f; // @[pic_ctrl.scala 141:139]
  wire  _T_128 = waddr_intpriority_base_match & _T_127; // @[pic_ctrl.scala 141:106]
  wire  intpriority_reg_we_31 = _T_128 & picm_wren_ff; // @[pic_ctrl.scala 141:153]
  wire  _T_130 = picm_raddr_ff[6:2] == 5'h1; // @[pic_ctrl.scala 142:139]
  wire  _T_131 = raddr_intpriority_base_match & _T_130; // @[pic_ctrl.scala 142:106]
  wire  intpriority_reg_re_1 = _T_131 & picm_rden_ff; // @[pic_ctrl.scala 142:153]
  wire  _T_133 = picm_raddr_ff[6:2] == 5'h2; // @[pic_ctrl.scala 142:139]
  wire  _T_134 = raddr_intpriority_base_match & _T_133; // @[pic_ctrl.scala 142:106]
  wire  intpriority_reg_re_2 = _T_134 & picm_rden_ff; // @[pic_ctrl.scala 142:153]
  wire  _T_136 = picm_raddr_ff[6:2] == 5'h3; // @[pic_ctrl.scala 142:139]
  wire  _T_137 = raddr_intpriority_base_match & _T_136; // @[pic_ctrl.scala 142:106]
  wire  intpriority_reg_re_3 = _T_137 & picm_rden_ff; // @[pic_ctrl.scala 142:153]
  wire  _T_139 = picm_raddr_ff[6:2] == 5'h4; // @[pic_ctrl.scala 142:139]
  wire  _T_140 = raddr_intpriority_base_match & _T_139; // @[pic_ctrl.scala 142:106]
  wire  intpriority_reg_re_4 = _T_140 & picm_rden_ff; // @[pic_ctrl.scala 142:153]
  wire  _T_142 = picm_raddr_ff[6:2] == 5'h5; // @[pic_ctrl.scala 142:139]
  wire  _T_143 = raddr_intpriority_base_match & _T_142; // @[pic_ctrl.scala 142:106]
  wire  intpriority_reg_re_5 = _T_143 & picm_rden_ff; // @[pic_ctrl.scala 142:153]
  wire  _T_145 = picm_raddr_ff[6:2] == 5'h6; // @[pic_ctrl.scala 142:139]
  wire  _T_146 = raddr_intpriority_base_match & _T_145; // @[pic_ctrl.scala 142:106]
  wire  intpriority_reg_re_6 = _T_146 & picm_rden_ff; // @[pic_ctrl.scala 142:153]
  wire  _T_148 = picm_raddr_ff[6:2] == 5'h7; // @[pic_ctrl.scala 142:139]
  wire  _T_149 = raddr_intpriority_base_match & _T_148; // @[pic_ctrl.scala 142:106]
  wire  intpriority_reg_re_7 = _T_149 & picm_rden_ff; // @[pic_ctrl.scala 142:153]
  wire  _T_151 = picm_raddr_ff[6:2] == 5'h8; // @[pic_ctrl.scala 142:139]
  wire  _T_152 = raddr_intpriority_base_match & _T_151; // @[pic_ctrl.scala 142:106]
  wire  intpriority_reg_re_8 = _T_152 & picm_rden_ff; // @[pic_ctrl.scala 142:153]
  wire  _T_154 = picm_raddr_ff[6:2] == 5'h9; // @[pic_ctrl.scala 142:139]
  wire  _T_155 = raddr_intpriority_base_match & _T_154; // @[pic_ctrl.scala 142:106]
  wire  intpriority_reg_re_9 = _T_155 & picm_rden_ff; // @[pic_ctrl.scala 142:153]
  wire  _T_157 = picm_raddr_ff[6:2] == 5'ha; // @[pic_ctrl.scala 142:139]
  wire  _T_158 = raddr_intpriority_base_match & _T_157; // @[pic_ctrl.scala 142:106]
  wire  intpriority_reg_re_10 = _T_158 & picm_rden_ff; // @[pic_ctrl.scala 142:153]
  wire  _T_160 = picm_raddr_ff[6:2] == 5'hb; // @[pic_ctrl.scala 142:139]
  wire  _T_161 = raddr_intpriority_base_match & _T_160; // @[pic_ctrl.scala 142:106]
  wire  intpriority_reg_re_11 = _T_161 & picm_rden_ff; // @[pic_ctrl.scala 142:153]
  wire  _T_163 = picm_raddr_ff[6:2] == 5'hc; // @[pic_ctrl.scala 142:139]
  wire  _T_164 = raddr_intpriority_base_match & _T_163; // @[pic_ctrl.scala 142:106]
  wire  intpriority_reg_re_12 = _T_164 & picm_rden_ff; // @[pic_ctrl.scala 142:153]
  wire  _T_166 = picm_raddr_ff[6:2] == 5'hd; // @[pic_ctrl.scala 142:139]
  wire  _T_167 = raddr_intpriority_base_match & _T_166; // @[pic_ctrl.scala 142:106]
  wire  intpriority_reg_re_13 = _T_167 & picm_rden_ff; // @[pic_ctrl.scala 142:153]
  wire  _T_169 = picm_raddr_ff[6:2] == 5'he; // @[pic_ctrl.scala 142:139]
  wire  _T_170 = raddr_intpriority_base_match & _T_169; // @[pic_ctrl.scala 142:106]
  wire  intpriority_reg_re_14 = _T_170 & picm_rden_ff; // @[pic_ctrl.scala 142:153]
  wire  _T_172 = picm_raddr_ff[6:2] == 5'hf; // @[pic_ctrl.scala 142:139]
  wire  _T_173 = raddr_intpriority_base_match & _T_172; // @[pic_ctrl.scala 142:106]
  wire  intpriority_reg_re_15 = _T_173 & picm_rden_ff; // @[pic_ctrl.scala 142:153]
  wire  _T_175 = picm_raddr_ff[6:2] == 5'h10; // @[pic_ctrl.scala 142:139]
  wire  _T_176 = raddr_intpriority_base_match & _T_175; // @[pic_ctrl.scala 142:106]
  wire  intpriority_reg_re_16 = _T_176 & picm_rden_ff; // @[pic_ctrl.scala 142:153]
  wire  _T_178 = picm_raddr_ff[6:2] == 5'h11; // @[pic_ctrl.scala 142:139]
  wire  _T_179 = raddr_intpriority_base_match & _T_178; // @[pic_ctrl.scala 142:106]
  wire  intpriority_reg_re_17 = _T_179 & picm_rden_ff; // @[pic_ctrl.scala 142:153]
  wire  _T_181 = picm_raddr_ff[6:2] == 5'h12; // @[pic_ctrl.scala 142:139]
  wire  _T_182 = raddr_intpriority_base_match & _T_181; // @[pic_ctrl.scala 142:106]
  wire  intpriority_reg_re_18 = _T_182 & picm_rden_ff; // @[pic_ctrl.scala 142:153]
  wire  _T_184 = picm_raddr_ff[6:2] == 5'h13; // @[pic_ctrl.scala 142:139]
  wire  _T_185 = raddr_intpriority_base_match & _T_184; // @[pic_ctrl.scala 142:106]
  wire  intpriority_reg_re_19 = _T_185 & picm_rden_ff; // @[pic_ctrl.scala 142:153]
  wire  _T_187 = picm_raddr_ff[6:2] == 5'h14; // @[pic_ctrl.scala 142:139]
  wire  _T_188 = raddr_intpriority_base_match & _T_187; // @[pic_ctrl.scala 142:106]
  wire  intpriority_reg_re_20 = _T_188 & picm_rden_ff; // @[pic_ctrl.scala 142:153]
  wire  _T_190 = picm_raddr_ff[6:2] == 5'h15; // @[pic_ctrl.scala 142:139]
  wire  _T_191 = raddr_intpriority_base_match & _T_190; // @[pic_ctrl.scala 142:106]
  wire  intpriority_reg_re_21 = _T_191 & picm_rden_ff; // @[pic_ctrl.scala 142:153]
  wire  _T_193 = picm_raddr_ff[6:2] == 5'h16; // @[pic_ctrl.scala 142:139]
  wire  _T_194 = raddr_intpriority_base_match & _T_193; // @[pic_ctrl.scala 142:106]
  wire  intpriority_reg_re_22 = _T_194 & picm_rden_ff; // @[pic_ctrl.scala 142:153]
  wire  _T_196 = picm_raddr_ff[6:2] == 5'h17; // @[pic_ctrl.scala 142:139]
  wire  _T_197 = raddr_intpriority_base_match & _T_196; // @[pic_ctrl.scala 142:106]
  wire  intpriority_reg_re_23 = _T_197 & picm_rden_ff; // @[pic_ctrl.scala 142:153]
  wire  _T_199 = picm_raddr_ff[6:2] == 5'h18; // @[pic_ctrl.scala 142:139]
  wire  _T_200 = raddr_intpriority_base_match & _T_199; // @[pic_ctrl.scala 142:106]
  wire  intpriority_reg_re_24 = _T_200 & picm_rden_ff; // @[pic_ctrl.scala 142:153]
  wire  _T_202 = picm_raddr_ff[6:2] == 5'h19; // @[pic_ctrl.scala 142:139]
  wire  _T_203 = raddr_intpriority_base_match & _T_202; // @[pic_ctrl.scala 142:106]
  wire  intpriority_reg_re_25 = _T_203 & picm_rden_ff; // @[pic_ctrl.scala 142:153]
  wire  _T_205 = picm_raddr_ff[6:2] == 5'h1a; // @[pic_ctrl.scala 142:139]
  wire  _T_206 = raddr_intpriority_base_match & _T_205; // @[pic_ctrl.scala 142:106]
  wire  intpriority_reg_re_26 = _T_206 & picm_rden_ff; // @[pic_ctrl.scala 142:153]
  wire  _T_208 = picm_raddr_ff[6:2] == 5'h1b; // @[pic_ctrl.scala 142:139]
  wire  _T_209 = raddr_intpriority_base_match & _T_208; // @[pic_ctrl.scala 142:106]
  wire  intpriority_reg_re_27 = _T_209 & picm_rden_ff; // @[pic_ctrl.scala 142:153]
  wire  _T_211 = picm_raddr_ff[6:2] == 5'h1c; // @[pic_ctrl.scala 142:139]
  wire  _T_212 = raddr_intpriority_base_match & _T_211; // @[pic_ctrl.scala 142:106]
  wire  intpriority_reg_re_28 = _T_212 & picm_rden_ff; // @[pic_ctrl.scala 142:153]
  wire  _T_214 = picm_raddr_ff[6:2] == 5'h1d; // @[pic_ctrl.scala 142:139]
  wire  _T_215 = raddr_intpriority_base_match & _T_214; // @[pic_ctrl.scala 142:106]
  wire  intpriority_reg_re_29 = _T_215 & picm_rden_ff; // @[pic_ctrl.scala 142:153]
  wire  _T_217 = picm_raddr_ff[6:2] == 5'h1e; // @[pic_ctrl.scala 142:139]
  wire  _T_218 = raddr_intpriority_base_match & _T_217; // @[pic_ctrl.scala 142:106]
  wire  intpriority_reg_re_30 = _T_218 & picm_rden_ff; // @[pic_ctrl.scala 142:153]
  wire  _T_220 = picm_raddr_ff[6:2] == 5'h1f; // @[pic_ctrl.scala 142:139]
  wire  _T_221 = raddr_intpriority_base_match & _T_220; // @[pic_ctrl.scala 142:106]
  wire  intpriority_reg_re_31 = _T_221 & picm_rden_ff; // @[pic_ctrl.scala 142:153]
  wire  _T_224 = waddr_intenable_base_match & _T_37; // @[pic_ctrl.scala 143:106]
  wire  intenable_reg_we_1 = _T_224 & picm_wren_ff; // @[pic_ctrl.scala 143:153]
  wire  _T_227 = waddr_intenable_base_match & _T_40; // @[pic_ctrl.scala 143:106]
  wire  intenable_reg_we_2 = _T_227 & picm_wren_ff; // @[pic_ctrl.scala 143:153]
  wire  _T_230 = waddr_intenable_base_match & _T_43; // @[pic_ctrl.scala 143:106]
  wire  intenable_reg_we_3 = _T_230 & picm_wren_ff; // @[pic_ctrl.scala 143:153]
  wire  _T_233 = waddr_intenable_base_match & _T_46; // @[pic_ctrl.scala 143:106]
  wire  intenable_reg_we_4 = _T_233 & picm_wren_ff; // @[pic_ctrl.scala 143:153]
  wire  _T_236 = waddr_intenable_base_match & _T_49; // @[pic_ctrl.scala 143:106]
  wire  intenable_reg_we_5 = _T_236 & picm_wren_ff; // @[pic_ctrl.scala 143:153]
  wire  _T_239 = waddr_intenable_base_match & _T_52; // @[pic_ctrl.scala 143:106]
  wire  intenable_reg_we_6 = _T_239 & picm_wren_ff; // @[pic_ctrl.scala 143:153]
  wire  _T_242 = waddr_intenable_base_match & _T_55; // @[pic_ctrl.scala 143:106]
  wire  intenable_reg_we_7 = _T_242 & picm_wren_ff; // @[pic_ctrl.scala 143:153]
  wire  _T_245 = waddr_intenable_base_match & _T_58; // @[pic_ctrl.scala 143:106]
  wire  intenable_reg_we_8 = _T_245 & picm_wren_ff; // @[pic_ctrl.scala 143:153]
  wire  _T_248 = waddr_intenable_base_match & _T_61; // @[pic_ctrl.scala 143:106]
  wire  intenable_reg_we_9 = _T_248 & picm_wren_ff; // @[pic_ctrl.scala 143:153]
  wire  _T_251 = waddr_intenable_base_match & _T_64; // @[pic_ctrl.scala 143:106]
  wire  intenable_reg_we_10 = _T_251 & picm_wren_ff; // @[pic_ctrl.scala 143:153]
  wire  _T_254 = waddr_intenable_base_match & _T_67; // @[pic_ctrl.scala 143:106]
  wire  intenable_reg_we_11 = _T_254 & picm_wren_ff; // @[pic_ctrl.scala 143:153]
  wire  _T_257 = waddr_intenable_base_match & _T_70; // @[pic_ctrl.scala 143:106]
  wire  intenable_reg_we_12 = _T_257 & picm_wren_ff; // @[pic_ctrl.scala 143:153]
  wire  _T_260 = waddr_intenable_base_match & _T_73; // @[pic_ctrl.scala 143:106]
  wire  intenable_reg_we_13 = _T_260 & picm_wren_ff; // @[pic_ctrl.scala 143:153]
  wire  _T_263 = waddr_intenable_base_match & _T_76; // @[pic_ctrl.scala 143:106]
  wire  intenable_reg_we_14 = _T_263 & picm_wren_ff; // @[pic_ctrl.scala 143:153]
  wire  _T_266 = waddr_intenable_base_match & _T_79; // @[pic_ctrl.scala 143:106]
  wire  intenable_reg_we_15 = _T_266 & picm_wren_ff; // @[pic_ctrl.scala 143:153]
  wire  _T_269 = waddr_intenable_base_match & _T_82; // @[pic_ctrl.scala 143:106]
  wire  intenable_reg_we_16 = _T_269 & picm_wren_ff; // @[pic_ctrl.scala 143:153]
  wire  _T_272 = waddr_intenable_base_match & _T_85; // @[pic_ctrl.scala 143:106]
  wire  intenable_reg_we_17 = _T_272 & picm_wren_ff; // @[pic_ctrl.scala 143:153]
  wire  _T_275 = waddr_intenable_base_match & _T_88; // @[pic_ctrl.scala 143:106]
  wire  intenable_reg_we_18 = _T_275 & picm_wren_ff; // @[pic_ctrl.scala 143:153]
  wire  _T_278 = waddr_intenable_base_match & _T_91; // @[pic_ctrl.scala 143:106]
  wire  intenable_reg_we_19 = _T_278 & picm_wren_ff; // @[pic_ctrl.scala 143:153]
  wire  _T_281 = waddr_intenable_base_match & _T_94; // @[pic_ctrl.scala 143:106]
  wire  intenable_reg_we_20 = _T_281 & picm_wren_ff; // @[pic_ctrl.scala 143:153]
  wire  _T_284 = waddr_intenable_base_match & _T_97; // @[pic_ctrl.scala 143:106]
  wire  intenable_reg_we_21 = _T_284 & picm_wren_ff; // @[pic_ctrl.scala 143:153]
  wire  _T_287 = waddr_intenable_base_match & _T_100; // @[pic_ctrl.scala 143:106]
  wire  intenable_reg_we_22 = _T_287 & picm_wren_ff; // @[pic_ctrl.scala 143:153]
  wire  _T_290 = waddr_intenable_base_match & _T_103; // @[pic_ctrl.scala 143:106]
  wire  intenable_reg_we_23 = _T_290 & picm_wren_ff; // @[pic_ctrl.scala 143:153]
  wire  _T_293 = waddr_intenable_base_match & _T_106; // @[pic_ctrl.scala 143:106]
  wire  intenable_reg_we_24 = _T_293 & picm_wren_ff; // @[pic_ctrl.scala 143:153]
  wire  _T_296 = waddr_intenable_base_match & _T_109; // @[pic_ctrl.scala 143:106]
  wire  intenable_reg_we_25 = _T_296 & picm_wren_ff; // @[pic_ctrl.scala 143:153]
  wire  _T_299 = waddr_intenable_base_match & _T_112; // @[pic_ctrl.scala 143:106]
  wire  intenable_reg_we_26 = _T_299 & picm_wren_ff; // @[pic_ctrl.scala 143:153]
  wire  _T_302 = waddr_intenable_base_match & _T_115; // @[pic_ctrl.scala 143:106]
  wire  intenable_reg_we_27 = _T_302 & picm_wren_ff; // @[pic_ctrl.scala 143:153]
  wire  _T_305 = waddr_intenable_base_match & _T_118; // @[pic_ctrl.scala 143:106]
  wire  intenable_reg_we_28 = _T_305 & picm_wren_ff; // @[pic_ctrl.scala 143:153]
  wire  _T_308 = waddr_intenable_base_match & _T_121; // @[pic_ctrl.scala 143:106]
  wire  intenable_reg_we_29 = _T_308 & picm_wren_ff; // @[pic_ctrl.scala 143:153]
  wire  _T_311 = waddr_intenable_base_match & _T_124; // @[pic_ctrl.scala 143:106]
  wire  intenable_reg_we_30 = _T_311 & picm_wren_ff; // @[pic_ctrl.scala 143:153]
  wire  _T_314 = waddr_intenable_base_match & _T_127; // @[pic_ctrl.scala 143:106]
  wire  intenable_reg_we_31 = _T_314 & picm_wren_ff; // @[pic_ctrl.scala 143:153]
  wire  _T_317 = raddr_intenable_base_match & _T_130; // @[pic_ctrl.scala 144:106]
  wire  intenable_reg_re_1 = _T_317 & picm_rden_ff; // @[pic_ctrl.scala 144:153]
  wire  _T_320 = raddr_intenable_base_match & _T_133; // @[pic_ctrl.scala 144:106]
  wire  intenable_reg_re_2 = _T_320 & picm_rden_ff; // @[pic_ctrl.scala 144:153]
  wire  _T_323 = raddr_intenable_base_match & _T_136; // @[pic_ctrl.scala 144:106]
  wire  intenable_reg_re_3 = _T_323 & picm_rden_ff; // @[pic_ctrl.scala 144:153]
  wire  _T_326 = raddr_intenable_base_match & _T_139; // @[pic_ctrl.scala 144:106]
  wire  intenable_reg_re_4 = _T_326 & picm_rden_ff; // @[pic_ctrl.scala 144:153]
  wire  _T_329 = raddr_intenable_base_match & _T_142; // @[pic_ctrl.scala 144:106]
  wire  intenable_reg_re_5 = _T_329 & picm_rden_ff; // @[pic_ctrl.scala 144:153]
  wire  _T_332 = raddr_intenable_base_match & _T_145; // @[pic_ctrl.scala 144:106]
  wire  intenable_reg_re_6 = _T_332 & picm_rden_ff; // @[pic_ctrl.scala 144:153]
  wire  _T_335 = raddr_intenable_base_match & _T_148; // @[pic_ctrl.scala 144:106]
  wire  intenable_reg_re_7 = _T_335 & picm_rden_ff; // @[pic_ctrl.scala 144:153]
  wire  _T_338 = raddr_intenable_base_match & _T_151; // @[pic_ctrl.scala 144:106]
  wire  intenable_reg_re_8 = _T_338 & picm_rden_ff; // @[pic_ctrl.scala 144:153]
  wire  _T_341 = raddr_intenable_base_match & _T_154; // @[pic_ctrl.scala 144:106]
  wire  intenable_reg_re_9 = _T_341 & picm_rden_ff; // @[pic_ctrl.scala 144:153]
  wire  _T_344 = raddr_intenable_base_match & _T_157; // @[pic_ctrl.scala 144:106]
  wire  intenable_reg_re_10 = _T_344 & picm_rden_ff; // @[pic_ctrl.scala 144:153]
  wire  _T_347 = raddr_intenable_base_match & _T_160; // @[pic_ctrl.scala 144:106]
  wire  intenable_reg_re_11 = _T_347 & picm_rden_ff; // @[pic_ctrl.scala 144:153]
  wire  _T_350 = raddr_intenable_base_match & _T_163; // @[pic_ctrl.scala 144:106]
  wire  intenable_reg_re_12 = _T_350 & picm_rden_ff; // @[pic_ctrl.scala 144:153]
  wire  _T_353 = raddr_intenable_base_match & _T_166; // @[pic_ctrl.scala 144:106]
  wire  intenable_reg_re_13 = _T_353 & picm_rden_ff; // @[pic_ctrl.scala 144:153]
  wire  _T_356 = raddr_intenable_base_match & _T_169; // @[pic_ctrl.scala 144:106]
  wire  intenable_reg_re_14 = _T_356 & picm_rden_ff; // @[pic_ctrl.scala 144:153]
  wire  _T_359 = raddr_intenable_base_match & _T_172; // @[pic_ctrl.scala 144:106]
  wire  intenable_reg_re_15 = _T_359 & picm_rden_ff; // @[pic_ctrl.scala 144:153]
  wire  _T_362 = raddr_intenable_base_match & _T_175; // @[pic_ctrl.scala 144:106]
  wire  intenable_reg_re_16 = _T_362 & picm_rden_ff; // @[pic_ctrl.scala 144:153]
  wire  _T_365 = raddr_intenable_base_match & _T_178; // @[pic_ctrl.scala 144:106]
  wire  intenable_reg_re_17 = _T_365 & picm_rden_ff; // @[pic_ctrl.scala 144:153]
  wire  _T_368 = raddr_intenable_base_match & _T_181; // @[pic_ctrl.scala 144:106]
  wire  intenable_reg_re_18 = _T_368 & picm_rden_ff; // @[pic_ctrl.scala 144:153]
  wire  _T_371 = raddr_intenable_base_match & _T_184; // @[pic_ctrl.scala 144:106]
  wire  intenable_reg_re_19 = _T_371 & picm_rden_ff; // @[pic_ctrl.scala 144:153]
  wire  _T_374 = raddr_intenable_base_match & _T_187; // @[pic_ctrl.scala 144:106]
  wire  intenable_reg_re_20 = _T_374 & picm_rden_ff; // @[pic_ctrl.scala 144:153]
  wire  _T_377 = raddr_intenable_base_match & _T_190; // @[pic_ctrl.scala 144:106]
  wire  intenable_reg_re_21 = _T_377 & picm_rden_ff; // @[pic_ctrl.scala 144:153]
  wire  _T_380 = raddr_intenable_base_match & _T_193; // @[pic_ctrl.scala 144:106]
  wire  intenable_reg_re_22 = _T_380 & picm_rden_ff; // @[pic_ctrl.scala 144:153]
  wire  _T_383 = raddr_intenable_base_match & _T_196; // @[pic_ctrl.scala 144:106]
  wire  intenable_reg_re_23 = _T_383 & picm_rden_ff; // @[pic_ctrl.scala 144:153]
  wire  _T_386 = raddr_intenable_base_match & _T_199; // @[pic_ctrl.scala 144:106]
  wire  intenable_reg_re_24 = _T_386 & picm_rden_ff; // @[pic_ctrl.scala 144:153]
  wire  _T_389 = raddr_intenable_base_match & _T_202; // @[pic_ctrl.scala 144:106]
  wire  intenable_reg_re_25 = _T_389 & picm_rden_ff; // @[pic_ctrl.scala 144:153]
  wire  _T_392 = raddr_intenable_base_match & _T_205; // @[pic_ctrl.scala 144:106]
  wire  intenable_reg_re_26 = _T_392 & picm_rden_ff; // @[pic_ctrl.scala 144:153]
  wire  _T_395 = raddr_intenable_base_match & _T_208; // @[pic_ctrl.scala 144:106]
  wire  intenable_reg_re_27 = _T_395 & picm_rden_ff; // @[pic_ctrl.scala 144:153]
  wire  _T_398 = raddr_intenable_base_match & _T_211; // @[pic_ctrl.scala 144:106]
  wire  intenable_reg_re_28 = _T_398 & picm_rden_ff; // @[pic_ctrl.scala 144:153]
  wire  _T_401 = raddr_intenable_base_match & _T_214; // @[pic_ctrl.scala 144:106]
  wire  intenable_reg_re_29 = _T_401 & picm_rden_ff; // @[pic_ctrl.scala 144:153]
  wire  _T_404 = raddr_intenable_base_match & _T_217; // @[pic_ctrl.scala 144:106]
  wire  intenable_reg_re_30 = _T_404 & picm_rden_ff; // @[pic_ctrl.scala 144:153]
  wire  _T_407 = raddr_intenable_base_match & _T_220; // @[pic_ctrl.scala 144:106]
  wire  intenable_reg_re_31 = _T_407 & picm_rden_ff; // @[pic_ctrl.scala 144:153]
  wire  _T_410 = waddr_config_gw_base_match & _T_37; // @[pic_ctrl.scala 145:106]
  wire  gw_config_reg_we_1 = _T_410 & picm_wren_ff; // @[pic_ctrl.scala 145:153]
  wire  _T_413 = waddr_config_gw_base_match & _T_40; // @[pic_ctrl.scala 145:106]
  wire  gw_config_reg_we_2 = _T_413 & picm_wren_ff; // @[pic_ctrl.scala 145:153]
  wire  _T_416 = waddr_config_gw_base_match & _T_43; // @[pic_ctrl.scala 145:106]
  wire  gw_config_reg_we_3 = _T_416 & picm_wren_ff; // @[pic_ctrl.scala 145:153]
  wire  _T_419 = waddr_config_gw_base_match & _T_46; // @[pic_ctrl.scala 145:106]
  wire  gw_config_reg_we_4 = _T_419 & picm_wren_ff; // @[pic_ctrl.scala 145:153]
  wire  _T_422 = waddr_config_gw_base_match & _T_49; // @[pic_ctrl.scala 145:106]
  wire  gw_config_reg_we_5 = _T_422 & picm_wren_ff; // @[pic_ctrl.scala 145:153]
  wire  _T_425 = waddr_config_gw_base_match & _T_52; // @[pic_ctrl.scala 145:106]
  wire  gw_config_reg_we_6 = _T_425 & picm_wren_ff; // @[pic_ctrl.scala 145:153]
  wire  _T_428 = waddr_config_gw_base_match & _T_55; // @[pic_ctrl.scala 145:106]
  wire  gw_config_reg_we_7 = _T_428 & picm_wren_ff; // @[pic_ctrl.scala 145:153]
  wire  _T_431 = waddr_config_gw_base_match & _T_58; // @[pic_ctrl.scala 145:106]
  wire  gw_config_reg_we_8 = _T_431 & picm_wren_ff; // @[pic_ctrl.scala 145:153]
  wire  _T_434 = waddr_config_gw_base_match & _T_61; // @[pic_ctrl.scala 145:106]
  wire  gw_config_reg_we_9 = _T_434 & picm_wren_ff; // @[pic_ctrl.scala 145:153]
  wire  _T_437 = waddr_config_gw_base_match & _T_64; // @[pic_ctrl.scala 145:106]
  wire  gw_config_reg_we_10 = _T_437 & picm_wren_ff; // @[pic_ctrl.scala 145:153]
  wire  _T_440 = waddr_config_gw_base_match & _T_67; // @[pic_ctrl.scala 145:106]
  wire  gw_config_reg_we_11 = _T_440 & picm_wren_ff; // @[pic_ctrl.scala 145:153]
  wire  _T_443 = waddr_config_gw_base_match & _T_70; // @[pic_ctrl.scala 145:106]
  wire  gw_config_reg_we_12 = _T_443 & picm_wren_ff; // @[pic_ctrl.scala 145:153]
  wire  _T_446 = waddr_config_gw_base_match & _T_73; // @[pic_ctrl.scala 145:106]
  wire  gw_config_reg_we_13 = _T_446 & picm_wren_ff; // @[pic_ctrl.scala 145:153]
  wire  _T_449 = waddr_config_gw_base_match & _T_76; // @[pic_ctrl.scala 145:106]
  wire  gw_config_reg_we_14 = _T_449 & picm_wren_ff; // @[pic_ctrl.scala 145:153]
  wire  _T_452 = waddr_config_gw_base_match & _T_79; // @[pic_ctrl.scala 145:106]
  wire  gw_config_reg_we_15 = _T_452 & picm_wren_ff; // @[pic_ctrl.scala 145:153]
  wire  _T_455 = waddr_config_gw_base_match & _T_82; // @[pic_ctrl.scala 145:106]
  wire  gw_config_reg_we_16 = _T_455 & picm_wren_ff; // @[pic_ctrl.scala 145:153]
  wire  _T_458 = waddr_config_gw_base_match & _T_85; // @[pic_ctrl.scala 145:106]
  wire  gw_config_reg_we_17 = _T_458 & picm_wren_ff; // @[pic_ctrl.scala 145:153]
  wire  _T_461 = waddr_config_gw_base_match & _T_88; // @[pic_ctrl.scala 145:106]
  wire  gw_config_reg_we_18 = _T_461 & picm_wren_ff; // @[pic_ctrl.scala 145:153]
  wire  _T_464 = waddr_config_gw_base_match & _T_91; // @[pic_ctrl.scala 145:106]
  wire  gw_config_reg_we_19 = _T_464 & picm_wren_ff; // @[pic_ctrl.scala 145:153]
  wire  _T_467 = waddr_config_gw_base_match & _T_94; // @[pic_ctrl.scala 145:106]
  wire  gw_config_reg_we_20 = _T_467 & picm_wren_ff; // @[pic_ctrl.scala 145:153]
  wire  _T_470 = waddr_config_gw_base_match & _T_97; // @[pic_ctrl.scala 145:106]
  wire  gw_config_reg_we_21 = _T_470 & picm_wren_ff; // @[pic_ctrl.scala 145:153]
  wire  _T_473 = waddr_config_gw_base_match & _T_100; // @[pic_ctrl.scala 145:106]
  wire  gw_config_reg_we_22 = _T_473 & picm_wren_ff; // @[pic_ctrl.scala 145:153]
  wire  _T_476 = waddr_config_gw_base_match & _T_103; // @[pic_ctrl.scala 145:106]
  wire  gw_config_reg_we_23 = _T_476 & picm_wren_ff; // @[pic_ctrl.scala 145:153]
  wire  _T_479 = waddr_config_gw_base_match & _T_106; // @[pic_ctrl.scala 145:106]
  wire  gw_config_reg_we_24 = _T_479 & picm_wren_ff; // @[pic_ctrl.scala 145:153]
  wire  _T_482 = waddr_config_gw_base_match & _T_109; // @[pic_ctrl.scala 145:106]
  wire  gw_config_reg_we_25 = _T_482 & picm_wren_ff; // @[pic_ctrl.scala 145:153]
  wire  _T_485 = waddr_config_gw_base_match & _T_112; // @[pic_ctrl.scala 145:106]
  wire  gw_config_reg_we_26 = _T_485 & picm_wren_ff; // @[pic_ctrl.scala 145:153]
  wire  _T_488 = waddr_config_gw_base_match & _T_115; // @[pic_ctrl.scala 145:106]
  wire  gw_config_reg_we_27 = _T_488 & picm_wren_ff; // @[pic_ctrl.scala 145:153]
  wire  _T_491 = waddr_config_gw_base_match & _T_118; // @[pic_ctrl.scala 145:106]
  wire  gw_config_reg_we_28 = _T_491 & picm_wren_ff; // @[pic_ctrl.scala 145:153]
  wire  _T_494 = waddr_config_gw_base_match & _T_121; // @[pic_ctrl.scala 145:106]
  wire  gw_config_reg_we_29 = _T_494 & picm_wren_ff; // @[pic_ctrl.scala 145:153]
  wire  _T_497 = waddr_config_gw_base_match & _T_124; // @[pic_ctrl.scala 145:106]
  wire  gw_config_reg_we_30 = _T_497 & picm_wren_ff; // @[pic_ctrl.scala 145:153]
  wire  _T_500 = waddr_config_gw_base_match & _T_127; // @[pic_ctrl.scala 145:106]
  wire  gw_config_reg_we_31 = _T_500 & picm_wren_ff; // @[pic_ctrl.scala 145:153]
  wire  _T_503 = raddr_config_gw_base_match & _T_130; // @[pic_ctrl.scala 146:106]
  wire  gw_config_reg_re_1 = _T_503 & picm_rden_ff; // @[pic_ctrl.scala 146:153]
  wire  _T_506 = raddr_config_gw_base_match & _T_133; // @[pic_ctrl.scala 146:106]
  wire  gw_config_reg_re_2 = _T_506 & picm_rden_ff; // @[pic_ctrl.scala 146:153]
  wire  _T_509 = raddr_config_gw_base_match & _T_136; // @[pic_ctrl.scala 146:106]
  wire  gw_config_reg_re_3 = _T_509 & picm_rden_ff; // @[pic_ctrl.scala 146:153]
  wire  _T_512 = raddr_config_gw_base_match & _T_139; // @[pic_ctrl.scala 146:106]
  wire  gw_config_reg_re_4 = _T_512 & picm_rden_ff; // @[pic_ctrl.scala 146:153]
  wire  _T_515 = raddr_config_gw_base_match & _T_142; // @[pic_ctrl.scala 146:106]
  wire  gw_config_reg_re_5 = _T_515 & picm_rden_ff; // @[pic_ctrl.scala 146:153]
  wire  _T_518 = raddr_config_gw_base_match & _T_145; // @[pic_ctrl.scala 146:106]
  wire  gw_config_reg_re_6 = _T_518 & picm_rden_ff; // @[pic_ctrl.scala 146:153]
  wire  _T_521 = raddr_config_gw_base_match & _T_148; // @[pic_ctrl.scala 146:106]
  wire  gw_config_reg_re_7 = _T_521 & picm_rden_ff; // @[pic_ctrl.scala 146:153]
  wire  _T_524 = raddr_config_gw_base_match & _T_151; // @[pic_ctrl.scala 146:106]
  wire  gw_config_reg_re_8 = _T_524 & picm_rden_ff; // @[pic_ctrl.scala 146:153]
  wire  _T_527 = raddr_config_gw_base_match & _T_154; // @[pic_ctrl.scala 146:106]
  wire  gw_config_reg_re_9 = _T_527 & picm_rden_ff; // @[pic_ctrl.scala 146:153]
  wire  _T_530 = raddr_config_gw_base_match & _T_157; // @[pic_ctrl.scala 146:106]
  wire  gw_config_reg_re_10 = _T_530 & picm_rden_ff; // @[pic_ctrl.scala 146:153]
  wire  _T_533 = raddr_config_gw_base_match & _T_160; // @[pic_ctrl.scala 146:106]
  wire  gw_config_reg_re_11 = _T_533 & picm_rden_ff; // @[pic_ctrl.scala 146:153]
  wire  _T_536 = raddr_config_gw_base_match & _T_163; // @[pic_ctrl.scala 146:106]
  wire  gw_config_reg_re_12 = _T_536 & picm_rden_ff; // @[pic_ctrl.scala 146:153]
  wire  _T_539 = raddr_config_gw_base_match & _T_166; // @[pic_ctrl.scala 146:106]
  wire  gw_config_reg_re_13 = _T_539 & picm_rden_ff; // @[pic_ctrl.scala 146:153]
  wire  _T_542 = raddr_config_gw_base_match & _T_169; // @[pic_ctrl.scala 146:106]
  wire  gw_config_reg_re_14 = _T_542 & picm_rden_ff; // @[pic_ctrl.scala 146:153]
  wire  _T_545 = raddr_config_gw_base_match & _T_172; // @[pic_ctrl.scala 146:106]
  wire  gw_config_reg_re_15 = _T_545 & picm_rden_ff; // @[pic_ctrl.scala 146:153]
  wire  _T_548 = raddr_config_gw_base_match & _T_175; // @[pic_ctrl.scala 146:106]
  wire  gw_config_reg_re_16 = _T_548 & picm_rden_ff; // @[pic_ctrl.scala 146:153]
  wire  _T_551 = raddr_config_gw_base_match & _T_178; // @[pic_ctrl.scala 146:106]
  wire  gw_config_reg_re_17 = _T_551 & picm_rden_ff; // @[pic_ctrl.scala 146:153]
  wire  _T_554 = raddr_config_gw_base_match & _T_181; // @[pic_ctrl.scala 146:106]
  wire  gw_config_reg_re_18 = _T_554 & picm_rden_ff; // @[pic_ctrl.scala 146:153]
  wire  _T_557 = raddr_config_gw_base_match & _T_184; // @[pic_ctrl.scala 146:106]
  wire  gw_config_reg_re_19 = _T_557 & picm_rden_ff; // @[pic_ctrl.scala 146:153]
  wire  _T_560 = raddr_config_gw_base_match & _T_187; // @[pic_ctrl.scala 146:106]
  wire  gw_config_reg_re_20 = _T_560 & picm_rden_ff; // @[pic_ctrl.scala 146:153]
  wire  _T_563 = raddr_config_gw_base_match & _T_190; // @[pic_ctrl.scala 146:106]
  wire  gw_config_reg_re_21 = _T_563 & picm_rden_ff; // @[pic_ctrl.scala 146:153]
  wire  _T_566 = raddr_config_gw_base_match & _T_193; // @[pic_ctrl.scala 146:106]
  wire  gw_config_reg_re_22 = _T_566 & picm_rden_ff; // @[pic_ctrl.scala 146:153]
  wire  _T_569 = raddr_config_gw_base_match & _T_196; // @[pic_ctrl.scala 146:106]
  wire  gw_config_reg_re_23 = _T_569 & picm_rden_ff; // @[pic_ctrl.scala 146:153]
  wire  _T_572 = raddr_config_gw_base_match & _T_199; // @[pic_ctrl.scala 146:106]
  wire  gw_config_reg_re_24 = _T_572 & picm_rden_ff; // @[pic_ctrl.scala 146:153]
  wire  _T_575 = raddr_config_gw_base_match & _T_202; // @[pic_ctrl.scala 146:106]
  wire  gw_config_reg_re_25 = _T_575 & picm_rden_ff; // @[pic_ctrl.scala 146:153]
  wire  _T_578 = raddr_config_gw_base_match & _T_205; // @[pic_ctrl.scala 146:106]
  wire  gw_config_reg_re_26 = _T_578 & picm_rden_ff; // @[pic_ctrl.scala 146:153]
  wire  _T_581 = raddr_config_gw_base_match & _T_208; // @[pic_ctrl.scala 146:106]
  wire  gw_config_reg_re_27 = _T_581 & picm_rden_ff; // @[pic_ctrl.scala 146:153]
  wire  _T_584 = raddr_config_gw_base_match & _T_211; // @[pic_ctrl.scala 146:106]
  wire  gw_config_reg_re_28 = _T_584 & picm_rden_ff; // @[pic_ctrl.scala 146:153]
  wire  _T_587 = raddr_config_gw_base_match & _T_214; // @[pic_ctrl.scala 146:106]
  wire  gw_config_reg_re_29 = _T_587 & picm_rden_ff; // @[pic_ctrl.scala 146:153]
  wire  _T_590 = raddr_config_gw_base_match & _T_217; // @[pic_ctrl.scala 146:106]
  wire  gw_config_reg_re_30 = _T_590 & picm_rden_ff; // @[pic_ctrl.scala 146:153]
  wire  _T_593 = raddr_config_gw_base_match & _T_220; // @[pic_ctrl.scala 146:106]
  wire  gw_config_reg_re_31 = _T_593 & picm_rden_ff; // @[pic_ctrl.scala 146:153]
  wire  _T_596 = addr_clear_gw_base_match & _T_37; // @[pic_ctrl.scala 147:106]
  wire  gw_clear_reg_we_1 = _T_596 & picm_wren_ff; // @[pic_ctrl.scala 147:153]
  wire  _T_599 = addr_clear_gw_base_match & _T_40; // @[pic_ctrl.scala 147:106]
  wire  gw_clear_reg_we_2 = _T_599 & picm_wren_ff; // @[pic_ctrl.scala 147:153]
  wire  _T_602 = addr_clear_gw_base_match & _T_43; // @[pic_ctrl.scala 147:106]
  wire  gw_clear_reg_we_3 = _T_602 & picm_wren_ff; // @[pic_ctrl.scala 147:153]
  wire  _T_605 = addr_clear_gw_base_match & _T_46; // @[pic_ctrl.scala 147:106]
  wire  gw_clear_reg_we_4 = _T_605 & picm_wren_ff; // @[pic_ctrl.scala 147:153]
  wire  _T_608 = addr_clear_gw_base_match & _T_49; // @[pic_ctrl.scala 147:106]
  wire  gw_clear_reg_we_5 = _T_608 & picm_wren_ff; // @[pic_ctrl.scala 147:153]
  wire  _T_611 = addr_clear_gw_base_match & _T_52; // @[pic_ctrl.scala 147:106]
  wire  gw_clear_reg_we_6 = _T_611 & picm_wren_ff; // @[pic_ctrl.scala 147:153]
  wire  _T_614 = addr_clear_gw_base_match & _T_55; // @[pic_ctrl.scala 147:106]
  wire  gw_clear_reg_we_7 = _T_614 & picm_wren_ff; // @[pic_ctrl.scala 147:153]
  wire  _T_617 = addr_clear_gw_base_match & _T_58; // @[pic_ctrl.scala 147:106]
  wire  gw_clear_reg_we_8 = _T_617 & picm_wren_ff; // @[pic_ctrl.scala 147:153]
  wire  _T_620 = addr_clear_gw_base_match & _T_61; // @[pic_ctrl.scala 147:106]
  wire  gw_clear_reg_we_9 = _T_620 & picm_wren_ff; // @[pic_ctrl.scala 147:153]
  wire  _T_623 = addr_clear_gw_base_match & _T_64; // @[pic_ctrl.scala 147:106]
  wire  gw_clear_reg_we_10 = _T_623 & picm_wren_ff; // @[pic_ctrl.scala 147:153]
  wire  _T_626 = addr_clear_gw_base_match & _T_67; // @[pic_ctrl.scala 147:106]
  wire  gw_clear_reg_we_11 = _T_626 & picm_wren_ff; // @[pic_ctrl.scala 147:153]
  wire  _T_629 = addr_clear_gw_base_match & _T_70; // @[pic_ctrl.scala 147:106]
  wire  gw_clear_reg_we_12 = _T_629 & picm_wren_ff; // @[pic_ctrl.scala 147:153]
  wire  _T_632 = addr_clear_gw_base_match & _T_73; // @[pic_ctrl.scala 147:106]
  wire  gw_clear_reg_we_13 = _T_632 & picm_wren_ff; // @[pic_ctrl.scala 147:153]
  wire  _T_635 = addr_clear_gw_base_match & _T_76; // @[pic_ctrl.scala 147:106]
  wire  gw_clear_reg_we_14 = _T_635 & picm_wren_ff; // @[pic_ctrl.scala 147:153]
  wire  _T_638 = addr_clear_gw_base_match & _T_79; // @[pic_ctrl.scala 147:106]
  wire  gw_clear_reg_we_15 = _T_638 & picm_wren_ff; // @[pic_ctrl.scala 147:153]
  wire  _T_641 = addr_clear_gw_base_match & _T_82; // @[pic_ctrl.scala 147:106]
  wire  gw_clear_reg_we_16 = _T_641 & picm_wren_ff; // @[pic_ctrl.scala 147:153]
  wire  _T_644 = addr_clear_gw_base_match & _T_85; // @[pic_ctrl.scala 147:106]
  wire  gw_clear_reg_we_17 = _T_644 & picm_wren_ff; // @[pic_ctrl.scala 147:153]
  wire  _T_647 = addr_clear_gw_base_match & _T_88; // @[pic_ctrl.scala 147:106]
  wire  gw_clear_reg_we_18 = _T_647 & picm_wren_ff; // @[pic_ctrl.scala 147:153]
  wire  _T_650 = addr_clear_gw_base_match & _T_91; // @[pic_ctrl.scala 147:106]
  wire  gw_clear_reg_we_19 = _T_650 & picm_wren_ff; // @[pic_ctrl.scala 147:153]
  wire  _T_653 = addr_clear_gw_base_match & _T_94; // @[pic_ctrl.scala 147:106]
  wire  gw_clear_reg_we_20 = _T_653 & picm_wren_ff; // @[pic_ctrl.scala 147:153]
  wire  _T_656 = addr_clear_gw_base_match & _T_97; // @[pic_ctrl.scala 147:106]
  wire  gw_clear_reg_we_21 = _T_656 & picm_wren_ff; // @[pic_ctrl.scala 147:153]
  wire  _T_659 = addr_clear_gw_base_match & _T_100; // @[pic_ctrl.scala 147:106]
  wire  gw_clear_reg_we_22 = _T_659 & picm_wren_ff; // @[pic_ctrl.scala 147:153]
  wire  _T_662 = addr_clear_gw_base_match & _T_103; // @[pic_ctrl.scala 147:106]
  wire  gw_clear_reg_we_23 = _T_662 & picm_wren_ff; // @[pic_ctrl.scala 147:153]
  wire  _T_665 = addr_clear_gw_base_match & _T_106; // @[pic_ctrl.scala 147:106]
  wire  gw_clear_reg_we_24 = _T_665 & picm_wren_ff; // @[pic_ctrl.scala 147:153]
  wire  _T_668 = addr_clear_gw_base_match & _T_109; // @[pic_ctrl.scala 147:106]
  wire  gw_clear_reg_we_25 = _T_668 & picm_wren_ff; // @[pic_ctrl.scala 147:153]
  wire  _T_671 = addr_clear_gw_base_match & _T_112; // @[pic_ctrl.scala 147:106]
  wire  gw_clear_reg_we_26 = _T_671 & picm_wren_ff; // @[pic_ctrl.scala 147:153]
  wire  _T_674 = addr_clear_gw_base_match & _T_115; // @[pic_ctrl.scala 147:106]
  wire  gw_clear_reg_we_27 = _T_674 & picm_wren_ff; // @[pic_ctrl.scala 147:153]
  wire  _T_677 = addr_clear_gw_base_match & _T_118; // @[pic_ctrl.scala 147:106]
  wire  gw_clear_reg_we_28 = _T_677 & picm_wren_ff; // @[pic_ctrl.scala 147:153]
  wire  _T_680 = addr_clear_gw_base_match & _T_121; // @[pic_ctrl.scala 147:106]
  wire  gw_clear_reg_we_29 = _T_680 & picm_wren_ff; // @[pic_ctrl.scala 147:153]
  wire  _T_683 = addr_clear_gw_base_match & _T_124; // @[pic_ctrl.scala 147:106]
  wire  gw_clear_reg_we_30 = _T_683 & picm_wren_ff; // @[pic_ctrl.scala 147:153]
  wire  _T_686 = addr_clear_gw_base_match & _T_127; // @[pic_ctrl.scala 147:106]
  wire  gw_clear_reg_we_31 = _T_686 & picm_wren_ff; // @[pic_ctrl.scala 147:153]
  wire  pic_pri_c1_clk = rvclkhdr_2_io_l1clk; // @[pic_ctrl.scala 97:42 pic_ctrl.scala 134:21]
  reg [3:0] intpriority_reg_1; // @[Reg.scala 27:20]
  reg [3:0] intpriority_reg_2; // @[Reg.scala 27:20]
  reg [3:0] intpriority_reg_3; // @[Reg.scala 27:20]
  reg [3:0] intpriority_reg_4; // @[Reg.scala 27:20]
  reg [3:0] intpriority_reg_5; // @[Reg.scala 27:20]
  reg [3:0] intpriority_reg_6; // @[Reg.scala 27:20]
  reg [3:0] intpriority_reg_7; // @[Reg.scala 27:20]
  reg [3:0] intpriority_reg_8; // @[Reg.scala 27:20]
  reg [3:0] intpriority_reg_9; // @[Reg.scala 27:20]
  reg [3:0] intpriority_reg_10; // @[Reg.scala 27:20]
  reg [3:0] intpriority_reg_11; // @[Reg.scala 27:20]
  reg [3:0] intpriority_reg_12; // @[Reg.scala 27:20]
  reg [3:0] intpriority_reg_13; // @[Reg.scala 27:20]
  reg [3:0] intpriority_reg_14; // @[Reg.scala 27:20]
  reg [3:0] intpriority_reg_15; // @[Reg.scala 27:20]
  reg [3:0] intpriority_reg_16; // @[Reg.scala 27:20]
  reg [3:0] intpriority_reg_17; // @[Reg.scala 27:20]
  reg [3:0] intpriority_reg_18; // @[Reg.scala 27:20]
  reg [3:0] intpriority_reg_19; // @[Reg.scala 27:20]
  reg [3:0] intpriority_reg_20; // @[Reg.scala 27:20]
  reg [3:0] intpriority_reg_21; // @[Reg.scala 27:20]
  reg [3:0] intpriority_reg_22; // @[Reg.scala 27:20]
  reg [3:0] intpriority_reg_23; // @[Reg.scala 27:20]
  reg [3:0] intpriority_reg_24; // @[Reg.scala 27:20]
  reg [3:0] intpriority_reg_25; // @[Reg.scala 27:20]
  reg [3:0] intpriority_reg_26; // @[Reg.scala 27:20]
  reg [3:0] intpriority_reg_27; // @[Reg.scala 27:20]
  reg [3:0] intpriority_reg_28; // @[Reg.scala 27:20]
  reg [3:0] intpriority_reg_29; // @[Reg.scala 27:20]
  reg [3:0] intpriority_reg_30; // @[Reg.scala 27:20]
  reg [3:0] intpriority_reg_31; // @[Reg.scala 27:20]
  wire  pic_int_c1_clk = rvclkhdr_3_io_l1clk; // @[pic_ctrl.scala 98:42 pic_ctrl.scala 135:21]
  reg  intenable_reg_1; // @[Reg.scala 27:20]
  reg  intenable_reg_2; // @[Reg.scala 27:20]
  reg  intenable_reg_3; // @[Reg.scala 27:20]
  reg  intenable_reg_4; // @[Reg.scala 27:20]
  reg  intenable_reg_5; // @[Reg.scala 27:20]
  reg  intenable_reg_6; // @[Reg.scala 27:20]
  reg  intenable_reg_7; // @[Reg.scala 27:20]
  reg  intenable_reg_8; // @[Reg.scala 27:20]
  reg  intenable_reg_9; // @[Reg.scala 27:20]
  reg  intenable_reg_10; // @[Reg.scala 27:20]
  reg  intenable_reg_11; // @[Reg.scala 27:20]
  reg  intenable_reg_12; // @[Reg.scala 27:20]
  reg  intenable_reg_13; // @[Reg.scala 27:20]
  reg  intenable_reg_14; // @[Reg.scala 27:20]
  reg  intenable_reg_15; // @[Reg.scala 27:20]
  reg  intenable_reg_16; // @[Reg.scala 27:20]
  reg  intenable_reg_17; // @[Reg.scala 27:20]
  reg  intenable_reg_18; // @[Reg.scala 27:20]
  reg  intenable_reg_19; // @[Reg.scala 27:20]
  reg  intenable_reg_20; // @[Reg.scala 27:20]
  reg  intenable_reg_21; // @[Reg.scala 27:20]
  reg  intenable_reg_22; // @[Reg.scala 27:20]
  reg  intenable_reg_23; // @[Reg.scala 27:20]
  reg  intenable_reg_24; // @[Reg.scala 27:20]
  reg  intenable_reg_25; // @[Reg.scala 27:20]
  reg  intenable_reg_26; // @[Reg.scala 27:20]
  reg  intenable_reg_27; // @[Reg.scala 27:20]
  reg  intenable_reg_28; // @[Reg.scala 27:20]
  reg  intenable_reg_29; // @[Reg.scala 27:20]
  reg  intenable_reg_30; // @[Reg.scala 27:20]
  reg  intenable_reg_31; // @[Reg.scala 27:20]
  wire  gw_config_c1_clk = rvclkhdr_4_io_l1clk; // @[pic_ctrl.scala 99:42 pic_ctrl.scala 136:21]
  reg [1:0] gw_config_reg_1; // @[Reg.scala 27:20]
  reg [1:0] gw_config_reg_2; // @[Reg.scala 27:20]
  reg [1:0] gw_config_reg_3; // @[Reg.scala 27:20]
  reg [1:0] gw_config_reg_4; // @[Reg.scala 27:20]
  reg [1:0] gw_config_reg_5; // @[Reg.scala 27:20]
  reg [1:0] gw_config_reg_6; // @[Reg.scala 27:20]
  reg [1:0] gw_config_reg_7; // @[Reg.scala 27:20]
  reg [1:0] gw_config_reg_8; // @[Reg.scala 27:20]
  reg [1:0] gw_config_reg_9; // @[Reg.scala 27:20]
  reg [1:0] gw_config_reg_10; // @[Reg.scala 27:20]
  reg [1:0] gw_config_reg_11; // @[Reg.scala 27:20]
  reg [1:0] gw_config_reg_12; // @[Reg.scala 27:20]
  reg [1:0] gw_config_reg_13; // @[Reg.scala 27:20]
  reg [1:0] gw_config_reg_14; // @[Reg.scala 27:20]
  reg [1:0] gw_config_reg_15; // @[Reg.scala 27:20]
  reg [1:0] gw_config_reg_16; // @[Reg.scala 27:20]
  reg [1:0] gw_config_reg_17; // @[Reg.scala 27:20]
  reg [1:0] gw_config_reg_18; // @[Reg.scala 27:20]
  reg [1:0] gw_config_reg_19; // @[Reg.scala 27:20]
  reg [1:0] gw_config_reg_20; // @[Reg.scala 27:20]
  reg [1:0] gw_config_reg_21; // @[Reg.scala 27:20]
  reg [1:0] gw_config_reg_22; // @[Reg.scala 27:20]
  reg [1:0] gw_config_reg_23; // @[Reg.scala 27:20]
  reg [1:0] gw_config_reg_24; // @[Reg.scala 27:20]
  reg [1:0] gw_config_reg_25; // @[Reg.scala 27:20]
  reg [1:0] gw_config_reg_26; // @[Reg.scala 27:20]
  reg [1:0] gw_config_reg_27; // @[Reg.scala 27:20]
  reg [1:0] gw_config_reg_28; // @[Reg.scala 27:20]
  reg [1:0] gw_config_reg_29; // @[Reg.scala 27:20]
  reg [1:0] gw_config_reg_30; // @[Reg.scala 27:20]
  reg [1:0] gw_config_reg_31; // @[Reg.scala 27:20]
  wire  _T_970 = extintsrc_req_sync[1] ^ gw_config_reg_1[0]; // @[pic_ctrl.scala 31:50]
  wire  _T_971 = ~gw_clear_reg_we_1; // @[pic_ctrl.scala 31:92]
  reg  gw_int_pending; // @[pic_ctrl.scala 32:45]
  wire  _T_972 = gw_int_pending & _T_971; // @[pic_ctrl.scala 31:90]
  wire  _T_976 = _T_970 | gw_int_pending; // @[pic_ctrl.scala 33:78]
  wire  extintsrc_req_gw_1 = gw_config_reg_1[1] ? _T_976 : _T_970; // @[pic_ctrl.scala 33:8]
  wire  _T_982 = extintsrc_req_sync[2] ^ gw_config_reg_2[0]; // @[pic_ctrl.scala 31:50]
  wire  _T_983 = ~gw_clear_reg_we_2; // @[pic_ctrl.scala 31:92]
  reg  gw_int_pending_1; // @[pic_ctrl.scala 32:45]
  wire  _T_984 = gw_int_pending_1 & _T_983; // @[pic_ctrl.scala 31:90]
  wire  _T_988 = _T_982 | gw_int_pending_1; // @[pic_ctrl.scala 33:78]
  wire  extintsrc_req_gw_2 = gw_config_reg_2[1] ? _T_988 : _T_982; // @[pic_ctrl.scala 33:8]
  wire  _T_994 = extintsrc_req_sync[3] ^ gw_config_reg_3[0]; // @[pic_ctrl.scala 31:50]
  wire  _T_995 = ~gw_clear_reg_we_3; // @[pic_ctrl.scala 31:92]
  reg  gw_int_pending_2; // @[pic_ctrl.scala 32:45]
  wire  _T_996 = gw_int_pending_2 & _T_995; // @[pic_ctrl.scala 31:90]
  wire  _T_1000 = _T_994 | gw_int_pending_2; // @[pic_ctrl.scala 33:78]
  wire  extintsrc_req_gw_3 = gw_config_reg_3[1] ? _T_1000 : _T_994; // @[pic_ctrl.scala 33:8]
  wire  _T_1006 = extintsrc_req_sync[4] ^ gw_config_reg_4[0]; // @[pic_ctrl.scala 31:50]
  wire  _T_1007 = ~gw_clear_reg_we_4; // @[pic_ctrl.scala 31:92]
  reg  gw_int_pending_3; // @[pic_ctrl.scala 32:45]
  wire  _T_1008 = gw_int_pending_3 & _T_1007; // @[pic_ctrl.scala 31:90]
  wire  _T_1012 = _T_1006 | gw_int_pending_3; // @[pic_ctrl.scala 33:78]
  wire  extintsrc_req_gw_4 = gw_config_reg_4[1] ? _T_1012 : _T_1006; // @[pic_ctrl.scala 33:8]
  wire  _T_1018 = extintsrc_req_sync[5] ^ gw_config_reg_5[0]; // @[pic_ctrl.scala 31:50]
  wire  _T_1019 = ~gw_clear_reg_we_5; // @[pic_ctrl.scala 31:92]
  reg  gw_int_pending_4; // @[pic_ctrl.scala 32:45]
  wire  _T_1020 = gw_int_pending_4 & _T_1019; // @[pic_ctrl.scala 31:90]
  wire  _T_1024 = _T_1018 | gw_int_pending_4; // @[pic_ctrl.scala 33:78]
  wire  extintsrc_req_gw_5 = gw_config_reg_5[1] ? _T_1024 : _T_1018; // @[pic_ctrl.scala 33:8]
  wire  _T_1030 = extintsrc_req_sync[6] ^ gw_config_reg_6[0]; // @[pic_ctrl.scala 31:50]
  wire  _T_1031 = ~gw_clear_reg_we_6; // @[pic_ctrl.scala 31:92]
  reg  gw_int_pending_5; // @[pic_ctrl.scala 32:45]
  wire  _T_1032 = gw_int_pending_5 & _T_1031; // @[pic_ctrl.scala 31:90]
  wire  _T_1036 = _T_1030 | gw_int_pending_5; // @[pic_ctrl.scala 33:78]
  wire  extintsrc_req_gw_6 = gw_config_reg_6[1] ? _T_1036 : _T_1030; // @[pic_ctrl.scala 33:8]
  wire  _T_1042 = extintsrc_req_sync[7] ^ gw_config_reg_7[0]; // @[pic_ctrl.scala 31:50]
  wire  _T_1043 = ~gw_clear_reg_we_7; // @[pic_ctrl.scala 31:92]
  reg  gw_int_pending_6; // @[pic_ctrl.scala 32:45]
  wire  _T_1044 = gw_int_pending_6 & _T_1043; // @[pic_ctrl.scala 31:90]
  wire  _T_1048 = _T_1042 | gw_int_pending_6; // @[pic_ctrl.scala 33:78]
  wire  extintsrc_req_gw_7 = gw_config_reg_7[1] ? _T_1048 : _T_1042; // @[pic_ctrl.scala 33:8]
  wire  _T_1054 = extintsrc_req_sync[8] ^ gw_config_reg_8[0]; // @[pic_ctrl.scala 31:50]
  wire  _T_1055 = ~gw_clear_reg_we_8; // @[pic_ctrl.scala 31:92]
  reg  gw_int_pending_7; // @[pic_ctrl.scala 32:45]
  wire  _T_1056 = gw_int_pending_7 & _T_1055; // @[pic_ctrl.scala 31:90]
  wire  _T_1060 = _T_1054 | gw_int_pending_7; // @[pic_ctrl.scala 33:78]
  wire  extintsrc_req_gw_8 = gw_config_reg_8[1] ? _T_1060 : _T_1054; // @[pic_ctrl.scala 33:8]
  wire  _T_1066 = extintsrc_req_sync[9] ^ gw_config_reg_9[0]; // @[pic_ctrl.scala 31:50]
  wire  _T_1067 = ~gw_clear_reg_we_9; // @[pic_ctrl.scala 31:92]
  reg  gw_int_pending_8; // @[pic_ctrl.scala 32:45]
  wire  _T_1068 = gw_int_pending_8 & _T_1067; // @[pic_ctrl.scala 31:90]
  wire  _T_1072 = _T_1066 | gw_int_pending_8; // @[pic_ctrl.scala 33:78]
  wire  extintsrc_req_gw_9 = gw_config_reg_9[1] ? _T_1072 : _T_1066; // @[pic_ctrl.scala 33:8]
  wire  _T_1078 = extintsrc_req_sync[10] ^ gw_config_reg_10[0]; // @[pic_ctrl.scala 31:50]
  wire  _T_1079 = ~gw_clear_reg_we_10; // @[pic_ctrl.scala 31:92]
  reg  gw_int_pending_9; // @[pic_ctrl.scala 32:45]
  wire  _T_1080 = gw_int_pending_9 & _T_1079; // @[pic_ctrl.scala 31:90]
  wire  _T_1084 = _T_1078 | gw_int_pending_9; // @[pic_ctrl.scala 33:78]
  wire  extintsrc_req_gw_10 = gw_config_reg_10[1] ? _T_1084 : _T_1078; // @[pic_ctrl.scala 33:8]
  wire  _T_1090 = extintsrc_req_sync[11] ^ gw_config_reg_11[0]; // @[pic_ctrl.scala 31:50]
  wire  _T_1091 = ~gw_clear_reg_we_11; // @[pic_ctrl.scala 31:92]
  reg  gw_int_pending_10; // @[pic_ctrl.scala 32:45]
  wire  _T_1092 = gw_int_pending_10 & _T_1091; // @[pic_ctrl.scala 31:90]
  wire  _T_1096 = _T_1090 | gw_int_pending_10; // @[pic_ctrl.scala 33:78]
  wire  extintsrc_req_gw_11 = gw_config_reg_11[1] ? _T_1096 : _T_1090; // @[pic_ctrl.scala 33:8]
  wire  _T_1102 = extintsrc_req_sync[12] ^ gw_config_reg_12[0]; // @[pic_ctrl.scala 31:50]
  wire  _T_1103 = ~gw_clear_reg_we_12; // @[pic_ctrl.scala 31:92]
  reg  gw_int_pending_11; // @[pic_ctrl.scala 32:45]
  wire  _T_1104 = gw_int_pending_11 & _T_1103; // @[pic_ctrl.scala 31:90]
  wire  _T_1108 = _T_1102 | gw_int_pending_11; // @[pic_ctrl.scala 33:78]
  wire  extintsrc_req_gw_12 = gw_config_reg_12[1] ? _T_1108 : _T_1102; // @[pic_ctrl.scala 33:8]
  wire  _T_1114 = extintsrc_req_sync[13] ^ gw_config_reg_13[0]; // @[pic_ctrl.scala 31:50]
  wire  _T_1115 = ~gw_clear_reg_we_13; // @[pic_ctrl.scala 31:92]
  reg  gw_int_pending_12; // @[pic_ctrl.scala 32:45]
  wire  _T_1116 = gw_int_pending_12 & _T_1115; // @[pic_ctrl.scala 31:90]
  wire  _T_1120 = _T_1114 | gw_int_pending_12; // @[pic_ctrl.scala 33:78]
  wire  extintsrc_req_gw_13 = gw_config_reg_13[1] ? _T_1120 : _T_1114; // @[pic_ctrl.scala 33:8]
  wire  _T_1126 = extintsrc_req_sync[14] ^ gw_config_reg_14[0]; // @[pic_ctrl.scala 31:50]
  wire  _T_1127 = ~gw_clear_reg_we_14; // @[pic_ctrl.scala 31:92]
  reg  gw_int_pending_13; // @[pic_ctrl.scala 32:45]
  wire  _T_1128 = gw_int_pending_13 & _T_1127; // @[pic_ctrl.scala 31:90]
  wire  _T_1132 = _T_1126 | gw_int_pending_13; // @[pic_ctrl.scala 33:78]
  wire  extintsrc_req_gw_14 = gw_config_reg_14[1] ? _T_1132 : _T_1126; // @[pic_ctrl.scala 33:8]
  wire  _T_1138 = extintsrc_req_sync[15] ^ gw_config_reg_15[0]; // @[pic_ctrl.scala 31:50]
  wire  _T_1139 = ~gw_clear_reg_we_15; // @[pic_ctrl.scala 31:92]
  reg  gw_int_pending_14; // @[pic_ctrl.scala 32:45]
  wire  _T_1140 = gw_int_pending_14 & _T_1139; // @[pic_ctrl.scala 31:90]
  wire  _T_1144 = _T_1138 | gw_int_pending_14; // @[pic_ctrl.scala 33:78]
  wire  extintsrc_req_gw_15 = gw_config_reg_15[1] ? _T_1144 : _T_1138; // @[pic_ctrl.scala 33:8]
  wire  _T_1150 = extintsrc_req_sync[16] ^ gw_config_reg_16[0]; // @[pic_ctrl.scala 31:50]
  wire  _T_1151 = ~gw_clear_reg_we_16; // @[pic_ctrl.scala 31:92]
  reg  gw_int_pending_15; // @[pic_ctrl.scala 32:45]
  wire  _T_1152 = gw_int_pending_15 & _T_1151; // @[pic_ctrl.scala 31:90]
  wire  _T_1156 = _T_1150 | gw_int_pending_15; // @[pic_ctrl.scala 33:78]
  wire  extintsrc_req_gw_16 = gw_config_reg_16[1] ? _T_1156 : _T_1150; // @[pic_ctrl.scala 33:8]
  wire  _T_1162 = extintsrc_req_sync[17] ^ gw_config_reg_17[0]; // @[pic_ctrl.scala 31:50]
  wire  _T_1163 = ~gw_clear_reg_we_17; // @[pic_ctrl.scala 31:92]
  reg  gw_int_pending_16; // @[pic_ctrl.scala 32:45]
  wire  _T_1164 = gw_int_pending_16 & _T_1163; // @[pic_ctrl.scala 31:90]
  wire  _T_1168 = _T_1162 | gw_int_pending_16; // @[pic_ctrl.scala 33:78]
  wire  extintsrc_req_gw_17 = gw_config_reg_17[1] ? _T_1168 : _T_1162; // @[pic_ctrl.scala 33:8]
  wire  _T_1174 = extintsrc_req_sync[18] ^ gw_config_reg_18[0]; // @[pic_ctrl.scala 31:50]
  wire  _T_1175 = ~gw_clear_reg_we_18; // @[pic_ctrl.scala 31:92]
  reg  gw_int_pending_17; // @[pic_ctrl.scala 32:45]
  wire  _T_1176 = gw_int_pending_17 & _T_1175; // @[pic_ctrl.scala 31:90]
  wire  _T_1180 = _T_1174 | gw_int_pending_17; // @[pic_ctrl.scala 33:78]
  wire  extintsrc_req_gw_18 = gw_config_reg_18[1] ? _T_1180 : _T_1174; // @[pic_ctrl.scala 33:8]
  wire  _T_1186 = extintsrc_req_sync[19] ^ gw_config_reg_19[0]; // @[pic_ctrl.scala 31:50]
  wire  _T_1187 = ~gw_clear_reg_we_19; // @[pic_ctrl.scala 31:92]
  reg  gw_int_pending_18; // @[pic_ctrl.scala 32:45]
  wire  _T_1188 = gw_int_pending_18 & _T_1187; // @[pic_ctrl.scala 31:90]
  wire  _T_1192 = _T_1186 | gw_int_pending_18; // @[pic_ctrl.scala 33:78]
  wire  extintsrc_req_gw_19 = gw_config_reg_19[1] ? _T_1192 : _T_1186; // @[pic_ctrl.scala 33:8]
  wire  _T_1198 = extintsrc_req_sync[20] ^ gw_config_reg_20[0]; // @[pic_ctrl.scala 31:50]
  wire  _T_1199 = ~gw_clear_reg_we_20; // @[pic_ctrl.scala 31:92]
  reg  gw_int_pending_19; // @[pic_ctrl.scala 32:45]
  wire  _T_1200 = gw_int_pending_19 & _T_1199; // @[pic_ctrl.scala 31:90]
  wire  _T_1204 = _T_1198 | gw_int_pending_19; // @[pic_ctrl.scala 33:78]
  wire  extintsrc_req_gw_20 = gw_config_reg_20[1] ? _T_1204 : _T_1198; // @[pic_ctrl.scala 33:8]
  wire  _T_1210 = extintsrc_req_sync[21] ^ gw_config_reg_21[0]; // @[pic_ctrl.scala 31:50]
  wire  _T_1211 = ~gw_clear_reg_we_21; // @[pic_ctrl.scala 31:92]
  reg  gw_int_pending_20; // @[pic_ctrl.scala 32:45]
  wire  _T_1212 = gw_int_pending_20 & _T_1211; // @[pic_ctrl.scala 31:90]
  wire  _T_1216 = _T_1210 | gw_int_pending_20; // @[pic_ctrl.scala 33:78]
  wire  extintsrc_req_gw_21 = gw_config_reg_21[1] ? _T_1216 : _T_1210; // @[pic_ctrl.scala 33:8]
  wire  _T_1222 = extintsrc_req_sync[22] ^ gw_config_reg_22[0]; // @[pic_ctrl.scala 31:50]
  wire  _T_1223 = ~gw_clear_reg_we_22; // @[pic_ctrl.scala 31:92]
  reg  gw_int_pending_21; // @[pic_ctrl.scala 32:45]
  wire  _T_1224 = gw_int_pending_21 & _T_1223; // @[pic_ctrl.scala 31:90]
  wire  _T_1228 = _T_1222 | gw_int_pending_21; // @[pic_ctrl.scala 33:78]
  wire  extintsrc_req_gw_22 = gw_config_reg_22[1] ? _T_1228 : _T_1222; // @[pic_ctrl.scala 33:8]
  wire  _T_1234 = extintsrc_req_sync[23] ^ gw_config_reg_23[0]; // @[pic_ctrl.scala 31:50]
  wire  _T_1235 = ~gw_clear_reg_we_23; // @[pic_ctrl.scala 31:92]
  reg  gw_int_pending_22; // @[pic_ctrl.scala 32:45]
  wire  _T_1236 = gw_int_pending_22 & _T_1235; // @[pic_ctrl.scala 31:90]
  wire  _T_1240 = _T_1234 | gw_int_pending_22; // @[pic_ctrl.scala 33:78]
  wire  extintsrc_req_gw_23 = gw_config_reg_23[1] ? _T_1240 : _T_1234; // @[pic_ctrl.scala 33:8]
  wire  _T_1246 = extintsrc_req_sync[24] ^ gw_config_reg_24[0]; // @[pic_ctrl.scala 31:50]
  wire  _T_1247 = ~gw_clear_reg_we_24; // @[pic_ctrl.scala 31:92]
  reg  gw_int_pending_23; // @[pic_ctrl.scala 32:45]
  wire  _T_1248 = gw_int_pending_23 & _T_1247; // @[pic_ctrl.scala 31:90]
  wire  _T_1252 = _T_1246 | gw_int_pending_23; // @[pic_ctrl.scala 33:78]
  wire  extintsrc_req_gw_24 = gw_config_reg_24[1] ? _T_1252 : _T_1246; // @[pic_ctrl.scala 33:8]
  wire  _T_1258 = extintsrc_req_sync[25] ^ gw_config_reg_25[0]; // @[pic_ctrl.scala 31:50]
  wire  _T_1259 = ~gw_clear_reg_we_25; // @[pic_ctrl.scala 31:92]
  reg  gw_int_pending_24; // @[pic_ctrl.scala 32:45]
  wire  _T_1260 = gw_int_pending_24 & _T_1259; // @[pic_ctrl.scala 31:90]
  wire  _T_1264 = _T_1258 | gw_int_pending_24; // @[pic_ctrl.scala 33:78]
  wire  extintsrc_req_gw_25 = gw_config_reg_25[1] ? _T_1264 : _T_1258; // @[pic_ctrl.scala 33:8]
  wire  _T_1270 = extintsrc_req_sync[26] ^ gw_config_reg_26[0]; // @[pic_ctrl.scala 31:50]
  wire  _T_1271 = ~gw_clear_reg_we_26; // @[pic_ctrl.scala 31:92]
  reg  gw_int_pending_25; // @[pic_ctrl.scala 32:45]
  wire  _T_1272 = gw_int_pending_25 & _T_1271; // @[pic_ctrl.scala 31:90]
  wire  _T_1276 = _T_1270 | gw_int_pending_25; // @[pic_ctrl.scala 33:78]
  wire  extintsrc_req_gw_26 = gw_config_reg_26[1] ? _T_1276 : _T_1270; // @[pic_ctrl.scala 33:8]
  wire  _T_1282 = extintsrc_req_sync[27] ^ gw_config_reg_27[0]; // @[pic_ctrl.scala 31:50]
  wire  _T_1283 = ~gw_clear_reg_we_27; // @[pic_ctrl.scala 31:92]
  reg  gw_int_pending_26; // @[pic_ctrl.scala 32:45]
  wire  _T_1284 = gw_int_pending_26 & _T_1283; // @[pic_ctrl.scala 31:90]
  wire  _T_1288 = _T_1282 | gw_int_pending_26; // @[pic_ctrl.scala 33:78]
  wire  extintsrc_req_gw_27 = gw_config_reg_27[1] ? _T_1288 : _T_1282; // @[pic_ctrl.scala 33:8]
  wire  _T_1294 = extintsrc_req_sync[28] ^ gw_config_reg_28[0]; // @[pic_ctrl.scala 31:50]
  wire  _T_1295 = ~gw_clear_reg_we_28; // @[pic_ctrl.scala 31:92]
  reg  gw_int_pending_27; // @[pic_ctrl.scala 32:45]
  wire  _T_1296 = gw_int_pending_27 & _T_1295; // @[pic_ctrl.scala 31:90]
  wire  _T_1300 = _T_1294 | gw_int_pending_27; // @[pic_ctrl.scala 33:78]
  wire  extintsrc_req_gw_28 = gw_config_reg_28[1] ? _T_1300 : _T_1294; // @[pic_ctrl.scala 33:8]
  wire  _T_1306 = extintsrc_req_sync[29] ^ gw_config_reg_29[0]; // @[pic_ctrl.scala 31:50]
  wire  _T_1307 = ~gw_clear_reg_we_29; // @[pic_ctrl.scala 31:92]
  reg  gw_int_pending_28; // @[pic_ctrl.scala 32:45]
  wire  _T_1308 = gw_int_pending_28 & _T_1307; // @[pic_ctrl.scala 31:90]
  wire  _T_1312 = _T_1306 | gw_int_pending_28; // @[pic_ctrl.scala 33:78]
  wire  extintsrc_req_gw_29 = gw_config_reg_29[1] ? _T_1312 : _T_1306; // @[pic_ctrl.scala 33:8]
  wire  _T_1318 = extintsrc_req_sync[30] ^ gw_config_reg_30[0]; // @[pic_ctrl.scala 31:50]
  wire  _T_1319 = ~gw_clear_reg_we_30; // @[pic_ctrl.scala 31:92]
  reg  gw_int_pending_29; // @[pic_ctrl.scala 32:45]
  wire  _T_1320 = gw_int_pending_29 & _T_1319; // @[pic_ctrl.scala 31:90]
  wire  _T_1324 = _T_1318 | gw_int_pending_29; // @[pic_ctrl.scala 33:78]
  wire  extintsrc_req_gw_30 = gw_config_reg_30[1] ? _T_1324 : _T_1318; // @[pic_ctrl.scala 33:8]
  wire  _T_1330 = extintsrc_req_sync[31] ^ gw_config_reg_31[0]; // @[pic_ctrl.scala 31:50]
  wire  _T_1331 = ~gw_clear_reg_we_31; // @[pic_ctrl.scala 31:92]
  reg  gw_int_pending_30; // @[pic_ctrl.scala 32:45]
  wire  _T_1332 = gw_int_pending_30 & _T_1331; // @[pic_ctrl.scala 31:90]
  wire  _T_1336 = _T_1330 | gw_int_pending_30; // @[pic_ctrl.scala 33:78]
  wire  extintsrc_req_gw_31 = gw_config_reg_31[1] ? _T_1336 : _T_1330; // @[pic_ctrl.scala 33:8]
  reg  config_reg; // @[Reg.scala 27:20]
  wire [3:0] intpriority_reg_0 = 4'h0; // @[pic_ctrl.scala 148:32 pic_ctrl.scala 149:208]
  wire [3:0] _T_1342 = ~intpriority_reg_1; // @[pic_ctrl.scala 160:90]
  wire [3:0] intpriority_reg_inv_1 = config_reg ? _T_1342 : intpriority_reg_1; // @[pic_ctrl.scala 160:71]
  wire [3:0] _T_1345 = ~intpriority_reg_2; // @[pic_ctrl.scala 160:90]
  wire [3:0] intpriority_reg_inv_2 = config_reg ? _T_1345 : intpriority_reg_2; // @[pic_ctrl.scala 160:71]
  wire [3:0] _T_1348 = ~intpriority_reg_3; // @[pic_ctrl.scala 160:90]
  wire [3:0] intpriority_reg_inv_3 = config_reg ? _T_1348 : intpriority_reg_3; // @[pic_ctrl.scala 160:71]
  wire [3:0] _T_1351 = ~intpriority_reg_4; // @[pic_ctrl.scala 160:90]
  wire [3:0] intpriority_reg_inv_4 = config_reg ? _T_1351 : intpriority_reg_4; // @[pic_ctrl.scala 160:71]
  wire [3:0] _T_1354 = ~intpriority_reg_5; // @[pic_ctrl.scala 160:90]
  wire [3:0] intpriority_reg_inv_5 = config_reg ? _T_1354 : intpriority_reg_5; // @[pic_ctrl.scala 160:71]
  wire [3:0] _T_1357 = ~intpriority_reg_6; // @[pic_ctrl.scala 160:90]
  wire [3:0] intpriority_reg_inv_6 = config_reg ? _T_1357 : intpriority_reg_6; // @[pic_ctrl.scala 160:71]
  wire [3:0] _T_1360 = ~intpriority_reg_7; // @[pic_ctrl.scala 160:90]
  wire [3:0] intpriority_reg_inv_7 = config_reg ? _T_1360 : intpriority_reg_7; // @[pic_ctrl.scala 160:71]
  wire [3:0] _T_1363 = ~intpriority_reg_8; // @[pic_ctrl.scala 160:90]
  wire [3:0] intpriority_reg_inv_8 = config_reg ? _T_1363 : intpriority_reg_8; // @[pic_ctrl.scala 160:71]
  wire [3:0] _T_1366 = ~intpriority_reg_9; // @[pic_ctrl.scala 160:90]
  wire [3:0] intpriority_reg_inv_9 = config_reg ? _T_1366 : intpriority_reg_9; // @[pic_ctrl.scala 160:71]
  wire [3:0] _T_1369 = ~intpriority_reg_10; // @[pic_ctrl.scala 160:90]
  wire [3:0] intpriority_reg_inv_10 = config_reg ? _T_1369 : intpriority_reg_10; // @[pic_ctrl.scala 160:71]
  wire [3:0] _T_1372 = ~intpriority_reg_11; // @[pic_ctrl.scala 160:90]
  wire [3:0] intpriority_reg_inv_11 = config_reg ? _T_1372 : intpriority_reg_11; // @[pic_ctrl.scala 160:71]
  wire [3:0] _T_1375 = ~intpriority_reg_12; // @[pic_ctrl.scala 160:90]
  wire [3:0] intpriority_reg_inv_12 = config_reg ? _T_1375 : intpriority_reg_12; // @[pic_ctrl.scala 160:71]
  wire [3:0] _T_1378 = ~intpriority_reg_13; // @[pic_ctrl.scala 160:90]
  wire [3:0] intpriority_reg_inv_13 = config_reg ? _T_1378 : intpriority_reg_13; // @[pic_ctrl.scala 160:71]
  wire [3:0] _T_1381 = ~intpriority_reg_14; // @[pic_ctrl.scala 160:90]
  wire [3:0] intpriority_reg_inv_14 = config_reg ? _T_1381 : intpriority_reg_14; // @[pic_ctrl.scala 160:71]
  wire [3:0] _T_1384 = ~intpriority_reg_15; // @[pic_ctrl.scala 160:90]
  wire [3:0] intpriority_reg_inv_15 = config_reg ? _T_1384 : intpriority_reg_15; // @[pic_ctrl.scala 160:71]
  wire [3:0] _T_1387 = ~intpriority_reg_16; // @[pic_ctrl.scala 160:90]
  wire [3:0] intpriority_reg_inv_16 = config_reg ? _T_1387 : intpriority_reg_16; // @[pic_ctrl.scala 160:71]
  wire [3:0] _T_1390 = ~intpriority_reg_17; // @[pic_ctrl.scala 160:90]
  wire [3:0] intpriority_reg_inv_17 = config_reg ? _T_1390 : intpriority_reg_17; // @[pic_ctrl.scala 160:71]
  wire [3:0] _T_1393 = ~intpriority_reg_18; // @[pic_ctrl.scala 160:90]
  wire [3:0] intpriority_reg_inv_18 = config_reg ? _T_1393 : intpriority_reg_18; // @[pic_ctrl.scala 160:71]
  wire [3:0] _T_1396 = ~intpriority_reg_19; // @[pic_ctrl.scala 160:90]
  wire [3:0] intpriority_reg_inv_19 = config_reg ? _T_1396 : intpriority_reg_19; // @[pic_ctrl.scala 160:71]
  wire [3:0] _T_1399 = ~intpriority_reg_20; // @[pic_ctrl.scala 160:90]
  wire [3:0] intpriority_reg_inv_20 = config_reg ? _T_1399 : intpriority_reg_20; // @[pic_ctrl.scala 160:71]
  wire [3:0] _T_1402 = ~intpriority_reg_21; // @[pic_ctrl.scala 160:90]
  wire [3:0] intpriority_reg_inv_21 = config_reg ? _T_1402 : intpriority_reg_21; // @[pic_ctrl.scala 160:71]
  wire [3:0] _T_1405 = ~intpriority_reg_22; // @[pic_ctrl.scala 160:90]
  wire [3:0] intpriority_reg_inv_22 = config_reg ? _T_1405 : intpriority_reg_22; // @[pic_ctrl.scala 160:71]
  wire [3:0] _T_1408 = ~intpriority_reg_23; // @[pic_ctrl.scala 160:90]
  wire [3:0] intpriority_reg_inv_23 = config_reg ? _T_1408 : intpriority_reg_23; // @[pic_ctrl.scala 160:71]
  wire [3:0] _T_1411 = ~intpriority_reg_24; // @[pic_ctrl.scala 160:90]
  wire [3:0] intpriority_reg_inv_24 = config_reg ? _T_1411 : intpriority_reg_24; // @[pic_ctrl.scala 160:71]
  wire [3:0] _T_1414 = ~intpriority_reg_25; // @[pic_ctrl.scala 160:90]
  wire [3:0] intpriority_reg_inv_25 = config_reg ? _T_1414 : intpriority_reg_25; // @[pic_ctrl.scala 160:71]
  wire [3:0] _T_1417 = ~intpriority_reg_26; // @[pic_ctrl.scala 160:90]
  wire [3:0] intpriority_reg_inv_26 = config_reg ? _T_1417 : intpriority_reg_26; // @[pic_ctrl.scala 160:71]
  wire [3:0] _T_1420 = ~intpriority_reg_27; // @[pic_ctrl.scala 160:90]
  wire [3:0] intpriority_reg_inv_27 = config_reg ? _T_1420 : intpriority_reg_27; // @[pic_ctrl.scala 160:71]
  wire [3:0] _T_1423 = ~intpriority_reg_28; // @[pic_ctrl.scala 160:90]
  wire [3:0] intpriority_reg_inv_28 = config_reg ? _T_1423 : intpriority_reg_28; // @[pic_ctrl.scala 160:71]
  wire [3:0] _T_1426 = ~intpriority_reg_29; // @[pic_ctrl.scala 160:90]
  wire [3:0] intpriority_reg_inv_29 = config_reg ? _T_1426 : intpriority_reg_29; // @[pic_ctrl.scala 160:71]
  wire [3:0] _T_1429 = ~intpriority_reg_30; // @[pic_ctrl.scala 160:90]
  wire [3:0] intpriority_reg_inv_30 = config_reg ? _T_1429 : intpriority_reg_30; // @[pic_ctrl.scala 160:71]
  wire [3:0] _T_1432 = ~intpriority_reg_31; // @[pic_ctrl.scala 160:90]
  wire [3:0] intpriority_reg_inv_31 = config_reg ? _T_1432 : intpriority_reg_31; // @[pic_ctrl.scala 160:71]
  wire  _T_1438 = extintsrc_req_gw_1 & intenable_reg_1; // @[pic_ctrl.scala 161:110]
  wire [3:0] _T_1440 = _T_1438 ? 4'hf : 4'h0; // @[Bitwise.scala 72:12]
  wire [3:0] intpend_w_prior_en_1 = _T_1440 & intpriority_reg_inv_1; // @[pic_ctrl.scala 161:130]
  wire  _T_1442 = extintsrc_req_gw_2 & intenable_reg_2; // @[pic_ctrl.scala 161:110]
  wire [3:0] _T_1444 = _T_1442 ? 4'hf : 4'h0; // @[Bitwise.scala 72:12]
  wire [3:0] intpend_w_prior_en_2 = _T_1444 & intpriority_reg_inv_2; // @[pic_ctrl.scala 161:130]
  wire  _T_1446 = extintsrc_req_gw_3 & intenable_reg_3; // @[pic_ctrl.scala 161:110]
  wire [3:0] _T_1448 = _T_1446 ? 4'hf : 4'h0; // @[Bitwise.scala 72:12]
  wire [3:0] intpend_w_prior_en_3 = _T_1448 & intpriority_reg_inv_3; // @[pic_ctrl.scala 161:130]
  wire  _T_1450 = extintsrc_req_gw_4 & intenable_reg_4; // @[pic_ctrl.scala 161:110]
  wire [3:0] _T_1452 = _T_1450 ? 4'hf : 4'h0; // @[Bitwise.scala 72:12]
  wire [3:0] intpend_w_prior_en_4 = _T_1452 & intpriority_reg_inv_4; // @[pic_ctrl.scala 161:130]
  wire  _T_1454 = extintsrc_req_gw_5 & intenable_reg_5; // @[pic_ctrl.scala 161:110]
  wire [3:0] _T_1456 = _T_1454 ? 4'hf : 4'h0; // @[Bitwise.scala 72:12]
  wire [3:0] intpend_w_prior_en_5 = _T_1456 & intpriority_reg_inv_5; // @[pic_ctrl.scala 161:130]
  wire  _T_1458 = extintsrc_req_gw_6 & intenable_reg_6; // @[pic_ctrl.scala 161:110]
  wire [3:0] _T_1460 = _T_1458 ? 4'hf : 4'h0; // @[Bitwise.scala 72:12]
  wire [3:0] intpend_w_prior_en_6 = _T_1460 & intpriority_reg_inv_6; // @[pic_ctrl.scala 161:130]
  wire  _T_1462 = extintsrc_req_gw_7 & intenable_reg_7; // @[pic_ctrl.scala 161:110]
  wire [3:0] _T_1464 = _T_1462 ? 4'hf : 4'h0; // @[Bitwise.scala 72:12]
  wire [3:0] intpend_w_prior_en_7 = _T_1464 & intpriority_reg_inv_7; // @[pic_ctrl.scala 161:130]
  wire  _T_1466 = extintsrc_req_gw_8 & intenable_reg_8; // @[pic_ctrl.scala 161:110]
  wire [3:0] _T_1468 = _T_1466 ? 4'hf : 4'h0; // @[Bitwise.scala 72:12]
  wire [3:0] intpend_w_prior_en_8 = _T_1468 & intpriority_reg_inv_8; // @[pic_ctrl.scala 161:130]
  wire  _T_1470 = extintsrc_req_gw_9 & intenable_reg_9; // @[pic_ctrl.scala 161:110]
  wire [3:0] _T_1472 = _T_1470 ? 4'hf : 4'h0; // @[Bitwise.scala 72:12]
  wire [3:0] intpend_w_prior_en_9 = _T_1472 & intpriority_reg_inv_9; // @[pic_ctrl.scala 161:130]
  wire  _T_1474 = extintsrc_req_gw_10 & intenable_reg_10; // @[pic_ctrl.scala 161:110]
  wire [3:0] _T_1476 = _T_1474 ? 4'hf : 4'h0; // @[Bitwise.scala 72:12]
  wire [3:0] intpend_w_prior_en_10 = _T_1476 & intpriority_reg_inv_10; // @[pic_ctrl.scala 161:130]
  wire  _T_1478 = extintsrc_req_gw_11 & intenable_reg_11; // @[pic_ctrl.scala 161:110]
  wire [3:0] _T_1480 = _T_1478 ? 4'hf : 4'h0; // @[Bitwise.scala 72:12]
  wire [3:0] intpend_w_prior_en_11 = _T_1480 & intpriority_reg_inv_11; // @[pic_ctrl.scala 161:130]
  wire  _T_1482 = extintsrc_req_gw_12 & intenable_reg_12; // @[pic_ctrl.scala 161:110]
  wire [3:0] _T_1484 = _T_1482 ? 4'hf : 4'h0; // @[Bitwise.scala 72:12]
  wire [3:0] intpend_w_prior_en_12 = _T_1484 & intpriority_reg_inv_12; // @[pic_ctrl.scala 161:130]
  wire  _T_1486 = extintsrc_req_gw_13 & intenable_reg_13; // @[pic_ctrl.scala 161:110]
  wire [3:0] _T_1488 = _T_1486 ? 4'hf : 4'h0; // @[Bitwise.scala 72:12]
  wire [3:0] intpend_w_prior_en_13 = _T_1488 & intpriority_reg_inv_13; // @[pic_ctrl.scala 161:130]
  wire  _T_1490 = extintsrc_req_gw_14 & intenable_reg_14; // @[pic_ctrl.scala 161:110]
  wire [3:0] _T_1492 = _T_1490 ? 4'hf : 4'h0; // @[Bitwise.scala 72:12]
  wire [3:0] intpend_w_prior_en_14 = _T_1492 & intpriority_reg_inv_14; // @[pic_ctrl.scala 161:130]
  wire  _T_1494 = extintsrc_req_gw_15 & intenable_reg_15; // @[pic_ctrl.scala 161:110]
  wire [3:0] _T_1496 = _T_1494 ? 4'hf : 4'h0; // @[Bitwise.scala 72:12]
  wire [3:0] intpend_w_prior_en_15 = _T_1496 & intpriority_reg_inv_15; // @[pic_ctrl.scala 161:130]
  wire  _T_1498 = extintsrc_req_gw_16 & intenable_reg_16; // @[pic_ctrl.scala 161:110]
  wire [3:0] _T_1500 = _T_1498 ? 4'hf : 4'h0; // @[Bitwise.scala 72:12]
  wire [3:0] intpend_w_prior_en_16 = _T_1500 & intpriority_reg_inv_16; // @[pic_ctrl.scala 161:130]
  wire  _T_1502 = extintsrc_req_gw_17 & intenable_reg_17; // @[pic_ctrl.scala 161:110]
  wire [3:0] _T_1504 = _T_1502 ? 4'hf : 4'h0; // @[Bitwise.scala 72:12]
  wire [3:0] intpend_w_prior_en_17 = _T_1504 & intpriority_reg_inv_17; // @[pic_ctrl.scala 161:130]
  wire  _T_1506 = extintsrc_req_gw_18 & intenable_reg_18; // @[pic_ctrl.scala 161:110]
  wire [3:0] _T_1508 = _T_1506 ? 4'hf : 4'h0; // @[Bitwise.scala 72:12]
  wire [3:0] intpend_w_prior_en_18 = _T_1508 & intpriority_reg_inv_18; // @[pic_ctrl.scala 161:130]
  wire  _T_1510 = extintsrc_req_gw_19 & intenable_reg_19; // @[pic_ctrl.scala 161:110]
  wire [3:0] _T_1512 = _T_1510 ? 4'hf : 4'h0; // @[Bitwise.scala 72:12]
  wire [3:0] intpend_w_prior_en_19 = _T_1512 & intpriority_reg_inv_19; // @[pic_ctrl.scala 161:130]
  wire  _T_1514 = extintsrc_req_gw_20 & intenable_reg_20; // @[pic_ctrl.scala 161:110]
  wire [3:0] _T_1516 = _T_1514 ? 4'hf : 4'h0; // @[Bitwise.scala 72:12]
  wire [3:0] intpend_w_prior_en_20 = _T_1516 & intpriority_reg_inv_20; // @[pic_ctrl.scala 161:130]
  wire  _T_1518 = extintsrc_req_gw_21 & intenable_reg_21; // @[pic_ctrl.scala 161:110]
  wire [3:0] _T_1520 = _T_1518 ? 4'hf : 4'h0; // @[Bitwise.scala 72:12]
  wire [3:0] intpend_w_prior_en_21 = _T_1520 & intpriority_reg_inv_21; // @[pic_ctrl.scala 161:130]
  wire  _T_1522 = extintsrc_req_gw_22 & intenable_reg_22; // @[pic_ctrl.scala 161:110]
  wire [3:0] _T_1524 = _T_1522 ? 4'hf : 4'h0; // @[Bitwise.scala 72:12]
  wire [3:0] intpend_w_prior_en_22 = _T_1524 & intpriority_reg_inv_22; // @[pic_ctrl.scala 161:130]
  wire  _T_1526 = extintsrc_req_gw_23 & intenable_reg_23; // @[pic_ctrl.scala 161:110]
  wire [3:0] _T_1528 = _T_1526 ? 4'hf : 4'h0; // @[Bitwise.scala 72:12]
  wire [3:0] intpend_w_prior_en_23 = _T_1528 & intpriority_reg_inv_23; // @[pic_ctrl.scala 161:130]
  wire  _T_1530 = extintsrc_req_gw_24 & intenable_reg_24; // @[pic_ctrl.scala 161:110]
  wire [3:0] _T_1532 = _T_1530 ? 4'hf : 4'h0; // @[Bitwise.scala 72:12]
  wire [3:0] intpend_w_prior_en_24 = _T_1532 & intpriority_reg_inv_24; // @[pic_ctrl.scala 161:130]
  wire  _T_1534 = extintsrc_req_gw_25 & intenable_reg_25; // @[pic_ctrl.scala 161:110]
  wire [3:0] _T_1536 = _T_1534 ? 4'hf : 4'h0; // @[Bitwise.scala 72:12]
  wire [3:0] intpend_w_prior_en_25 = _T_1536 & intpriority_reg_inv_25; // @[pic_ctrl.scala 161:130]
  wire  _T_1538 = extintsrc_req_gw_26 & intenable_reg_26; // @[pic_ctrl.scala 161:110]
  wire [3:0] _T_1540 = _T_1538 ? 4'hf : 4'h0; // @[Bitwise.scala 72:12]
  wire [3:0] intpend_w_prior_en_26 = _T_1540 & intpriority_reg_inv_26; // @[pic_ctrl.scala 161:130]
  wire  _T_1542 = extintsrc_req_gw_27 & intenable_reg_27; // @[pic_ctrl.scala 161:110]
  wire [3:0] _T_1544 = _T_1542 ? 4'hf : 4'h0; // @[Bitwise.scala 72:12]
  wire [3:0] intpend_w_prior_en_27 = _T_1544 & intpriority_reg_inv_27; // @[pic_ctrl.scala 161:130]
  wire  _T_1546 = extintsrc_req_gw_28 & intenable_reg_28; // @[pic_ctrl.scala 161:110]
  wire [3:0] _T_1548 = _T_1546 ? 4'hf : 4'h0; // @[Bitwise.scala 72:12]
  wire [3:0] intpend_w_prior_en_28 = _T_1548 & intpriority_reg_inv_28; // @[pic_ctrl.scala 161:130]
  wire  _T_1550 = extintsrc_req_gw_29 & intenable_reg_29; // @[pic_ctrl.scala 161:110]
  wire [3:0] _T_1552 = _T_1550 ? 4'hf : 4'h0; // @[Bitwise.scala 72:12]
  wire [3:0] intpend_w_prior_en_29 = _T_1552 & intpriority_reg_inv_29; // @[pic_ctrl.scala 161:130]
  wire  _T_1554 = extintsrc_req_gw_30 & intenable_reg_30; // @[pic_ctrl.scala 161:110]
  wire [3:0] _T_1556 = _T_1554 ? 4'hf : 4'h0; // @[Bitwise.scala 72:12]
  wire [3:0] intpend_w_prior_en_30 = _T_1556 & intpriority_reg_inv_30; // @[pic_ctrl.scala 161:130]
  wire  _T_1558 = extintsrc_req_gw_31 & intenable_reg_31; // @[pic_ctrl.scala 161:110]
  wire [3:0] _T_1560 = _T_1558 ? 4'hf : 4'h0; // @[Bitwise.scala 72:12]
  wire [3:0] intpend_w_prior_en_31 = _T_1560 & intpriority_reg_inv_31; // @[pic_ctrl.scala 161:130]
  wire [7:0] _T_1564 = 8'hff; // @[Bitwise.scala 72:12]
  wire [3:0] level_intpend_w_prior_en_0_0 = 4'h0; // @[pic_ctrl.scala 213:40 pic_ctrl.scala 217:38 pic_ctrl.scala 220:33]
  wire [3:0] _T_1441 = intpend_w_prior_en_1; // @[pic_ctrl.scala 70:42 pic_ctrl.scala 161:64]
  wire [3:0] level_intpend_w_prior_en_0_1 = intpend_w_prior_en_1; // @[pic_ctrl.scala 213:40 pic_ctrl.scala 217:38 pic_ctrl.scala 220:33]
  wire  _T_1566 = intpriority_reg_0 < _T_1441; // @[pic_ctrl.scala 27:20]
  wire [7:0] intpend_id_1 = 8'h1; // @[pic_ctrl.scala 71:42 pic_ctrl.scala 162:56]
  wire [7:0] level_intpend_id_0_1 = 8'h1; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30 pic_ctrl.scala 221:33]
  wire [7:0] intpend_id_0 = 8'h0; // @[pic_ctrl.scala 71:42 pic_ctrl.scala 162:56]
  wire [7:0] level_intpend_id_0_0 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30 pic_ctrl.scala 221:33]
  wire [7:0] out_id = _T_1566 ? intpend_id_1 : intpend_id_0; // @[pic_ctrl.scala 27:9]
  wire [3:0] out_priority = _T_1566 ? _T_1441 : intpriority_reg_0; // @[pic_ctrl.scala 27:49]
  wire [3:0] _T_1445 = intpend_w_prior_en_2; // @[pic_ctrl.scala 70:42 pic_ctrl.scala 161:64]
  wire [3:0] level_intpend_w_prior_en_0_2 = intpend_w_prior_en_2; // @[pic_ctrl.scala 213:40 pic_ctrl.scala 217:38 pic_ctrl.scala 220:33]
  wire [3:0] _T_1449 = intpend_w_prior_en_3; // @[pic_ctrl.scala 70:42 pic_ctrl.scala 161:64]
  wire [3:0] level_intpend_w_prior_en_0_3 = intpend_w_prior_en_3; // @[pic_ctrl.scala 213:40 pic_ctrl.scala 217:38 pic_ctrl.scala 220:33]
  wire  _T_1568 = _T_1445 < _T_1449; // @[pic_ctrl.scala 27:20]
  wire [7:0] intpend_id_3 = 8'h3; // @[pic_ctrl.scala 71:42 pic_ctrl.scala 162:56]
  wire [7:0] level_intpend_id_0_3 = 8'h3; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30 pic_ctrl.scala 221:33]
  wire [7:0] intpend_id_2 = 8'h2; // @[pic_ctrl.scala 71:42 pic_ctrl.scala 162:56]
  wire [7:0] level_intpend_id_0_2 = 8'h2; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30 pic_ctrl.scala 221:33]
  wire [7:0] out_id_1 = _T_1568 ? intpend_id_3 : intpend_id_2; // @[pic_ctrl.scala 27:9]
  wire [3:0] out_priority_1 = _T_1568 ? _T_1449 : _T_1445; // @[pic_ctrl.scala 27:49]
  wire [3:0] _T_1453 = intpend_w_prior_en_4; // @[pic_ctrl.scala 70:42 pic_ctrl.scala 161:64]
  wire [3:0] level_intpend_w_prior_en_0_4 = intpend_w_prior_en_4; // @[pic_ctrl.scala 213:40 pic_ctrl.scala 217:38 pic_ctrl.scala 220:33]
  wire [3:0] _T_1457 = intpend_w_prior_en_5; // @[pic_ctrl.scala 70:42 pic_ctrl.scala 161:64]
  wire [3:0] level_intpend_w_prior_en_0_5 = intpend_w_prior_en_5; // @[pic_ctrl.scala 213:40 pic_ctrl.scala 217:38 pic_ctrl.scala 220:33]
  wire  _T_1570 = _T_1453 < _T_1457; // @[pic_ctrl.scala 27:20]
  wire [7:0] intpend_id_5 = 8'h5; // @[pic_ctrl.scala 71:42 pic_ctrl.scala 162:56]
  wire [7:0] level_intpend_id_0_5 = 8'h5; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30 pic_ctrl.scala 221:33]
  wire [7:0] intpend_id_4 = 8'h4; // @[pic_ctrl.scala 71:42 pic_ctrl.scala 162:56]
  wire [7:0] level_intpend_id_0_4 = 8'h4; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30 pic_ctrl.scala 221:33]
  wire [7:0] out_id_2 = _T_1570 ? intpend_id_5 : intpend_id_4; // @[pic_ctrl.scala 27:9]
  wire [3:0] out_priority_2 = _T_1570 ? _T_1457 : _T_1453; // @[pic_ctrl.scala 27:49]
  wire [3:0] _T_1461 = intpend_w_prior_en_6; // @[pic_ctrl.scala 70:42 pic_ctrl.scala 161:64]
  wire [3:0] level_intpend_w_prior_en_0_6 = intpend_w_prior_en_6; // @[pic_ctrl.scala 213:40 pic_ctrl.scala 217:38 pic_ctrl.scala 220:33]
  wire [3:0] _T_1465 = intpend_w_prior_en_7; // @[pic_ctrl.scala 70:42 pic_ctrl.scala 161:64]
  wire [3:0] level_intpend_w_prior_en_0_7 = intpend_w_prior_en_7; // @[pic_ctrl.scala 213:40 pic_ctrl.scala 217:38 pic_ctrl.scala 220:33]
  wire  _T_1572 = _T_1461 < _T_1465; // @[pic_ctrl.scala 27:20]
  wire [7:0] intpend_id_7 = 8'h7; // @[pic_ctrl.scala 71:42 pic_ctrl.scala 162:56]
  wire [7:0] level_intpend_id_0_7 = 8'h7; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30 pic_ctrl.scala 221:33]
  wire [7:0] intpend_id_6 = 8'h6; // @[pic_ctrl.scala 71:42 pic_ctrl.scala 162:56]
  wire [7:0] level_intpend_id_0_6 = 8'h6; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30 pic_ctrl.scala 221:33]
  wire [7:0] out_id_3 = _T_1572 ? intpend_id_7 : intpend_id_6; // @[pic_ctrl.scala 27:9]
  wire [3:0] out_priority_3 = _T_1572 ? _T_1465 : _T_1461; // @[pic_ctrl.scala 27:49]
  wire [3:0] _T_1469 = intpend_w_prior_en_8; // @[pic_ctrl.scala 70:42 pic_ctrl.scala 161:64]
  wire [3:0] level_intpend_w_prior_en_0_8 = intpend_w_prior_en_8; // @[pic_ctrl.scala 213:40 pic_ctrl.scala 217:38 pic_ctrl.scala 220:33]
  wire [3:0] _T_1473 = intpend_w_prior_en_9; // @[pic_ctrl.scala 70:42 pic_ctrl.scala 161:64]
  wire [3:0] level_intpend_w_prior_en_0_9 = intpend_w_prior_en_9; // @[pic_ctrl.scala 213:40 pic_ctrl.scala 217:38 pic_ctrl.scala 220:33]
  wire  _T_1574 = _T_1469 < _T_1473; // @[pic_ctrl.scala 27:20]
  wire [7:0] intpend_id_9 = 8'h9; // @[pic_ctrl.scala 71:42 pic_ctrl.scala 162:56]
  wire [7:0] level_intpend_id_0_9 = 8'h9; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30 pic_ctrl.scala 221:33]
  wire [7:0] intpend_id_8 = 8'h8; // @[pic_ctrl.scala 71:42 pic_ctrl.scala 162:56]
  wire [7:0] level_intpend_id_0_8 = 8'h8; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30 pic_ctrl.scala 221:33]
  wire [7:0] out_id_4 = _T_1574 ? intpend_id_9 : intpend_id_8; // @[pic_ctrl.scala 27:9]
  wire [3:0] out_priority_4 = _T_1574 ? _T_1473 : _T_1469; // @[pic_ctrl.scala 27:49]
  wire [3:0] _T_1477 = intpend_w_prior_en_10; // @[pic_ctrl.scala 70:42 pic_ctrl.scala 161:64]
  wire [3:0] level_intpend_w_prior_en_0_10 = intpend_w_prior_en_10; // @[pic_ctrl.scala 213:40 pic_ctrl.scala 217:38 pic_ctrl.scala 220:33]
  wire [3:0] _T_1481 = intpend_w_prior_en_11; // @[pic_ctrl.scala 70:42 pic_ctrl.scala 161:64]
  wire [3:0] level_intpend_w_prior_en_0_11 = intpend_w_prior_en_11; // @[pic_ctrl.scala 213:40 pic_ctrl.scala 217:38 pic_ctrl.scala 220:33]
  wire  _T_1576 = _T_1477 < _T_1481; // @[pic_ctrl.scala 27:20]
  wire [7:0] intpend_id_11 = 8'hb; // @[pic_ctrl.scala 71:42 pic_ctrl.scala 162:56]
  wire [7:0] level_intpend_id_0_11 = 8'hb; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30 pic_ctrl.scala 221:33]
  wire [7:0] intpend_id_10 = 8'ha; // @[pic_ctrl.scala 71:42 pic_ctrl.scala 162:56]
  wire [7:0] level_intpend_id_0_10 = 8'ha; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30 pic_ctrl.scala 221:33]
  wire [7:0] out_id_5 = _T_1576 ? intpend_id_11 : intpend_id_10; // @[pic_ctrl.scala 27:9]
  wire [3:0] out_priority_5 = _T_1576 ? _T_1481 : _T_1477; // @[pic_ctrl.scala 27:49]
  wire [3:0] _T_1485 = intpend_w_prior_en_12; // @[pic_ctrl.scala 70:42 pic_ctrl.scala 161:64]
  wire [3:0] level_intpend_w_prior_en_0_12 = intpend_w_prior_en_12; // @[pic_ctrl.scala 213:40 pic_ctrl.scala 217:38 pic_ctrl.scala 220:33]
  wire [3:0] _T_1489 = intpend_w_prior_en_13; // @[pic_ctrl.scala 70:42 pic_ctrl.scala 161:64]
  wire [3:0] level_intpend_w_prior_en_0_13 = intpend_w_prior_en_13; // @[pic_ctrl.scala 213:40 pic_ctrl.scala 217:38 pic_ctrl.scala 220:33]
  wire  _T_1578 = _T_1485 < _T_1489; // @[pic_ctrl.scala 27:20]
  wire [7:0] intpend_id_13 = 8'hd; // @[pic_ctrl.scala 71:42 pic_ctrl.scala 162:56]
  wire [7:0] level_intpend_id_0_13 = 8'hd; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30 pic_ctrl.scala 221:33]
  wire [7:0] intpend_id_12 = 8'hc; // @[pic_ctrl.scala 71:42 pic_ctrl.scala 162:56]
  wire [7:0] level_intpend_id_0_12 = 8'hc; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30 pic_ctrl.scala 221:33]
  wire [7:0] out_id_6 = _T_1578 ? intpend_id_13 : intpend_id_12; // @[pic_ctrl.scala 27:9]
  wire [3:0] out_priority_6 = _T_1578 ? _T_1489 : _T_1485; // @[pic_ctrl.scala 27:49]
  wire [3:0] _T_1493 = intpend_w_prior_en_14; // @[pic_ctrl.scala 70:42 pic_ctrl.scala 161:64]
  wire [3:0] level_intpend_w_prior_en_0_14 = intpend_w_prior_en_14; // @[pic_ctrl.scala 213:40 pic_ctrl.scala 217:38 pic_ctrl.scala 220:33]
  wire [3:0] _T_1497 = intpend_w_prior_en_15; // @[pic_ctrl.scala 70:42 pic_ctrl.scala 161:64]
  wire [3:0] level_intpend_w_prior_en_0_15 = intpend_w_prior_en_15; // @[pic_ctrl.scala 213:40 pic_ctrl.scala 217:38 pic_ctrl.scala 220:33]
  wire  _T_1580 = _T_1493 < _T_1497; // @[pic_ctrl.scala 27:20]
  wire [7:0] intpend_id_15 = 8'hf; // @[pic_ctrl.scala 71:42 pic_ctrl.scala 162:56]
  wire [7:0] level_intpend_id_0_15 = 8'hf; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30 pic_ctrl.scala 221:33]
  wire [7:0] intpend_id_14 = 8'he; // @[pic_ctrl.scala 71:42 pic_ctrl.scala 162:56]
  wire [7:0] level_intpend_id_0_14 = 8'he; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30 pic_ctrl.scala 221:33]
  wire [7:0] out_id_7 = _T_1580 ? intpend_id_15 : intpend_id_14; // @[pic_ctrl.scala 27:9]
  wire [3:0] out_priority_7 = _T_1580 ? _T_1497 : _T_1493; // @[pic_ctrl.scala 27:49]
  wire [3:0] _T_1501 = intpend_w_prior_en_16; // @[pic_ctrl.scala 70:42 pic_ctrl.scala 161:64]
  wire [3:0] level_intpend_w_prior_en_0_16 = intpend_w_prior_en_16; // @[pic_ctrl.scala 213:40 pic_ctrl.scala 217:38 pic_ctrl.scala 220:33]
  wire [3:0] _T_1505 = intpend_w_prior_en_17; // @[pic_ctrl.scala 70:42 pic_ctrl.scala 161:64]
  wire [3:0] level_intpend_w_prior_en_0_17 = intpend_w_prior_en_17; // @[pic_ctrl.scala 213:40 pic_ctrl.scala 217:38 pic_ctrl.scala 220:33]
  wire  _T_1582 = _T_1501 < _T_1505; // @[pic_ctrl.scala 27:20]
  wire [7:0] intpend_id_17 = 8'h11; // @[pic_ctrl.scala 71:42 pic_ctrl.scala 162:56]
  wire [7:0] level_intpend_id_0_17 = 8'h11; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30 pic_ctrl.scala 221:33]
  wire [7:0] intpend_id_16 = 8'h10; // @[pic_ctrl.scala 71:42 pic_ctrl.scala 162:56]
  wire [7:0] level_intpend_id_0_16 = 8'h10; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30 pic_ctrl.scala 221:33]
  wire [7:0] out_id_8 = _T_1582 ? intpend_id_17 : intpend_id_16; // @[pic_ctrl.scala 27:9]
  wire [3:0] out_priority_8 = _T_1582 ? _T_1505 : _T_1501; // @[pic_ctrl.scala 27:49]
  wire [3:0] _T_1509 = intpend_w_prior_en_18; // @[pic_ctrl.scala 70:42 pic_ctrl.scala 161:64]
  wire [3:0] level_intpend_w_prior_en_0_18 = intpend_w_prior_en_18; // @[pic_ctrl.scala 213:40 pic_ctrl.scala 217:38 pic_ctrl.scala 220:33]
  wire [3:0] _T_1513 = intpend_w_prior_en_19; // @[pic_ctrl.scala 70:42 pic_ctrl.scala 161:64]
  wire [3:0] level_intpend_w_prior_en_0_19 = intpend_w_prior_en_19; // @[pic_ctrl.scala 213:40 pic_ctrl.scala 217:38 pic_ctrl.scala 220:33]
  wire  _T_1584 = _T_1509 < _T_1513; // @[pic_ctrl.scala 27:20]
  wire [7:0] intpend_id_19 = 8'h13; // @[pic_ctrl.scala 71:42 pic_ctrl.scala 162:56]
  wire [7:0] level_intpend_id_0_19 = 8'h13; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30 pic_ctrl.scala 221:33]
  wire [7:0] intpend_id_18 = 8'h12; // @[pic_ctrl.scala 71:42 pic_ctrl.scala 162:56]
  wire [7:0] level_intpend_id_0_18 = 8'h12; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30 pic_ctrl.scala 221:33]
  wire [7:0] out_id_9 = _T_1584 ? intpend_id_19 : intpend_id_18; // @[pic_ctrl.scala 27:9]
  wire [3:0] out_priority_9 = _T_1584 ? _T_1513 : _T_1509; // @[pic_ctrl.scala 27:49]
  wire [3:0] _T_1517 = intpend_w_prior_en_20; // @[pic_ctrl.scala 70:42 pic_ctrl.scala 161:64]
  wire [3:0] level_intpend_w_prior_en_0_20 = intpend_w_prior_en_20; // @[pic_ctrl.scala 213:40 pic_ctrl.scala 217:38 pic_ctrl.scala 220:33]
  wire [3:0] _T_1521 = intpend_w_prior_en_21; // @[pic_ctrl.scala 70:42 pic_ctrl.scala 161:64]
  wire [3:0] level_intpend_w_prior_en_0_21 = intpend_w_prior_en_21; // @[pic_ctrl.scala 213:40 pic_ctrl.scala 217:38 pic_ctrl.scala 220:33]
  wire  _T_1586 = _T_1517 < _T_1521; // @[pic_ctrl.scala 27:20]
  wire [7:0] intpend_id_21 = 8'h15; // @[pic_ctrl.scala 71:42 pic_ctrl.scala 162:56]
  wire [7:0] level_intpend_id_0_21 = 8'h15; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30 pic_ctrl.scala 221:33]
  wire [7:0] intpend_id_20 = 8'h14; // @[pic_ctrl.scala 71:42 pic_ctrl.scala 162:56]
  wire [7:0] level_intpend_id_0_20 = 8'h14; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30 pic_ctrl.scala 221:33]
  wire [7:0] out_id_10 = _T_1586 ? intpend_id_21 : intpend_id_20; // @[pic_ctrl.scala 27:9]
  wire [3:0] out_priority_10 = _T_1586 ? _T_1521 : _T_1517; // @[pic_ctrl.scala 27:49]
  wire [3:0] _T_1525 = intpend_w_prior_en_22; // @[pic_ctrl.scala 70:42 pic_ctrl.scala 161:64]
  wire [3:0] level_intpend_w_prior_en_0_22 = intpend_w_prior_en_22; // @[pic_ctrl.scala 213:40 pic_ctrl.scala 217:38 pic_ctrl.scala 220:33]
  wire [3:0] _T_1529 = intpend_w_prior_en_23; // @[pic_ctrl.scala 70:42 pic_ctrl.scala 161:64]
  wire [3:0] level_intpend_w_prior_en_0_23 = intpend_w_prior_en_23; // @[pic_ctrl.scala 213:40 pic_ctrl.scala 217:38 pic_ctrl.scala 220:33]
  wire  _T_1588 = _T_1525 < _T_1529; // @[pic_ctrl.scala 27:20]
  wire [7:0] intpend_id_23 = 8'h17; // @[pic_ctrl.scala 71:42 pic_ctrl.scala 162:56]
  wire [7:0] level_intpend_id_0_23 = 8'h17; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30 pic_ctrl.scala 221:33]
  wire [7:0] intpend_id_22 = 8'h16; // @[pic_ctrl.scala 71:42 pic_ctrl.scala 162:56]
  wire [7:0] level_intpend_id_0_22 = 8'h16; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30 pic_ctrl.scala 221:33]
  wire [7:0] out_id_11 = _T_1588 ? intpend_id_23 : intpend_id_22; // @[pic_ctrl.scala 27:9]
  wire [3:0] out_priority_11 = _T_1588 ? _T_1529 : _T_1525; // @[pic_ctrl.scala 27:49]
  wire [3:0] _T_1533 = intpend_w_prior_en_24; // @[pic_ctrl.scala 70:42 pic_ctrl.scala 161:64]
  wire [3:0] level_intpend_w_prior_en_0_24 = intpend_w_prior_en_24; // @[pic_ctrl.scala 213:40 pic_ctrl.scala 217:38 pic_ctrl.scala 220:33]
  wire [3:0] _T_1537 = intpend_w_prior_en_25; // @[pic_ctrl.scala 70:42 pic_ctrl.scala 161:64]
  wire [3:0] level_intpend_w_prior_en_0_25 = intpend_w_prior_en_25; // @[pic_ctrl.scala 213:40 pic_ctrl.scala 217:38 pic_ctrl.scala 220:33]
  wire  _T_1590 = _T_1533 < _T_1537; // @[pic_ctrl.scala 27:20]
  wire [7:0] intpend_id_25 = 8'h19; // @[pic_ctrl.scala 71:42 pic_ctrl.scala 162:56]
  wire [7:0] level_intpend_id_0_25 = 8'h19; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30 pic_ctrl.scala 221:33]
  wire [7:0] intpend_id_24 = 8'h18; // @[pic_ctrl.scala 71:42 pic_ctrl.scala 162:56]
  wire [7:0] level_intpend_id_0_24 = 8'h18; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30 pic_ctrl.scala 221:33]
  wire [7:0] out_id_12 = _T_1590 ? intpend_id_25 : intpend_id_24; // @[pic_ctrl.scala 27:9]
  wire [3:0] out_priority_12 = _T_1590 ? _T_1537 : _T_1533; // @[pic_ctrl.scala 27:49]
  wire [3:0] _T_1541 = intpend_w_prior_en_26; // @[pic_ctrl.scala 70:42 pic_ctrl.scala 161:64]
  wire [3:0] level_intpend_w_prior_en_0_26 = intpend_w_prior_en_26; // @[pic_ctrl.scala 213:40 pic_ctrl.scala 217:38 pic_ctrl.scala 220:33]
  wire [3:0] _T_1545 = intpend_w_prior_en_27; // @[pic_ctrl.scala 70:42 pic_ctrl.scala 161:64]
  wire [3:0] level_intpend_w_prior_en_0_27 = intpend_w_prior_en_27; // @[pic_ctrl.scala 213:40 pic_ctrl.scala 217:38 pic_ctrl.scala 220:33]
  wire  _T_1592 = _T_1541 < _T_1545; // @[pic_ctrl.scala 27:20]
  wire [7:0] intpend_id_27 = 8'h1b; // @[pic_ctrl.scala 71:42 pic_ctrl.scala 162:56]
  wire [7:0] level_intpend_id_0_27 = 8'h1b; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30 pic_ctrl.scala 221:33]
  wire [7:0] intpend_id_26 = 8'h1a; // @[pic_ctrl.scala 71:42 pic_ctrl.scala 162:56]
  wire [7:0] level_intpend_id_0_26 = 8'h1a; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30 pic_ctrl.scala 221:33]
  wire [7:0] out_id_13 = _T_1592 ? intpend_id_27 : intpend_id_26; // @[pic_ctrl.scala 27:9]
  wire [3:0] out_priority_13 = _T_1592 ? _T_1545 : _T_1541; // @[pic_ctrl.scala 27:49]
  wire [3:0] _T_1549 = intpend_w_prior_en_28; // @[pic_ctrl.scala 70:42 pic_ctrl.scala 161:64]
  wire [3:0] level_intpend_w_prior_en_0_28 = intpend_w_prior_en_28; // @[pic_ctrl.scala 213:40 pic_ctrl.scala 217:38 pic_ctrl.scala 220:33]
  wire [3:0] _T_1553 = intpend_w_prior_en_29; // @[pic_ctrl.scala 70:42 pic_ctrl.scala 161:64]
  wire [3:0] level_intpend_w_prior_en_0_29 = intpend_w_prior_en_29; // @[pic_ctrl.scala 213:40 pic_ctrl.scala 217:38 pic_ctrl.scala 220:33]
  wire  _T_1594 = _T_1549 < _T_1553; // @[pic_ctrl.scala 27:20]
  wire [7:0] intpend_id_29 = 8'h1d; // @[pic_ctrl.scala 71:42 pic_ctrl.scala 162:56]
  wire [7:0] level_intpend_id_0_29 = 8'h1d; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30 pic_ctrl.scala 221:33]
  wire [7:0] intpend_id_28 = 8'h1c; // @[pic_ctrl.scala 71:42 pic_ctrl.scala 162:56]
  wire [7:0] level_intpend_id_0_28 = 8'h1c; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30 pic_ctrl.scala 221:33]
  wire [7:0] out_id_14 = _T_1594 ? intpend_id_29 : intpend_id_28; // @[pic_ctrl.scala 27:9]
  wire [3:0] out_priority_14 = _T_1594 ? _T_1553 : _T_1549; // @[pic_ctrl.scala 27:49]
  wire [3:0] _T_1557 = intpend_w_prior_en_30; // @[pic_ctrl.scala 70:42 pic_ctrl.scala 161:64]
  wire [3:0] level_intpend_w_prior_en_0_30 = intpend_w_prior_en_30; // @[pic_ctrl.scala 213:40 pic_ctrl.scala 217:38 pic_ctrl.scala 220:33]
  wire [3:0] _T_1561 = intpend_w_prior_en_31; // @[pic_ctrl.scala 70:42 pic_ctrl.scala 161:64]
  wire [3:0] level_intpend_w_prior_en_0_31 = intpend_w_prior_en_31; // @[pic_ctrl.scala 213:40 pic_ctrl.scala 217:38 pic_ctrl.scala 220:33]
  wire  _T_1596 = _T_1557 < _T_1561; // @[pic_ctrl.scala 27:20]
  wire [7:0] intpend_id_31 = 8'h1f; // @[pic_ctrl.scala 71:42 pic_ctrl.scala 162:56]
  wire [7:0] level_intpend_id_0_31 = 8'h1f; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30 pic_ctrl.scala 221:33]
  wire [7:0] intpend_id_30 = 8'h1e; // @[pic_ctrl.scala 71:42 pic_ctrl.scala 162:56]
  wire [7:0] level_intpend_id_0_30 = 8'h1e; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30 pic_ctrl.scala 221:33]
  wire [7:0] out_id_15 = _T_1596 ? intpend_id_31 : intpend_id_30; // @[pic_ctrl.scala 27:9]
  wire [3:0] out_priority_15 = _T_1596 ? _T_1561 : _T_1557; // @[pic_ctrl.scala 27:49]
  wire [3:0] level_intpend_w_prior_en_0_32 = 4'h0; // @[pic_ctrl.scala 213:40 pic_ctrl.scala 217:38 pic_ctrl.scala 220:33]
  wire [3:0] level_intpend_w_prior_en_0_33 = 4'h0; // @[pic_ctrl.scala 213:40 pic_ctrl.scala 217:38 pic_ctrl.scala 220:33]
  wire  _T_1598 = intpriority_reg_0 < intpriority_reg_0; // @[pic_ctrl.scala 27:20]
  wire [7:0] level_intpend_id_0_33 = 8'hff; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30 pic_ctrl.scala 221:33]
  wire [7:0] level_intpend_id_0_32 = 8'hff; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30 pic_ctrl.scala 221:33]
  wire [7:0] out_id_16 = _T_1598 ? _T_1564 : _T_1564; // @[pic_ctrl.scala 27:9]
  wire  _T_1600 = out_priority < out_priority_1; // @[pic_ctrl.scala 27:20]
  wire [7:0] level_intpend_id_1_1 = out_id_1; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30 pic_ctrl.scala 232:41]
  wire [7:0] level_intpend_id_1_0 = out_id; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30 pic_ctrl.scala 232:41]
  wire [7:0] out_id_17 = _T_1600 ? level_intpend_id_1_1 : level_intpend_id_1_0; // @[pic_ctrl.scala 27:9]
  wire [3:0] out_priority_17 = _T_1600 ? out_priority_1 : out_priority; // @[pic_ctrl.scala 27:49]
  wire  _T_1602 = out_priority_2 < out_priority_3; // @[pic_ctrl.scala 27:20]
  wire [7:0] level_intpend_id_1_3 = out_id_3; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30 pic_ctrl.scala 232:41]
  wire [7:0] level_intpend_id_1_2 = out_id_2; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30 pic_ctrl.scala 232:41]
  wire [7:0] out_id_18 = _T_1602 ? level_intpend_id_1_3 : level_intpend_id_1_2; // @[pic_ctrl.scala 27:9]
  wire [3:0] out_priority_18 = _T_1602 ? out_priority_3 : out_priority_2; // @[pic_ctrl.scala 27:49]
  wire  _T_1604 = out_priority_4 < out_priority_5; // @[pic_ctrl.scala 27:20]
  wire [7:0] level_intpend_id_1_5 = out_id_5; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30 pic_ctrl.scala 232:41]
  wire [7:0] level_intpend_id_1_4 = out_id_4; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30 pic_ctrl.scala 232:41]
  wire [7:0] out_id_19 = _T_1604 ? level_intpend_id_1_5 : level_intpend_id_1_4; // @[pic_ctrl.scala 27:9]
  wire [3:0] out_priority_19 = _T_1604 ? out_priority_5 : out_priority_4; // @[pic_ctrl.scala 27:49]
  wire  _T_1606 = out_priority_6 < out_priority_7; // @[pic_ctrl.scala 27:20]
  wire [7:0] level_intpend_id_1_7 = out_id_7; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30 pic_ctrl.scala 232:41]
  wire [7:0] level_intpend_id_1_6 = out_id_6; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30 pic_ctrl.scala 232:41]
  wire [7:0] out_id_20 = _T_1606 ? level_intpend_id_1_7 : level_intpend_id_1_6; // @[pic_ctrl.scala 27:9]
  wire [3:0] out_priority_20 = _T_1606 ? out_priority_7 : out_priority_6; // @[pic_ctrl.scala 27:49]
  wire  _T_1608 = out_priority_8 < out_priority_9; // @[pic_ctrl.scala 27:20]
  wire [7:0] level_intpend_id_1_9 = out_id_9; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30 pic_ctrl.scala 232:41]
  wire [7:0] level_intpend_id_1_8 = out_id_8; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30 pic_ctrl.scala 232:41]
  wire [7:0] out_id_21 = _T_1608 ? level_intpend_id_1_9 : level_intpend_id_1_8; // @[pic_ctrl.scala 27:9]
  wire [3:0] out_priority_21 = _T_1608 ? out_priority_9 : out_priority_8; // @[pic_ctrl.scala 27:49]
  wire  _T_1610 = out_priority_10 < out_priority_11; // @[pic_ctrl.scala 27:20]
  wire [7:0] level_intpend_id_1_11 = out_id_11; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30 pic_ctrl.scala 232:41]
  wire [7:0] level_intpend_id_1_10 = out_id_10; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30 pic_ctrl.scala 232:41]
  wire [7:0] out_id_22 = _T_1610 ? level_intpend_id_1_11 : level_intpend_id_1_10; // @[pic_ctrl.scala 27:9]
  wire [3:0] out_priority_22 = _T_1610 ? out_priority_11 : out_priority_10; // @[pic_ctrl.scala 27:49]
  wire  _T_1612 = out_priority_12 < out_priority_13; // @[pic_ctrl.scala 27:20]
  wire [7:0] level_intpend_id_1_13 = out_id_13; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30 pic_ctrl.scala 232:41]
  wire [7:0] level_intpend_id_1_12 = out_id_12; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30 pic_ctrl.scala 232:41]
  wire [7:0] out_id_23 = _T_1612 ? level_intpend_id_1_13 : level_intpend_id_1_12; // @[pic_ctrl.scala 27:9]
  wire [3:0] out_priority_23 = _T_1612 ? out_priority_13 : out_priority_12; // @[pic_ctrl.scala 27:49]
  wire  _T_1614 = out_priority_14 < out_priority_15; // @[pic_ctrl.scala 27:20]
  wire [7:0] level_intpend_id_1_15 = out_id_15; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30 pic_ctrl.scala 232:41]
  wire [7:0] level_intpend_id_1_14 = out_id_14; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30 pic_ctrl.scala 232:41]
  wire [7:0] out_id_24 = _T_1614 ? level_intpend_id_1_15 : level_intpend_id_1_14; // @[pic_ctrl.scala 27:9]
  wire [3:0] out_priority_24 = _T_1614 ? out_priority_15 : out_priority_14; // @[pic_ctrl.scala 27:49]
  wire [7:0] level_intpend_id_1_17 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30 pic_ctrl.scala 229:44]
  wire [7:0] level_intpend_id_1_16 = out_id_16; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30 pic_ctrl.scala 232:41]
  wire [7:0] out_id_25 = level_intpend_id_1_16; // @[pic_ctrl.scala 27:9]
  wire  _T_1618 = out_priority_17 < out_priority_18; // @[pic_ctrl.scala 27:20]
  wire [7:0] level_intpend_id_2_1 = out_id_18; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30 pic_ctrl.scala 232:41]
  wire [7:0] level_intpend_id_2_0 = out_id_17; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30 pic_ctrl.scala 232:41]
  wire [7:0] out_id_26 = _T_1618 ? level_intpend_id_2_1 : level_intpend_id_2_0; // @[pic_ctrl.scala 27:9]
  wire [3:0] out_priority_26 = _T_1618 ? out_priority_18 : out_priority_17; // @[pic_ctrl.scala 27:49]
  wire  _T_1620 = out_priority_19 < out_priority_20; // @[pic_ctrl.scala 27:20]
  wire [7:0] level_intpend_id_2_3 = out_id_20; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30 pic_ctrl.scala 232:41]
  wire [7:0] level_intpend_id_2_2 = out_id_19; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30 pic_ctrl.scala 232:41]
  wire [7:0] out_id_27 = _T_1620 ? level_intpend_id_2_3 : level_intpend_id_2_2; // @[pic_ctrl.scala 27:9]
  wire [3:0] out_priority_27 = _T_1620 ? out_priority_20 : out_priority_19; // @[pic_ctrl.scala 27:49]
  wire  _T_1622 = out_priority_21 < out_priority_22; // @[pic_ctrl.scala 27:20]
  wire [7:0] level_intpend_id_2_5 = out_id_22; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30 pic_ctrl.scala 232:41]
  wire [7:0] level_intpend_id_2_4 = out_id_21; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30 pic_ctrl.scala 232:41]
  wire [7:0] out_id_28 = _T_1622 ? level_intpend_id_2_5 : level_intpend_id_2_4; // @[pic_ctrl.scala 27:9]
  wire [3:0] out_priority_28 = _T_1622 ? out_priority_22 : out_priority_21; // @[pic_ctrl.scala 27:49]
  wire  _T_1624 = out_priority_23 < out_priority_24; // @[pic_ctrl.scala 27:20]
  wire [7:0] level_intpend_id_2_7 = out_id_24; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30 pic_ctrl.scala 232:41]
  wire [7:0] level_intpend_id_2_6 = out_id_23; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30 pic_ctrl.scala 232:41]
  wire [7:0] out_id_29 = _T_1624 ? level_intpend_id_2_7 : level_intpend_id_2_6; // @[pic_ctrl.scala 27:9]
  wire [3:0] out_priority_29 = _T_1624 ? out_priority_24 : out_priority_23; // @[pic_ctrl.scala 27:49]
  wire [7:0] level_intpend_id_2_9 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30 pic_ctrl.scala 229:44]
  wire [7:0] level_intpend_id_2_8 = level_intpend_id_1_16; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30 pic_ctrl.scala 232:41]
  wire [7:0] out_id_30 = out_id_25; // @[pic_ctrl.scala 27:9]
  wire  _T_1628 = out_priority_26 < out_priority_27; // @[pic_ctrl.scala 27:20]
  wire [7:0] level_intpend_id_3_1 = out_id_27; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30 pic_ctrl.scala 232:41]
  wire [7:0] level_intpend_id_3_0 = out_id_26; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30 pic_ctrl.scala 232:41]
  wire [7:0] out_id_31 = _T_1628 ? level_intpend_id_3_1 : level_intpend_id_3_0; // @[pic_ctrl.scala 27:9]
  wire [3:0] out_priority_31 = _T_1628 ? out_priority_27 : out_priority_26; // @[pic_ctrl.scala 27:49]
  wire  _T_1630 = out_priority_28 < out_priority_29; // @[pic_ctrl.scala 27:20]
  wire [7:0] level_intpend_id_3_3 = out_id_29; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30 pic_ctrl.scala 232:41]
  wire [7:0] level_intpend_id_3_2 = out_id_28; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30 pic_ctrl.scala 232:41]
  wire [7:0] out_id_32 = _T_1630 ? level_intpend_id_3_3 : level_intpend_id_3_2; // @[pic_ctrl.scala 27:9]
  wire [3:0] out_priority_32 = _T_1630 ? out_priority_29 : out_priority_28; // @[pic_ctrl.scala 27:49]
  wire [7:0] level_intpend_id_3_5 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30 pic_ctrl.scala 229:44]
  wire [7:0] level_intpend_id_3_4 = out_id_25; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30 pic_ctrl.scala 232:41]
  wire [7:0] out_id_33 = out_id_30; // @[pic_ctrl.scala 27:9]
  wire  _T_1634 = out_priority_31 < out_priority_32; // @[pic_ctrl.scala 27:20]
  wire [7:0] level_intpend_id_4_1 = out_id_32; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30 pic_ctrl.scala 232:41]
  wire [7:0] level_intpend_id_4_0 = out_id_31; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30 pic_ctrl.scala 232:41]
  wire [7:0] out_id_34 = _T_1634 ? level_intpend_id_4_1 : level_intpend_id_4_0; // @[pic_ctrl.scala 27:9]
  wire [3:0] out_priority_34 = _T_1634 ? out_priority_32 : out_priority_31; // @[pic_ctrl.scala 27:49]
  wire [7:0] level_intpend_id_4_3 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30 pic_ctrl.scala 229:44]
  wire [7:0] level_intpend_id_4_2 = out_id_30; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30 pic_ctrl.scala 232:41]
  wire  config_reg_we = waddr_config_pic_match & picm_wren_ff; // @[pic_ctrl.scala 249:47]
  wire  config_reg_re = raddr_config_pic_match & picm_rden_ff; // @[pic_ctrl.scala 250:47]
  wire [3:0] level_intpend_w_prior_en_5_0 = out_priority_34; // @[pic_ctrl.scala 213:40 pic_ctrl.scala 217:38 pic_ctrl.scala 233:41]
  wire [3:0] selected_int_priority = out_priority_34; // @[pic_ctrl.scala 237:29]
  wire [3:0] _T_1641 = ~level_intpend_w_prior_en_5_0; // @[pic_ctrl.scala 261:38]
  wire [3:0] pl_in_q = config_reg ? _T_1641 : level_intpend_w_prior_en_5_0; // @[pic_ctrl.scala 261:20]
  reg [7:0] _T_1642; // @[pic_ctrl.scala 262:59]
  reg [3:0] _T_1643; // @[pic_ctrl.scala 263:54]
  wire [3:0] _T_1645 = ~io_dec_pic_dec_tlu_meipt; // @[pic_ctrl.scala 264:40]
  wire [3:0] meipt_inv = config_reg ? _T_1645 : io_dec_pic_dec_tlu_meipt; // @[pic_ctrl.scala 264:22]
  wire [3:0] _T_1647 = ~io_dec_pic_dec_tlu_meicurpl; // @[pic_ctrl.scala 265:43]
  wire [3:0] meicurpl_inv = config_reg ? _T_1647 : io_dec_pic_dec_tlu_meicurpl; // @[pic_ctrl.scala 265:25]
  wire  _T_1648 = level_intpend_w_prior_en_5_0 > meipt_inv; // @[pic_ctrl.scala 266:47]
  wire  _T_1649 = level_intpend_w_prior_en_5_0 > meicurpl_inv; // @[pic_ctrl.scala 266:86]
  reg  _T_1650; // @[pic_ctrl.scala 267:58]
  wire [3:0] maxint = config_reg ? 4'h0 : 4'hf; // @[pic_ctrl.scala 268:19]
  reg  _T_1652; // @[pic_ctrl.scala 270:56]
  wire  intpend_reg_read = addr_intpend_base_match & picm_rden_ff; // @[pic_ctrl.scala 276:60]
  wire [9:0] _T_1662 = {extintsrc_req_gw_31,extintsrc_req_gw_30,extintsrc_req_gw_29,extintsrc_req_gw_28,extintsrc_req_gw_27,extintsrc_req_gw_26,extintsrc_req_gw_25,extintsrc_req_gw_24,extintsrc_req_gw_23,extintsrc_req_gw_22}; // @[Cat.scala 29:58]
  wire [18:0] _T_1671 = {_T_1662,extintsrc_req_gw_21,extintsrc_req_gw_20,extintsrc_req_gw_19,extintsrc_req_gw_18,extintsrc_req_gw_17,extintsrc_req_gw_16,extintsrc_req_gw_15,extintsrc_req_gw_14,extintsrc_req_gw_13}; // @[Cat.scala 29:58]
  wire [27:0] _T_1680 = {_T_1671,extintsrc_req_gw_12,extintsrc_req_gw_11,extintsrc_req_gw_10,extintsrc_req_gw_9,extintsrc_req_gw_8,extintsrc_req_gw_7,extintsrc_req_gw_6,extintsrc_req_gw_5,extintsrc_req_gw_4}; // @[Cat.scala 29:58]
  wire [63:0] intpend_reg_extended = {32'h0,_T_1680,extintsrc_req_gw_3,extintsrc_req_gw_2,extintsrc_req_gw_1,1'h0}; // @[Cat.scala 29:58]
  wire  _T_1687 = picm_raddr_ff[5:2] == 4'h0; // @[pic_ctrl.scala 284:107]
  wire  _T_1688 = intpend_reg_read & _T_1687; // @[pic_ctrl.scala 284:85]
  wire [31:0] _T_1690 = _T_1688 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] intpend_rd_part_out_0 = _T_1690 & intpend_reg_extended[31:0]; // @[pic_ctrl.scala 284:123]
  wire  _T_1694 = picm_raddr_ff[5:2] == 4'h1; // @[pic_ctrl.scala 284:107]
  wire  _T_1695 = intpend_reg_read & _T_1694; // @[pic_ctrl.scala 284:85]
  wire [31:0] _T_1697 = _T_1695 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] intpend_rd_part_out_1 = _T_1697 & intpend_reg_extended[63:32]; // @[pic_ctrl.scala 284:123]
  wire [31:0] intpend_rd_out = intpend_rd_part_out_0 | intpend_rd_part_out_1; // @[pic_ctrl.scala 285:58]
  wire  _T_1732 = intenable_reg_re_31 & intenable_reg_31; // @[Mux.scala 98:16]
  wire  _T_1733 = intenable_reg_re_30 ? intenable_reg_30 : _T_1732; // @[Mux.scala 98:16]
  wire  _T_1734 = intenable_reg_re_29 ? intenable_reg_29 : _T_1733; // @[Mux.scala 98:16]
  wire  _T_1735 = intenable_reg_re_28 ? intenable_reg_28 : _T_1734; // @[Mux.scala 98:16]
  wire  _T_1736 = intenable_reg_re_27 ? intenable_reg_27 : _T_1735; // @[Mux.scala 98:16]
  wire  _T_1737 = intenable_reg_re_26 ? intenable_reg_26 : _T_1736; // @[Mux.scala 98:16]
  wire  _T_1738 = intenable_reg_re_25 ? intenable_reg_25 : _T_1737; // @[Mux.scala 98:16]
  wire  _T_1739 = intenable_reg_re_24 ? intenable_reg_24 : _T_1738; // @[Mux.scala 98:16]
  wire  _T_1740 = intenable_reg_re_23 ? intenable_reg_23 : _T_1739; // @[Mux.scala 98:16]
  wire  _T_1741 = intenable_reg_re_22 ? intenable_reg_22 : _T_1740; // @[Mux.scala 98:16]
  wire  _T_1742 = intenable_reg_re_21 ? intenable_reg_21 : _T_1741; // @[Mux.scala 98:16]
  wire  _T_1743 = intenable_reg_re_20 ? intenable_reg_20 : _T_1742; // @[Mux.scala 98:16]
  wire  _T_1744 = intenable_reg_re_19 ? intenable_reg_19 : _T_1743; // @[Mux.scala 98:16]
  wire  _T_1745 = intenable_reg_re_18 ? intenable_reg_18 : _T_1744; // @[Mux.scala 98:16]
  wire  _T_1746 = intenable_reg_re_17 ? intenable_reg_17 : _T_1745; // @[Mux.scala 98:16]
  wire  _T_1747 = intenable_reg_re_16 ? intenable_reg_16 : _T_1746; // @[Mux.scala 98:16]
  wire  _T_1748 = intenable_reg_re_15 ? intenable_reg_15 : _T_1747; // @[Mux.scala 98:16]
  wire  _T_1749 = intenable_reg_re_14 ? intenable_reg_14 : _T_1748; // @[Mux.scala 98:16]
  wire  _T_1750 = intenable_reg_re_13 ? intenable_reg_13 : _T_1749; // @[Mux.scala 98:16]
  wire  _T_1751 = intenable_reg_re_12 ? intenable_reg_12 : _T_1750; // @[Mux.scala 98:16]
  wire  _T_1752 = intenable_reg_re_11 ? intenable_reg_11 : _T_1751; // @[Mux.scala 98:16]
  wire  _T_1753 = intenable_reg_re_10 ? intenable_reg_10 : _T_1752; // @[Mux.scala 98:16]
  wire  _T_1754 = intenable_reg_re_9 ? intenable_reg_9 : _T_1753; // @[Mux.scala 98:16]
  wire  _T_1755 = intenable_reg_re_8 ? intenable_reg_8 : _T_1754; // @[Mux.scala 98:16]
  wire  _T_1756 = intenable_reg_re_7 ? intenable_reg_7 : _T_1755; // @[Mux.scala 98:16]
  wire  _T_1757 = intenable_reg_re_6 ? intenable_reg_6 : _T_1756; // @[Mux.scala 98:16]
  wire  _T_1758 = intenable_reg_re_5 ? intenable_reg_5 : _T_1757; // @[Mux.scala 98:16]
  wire  _T_1759 = intenable_reg_re_4 ? intenable_reg_4 : _T_1758; // @[Mux.scala 98:16]
  wire  _T_1760 = intenable_reg_re_3 ? intenable_reg_3 : _T_1759; // @[Mux.scala 98:16]
  wire  _T_1761 = intenable_reg_re_2 ? intenable_reg_2 : _T_1760; // @[Mux.scala 98:16]
  wire  intenable_rd_out = intenable_reg_re_1 ? intenable_reg_1 : _T_1761; // @[Mux.scala 98:16]
  wire [3:0] _T_1794 = intpriority_reg_re_31 ? intpriority_reg_31 : 4'h0; // @[Mux.scala 98:16]
  wire [3:0] _T_1795 = intpriority_reg_re_30 ? intpriority_reg_30 : _T_1794; // @[Mux.scala 98:16]
  wire [3:0] _T_1796 = intpriority_reg_re_29 ? intpriority_reg_29 : _T_1795; // @[Mux.scala 98:16]
  wire [3:0] _T_1797 = intpriority_reg_re_28 ? intpriority_reg_28 : _T_1796; // @[Mux.scala 98:16]
  wire [3:0] _T_1798 = intpriority_reg_re_27 ? intpriority_reg_27 : _T_1797; // @[Mux.scala 98:16]
  wire [3:0] _T_1799 = intpriority_reg_re_26 ? intpriority_reg_26 : _T_1798; // @[Mux.scala 98:16]
  wire [3:0] _T_1800 = intpriority_reg_re_25 ? intpriority_reg_25 : _T_1799; // @[Mux.scala 98:16]
  wire [3:0] _T_1801 = intpriority_reg_re_24 ? intpriority_reg_24 : _T_1800; // @[Mux.scala 98:16]
  wire [3:0] _T_1802 = intpriority_reg_re_23 ? intpriority_reg_23 : _T_1801; // @[Mux.scala 98:16]
  wire [3:0] _T_1803 = intpriority_reg_re_22 ? intpriority_reg_22 : _T_1802; // @[Mux.scala 98:16]
  wire [3:0] _T_1804 = intpriority_reg_re_21 ? intpriority_reg_21 : _T_1803; // @[Mux.scala 98:16]
  wire [3:0] _T_1805 = intpriority_reg_re_20 ? intpriority_reg_20 : _T_1804; // @[Mux.scala 98:16]
  wire [3:0] _T_1806 = intpriority_reg_re_19 ? intpriority_reg_19 : _T_1805; // @[Mux.scala 98:16]
  wire [3:0] _T_1807 = intpriority_reg_re_18 ? intpriority_reg_18 : _T_1806; // @[Mux.scala 98:16]
  wire [3:0] _T_1808 = intpriority_reg_re_17 ? intpriority_reg_17 : _T_1807; // @[Mux.scala 98:16]
  wire [3:0] _T_1809 = intpriority_reg_re_16 ? intpriority_reg_16 : _T_1808; // @[Mux.scala 98:16]
  wire [3:0] _T_1810 = intpriority_reg_re_15 ? intpriority_reg_15 : _T_1809; // @[Mux.scala 98:16]
  wire [3:0] _T_1811 = intpriority_reg_re_14 ? intpriority_reg_14 : _T_1810; // @[Mux.scala 98:16]
  wire [3:0] _T_1812 = intpriority_reg_re_13 ? intpriority_reg_13 : _T_1811; // @[Mux.scala 98:16]
  wire [3:0] _T_1813 = intpriority_reg_re_12 ? intpriority_reg_12 : _T_1812; // @[Mux.scala 98:16]
  wire [3:0] _T_1814 = intpriority_reg_re_11 ? intpriority_reg_11 : _T_1813; // @[Mux.scala 98:16]
  wire [3:0] _T_1815 = intpriority_reg_re_10 ? intpriority_reg_10 : _T_1814; // @[Mux.scala 98:16]
  wire [3:0] _T_1816 = intpriority_reg_re_9 ? intpriority_reg_9 : _T_1815; // @[Mux.scala 98:16]
  wire [3:0] _T_1817 = intpriority_reg_re_8 ? intpriority_reg_8 : _T_1816; // @[Mux.scala 98:16]
  wire [3:0] _T_1818 = intpriority_reg_re_7 ? intpriority_reg_7 : _T_1817; // @[Mux.scala 98:16]
  wire [3:0] _T_1819 = intpriority_reg_re_6 ? intpriority_reg_6 : _T_1818; // @[Mux.scala 98:16]
  wire [3:0] _T_1820 = intpriority_reg_re_5 ? intpriority_reg_5 : _T_1819; // @[Mux.scala 98:16]
  wire [3:0] _T_1821 = intpriority_reg_re_4 ? intpriority_reg_4 : _T_1820; // @[Mux.scala 98:16]
  wire [3:0] _T_1822 = intpriority_reg_re_3 ? intpriority_reg_3 : _T_1821; // @[Mux.scala 98:16]
  wire [3:0] _T_1823 = intpriority_reg_re_2 ? intpriority_reg_2 : _T_1822; // @[Mux.scala 98:16]
  wire [3:0] intpriority_rd_out = intpriority_reg_re_1 ? intpriority_reg_1 : _T_1823; // @[Mux.scala 98:16]
  wire [1:0] _T_1856 = gw_config_reg_re_31 ? gw_config_reg_31 : 2'h0; // @[Mux.scala 98:16]
  wire [1:0] _T_1857 = gw_config_reg_re_30 ? gw_config_reg_30 : _T_1856; // @[Mux.scala 98:16]
  wire [1:0] _T_1858 = gw_config_reg_re_29 ? gw_config_reg_29 : _T_1857; // @[Mux.scala 98:16]
  wire [1:0] _T_1859 = gw_config_reg_re_28 ? gw_config_reg_28 : _T_1858; // @[Mux.scala 98:16]
  wire [1:0] _T_1860 = gw_config_reg_re_27 ? gw_config_reg_27 : _T_1859; // @[Mux.scala 98:16]
  wire [1:0] _T_1861 = gw_config_reg_re_26 ? gw_config_reg_26 : _T_1860; // @[Mux.scala 98:16]
  wire [1:0] _T_1862 = gw_config_reg_re_25 ? gw_config_reg_25 : _T_1861; // @[Mux.scala 98:16]
  wire [1:0] _T_1863 = gw_config_reg_re_24 ? gw_config_reg_24 : _T_1862; // @[Mux.scala 98:16]
  wire [1:0] _T_1864 = gw_config_reg_re_23 ? gw_config_reg_23 : _T_1863; // @[Mux.scala 98:16]
  wire [1:0] _T_1865 = gw_config_reg_re_22 ? gw_config_reg_22 : _T_1864; // @[Mux.scala 98:16]
  wire [1:0] _T_1866 = gw_config_reg_re_21 ? gw_config_reg_21 : _T_1865; // @[Mux.scala 98:16]
  wire [1:0] _T_1867 = gw_config_reg_re_20 ? gw_config_reg_20 : _T_1866; // @[Mux.scala 98:16]
  wire [1:0] _T_1868 = gw_config_reg_re_19 ? gw_config_reg_19 : _T_1867; // @[Mux.scala 98:16]
  wire [1:0] _T_1869 = gw_config_reg_re_18 ? gw_config_reg_18 : _T_1868; // @[Mux.scala 98:16]
  wire [1:0] _T_1870 = gw_config_reg_re_17 ? gw_config_reg_17 : _T_1869; // @[Mux.scala 98:16]
  wire [1:0] _T_1871 = gw_config_reg_re_16 ? gw_config_reg_16 : _T_1870; // @[Mux.scala 98:16]
  wire [1:0] _T_1872 = gw_config_reg_re_15 ? gw_config_reg_15 : _T_1871; // @[Mux.scala 98:16]
  wire [1:0] _T_1873 = gw_config_reg_re_14 ? gw_config_reg_14 : _T_1872; // @[Mux.scala 98:16]
  wire [1:0] _T_1874 = gw_config_reg_re_13 ? gw_config_reg_13 : _T_1873; // @[Mux.scala 98:16]
  wire [1:0] _T_1875 = gw_config_reg_re_12 ? gw_config_reg_12 : _T_1874; // @[Mux.scala 98:16]
  wire [1:0] _T_1876 = gw_config_reg_re_11 ? gw_config_reg_11 : _T_1875; // @[Mux.scala 98:16]
  wire [1:0] _T_1877 = gw_config_reg_re_10 ? gw_config_reg_10 : _T_1876; // @[Mux.scala 98:16]
  wire [1:0] _T_1878 = gw_config_reg_re_9 ? gw_config_reg_9 : _T_1877; // @[Mux.scala 98:16]
  wire [1:0] _T_1879 = gw_config_reg_re_8 ? gw_config_reg_8 : _T_1878; // @[Mux.scala 98:16]
  wire [1:0] _T_1880 = gw_config_reg_re_7 ? gw_config_reg_7 : _T_1879; // @[Mux.scala 98:16]
  wire [1:0] _T_1881 = gw_config_reg_re_6 ? gw_config_reg_6 : _T_1880; // @[Mux.scala 98:16]
  wire [1:0] _T_1882 = gw_config_reg_re_5 ? gw_config_reg_5 : _T_1881; // @[Mux.scala 98:16]
  wire [1:0] _T_1883 = gw_config_reg_re_4 ? gw_config_reg_4 : _T_1882; // @[Mux.scala 98:16]
  wire [1:0] _T_1884 = gw_config_reg_re_3 ? gw_config_reg_3 : _T_1883; // @[Mux.scala 98:16]
  wire [1:0] _T_1885 = gw_config_reg_re_2 ? gw_config_reg_2 : _T_1884; // @[Mux.scala 98:16]
  wire [1:0] gw_config_rd_out = gw_config_reg_re_1 ? gw_config_reg_1 : _T_1885; // @[Mux.scala 98:16]
  wire [31:0] _T_1890 = {28'h0,intpriority_rd_out}; // @[Cat.scala 29:58]
  wire [31:0] _T_1893 = {31'h0,intenable_rd_out}; // @[Cat.scala 29:58]
  wire [31:0] _T_1896 = {30'h0,gw_config_rd_out}; // @[Cat.scala 29:58]
  wire [31:0] _T_1899 = {31'h0,config_reg}; // @[Cat.scala 29:58]
  wire [14:0] address = picm_raddr_ff[14:0]; // @[pic_ctrl.scala 306:30]
  wire  _T_1939 = 15'h3000 == address; // @[Conditional.scala 37:30]
  wire  _T_1940 = 15'h4004 == address; // @[Conditional.scala 37:30]
  wire  _T_1941 = 15'h4008 == address; // @[Conditional.scala 37:30]
  wire  _T_1942 = 15'h400c == address; // @[Conditional.scala 37:30]
  wire  _T_1943 = 15'h4010 == address; // @[Conditional.scala 37:30]
  wire  _T_1944 = 15'h4014 == address; // @[Conditional.scala 37:30]
  wire  _T_1945 = 15'h4018 == address; // @[Conditional.scala 37:30]
  wire  _T_1946 = 15'h401c == address; // @[Conditional.scala 37:30]
  wire  _T_1947 = 15'h4020 == address; // @[Conditional.scala 37:30]
  wire  _T_1948 = 15'h4024 == address; // @[Conditional.scala 37:30]
  wire  _T_1949 = 15'h4028 == address; // @[Conditional.scala 37:30]
  wire  _T_1950 = 15'h402c == address; // @[Conditional.scala 37:30]
  wire  _T_1951 = 15'h4030 == address; // @[Conditional.scala 37:30]
  wire  _T_1952 = 15'h4034 == address; // @[Conditional.scala 37:30]
  wire  _T_1953 = 15'h4038 == address; // @[Conditional.scala 37:30]
  wire  _T_1954 = 15'h403c == address; // @[Conditional.scala 37:30]
  wire  _T_1955 = 15'h4040 == address; // @[Conditional.scala 37:30]
  wire  _T_1956 = 15'h4044 == address; // @[Conditional.scala 37:30]
  wire  _T_1957 = 15'h4048 == address; // @[Conditional.scala 37:30]
  wire  _T_1958 = 15'h404c == address; // @[Conditional.scala 37:30]
  wire  _T_1959 = 15'h4050 == address; // @[Conditional.scala 37:30]
  wire  _T_1960 = 15'h4054 == address; // @[Conditional.scala 37:30]
  wire  _T_1961 = 15'h4058 == address; // @[Conditional.scala 37:30]
  wire  _T_1962 = 15'h405c == address; // @[Conditional.scala 37:30]
  wire  _T_1963 = 15'h4060 == address; // @[Conditional.scala 37:30]
  wire  _T_1964 = 15'h4064 == address; // @[Conditional.scala 37:30]
  wire  _T_1965 = 15'h4068 == address; // @[Conditional.scala 37:30]
  wire  _T_1966 = 15'h406c == address; // @[Conditional.scala 37:30]
  wire  _T_1967 = 15'h4070 == address; // @[Conditional.scala 37:30]
  wire  _T_1968 = 15'h4074 == address; // @[Conditional.scala 37:30]
  wire  _T_1969 = 15'h4078 == address; // @[Conditional.scala 37:30]
  wire  _T_1970 = 15'h407c == address; // @[Conditional.scala 37:30]
  wire  _T_1971 = 15'h2004 == address; // @[Conditional.scala 37:30]
  wire  _T_1972 = 15'h2008 == address; // @[Conditional.scala 37:30]
  wire  _T_1973 = 15'h200c == address; // @[Conditional.scala 37:30]
  wire  _T_1974 = 15'h2010 == address; // @[Conditional.scala 37:30]
  wire  _T_1975 = 15'h2014 == address; // @[Conditional.scala 37:30]
  wire  _T_1976 = 15'h2018 == address; // @[Conditional.scala 37:30]
  wire  _T_1977 = 15'h201c == address; // @[Conditional.scala 37:30]
  wire  _T_1978 = 15'h2020 == address; // @[Conditional.scala 37:30]
  wire  _T_1979 = 15'h2024 == address; // @[Conditional.scala 37:30]
  wire  _T_1980 = 15'h2028 == address; // @[Conditional.scala 37:30]
  wire  _T_1981 = 15'h202c == address; // @[Conditional.scala 37:30]
  wire  _T_1982 = 15'h2030 == address; // @[Conditional.scala 37:30]
  wire  _T_1983 = 15'h2034 == address; // @[Conditional.scala 37:30]
  wire  _T_1984 = 15'h2038 == address; // @[Conditional.scala 37:30]
  wire  _T_1985 = 15'h203c == address; // @[Conditional.scala 37:30]
  wire  _T_1986 = 15'h2040 == address; // @[Conditional.scala 37:30]
  wire  _T_1987 = 15'h2044 == address; // @[Conditional.scala 37:30]
  wire  _T_1988 = 15'h2048 == address; // @[Conditional.scala 37:30]
  wire  _T_1989 = 15'h204c == address; // @[Conditional.scala 37:30]
  wire  _T_1990 = 15'h2050 == address; // @[Conditional.scala 37:30]
  wire  _T_1991 = 15'h2054 == address; // @[Conditional.scala 37:30]
  wire  _T_1992 = 15'h2058 == address; // @[Conditional.scala 37:30]
  wire  _T_1993 = 15'h205c == address; // @[Conditional.scala 37:30]
  wire  _T_1994 = 15'h2060 == address; // @[Conditional.scala 37:30]
  wire  _T_1995 = 15'h2064 == address; // @[Conditional.scala 37:30]
  wire  _T_1996 = 15'h2068 == address; // @[Conditional.scala 37:30]
  wire  _T_1997 = 15'h206c == address; // @[Conditional.scala 37:30]
  wire  _T_1998 = 15'h2070 == address; // @[Conditional.scala 37:30]
  wire  _T_1999 = 15'h2074 == address; // @[Conditional.scala 37:30]
  wire  _T_2000 = 15'h2078 == address; // @[Conditional.scala 37:30]
  wire  _T_2001 = 15'h207c == address; // @[Conditional.scala 37:30]
  wire  _T_2002 = 15'h4 == address; // @[Conditional.scala 37:30]
  wire  _T_2003 = 15'h8 == address; // @[Conditional.scala 37:30]
  wire  _T_2004 = 15'hc == address; // @[Conditional.scala 37:30]
  wire  _T_2005 = 15'h10 == address; // @[Conditional.scala 37:30]
  wire  _T_2006 = 15'h14 == address; // @[Conditional.scala 37:30]
  wire  _T_2007 = 15'h18 == address; // @[Conditional.scala 37:30]
  wire  _T_2008 = 15'h1c == address; // @[Conditional.scala 37:30]
  wire  _T_2009 = 15'h20 == address; // @[Conditional.scala 37:30]
  wire  _T_2010 = 15'h24 == address; // @[Conditional.scala 37:30]
  wire  _T_2011 = 15'h28 == address; // @[Conditional.scala 37:30]
  wire  _T_2012 = 15'h2c == address; // @[Conditional.scala 37:30]
  wire  _T_2013 = 15'h30 == address; // @[Conditional.scala 37:30]
  wire  _T_2014 = 15'h34 == address; // @[Conditional.scala 37:30]
  wire  _T_2015 = 15'h38 == address; // @[Conditional.scala 37:30]
  wire  _T_2016 = 15'h3c == address; // @[Conditional.scala 37:30]
  wire  _T_2017 = 15'h40 == address; // @[Conditional.scala 37:30]
  wire  _T_2018 = 15'h44 == address; // @[Conditional.scala 37:30]
  wire  _T_2019 = 15'h48 == address; // @[Conditional.scala 37:30]
  wire  _T_2020 = 15'h4c == address; // @[Conditional.scala 37:30]
  wire  _T_2021 = 15'h50 == address; // @[Conditional.scala 37:30]
  wire  _T_2022 = 15'h54 == address; // @[Conditional.scala 37:30]
  wire  _T_2023 = 15'h58 == address; // @[Conditional.scala 37:30]
  wire  _T_2024 = 15'h5c == address; // @[Conditional.scala 37:30]
  wire  _T_2025 = 15'h60 == address; // @[Conditional.scala 37:30]
  wire  _T_2026 = 15'h64 == address; // @[Conditional.scala 37:30]
  wire  _T_2027 = 15'h68 == address; // @[Conditional.scala 37:30]
  wire  _T_2028 = 15'h6c == address; // @[Conditional.scala 37:30]
  wire  _T_2029 = 15'h70 == address; // @[Conditional.scala 37:30]
  wire  _T_2030 = 15'h74 == address; // @[Conditional.scala 37:30]
  wire  _T_2031 = 15'h78 == address; // @[Conditional.scala 37:30]
  wire  _T_2032 = 15'h7c == address; // @[Conditional.scala 37:30]
  wire [3:0] _GEN_94 = _T_2032 ? 4'h2 : 4'h1; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_95 = _T_2031 ? 4'h2 : _GEN_94; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_96 = _T_2030 ? 4'h2 : _GEN_95; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_97 = _T_2029 ? 4'h2 : _GEN_96; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_98 = _T_2028 ? 4'h2 : _GEN_97; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_99 = _T_2027 ? 4'h2 : _GEN_98; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_100 = _T_2026 ? 4'h2 : _GEN_99; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_101 = _T_2025 ? 4'h2 : _GEN_100; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_102 = _T_2024 ? 4'h2 : _GEN_101; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_103 = _T_2023 ? 4'h2 : _GEN_102; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_104 = _T_2022 ? 4'h2 : _GEN_103; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_105 = _T_2021 ? 4'h2 : _GEN_104; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_106 = _T_2020 ? 4'h2 : _GEN_105; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_107 = _T_2019 ? 4'h2 : _GEN_106; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_108 = _T_2018 ? 4'h2 : _GEN_107; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_109 = _T_2017 ? 4'h2 : _GEN_108; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_110 = _T_2016 ? 4'h2 : _GEN_109; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_111 = _T_2015 ? 4'h2 : _GEN_110; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_112 = _T_2014 ? 4'h2 : _GEN_111; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_113 = _T_2013 ? 4'h2 : _GEN_112; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_114 = _T_2012 ? 4'h2 : _GEN_113; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_115 = _T_2011 ? 4'h2 : _GEN_114; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_116 = _T_2010 ? 4'h2 : _GEN_115; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_117 = _T_2009 ? 4'h2 : _GEN_116; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_118 = _T_2008 ? 4'h2 : _GEN_117; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_119 = _T_2007 ? 4'h2 : _GEN_118; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_120 = _T_2006 ? 4'h2 : _GEN_119; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_121 = _T_2005 ? 4'h2 : _GEN_120; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_122 = _T_2004 ? 4'h2 : _GEN_121; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_123 = _T_2003 ? 4'h2 : _GEN_122; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_124 = _T_2002 ? 4'h2 : _GEN_123; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_125 = _T_2001 ? 4'h4 : _GEN_124; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_126 = _T_2000 ? 4'h4 : _GEN_125; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_127 = _T_1999 ? 4'h4 : _GEN_126; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_128 = _T_1998 ? 4'h4 : _GEN_127; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_129 = _T_1997 ? 4'h4 : _GEN_128; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_130 = _T_1996 ? 4'h4 : _GEN_129; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_131 = _T_1995 ? 4'h4 : _GEN_130; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_132 = _T_1994 ? 4'h4 : _GEN_131; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_133 = _T_1993 ? 4'h4 : _GEN_132; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_134 = _T_1992 ? 4'h4 : _GEN_133; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_135 = _T_1991 ? 4'h4 : _GEN_134; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_136 = _T_1990 ? 4'h4 : _GEN_135; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_137 = _T_1989 ? 4'h4 : _GEN_136; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_138 = _T_1988 ? 4'h4 : _GEN_137; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_139 = _T_1987 ? 4'h4 : _GEN_138; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_140 = _T_1986 ? 4'h4 : _GEN_139; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_141 = _T_1985 ? 4'h4 : _GEN_140; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_142 = _T_1984 ? 4'h4 : _GEN_141; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_143 = _T_1983 ? 4'h4 : _GEN_142; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_144 = _T_1982 ? 4'h4 : _GEN_143; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_145 = _T_1981 ? 4'h4 : _GEN_144; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_146 = _T_1980 ? 4'h4 : _GEN_145; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_147 = _T_1979 ? 4'h4 : _GEN_146; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_148 = _T_1978 ? 4'h4 : _GEN_147; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_149 = _T_1977 ? 4'h4 : _GEN_148; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_150 = _T_1976 ? 4'h4 : _GEN_149; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_151 = _T_1975 ? 4'h4 : _GEN_150; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_152 = _T_1974 ? 4'h4 : _GEN_151; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_153 = _T_1973 ? 4'h4 : _GEN_152; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_154 = _T_1972 ? 4'h4 : _GEN_153; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_155 = _T_1971 ? 4'h4 : _GEN_154; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_156 = _T_1970 ? 4'h8 : _GEN_155; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_157 = _T_1969 ? 4'h8 : _GEN_156; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_158 = _T_1968 ? 4'h8 : _GEN_157; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_159 = _T_1967 ? 4'h8 : _GEN_158; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_160 = _T_1966 ? 4'h8 : _GEN_159; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_161 = _T_1965 ? 4'h8 : _GEN_160; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_162 = _T_1964 ? 4'h8 : _GEN_161; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_163 = _T_1963 ? 4'h8 : _GEN_162; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_164 = _T_1962 ? 4'h8 : _GEN_163; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_165 = _T_1961 ? 4'h8 : _GEN_164; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_166 = _T_1960 ? 4'h8 : _GEN_165; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_167 = _T_1959 ? 4'h8 : _GEN_166; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_168 = _T_1958 ? 4'h8 : _GEN_167; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_169 = _T_1957 ? 4'h8 : _GEN_168; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_170 = _T_1956 ? 4'h8 : _GEN_169; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_171 = _T_1955 ? 4'h8 : _GEN_170; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_172 = _T_1954 ? 4'h8 : _GEN_171; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_173 = _T_1953 ? 4'h8 : _GEN_172; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_174 = _T_1952 ? 4'h8 : _GEN_173; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_175 = _T_1951 ? 4'h8 : _GEN_174; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_176 = _T_1950 ? 4'h8 : _GEN_175; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_177 = _T_1949 ? 4'h8 : _GEN_176; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_178 = _T_1948 ? 4'h8 : _GEN_177; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_179 = _T_1947 ? 4'h8 : _GEN_178; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_180 = _T_1946 ? 4'h8 : _GEN_179; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_181 = _T_1945 ? 4'h8 : _GEN_180; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_182 = _T_1944 ? 4'h8 : _GEN_181; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_183 = _T_1943 ? 4'h8 : _GEN_182; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_184 = _T_1942 ? 4'h8 : _GEN_183; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_185 = _T_1941 ? 4'h8 : _GEN_184; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_186 = _T_1940 ? 4'h8 : _GEN_185; // @[Conditional.scala 39:67]
  wire [3:0] mask = _T_1939 ? 4'h4 : _GEN_186; // @[Conditional.scala 40:58]
  wire  _T_1901 = picm_mken_ff & mask[3]; // @[pic_ctrl.scala 299:19]
  wire  _T_1906 = picm_mken_ff & mask[2]; // @[pic_ctrl.scala 300:19]
  wire  _T_1911 = picm_mken_ff & mask[1]; // @[pic_ctrl.scala 301:19]
  wire [31:0] _T_1919 = intpend_reg_read ? intpend_rd_out : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1920 = _T_21 ? _T_1890 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1921 = _T_24 ? _T_1893 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1922 = _T_27 ? _T_1896 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1923 = config_reg_re ? _T_1899 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1924 = _T_1901 ? 32'h3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1925 = _T_1906 ? 32'h1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1926 = _T_1911 ? 32'hf : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1928 = _T_1919 | _T_1920; // @[Mux.scala 27:72]
  wire [31:0] _T_1929 = _T_1928 | _T_1921; // @[Mux.scala 27:72]
  wire [31:0] _T_1930 = _T_1929 | _T_1922; // @[Mux.scala 27:72]
  wire [31:0] _T_1931 = _T_1930 | _T_1923; // @[Mux.scala 27:72]
  wire [31:0] _T_1932 = _T_1931 | _T_1924; // @[Mux.scala 27:72]
  wire [31:0] _T_1933 = _T_1932 | _T_1925; // @[Mux.scala 27:72]
  wire [31:0] picm_rd_data_in = _T_1933 | _T_1926; // @[Mux.scala 27:72]
  wire [7:0] level_intpend_id_5_0 = out_id_34; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30 pic_ctrl.scala 232:41]
  wire [7:0] level_intpend_id_1_18 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_1_19 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_1_20 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_1_21 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_1_22 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_1_23 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_1_24 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_1_25 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_1_26 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_1_27 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_1_28 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_1_29 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_1_30 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_1_31 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_1_32 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_1_33 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_2_10 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_2_11 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_2_12 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_2_13 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_2_14 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_2_15 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_2_16 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_2_17 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_2_18 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_2_19 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_2_20 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_2_21 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_2_22 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_2_23 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_2_24 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_2_25 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_2_26 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_2_27 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_2_28 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_2_29 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_2_30 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_2_31 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_2_32 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_2_33 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_3_6 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_3_7 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_3_8 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_3_9 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_3_10 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_3_11 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_3_12 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_3_13 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_3_14 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_3_15 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_3_16 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_3_17 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_3_18 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_3_19 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_3_20 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_3_21 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_3_22 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_3_23 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_3_24 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_3_25 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_3_26 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_3_27 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_3_28 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_3_29 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_3_30 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_3_31 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_3_32 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_3_33 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_4_4 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_4_5 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_4_6 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_4_7 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_4_8 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_4_9 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_4_10 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_4_11 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_4_12 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_4_13 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_4_14 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_4_15 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_4_16 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_4_17 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_4_18 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_4_19 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_4_20 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_4_21 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_4_22 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_4_23 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_4_24 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_4_25 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_4_26 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_4_27 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_4_28 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_4_29 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_4_30 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_4_31 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_4_32 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_4_33 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_5_1 = out_id_33; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30 pic_ctrl.scala 232:41]
  wire [7:0] level_intpend_id_5_2 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30 pic_ctrl.scala 229:44]
  wire [7:0] level_intpend_id_5_3 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_5_4 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_5_5 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_5_6 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_5_7 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_5_8 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_5_9 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_5_10 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_5_11 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_5_12 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_5_13 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_5_14 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_5_15 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_5_16 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_5_17 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_5_18 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_5_19 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_5_20 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_5_21 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_5_22 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_5_23 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_5_24 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_5_25 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_5_26 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_5_27 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_5_28 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_5_29 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_5_30 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_5_31 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_5_32 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  wire [7:0] level_intpend_id_5_33 = 8'h0; // @[pic_ctrl.scala 214:32 pic_ctrl.scala 218:30]
  rvclkhdr rvclkhdr ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_io_l1clk),
    .io_clk(rvclkhdr_io_clk),
    .io_en(rvclkhdr_io_en),
    .io_scan_mode(rvclkhdr_io_scan_mode)
  );
  rvclkhdr rvclkhdr_1 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_1_io_l1clk),
    .io_clk(rvclkhdr_1_io_clk),
    .io_en(rvclkhdr_1_io_en),
    .io_scan_mode(rvclkhdr_1_io_scan_mode)
  );
  rvclkhdr rvclkhdr_2 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_2_io_l1clk),
    .io_clk(rvclkhdr_2_io_clk),
    .io_en(rvclkhdr_2_io_en),
    .io_scan_mode(rvclkhdr_2_io_scan_mode)
  );
  rvclkhdr rvclkhdr_3 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_3_io_l1clk),
    .io_clk(rvclkhdr_3_io_clk),
    .io_en(rvclkhdr_3_io_en),
    .io_scan_mode(rvclkhdr_3_io_scan_mode)
  );
  rvclkhdr rvclkhdr_4 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_4_io_l1clk),
    .io_clk(rvclkhdr_4_io_clk),
    .io_en(rvclkhdr_4_io_en),
    .io_scan_mode(rvclkhdr_4_io_scan_mode)
  );
  assign io_lsu_pic_picm_rd_data = picm_bypass_ff ? picm_wr_data_ff : picm_rd_data_in; // @[pic_ctrl.scala 305:27]
  assign io_dec_pic_pic_claimid = _T_1642; // @[pic_ctrl.scala 262:49]
  assign io_dec_pic_pic_pl = _T_1643; // @[pic_ctrl.scala 263:44]
  assign io_dec_pic_mhwakeup = _T_1652; // @[pic_ctrl.scala 270:23]
  assign io_dec_pic_mexintpend = _T_1650; // @[pic_ctrl.scala 267:25]
  assign rvclkhdr_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_io_en = _T_19 | io_clk_override; // @[lib.scala 345:16]
  assign rvclkhdr_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_1_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_1_io_en = io_lsu_pic_picm_wren | io_clk_override; // @[lib.scala 345:16]
  assign rvclkhdr_1_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_2_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_2_io_en = _T_22 | io_clk_override; // @[lib.scala 345:16]
  assign rvclkhdr_2_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_3_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_3_io_en = _T_25 | io_clk_override; // @[lib.scala 345:16]
  assign rvclkhdr_3_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_4_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_4_io_en = _T_28 | io_clk_override; // @[lib.scala 345:16]
  assign rvclkhdr_4_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  picm_raddr_ff = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  picm_waddr_ff = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  picm_wren_ff = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  picm_rden_ff = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  picm_mken_ff = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  picm_wr_data_ff = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  _T_33 = _RAND_6[30:0];
  _RAND_7 = {1{`RANDOM}};
  _T_34 = _RAND_7[30:0];
  _RAND_8 = {1{`RANDOM}};
  intpriority_reg_1 = _RAND_8[3:0];
  _RAND_9 = {1{`RANDOM}};
  intpriority_reg_2 = _RAND_9[3:0];
  _RAND_10 = {1{`RANDOM}};
  intpriority_reg_3 = _RAND_10[3:0];
  _RAND_11 = {1{`RANDOM}};
  intpriority_reg_4 = _RAND_11[3:0];
  _RAND_12 = {1{`RANDOM}};
  intpriority_reg_5 = _RAND_12[3:0];
  _RAND_13 = {1{`RANDOM}};
  intpriority_reg_6 = _RAND_13[3:0];
  _RAND_14 = {1{`RANDOM}};
  intpriority_reg_7 = _RAND_14[3:0];
  _RAND_15 = {1{`RANDOM}};
  intpriority_reg_8 = _RAND_15[3:0];
  _RAND_16 = {1{`RANDOM}};
  intpriority_reg_9 = _RAND_16[3:0];
  _RAND_17 = {1{`RANDOM}};
  intpriority_reg_10 = _RAND_17[3:0];
  _RAND_18 = {1{`RANDOM}};
  intpriority_reg_11 = _RAND_18[3:0];
  _RAND_19 = {1{`RANDOM}};
  intpriority_reg_12 = _RAND_19[3:0];
  _RAND_20 = {1{`RANDOM}};
  intpriority_reg_13 = _RAND_20[3:0];
  _RAND_21 = {1{`RANDOM}};
  intpriority_reg_14 = _RAND_21[3:0];
  _RAND_22 = {1{`RANDOM}};
  intpriority_reg_15 = _RAND_22[3:0];
  _RAND_23 = {1{`RANDOM}};
  intpriority_reg_16 = _RAND_23[3:0];
  _RAND_24 = {1{`RANDOM}};
  intpriority_reg_17 = _RAND_24[3:0];
  _RAND_25 = {1{`RANDOM}};
  intpriority_reg_18 = _RAND_25[3:0];
  _RAND_26 = {1{`RANDOM}};
  intpriority_reg_19 = _RAND_26[3:0];
  _RAND_27 = {1{`RANDOM}};
  intpriority_reg_20 = _RAND_27[3:0];
  _RAND_28 = {1{`RANDOM}};
  intpriority_reg_21 = _RAND_28[3:0];
  _RAND_29 = {1{`RANDOM}};
  intpriority_reg_22 = _RAND_29[3:0];
  _RAND_30 = {1{`RANDOM}};
  intpriority_reg_23 = _RAND_30[3:0];
  _RAND_31 = {1{`RANDOM}};
  intpriority_reg_24 = _RAND_31[3:0];
  _RAND_32 = {1{`RANDOM}};
  intpriority_reg_25 = _RAND_32[3:0];
  _RAND_33 = {1{`RANDOM}};
  intpriority_reg_26 = _RAND_33[3:0];
  _RAND_34 = {1{`RANDOM}};
  intpriority_reg_27 = _RAND_34[3:0];
  _RAND_35 = {1{`RANDOM}};
  intpriority_reg_28 = _RAND_35[3:0];
  _RAND_36 = {1{`RANDOM}};
  intpriority_reg_29 = _RAND_36[3:0];
  _RAND_37 = {1{`RANDOM}};
  intpriority_reg_30 = _RAND_37[3:0];
  _RAND_38 = {1{`RANDOM}};
  intpriority_reg_31 = _RAND_38[3:0];
  _RAND_39 = {1{`RANDOM}};
  intenable_reg_1 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  intenable_reg_2 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  intenable_reg_3 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  intenable_reg_4 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  intenable_reg_5 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  intenable_reg_6 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  intenable_reg_7 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  intenable_reg_8 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  intenable_reg_9 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  intenable_reg_10 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  intenable_reg_11 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  intenable_reg_12 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  intenable_reg_13 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  intenable_reg_14 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  intenable_reg_15 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  intenable_reg_16 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  intenable_reg_17 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  intenable_reg_18 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  intenable_reg_19 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  intenable_reg_20 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  intenable_reg_21 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  intenable_reg_22 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  intenable_reg_23 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  intenable_reg_24 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  intenable_reg_25 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  intenable_reg_26 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  intenable_reg_27 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  intenable_reg_28 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  intenable_reg_29 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  intenable_reg_30 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  intenable_reg_31 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  gw_config_reg_1 = _RAND_70[1:0];
  _RAND_71 = {1{`RANDOM}};
  gw_config_reg_2 = _RAND_71[1:0];
  _RAND_72 = {1{`RANDOM}};
  gw_config_reg_3 = _RAND_72[1:0];
  _RAND_73 = {1{`RANDOM}};
  gw_config_reg_4 = _RAND_73[1:0];
  _RAND_74 = {1{`RANDOM}};
  gw_config_reg_5 = _RAND_74[1:0];
  _RAND_75 = {1{`RANDOM}};
  gw_config_reg_6 = _RAND_75[1:0];
  _RAND_76 = {1{`RANDOM}};
  gw_config_reg_7 = _RAND_76[1:0];
  _RAND_77 = {1{`RANDOM}};
  gw_config_reg_8 = _RAND_77[1:0];
  _RAND_78 = {1{`RANDOM}};
  gw_config_reg_9 = _RAND_78[1:0];
  _RAND_79 = {1{`RANDOM}};
  gw_config_reg_10 = _RAND_79[1:0];
  _RAND_80 = {1{`RANDOM}};
  gw_config_reg_11 = _RAND_80[1:0];
  _RAND_81 = {1{`RANDOM}};
  gw_config_reg_12 = _RAND_81[1:0];
  _RAND_82 = {1{`RANDOM}};
  gw_config_reg_13 = _RAND_82[1:0];
  _RAND_83 = {1{`RANDOM}};
  gw_config_reg_14 = _RAND_83[1:0];
  _RAND_84 = {1{`RANDOM}};
  gw_config_reg_15 = _RAND_84[1:0];
  _RAND_85 = {1{`RANDOM}};
  gw_config_reg_16 = _RAND_85[1:0];
  _RAND_86 = {1{`RANDOM}};
  gw_config_reg_17 = _RAND_86[1:0];
  _RAND_87 = {1{`RANDOM}};
  gw_config_reg_18 = _RAND_87[1:0];
  _RAND_88 = {1{`RANDOM}};
  gw_config_reg_19 = _RAND_88[1:0];
  _RAND_89 = {1{`RANDOM}};
  gw_config_reg_20 = _RAND_89[1:0];
  _RAND_90 = {1{`RANDOM}};
  gw_config_reg_21 = _RAND_90[1:0];
  _RAND_91 = {1{`RANDOM}};
  gw_config_reg_22 = _RAND_91[1:0];
  _RAND_92 = {1{`RANDOM}};
  gw_config_reg_23 = _RAND_92[1:0];
  _RAND_93 = {1{`RANDOM}};
  gw_config_reg_24 = _RAND_93[1:0];
  _RAND_94 = {1{`RANDOM}};
  gw_config_reg_25 = _RAND_94[1:0];
  _RAND_95 = {1{`RANDOM}};
  gw_config_reg_26 = _RAND_95[1:0];
  _RAND_96 = {1{`RANDOM}};
  gw_config_reg_27 = _RAND_96[1:0];
  _RAND_97 = {1{`RANDOM}};
  gw_config_reg_28 = _RAND_97[1:0];
  _RAND_98 = {1{`RANDOM}};
  gw_config_reg_29 = _RAND_98[1:0];
  _RAND_99 = {1{`RANDOM}};
  gw_config_reg_30 = _RAND_99[1:0];
  _RAND_100 = {1{`RANDOM}};
  gw_config_reg_31 = _RAND_100[1:0];
  _RAND_101 = {1{`RANDOM}};
  gw_int_pending = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  gw_int_pending_1 = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  gw_int_pending_2 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  gw_int_pending_3 = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  gw_int_pending_4 = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  gw_int_pending_5 = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  gw_int_pending_6 = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  gw_int_pending_7 = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  gw_int_pending_8 = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  gw_int_pending_9 = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  gw_int_pending_10 = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  gw_int_pending_11 = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  gw_int_pending_12 = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  gw_int_pending_13 = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  gw_int_pending_14 = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  gw_int_pending_15 = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  gw_int_pending_16 = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  gw_int_pending_17 = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  gw_int_pending_18 = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  gw_int_pending_19 = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  gw_int_pending_20 = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  gw_int_pending_21 = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  gw_int_pending_22 = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  gw_int_pending_23 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  gw_int_pending_24 = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  gw_int_pending_25 = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  gw_int_pending_26 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  gw_int_pending_27 = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  gw_int_pending_28 = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  gw_int_pending_29 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  gw_int_pending_30 = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  config_reg = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  _T_1642 = _RAND_133[7:0];
  _RAND_134 = {1{`RANDOM}};
  _T_1643 = _RAND_134[3:0];
  _RAND_135 = {1{`RANDOM}};
  _T_1650 = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  _T_1652 = _RAND_136[0:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    picm_raddr_ff = 32'h0;
  end
  if (reset) begin
    picm_waddr_ff = 32'h0;
  end
  if (reset) begin
    picm_wren_ff = 1'h0;
  end
  if (reset) begin
    picm_rden_ff = 1'h0;
  end
  if (reset) begin
    picm_mken_ff = 1'h0;
  end
  if (reset) begin
    picm_wr_data_ff = 32'h0;
  end
  if (reset) begin
    _T_33 = 31'h0;
  end
  if (reset) begin
    _T_34 = 31'h0;
  end
  if (reset) begin
    intpriority_reg_1 = 4'h0;
  end
  if (reset) begin
    intpriority_reg_2 = 4'h0;
  end
  if (reset) begin
    intpriority_reg_3 = 4'h0;
  end
  if (reset) begin
    intpriority_reg_4 = 4'h0;
  end
  if (reset) begin
    intpriority_reg_5 = 4'h0;
  end
  if (reset) begin
    intpriority_reg_6 = 4'h0;
  end
  if (reset) begin
    intpriority_reg_7 = 4'h0;
  end
  if (reset) begin
    intpriority_reg_8 = 4'h0;
  end
  if (reset) begin
    intpriority_reg_9 = 4'h0;
  end
  if (reset) begin
    intpriority_reg_10 = 4'h0;
  end
  if (reset) begin
    intpriority_reg_11 = 4'h0;
  end
  if (reset) begin
    intpriority_reg_12 = 4'h0;
  end
  if (reset) begin
    intpriority_reg_13 = 4'h0;
  end
  if (reset) begin
    intpriority_reg_14 = 4'h0;
  end
  if (reset) begin
    intpriority_reg_15 = 4'h0;
  end
  if (reset) begin
    intpriority_reg_16 = 4'h0;
  end
  if (reset) begin
    intpriority_reg_17 = 4'h0;
  end
  if (reset) begin
    intpriority_reg_18 = 4'h0;
  end
  if (reset) begin
    intpriority_reg_19 = 4'h0;
  end
  if (reset) begin
    intpriority_reg_20 = 4'h0;
  end
  if (reset) begin
    intpriority_reg_21 = 4'h0;
  end
  if (reset) begin
    intpriority_reg_22 = 4'h0;
  end
  if (reset) begin
    intpriority_reg_23 = 4'h0;
  end
  if (reset) begin
    intpriority_reg_24 = 4'h0;
  end
  if (reset) begin
    intpriority_reg_25 = 4'h0;
  end
  if (reset) begin
    intpriority_reg_26 = 4'h0;
  end
  if (reset) begin
    intpriority_reg_27 = 4'h0;
  end
  if (reset) begin
    intpriority_reg_28 = 4'h0;
  end
  if (reset) begin
    intpriority_reg_29 = 4'h0;
  end
  if (reset) begin
    intpriority_reg_30 = 4'h0;
  end
  if (reset) begin
    intpriority_reg_31 = 4'h0;
  end
  if (reset) begin
    intenable_reg_1 = 1'h0;
  end
  if (reset) begin
    intenable_reg_2 = 1'h0;
  end
  if (reset) begin
    intenable_reg_3 = 1'h0;
  end
  if (reset) begin
    intenable_reg_4 = 1'h0;
  end
  if (reset) begin
    intenable_reg_5 = 1'h0;
  end
  if (reset) begin
    intenable_reg_6 = 1'h0;
  end
  if (reset) begin
    intenable_reg_7 = 1'h0;
  end
  if (reset) begin
    intenable_reg_8 = 1'h0;
  end
  if (reset) begin
    intenable_reg_9 = 1'h0;
  end
  if (reset) begin
    intenable_reg_10 = 1'h0;
  end
  if (reset) begin
    intenable_reg_11 = 1'h0;
  end
  if (reset) begin
    intenable_reg_12 = 1'h0;
  end
  if (reset) begin
    intenable_reg_13 = 1'h0;
  end
  if (reset) begin
    intenable_reg_14 = 1'h0;
  end
  if (reset) begin
    intenable_reg_15 = 1'h0;
  end
  if (reset) begin
    intenable_reg_16 = 1'h0;
  end
  if (reset) begin
    intenable_reg_17 = 1'h0;
  end
  if (reset) begin
    intenable_reg_18 = 1'h0;
  end
  if (reset) begin
    intenable_reg_19 = 1'h0;
  end
  if (reset) begin
    intenable_reg_20 = 1'h0;
  end
  if (reset) begin
    intenable_reg_21 = 1'h0;
  end
  if (reset) begin
    intenable_reg_22 = 1'h0;
  end
  if (reset) begin
    intenable_reg_23 = 1'h0;
  end
  if (reset) begin
    intenable_reg_24 = 1'h0;
  end
  if (reset) begin
    intenable_reg_25 = 1'h0;
  end
  if (reset) begin
    intenable_reg_26 = 1'h0;
  end
  if (reset) begin
    intenable_reg_27 = 1'h0;
  end
  if (reset) begin
    intenable_reg_28 = 1'h0;
  end
  if (reset) begin
    intenable_reg_29 = 1'h0;
  end
  if (reset) begin
    intenable_reg_30 = 1'h0;
  end
  if (reset) begin
    intenable_reg_31 = 1'h0;
  end
  if (reset) begin
    gw_config_reg_1 = 2'h0;
  end
  if (reset) begin
    gw_config_reg_2 = 2'h0;
  end
  if (reset) begin
    gw_config_reg_3 = 2'h0;
  end
  if (reset) begin
    gw_config_reg_4 = 2'h0;
  end
  if (reset) begin
    gw_config_reg_5 = 2'h0;
  end
  if (reset) begin
    gw_config_reg_6 = 2'h0;
  end
  if (reset) begin
    gw_config_reg_7 = 2'h0;
  end
  if (reset) begin
    gw_config_reg_8 = 2'h0;
  end
  if (reset) begin
    gw_config_reg_9 = 2'h0;
  end
  if (reset) begin
    gw_config_reg_10 = 2'h0;
  end
  if (reset) begin
    gw_config_reg_11 = 2'h0;
  end
  if (reset) begin
    gw_config_reg_12 = 2'h0;
  end
  if (reset) begin
    gw_config_reg_13 = 2'h0;
  end
  if (reset) begin
    gw_config_reg_14 = 2'h0;
  end
  if (reset) begin
    gw_config_reg_15 = 2'h0;
  end
  if (reset) begin
    gw_config_reg_16 = 2'h0;
  end
  if (reset) begin
    gw_config_reg_17 = 2'h0;
  end
  if (reset) begin
    gw_config_reg_18 = 2'h0;
  end
  if (reset) begin
    gw_config_reg_19 = 2'h0;
  end
  if (reset) begin
    gw_config_reg_20 = 2'h0;
  end
  if (reset) begin
    gw_config_reg_21 = 2'h0;
  end
  if (reset) begin
    gw_config_reg_22 = 2'h0;
  end
  if (reset) begin
    gw_config_reg_23 = 2'h0;
  end
  if (reset) begin
    gw_config_reg_24 = 2'h0;
  end
  if (reset) begin
    gw_config_reg_25 = 2'h0;
  end
  if (reset) begin
    gw_config_reg_26 = 2'h0;
  end
  if (reset) begin
    gw_config_reg_27 = 2'h0;
  end
  if (reset) begin
    gw_config_reg_28 = 2'h0;
  end
  if (reset) begin
    gw_config_reg_29 = 2'h0;
  end
  if (reset) begin
    gw_config_reg_30 = 2'h0;
  end
  if (reset) begin
    gw_config_reg_31 = 2'h0;
  end
  if (reset) begin
    gw_int_pending = 1'h0;
  end
  if (reset) begin
    gw_int_pending_1 = 1'h0;
  end
  if (reset) begin
    gw_int_pending_2 = 1'h0;
  end
  if (reset) begin
    gw_int_pending_3 = 1'h0;
  end
  if (reset) begin
    gw_int_pending_4 = 1'h0;
  end
  if (reset) begin
    gw_int_pending_5 = 1'h0;
  end
  if (reset) begin
    gw_int_pending_6 = 1'h0;
  end
  if (reset) begin
    gw_int_pending_7 = 1'h0;
  end
  if (reset) begin
    gw_int_pending_8 = 1'h0;
  end
  if (reset) begin
    gw_int_pending_9 = 1'h0;
  end
  if (reset) begin
    gw_int_pending_10 = 1'h0;
  end
  if (reset) begin
    gw_int_pending_11 = 1'h0;
  end
  if (reset) begin
    gw_int_pending_12 = 1'h0;
  end
  if (reset) begin
    gw_int_pending_13 = 1'h0;
  end
  if (reset) begin
    gw_int_pending_14 = 1'h0;
  end
  if (reset) begin
    gw_int_pending_15 = 1'h0;
  end
  if (reset) begin
    gw_int_pending_16 = 1'h0;
  end
  if (reset) begin
    gw_int_pending_17 = 1'h0;
  end
  if (reset) begin
    gw_int_pending_18 = 1'h0;
  end
  if (reset) begin
    gw_int_pending_19 = 1'h0;
  end
  if (reset) begin
    gw_int_pending_20 = 1'h0;
  end
  if (reset) begin
    gw_int_pending_21 = 1'h0;
  end
  if (reset) begin
    gw_int_pending_22 = 1'h0;
  end
  if (reset) begin
    gw_int_pending_23 = 1'h0;
  end
  if (reset) begin
    gw_int_pending_24 = 1'h0;
  end
  if (reset) begin
    gw_int_pending_25 = 1'h0;
  end
  if (reset) begin
    gw_int_pending_26 = 1'h0;
  end
  if (reset) begin
    gw_int_pending_27 = 1'h0;
  end
  if (reset) begin
    gw_int_pending_28 = 1'h0;
  end
  if (reset) begin
    gw_int_pending_29 = 1'h0;
  end
  if (reset) begin
    gw_int_pending_30 = 1'h0;
  end
  if (reset) begin
    config_reg = 1'h0;
  end
  if (reset) begin
    _T_1642 = 8'h0;
  end
  if (reset) begin
    _T_1643 = 4'h0;
  end
  if (reset) begin
    _T_1650 = 1'h0;
  end
  if (reset) begin
    _T_1652 = 1'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge pic_raddr_c1_clk or posedge reset) begin
    if (reset) begin
      picm_raddr_ff <= 32'h0;
    end else begin
      picm_raddr_ff <= io_lsu_pic_picm_rdaddr;
    end
  end
  always @(posedge pic_data_c1_clk or posedge reset) begin
    if (reset) begin
      picm_waddr_ff <= 32'h0;
    end else begin
      picm_waddr_ff <= io_lsu_pic_picm_wraddr;
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      picm_wren_ff <= 1'h0;
    end else begin
      picm_wren_ff <= io_lsu_pic_picm_wren;
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      picm_rden_ff <= 1'h0;
    end else begin
      picm_rden_ff <= io_lsu_pic_picm_rden;
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      picm_mken_ff <= 1'h0;
    end else begin
      picm_mken_ff <= io_lsu_pic_picm_mken;
    end
  end
  always @(posedge pic_data_c1_clk or posedge reset) begin
    if (reset) begin
      picm_wr_data_ff <= 32'h0;
    end else begin
      picm_wr_data_ff <= io_lsu_pic_picm_wr_data;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      _T_33 <= 31'h0;
    end else begin
      _T_33 <= io_extintsrc_req[31:1];
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      _T_34 <= 31'h0;
    end else begin
      _T_34 <= _T_33;
    end
  end
  always @(posedge pic_pri_c1_clk or posedge reset) begin
    if (reset) begin
      intpriority_reg_1 <= 4'h0;
    end else if (intpriority_reg_we_1) begin
      intpriority_reg_1 <= picm_wr_data_ff[3:0];
    end
  end
  always @(posedge pic_pri_c1_clk or posedge reset) begin
    if (reset) begin
      intpriority_reg_2 <= 4'h0;
    end else if (intpriority_reg_we_2) begin
      intpriority_reg_2 <= picm_wr_data_ff[3:0];
    end
  end
  always @(posedge pic_pri_c1_clk or posedge reset) begin
    if (reset) begin
      intpriority_reg_3 <= 4'h0;
    end else if (intpriority_reg_we_3) begin
      intpriority_reg_3 <= picm_wr_data_ff[3:0];
    end
  end
  always @(posedge pic_pri_c1_clk or posedge reset) begin
    if (reset) begin
      intpriority_reg_4 <= 4'h0;
    end else if (intpriority_reg_we_4) begin
      intpriority_reg_4 <= picm_wr_data_ff[3:0];
    end
  end
  always @(posedge pic_pri_c1_clk or posedge reset) begin
    if (reset) begin
      intpriority_reg_5 <= 4'h0;
    end else if (intpriority_reg_we_5) begin
      intpriority_reg_5 <= picm_wr_data_ff[3:0];
    end
  end
  always @(posedge pic_pri_c1_clk or posedge reset) begin
    if (reset) begin
      intpriority_reg_6 <= 4'h0;
    end else if (intpriority_reg_we_6) begin
      intpriority_reg_6 <= picm_wr_data_ff[3:0];
    end
  end
  always @(posedge pic_pri_c1_clk or posedge reset) begin
    if (reset) begin
      intpriority_reg_7 <= 4'h0;
    end else if (intpriority_reg_we_7) begin
      intpriority_reg_7 <= picm_wr_data_ff[3:0];
    end
  end
  always @(posedge pic_pri_c1_clk or posedge reset) begin
    if (reset) begin
      intpriority_reg_8 <= 4'h0;
    end else if (intpriority_reg_we_8) begin
      intpriority_reg_8 <= picm_wr_data_ff[3:0];
    end
  end
  always @(posedge pic_pri_c1_clk or posedge reset) begin
    if (reset) begin
      intpriority_reg_9 <= 4'h0;
    end else if (intpriority_reg_we_9) begin
      intpriority_reg_9 <= picm_wr_data_ff[3:0];
    end
  end
  always @(posedge pic_pri_c1_clk or posedge reset) begin
    if (reset) begin
      intpriority_reg_10 <= 4'h0;
    end else if (intpriority_reg_we_10) begin
      intpriority_reg_10 <= picm_wr_data_ff[3:0];
    end
  end
  always @(posedge pic_pri_c1_clk or posedge reset) begin
    if (reset) begin
      intpriority_reg_11 <= 4'h0;
    end else if (intpriority_reg_we_11) begin
      intpriority_reg_11 <= picm_wr_data_ff[3:0];
    end
  end
  always @(posedge pic_pri_c1_clk or posedge reset) begin
    if (reset) begin
      intpriority_reg_12 <= 4'h0;
    end else if (intpriority_reg_we_12) begin
      intpriority_reg_12 <= picm_wr_data_ff[3:0];
    end
  end
  always @(posedge pic_pri_c1_clk or posedge reset) begin
    if (reset) begin
      intpriority_reg_13 <= 4'h0;
    end else if (intpriority_reg_we_13) begin
      intpriority_reg_13 <= picm_wr_data_ff[3:0];
    end
  end
  always @(posedge pic_pri_c1_clk or posedge reset) begin
    if (reset) begin
      intpriority_reg_14 <= 4'h0;
    end else if (intpriority_reg_we_14) begin
      intpriority_reg_14 <= picm_wr_data_ff[3:0];
    end
  end
  always @(posedge pic_pri_c1_clk or posedge reset) begin
    if (reset) begin
      intpriority_reg_15 <= 4'h0;
    end else if (intpriority_reg_we_15) begin
      intpriority_reg_15 <= picm_wr_data_ff[3:0];
    end
  end
  always @(posedge pic_pri_c1_clk or posedge reset) begin
    if (reset) begin
      intpriority_reg_16 <= 4'h0;
    end else if (intpriority_reg_we_16) begin
      intpriority_reg_16 <= picm_wr_data_ff[3:0];
    end
  end
  always @(posedge pic_pri_c1_clk or posedge reset) begin
    if (reset) begin
      intpriority_reg_17 <= 4'h0;
    end else if (intpriority_reg_we_17) begin
      intpriority_reg_17 <= picm_wr_data_ff[3:0];
    end
  end
  always @(posedge pic_pri_c1_clk or posedge reset) begin
    if (reset) begin
      intpriority_reg_18 <= 4'h0;
    end else if (intpriority_reg_we_18) begin
      intpriority_reg_18 <= picm_wr_data_ff[3:0];
    end
  end
  always @(posedge pic_pri_c1_clk or posedge reset) begin
    if (reset) begin
      intpriority_reg_19 <= 4'h0;
    end else if (intpriority_reg_we_19) begin
      intpriority_reg_19 <= picm_wr_data_ff[3:0];
    end
  end
  always @(posedge pic_pri_c1_clk or posedge reset) begin
    if (reset) begin
      intpriority_reg_20 <= 4'h0;
    end else if (intpriority_reg_we_20) begin
      intpriority_reg_20 <= picm_wr_data_ff[3:0];
    end
  end
  always @(posedge pic_pri_c1_clk or posedge reset) begin
    if (reset) begin
      intpriority_reg_21 <= 4'h0;
    end else if (intpriority_reg_we_21) begin
      intpriority_reg_21 <= picm_wr_data_ff[3:0];
    end
  end
  always @(posedge pic_pri_c1_clk or posedge reset) begin
    if (reset) begin
      intpriority_reg_22 <= 4'h0;
    end else if (intpriority_reg_we_22) begin
      intpriority_reg_22 <= picm_wr_data_ff[3:0];
    end
  end
  always @(posedge pic_pri_c1_clk or posedge reset) begin
    if (reset) begin
      intpriority_reg_23 <= 4'h0;
    end else if (intpriority_reg_we_23) begin
      intpriority_reg_23 <= picm_wr_data_ff[3:0];
    end
  end
  always @(posedge pic_pri_c1_clk or posedge reset) begin
    if (reset) begin
      intpriority_reg_24 <= 4'h0;
    end else if (intpriority_reg_we_24) begin
      intpriority_reg_24 <= picm_wr_data_ff[3:0];
    end
  end
  always @(posedge pic_pri_c1_clk or posedge reset) begin
    if (reset) begin
      intpriority_reg_25 <= 4'h0;
    end else if (intpriority_reg_we_25) begin
      intpriority_reg_25 <= picm_wr_data_ff[3:0];
    end
  end
  always @(posedge pic_pri_c1_clk or posedge reset) begin
    if (reset) begin
      intpriority_reg_26 <= 4'h0;
    end else if (intpriority_reg_we_26) begin
      intpriority_reg_26 <= picm_wr_data_ff[3:0];
    end
  end
  always @(posedge pic_pri_c1_clk or posedge reset) begin
    if (reset) begin
      intpriority_reg_27 <= 4'h0;
    end else if (intpriority_reg_we_27) begin
      intpriority_reg_27 <= picm_wr_data_ff[3:0];
    end
  end
  always @(posedge pic_pri_c1_clk or posedge reset) begin
    if (reset) begin
      intpriority_reg_28 <= 4'h0;
    end else if (intpriority_reg_we_28) begin
      intpriority_reg_28 <= picm_wr_data_ff[3:0];
    end
  end
  always @(posedge pic_pri_c1_clk or posedge reset) begin
    if (reset) begin
      intpriority_reg_29 <= 4'h0;
    end else if (intpriority_reg_we_29) begin
      intpriority_reg_29 <= picm_wr_data_ff[3:0];
    end
  end
  always @(posedge pic_pri_c1_clk or posedge reset) begin
    if (reset) begin
      intpriority_reg_30 <= 4'h0;
    end else if (intpriority_reg_we_30) begin
      intpriority_reg_30 <= picm_wr_data_ff[3:0];
    end
  end
  always @(posedge pic_pri_c1_clk or posedge reset) begin
    if (reset) begin
      intpriority_reg_31 <= 4'h0;
    end else if (intpriority_reg_we_31) begin
      intpriority_reg_31 <= picm_wr_data_ff[3:0];
    end
  end
  always @(posedge pic_int_c1_clk or posedge reset) begin
    if (reset) begin
      intenable_reg_1 <= 1'h0;
    end else if (intenable_reg_we_1) begin
      intenable_reg_1 <= picm_wr_data_ff[0];
    end
  end
  always @(posedge pic_int_c1_clk or posedge reset) begin
    if (reset) begin
      intenable_reg_2 <= 1'h0;
    end else if (intenable_reg_we_2) begin
      intenable_reg_2 <= picm_wr_data_ff[0];
    end
  end
  always @(posedge pic_int_c1_clk or posedge reset) begin
    if (reset) begin
      intenable_reg_3 <= 1'h0;
    end else if (intenable_reg_we_3) begin
      intenable_reg_3 <= picm_wr_data_ff[0];
    end
  end
  always @(posedge pic_int_c1_clk or posedge reset) begin
    if (reset) begin
      intenable_reg_4 <= 1'h0;
    end else if (intenable_reg_we_4) begin
      intenable_reg_4 <= picm_wr_data_ff[0];
    end
  end
  always @(posedge pic_int_c1_clk or posedge reset) begin
    if (reset) begin
      intenable_reg_5 <= 1'h0;
    end else if (intenable_reg_we_5) begin
      intenable_reg_5 <= picm_wr_data_ff[0];
    end
  end
  always @(posedge pic_int_c1_clk or posedge reset) begin
    if (reset) begin
      intenable_reg_6 <= 1'h0;
    end else if (intenable_reg_we_6) begin
      intenable_reg_6 <= picm_wr_data_ff[0];
    end
  end
  always @(posedge pic_int_c1_clk or posedge reset) begin
    if (reset) begin
      intenable_reg_7 <= 1'h0;
    end else if (intenable_reg_we_7) begin
      intenable_reg_7 <= picm_wr_data_ff[0];
    end
  end
  always @(posedge pic_int_c1_clk or posedge reset) begin
    if (reset) begin
      intenable_reg_8 <= 1'h0;
    end else if (intenable_reg_we_8) begin
      intenable_reg_8 <= picm_wr_data_ff[0];
    end
  end
  always @(posedge pic_int_c1_clk or posedge reset) begin
    if (reset) begin
      intenable_reg_9 <= 1'h0;
    end else if (intenable_reg_we_9) begin
      intenable_reg_9 <= picm_wr_data_ff[0];
    end
  end
  always @(posedge pic_int_c1_clk or posedge reset) begin
    if (reset) begin
      intenable_reg_10 <= 1'h0;
    end else if (intenable_reg_we_10) begin
      intenable_reg_10 <= picm_wr_data_ff[0];
    end
  end
  always @(posedge pic_int_c1_clk or posedge reset) begin
    if (reset) begin
      intenable_reg_11 <= 1'h0;
    end else if (intenable_reg_we_11) begin
      intenable_reg_11 <= picm_wr_data_ff[0];
    end
  end
  always @(posedge pic_int_c1_clk or posedge reset) begin
    if (reset) begin
      intenable_reg_12 <= 1'h0;
    end else if (intenable_reg_we_12) begin
      intenable_reg_12 <= picm_wr_data_ff[0];
    end
  end
  always @(posedge pic_int_c1_clk or posedge reset) begin
    if (reset) begin
      intenable_reg_13 <= 1'h0;
    end else if (intenable_reg_we_13) begin
      intenable_reg_13 <= picm_wr_data_ff[0];
    end
  end
  always @(posedge pic_int_c1_clk or posedge reset) begin
    if (reset) begin
      intenable_reg_14 <= 1'h0;
    end else if (intenable_reg_we_14) begin
      intenable_reg_14 <= picm_wr_data_ff[0];
    end
  end
  always @(posedge pic_int_c1_clk or posedge reset) begin
    if (reset) begin
      intenable_reg_15 <= 1'h0;
    end else if (intenable_reg_we_15) begin
      intenable_reg_15 <= picm_wr_data_ff[0];
    end
  end
  always @(posedge pic_int_c1_clk or posedge reset) begin
    if (reset) begin
      intenable_reg_16 <= 1'h0;
    end else if (intenable_reg_we_16) begin
      intenable_reg_16 <= picm_wr_data_ff[0];
    end
  end
  always @(posedge pic_int_c1_clk or posedge reset) begin
    if (reset) begin
      intenable_reg_17 <= 1'h0;
    end else if (intenable_reg_we_17) begin
      intenable_reg_17 <= picm_wr_data_ff[0];
    end
  end
  always @(posedge pic_int_c1_clk or posedge reset) begin
    if (reset) begin
      intenable_reg_18 <= 1'h0;
    end else if (intenable_reg_we_18) begin
      intenable_reg_18 <= picm_wr_data_ff[0];
    end
  end
  always @(posedge pic_int_c1_clk or posedge reset) begin
    if (reset) begin
      intenable_reg_19 <= 1'h0;
    end else if (intenable_reg_we_19) begin
      intenable_reg_19 <= picm_wr_data_ff[0];
    end
  end
  always @(posedge pic_int_c1_clk or posedge reset) begin
    if (reset) begin
      intenable_reg_20 <= 1'h0;
    end else if (intenable_reg_we_20) begin
      intenable_reg_20 <= picm_wr_data_ff[0];
    end
  end
  always @(posedge pic_int_c1_clk or posedge reset) begin
    if (reset) begin
      intenable_reg_21 <= 1'h0;
    end else if (intenable_reg_we_21) begin
      intenable_reg_21 <= picm_wr_data_ff[0];
    end
  end
  always @(posedge pic_int_c1_clk or posedge reset) begin
    if (reset) begin
      intenable_reg_22 <= 1'h0;
    end else if (intenable_reg_we_22) begin
      intenable_reg_22 <= picm_wr_data_ff[0];
    end
  end
  always @(posedge pic_int_c1_clk or posedge reset) begin
    if (reset) begin
      intenable_reg_23 <= 1'h0;
    end else if (intenable_reg_we_23) begin
      intenable_reg_23 <= picm_wr_data_ff[0];
    end
  end
  always @(posedge pic_int_c1_clk or posedge reset) begin
    if (reset) begin
      intenable_reg_24 <= 1'h0;
    end else if (intenable_reg_we_24) begin
      intenable_reg_24 <= picm_wr_data_ff[0];
    end
  end
  always @(posedge pic_int_c1_clk or posedge reset) begin
    if (reset) begin
      intenable_reg_25 <= 1'h0;
    end else if (intenable_reg_we_25) begin
      intenable_reg_25 <= picm_wr_data_ff[0];
    end
  end
  always @(posedge pic_int_c1_clk or posedge reset) begin
    if (reset) begin
      intenable_reg_26 <= 1'h0;
    end else if (intenable_reg_we_26) begin
      intenable_reg_26 <= picm_wr_data_ff[0];
    end
  end
  always @(posedge pic_int_c1_clk or posedge reset) begin
    if (reset) begin
      intenable_reg_27 <= 1'h0;
    end else if (intenable_reg_we_27) begin
      intenable_reg_27 <= picm_wr_data_ff[0];
    end
  end
  always @(posedge pic_int_c1_clk or posedge reset) begin
    if (reset) begin
      intenable_reg_28 <= 1'h0;
    end else if (intenable_reg_we_28) begin
      intenable_reg_28 <= picm_wr_data_ff[0];
    end
  end
  always @(posedge pic_int_c1_clk or posedge reset) begin
    if (reset) begin
      intenable_reg_29 <= 1'h0;
    end else if (intenable_reg_we_29) begin
      intenable_reg_29 <= picm_wr_data_ff[0];
    end
  end
  always @(posedge pic_int_c1_clk or posedge reset) begin
    if (reset) begin
      intenable_reg_30 <= 1'h0;
    end else if (intenable_reg_we_30) begin
      intenable_reg_30 <= picm_wr_data_ff[0];
    end
  end
  always @(posedge pic_int_c1_clk or posedge reset) begin
    if (reset) begin
      intenable_reg_31 <= 1'h0;
    end else if (intenable_reg_we_31) begin
      intenable_reg_31 <= picm_wr_data_ff[0];
    end
  end
  always @(posedge gw_config_c1_clk or posedge reset) begin
    if (reset) begin
      gw_config_reg_1 <= 2'h0;
    end else if (gw_config_reg_we_1) begin
      gw_config_reg_1 <= picm_wr_data_ff[1:0];
    end
  end
  always @(posedge gw_config_c1_clk or posedge reset) begin
    if (reset) begin
      gw_config_reg_2 <= 2'h0;
    end else if (gw_config_reg_we_2) begin
      gw_config_reg_2 <= picm_wr_data_ff[1:0];
    end
  end
  always @(posedge gw_config_c1_clk or posedge reset) begin
    if (reset) begin
      gw_config_reg_3 <= 2'h0;
    end else if (gw_config_reg_we_3) begin
      gw_config_reg_3 <= picm_wr_data_ff[1:0];
    end
  end
  always @(posedge gw_config_c1_clk or posedge reset) begin
    if (reset) begin
      gw_config_reg_4 <= 2'h0;
    end else if (gw_config_reg_we_4) begin
      gw_config_reg_4 <= picm_wr_data_ff[1:0];
    end
  end
  always @(posedge gw_config_c1_clk or posedge reset) begin
    if (reset) begin
      gw_config_reg_5 <= 2'h0;
    end else if (gw_config_reg_we_5) begin
      gw_config_reg_5 <= picm_wr_data_ff[1:0];
    end
  end
  always @(posedge gw_config_c1_clk or posedge reset) begin
    if (reset) begin
      gw_config_reg_6 <= 2'h0;
    end else if (gw_config_reg_we_6) begin
      gw_config_reg_6 <= picm_wr_data_ff[1:0];
    end
  end
  always @(posedge gw_config_c1_clk or posedge reset) begin
    if (reset) begin
      gw_config_reg_7 <= 2'h0;
    end else if (gw_config_reg_we_7) begin
      gw_config_reg_7 <= picm_wr_data_ff[1:0];
    end
  end
  always @(posedge gw_config_c1_clk or posedge reset) begin
    if (reset) begin
      gw_config_reg_8 <= 2'h0;
    end else if (gw_config_reg_we_8) begin
      gw_config_reg_8 <= picm_wr_data_ff[1:0];
    end
  end
  always @(posedge gw_config_c1_clk or posedge reset) begin
    if (reset) begin
      gw_config_reg_9 <= 2'h0;
    end else if (gw_config_reg_we_9) begin
      gw_config_reg_9 <= picm_wr_data_ff[1:0];
    end
  end
  always @(posedge gw_config_c1_clk or posedge reset) begin
    if (reset) begin
      gw_config_reg_10 <= 2'h0;
    end else if (gw_config_reg_we_10) begin
      gw_config_reg_10 <= picm_wr_data_ff[1:0];
    end
  end
  always @(posedge gw_config_c1_clk or posedge reset) begin
    if (reset) begin
      gw_config_reg_11 <= 2'h0;
    end else if (gw_config_reg_we_11) begin
      gw_config_reg_11 <= picm_wr_data_ff[1:0];
    end
  end
  always @(posedge gw_config_c1_clk or posedge reset) begin
    if (reset) begin
      gw_config_reg_12 <= 2'h0;
    end else if (gw_config_reg_we_12) begin
      gw_config_reg_12 <= picm_wr_data_ff[1:0];
    end
  end
  always @(posedge gw_config_c1_clk or posedge reset) begin
    if (reset) begin
      gw_config_reg_13 <= 2'h0;
    end else if (gw_config_reg_we_13) begin
      gw_config_reg_13 <= picm_wr_data_ff[1:0];
    end
  end
  always @(posedge gw_config_c1_clk or posedge reset) begin
    if (reset) begin
      gw_config_reg_14 <= 2'h0;
    end else if (gw_config_reg_we_14) begin
      gw_config_reg_14 <= picm_wr_data_ff[1:0];
    end
  end
  always @(posedge gw_config_c1_clk or posedge reset) begin
    if (reset) begin
      gw_config_reg_15 <= 2'h0;
    end else if (gw_config_reg_we_15) begin
      gw_config_reg_15 <= picm_wr_data_ff[1:0];
    end
  end
  always @(posedge gw_config_c1_clk or posedge reset) begin
    if (reset) begin
      gw_config_reg_16 <= 2'h0;
    end else if (gw_config_reg_we_16) begin
      gw_config_reg_16 <= picm_wr_data_ff[1:0];
    end
  end
  always @(posedge gw_config_c1_clk or posedge reset) begin
    if (reset) begin
      gw_config_reg_17 <= 2'h0;
    end else if (gw_config_reg_we_17) begin
      gw_config_reg_17 <= picm_wr_data_ff[1:0];
    end
  end
  always @(posedge gw_config_c1_clk or posedge reset) begin
    if (reset) begin
      gw_config_reg_18 <= 2'h0;
    end else if (gw_config_reg_we_18) begin
      gw_config_reg_18 <= picm_wr_data_ff[1:0];
    end
  end
  always @(posedge gw_config_c1_clk or posedge reset) begin
    if (reset) begin
      gw_config_reg_19 <= 2'h0;
    end else if (gw_config_reg_we_19) begin
      gw_config_reg_19 <= picm_wr_data_ff[1:0];
    end
  end
  always @(posedge gw_config_c1_clk or posedge reset) begin
    if (reset) begin
      gw_config_reg_20 <= 2'h0;
    end else if (gw_config_reg_we_20) begin
      gw_config_reg_20 <= picm_wr_data_ff[1:0];
    end
  end
  always @(posedge gw_config_c1_clk or posedge reset) begin
    if (reset) begin
      gw_config_reg_21 <= 2'h0;
    end else if (gw_config_reg_we_21) begin
      gw_config_reg_21 <= picm_wr_data_ff[1:0];
    end
  end
  always @(posedge gw_config_c1_clk or posedge reset) begin
    if (reset) begin
      gw_config_reg_22 <= 2'h0;
    end else if (gw_config_reg_we_22) begin
      gw_config_reg_22 <= picm_wr_data_ff[1:0];
    end
  end
  always @(posedge gw_config_c1_clk or posedge reset) begin
    if (reset) begin
      gw_config_reg_23 <= 2'h0;
    end else if (gw_config_reg_we_23) begin
      gw_config_reg_23 <= picm_wr_data_ff[1:0];
    end
  end
  always @(posedge gw_config_c1_clk or posedge reset) begin
    if (reset) begin
      gw_config_reg_24 <= 2'h0;
    end else if (gw_config_reg_we_24) begin
      gw_config_reg_24 <= picm_wr_data_ff[1:0];
    end
  end
  always @(posedge gw_config_c1_clk or posedge reset) begin
    if (reset) begin
      gw_config_reg_25 <= 2'h0;
    end else if (gw_config_reg_we_25) begin
      gw_config_reg_25 <= picm_wr_data_ff[1:0];
    end
  end
  always @(posedge gw_config_c1_clk or posedge reset) begin
    if (reset) begin
      gw_config_reg_26 <= 2'h0;
    end else if (gw_config_reg_we_26) begin
      gw_config_reg_26 <= picm_wr_data_ff[1:0];
    end
  end
  always @(posedge gw_config_c1_clk or posedge reset) begin
    if (reset) begin
      gw_config_reg_27 <= 2'h0;
    end else if (gw_config_reg_we_27) begin
      gw_config_reg_27 <= picm_wr_data_ff[1:0];
    end
  end
  always @(posedge gw_config_c1_clk or posedge reset) begin
    if (reset) begin
      gw_config_reg_28 <= 2'h0;
    end else if (gw_config_reg_we_28) begin
      gw_config_reg_28 <= picm_wr_data_ff[1:0];
    end
  end
  always @(posedge gw_config_c1_clk or posedge reset) begin
    if (reset) begin
      gw_config_reg_29 <= 2'h0;
    end else if (gw_config_reg_we_29) begin
      gw_config_reg_29 <= picm_wr_data_ff[1:0];
    end
  end
  always @(posedge gw_config_c1_clk or posedge reset) begin
    if (reset) begin
      gw_config_reg_30 <= 2'h0;
    end else if (gw_config_reg_we_30) begin
      gw_config_reg_30 <= picm_wr_data_ff[1:0];
    end
  end
  always @(posedge gw_config_c1_clk or posedge reset) begin
    if (reset) begin
      gw_config_reg_31 <= 2'h0;
    end else if (gw_config_reg_we_31) begin
      gw_config_reg_31 <= picm_wr_data_ff[1:0];
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      gw_int_pending <= 1'h0;
    end else begin
      gw_int_pending <= _T_970 | _T_972;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      gw_int_pending_1 <= 1'h0;
    end else begin
      gw_int_pending_1 <= _T_982 | _T_984;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      gw_int_pending_2 <= 1'h0;
    end else begin
      gw_int_pending_2 <= _T_994 | _T_996;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      gw_int_pending_3 <= 1'h0;
    end else begin
      gw_int_pending_3 <= _T_1006 | _T_1008;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      gw_int_pending_4 <= 1'h0;
    end else begin
      gw_int_pending_4 <= _T_1018 | _T_1020;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      gw_int_pending_5 <= 1'h0;
    end else begin
      gw_int_pending_5 <= _T_1030 | _T_1032;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      gw_int_pending_6 <= 1'h0;
    end else begin
      gw_int_pending_6 <= _T_1042 | _T_1044;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      gw_int_pending_7 <= 1'h0;
    end else begin
      gw_int_pending_7 <= _T_1054 | _T_1056;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      gw_int_pending_8 <= 1'h0;
    end else begin
      gw_int_pending_8 <= _T_1066 | _T_1068;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      gw_int_pending_9 <= 1'h0;
    end else begin
      gw_int_pending_9 <= _T_1078 | _T_1080;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      gw_int_pending_10 <= 1'h0;
    end else begin
      gw_int_pending_10 <= _T_1090 | _T_1092;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      gw_int_pending_11 <= 1'h0;
    end else begin
      gw_int_pending_11 <= _T_1102 | _T_1104;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      gw_int_pending_12 <= 1'h0;
    end else begin
      gw_int_pending_12 <= _T_1114 | _T_1116;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      gw_int_pending_13 <= 1'h0;
    end else begin
      gw_int_pending_13 <= _T_1126 | _T_1128;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      gw_int_pending_14 <= 1'h0;
    end else begin
      gw_int_pending_14 <= _T_1138 | _T_1140;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      gw_int_pending_15 <= 1'h0;
    end else begin
      gw_int_pending_15 <= _T_1150 | _T_1152;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      gw_int_pending_16 <= 1'h0;
    end else begin
      gw_int_pending_16 <= _T_1162 | _T_1164;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      gw_int_pending_17 <= 1'h0;
    end else begin
      gw_int_pending_17 <= _T_1174 | _T_1176;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      gw_int_pending_18 <= 1'h0;
    end else begin
      gw_int_pending_18 <= _T_1186 | _T_1188;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      gw_int_pending_19 <= 1'h0;
    end else begin
      gw_int_pending_19 <= _T_1198 | _T_1200;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      gw_int_pending_20 <= 1'h0;
    end else begin
      gw_int_pending_20 <= _T_1210 | _T_1212;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      gw_int_pending_21 <= 1'h0;
    end else begin
      gw_int_pending_21 <= _T_1222 | _T_1224;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      gw_int_pending_22 <= 1'h0;
    end else begin
      gw_int_pending_22 <= _T_1234 | _T_1236;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      gw_int_pending_23 <= 1'h0;
    end else begin
      gw_int_pending_23 <= _T_1246 | _T_1248;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      gw_int_pending_24 <= 1'h0;
    end else begin
      gw_int_pending_24 <= _T_1258 | _T_1260;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      gw_int_pending_25 <= 1'h0;
    end else begin
      gw_int_pending_25 <= _T_1270 | _T_1272;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      gw_int_pending_26 <= 1'h0;
    end else begin
      gw_int_pending_26 <= _T_1282 | _T_1284;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      gw_int_pending_27 <= 1'h0;
    end else begin
      gw_int_pending_27 <= _T_1294 | _T_1296;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      gw_int_pending_28 <= 1'h0;
    end else begin
      gw_int_pending_28 <= _T_1306 | _T_1308;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      gw_int_pending_29 <= 1'h0;
    end else begin
      gw_int_pending_29 <= _T_1318 | _T_1320;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      gw_int_pending_30 <= 1'h0;
    end else begin
      gw_int_pending_30 <= _T_1330 | _T_1332;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      config_reg <= 1'h0;
    end else if (config_reg_we) begin
      config_reg <= picm_wr_data_ff[0];
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      _T_1642 <= 8'h0;
    end else begin
      _T_1642 <= level_intpend_id_5_0;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      _T_1643 <= 4'h0;
    end else if (config_reg) begin
      _T_1643 <= _T_1641;
    end else begin
      _T_1643 <= level_intpend_w_prior_en_5_0;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      _T_1650 <= 1'h0;
    end else begin
      _T_1650 <= _T_1648 & _T_1649;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      _T_1652 <= 1'h0;
    end else begin
      _T_1652 <= pl_in_q == maxint;
    end
  end
endmodule
module dma_ctrl(
  input         clock,
  input         reset,
  input         io_free_clk,
  input         io_dma_bus_clk_en,
  input         io_clk_override,
  input         io_scan_mode,
  input  [1:0]  io_dbg_cmd_size,
  output [31:0] io_dma_dbg_rddata,
  output        io_dma_dbg_cmd_done,
  output        io_dma_dbg_cmd_fail,
  input         io_dbg_dma_dbg_ib_dbg_cmd_valid,
  input         io_dbg_dma_dbg_ib_dbg_cmd_write,
  input  [1:0]  io_dbg_dma_dbg_ib_dbg_cmd_type,
  input  [31:0] io_dbg_dma_dbg_ib_dbg_cmd_addr,
  input  [31:0] io_dbg_dma_dbg_dctl_dbg_cmd_wrdata,
  input         io_dbg_dma_io_dbg_dma_bubble,
  output        io_dbg_dma_io_dma_dbg_ready,
  output        io_dec_dma_dctl_dma_dma_dccm_stall_any,
  output        io_dec_dma_tlu_dma_dma_pmu_dccm_read,
  output        io_dec_dma_tlu_dma_dma_pmu_dccm_write,
  output        io_dec_dma_tlu_dma_dma_pmu_any_read,
  output        io_dec_dma_tlu_dma_dma_pmu_any_write,
  input  [2:0]  io_dec_dma_tlu_dma_dec_tlu_dma_qos_prty,
  output        io_dec_dma_tlu_dma_dma_dccm_stall_any,
  output        io_dec_dma_tlu_dma_dma_iccm_stall_any,
  input         io_iccm_dma_rvalid,
  input         io_iccm_dma_ecc_error,
  input  [2:0]  io_iccm_dma_rtag,
  input  [63:0] io_iccm_dma_rdata,
  input         io_iccm_ready,
  output        io_dma_axi_b_valid,
  output        io_dma_axi_r_valid,
  output [1:0]  io_dma_axi_r_bits_resp,
  output        io_lsu_dma_dma_lsc_ctl_dma_dccm_req,
  output [31:0] io_lsu_dma_dma_lsc_ctl_dma_mem_addr,
  output [2:0]  io_lsu_dma_dma_lsc_ctl_dma_mem_sz,
  output        io_lsu_dma_dma_lsc_ctl_dma_mem_write,
  output [63:0] io_lsu_dma_dma_lsc_ctl_dma_mem_wdata,
  output [31:0] io_lsu_dma_dma_dccm_ctl_dma_mem_addr,
  output [63:0] io_lsu_dma_dma_dccm_ctl_dma_mem_wdata,
  input         io_lsu_dma_dma_dccm_ctl_dccm_dma_rvalid,
  input         io_lsu_dma_dma_dccm_ctl_dccm_dma_ecc_error,
  input  [2:0]  io_lsu_dma_dma_dccm_ctl_dccm_dma_rtag,
  input  [63:0] io_lsu_dma_dma_dccm_ctl_dccm_dma_rdata,
  input         io_lsu_dma_dccm_ready,
  output [2:0]  io_lsu_dma_dma_mem_tag,
  output        io_ifu_dma_dma_ifc_dma_iccm_stall_any,
  output        io_ifu_dma_dma_mem_ctl_dma_iccm_req,
  output [31:0] io_ifu_dma_dma_mem_ctl_dma_mem_addr,
  output [2:0]  io_ifu_dma_dma_mem_ctl_dma_mem_sz,
  output        io_ifu_dma_dma_mem_ctl_dma_mem_write,
  output [63:0] io_ifu_dma_dma_mem_ctl_dma_mem_wdata,
  output [2:0]  io_ifu_dma_dma_mem_ctl_dma_mem_tag
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [63:0] _RAND_54;
  reg [63:0] _RAND_55;
  reg [63:0] _RAND_56;
  reg [63:0] _RAND_57;
  reg [63:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
`endif // RANDOMIZE_REG_INIT
  wire  rvclkhdr_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_1_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_1_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_1_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_1_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_2_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_2_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_2_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_2_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_3_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_3_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_3_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_3_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_4_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_4_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_4_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_4_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_5_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_5_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_5_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_5_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_6_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_6_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_6_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_6_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_7_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_7_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_7_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_7_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_8_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_8_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_8_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_8_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_9_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_9_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_9_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_9_io_scan_mode; // @[lib.scala 368:23]
  wire  dma_buffer_c1cgc_io_l1clk; // @[dma_ctrl.scala 389:32]
  wire  dma_buffer_c1cgc_io_clk; // @[dma_ctrl.scala 389:32]
  wire  dma_buffer_c1cgc_io_en; // @[dma_ctrl.scala 389:32]
  wire  dma_buffer_c1cgc_io_scan_mode; // @[dma_ctrl.scala 389:32]
  wire  dma_free_cgc_io_l1clk; // @[dma_ctrl.scala 395:28]
  wire  dma_free_cgc_io_clk; // @[dma_ctrl.scala 395:28]
  wire  dma_free_cgc_io_en; // @[dma_ctrl.scala 395:28]
  wire  dma_free_cgc_io_scan_mode; // @[dma_ctrl.scala 395:28]
  wire  dma_bus_cgc_io_l1clk; // @[dma_ctrl.scala 401:27]
  wire  dma_bus_cgc_io_clk; // @[dma_ctrl.scala 401:27]
  wire  dma_bus_cgc_io_en; // @[dma_ctrl.scala 401:27]
  wire  dma_bus_cgc_io_scan_mode; // @[dma_ctrl.scala 401:27]
  wire  rvclkhdr_10_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_10_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_10_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_10_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_11_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_11_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_11_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_11_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_12_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_12_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_12_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_12_io_scan_mode; // @[lib.scala 368:23]
  wire  dma_free_clk = dma_free_cgc_io_l1clk; // @[dma_ctrl.scala 168:26 dma_ctrl.scala 399:29]
  reg [2:0] RdPtr; // @[Reg.scala 27:20]
  reg [31:0] fifo_addr_4; // @[lib.scala 374:16]
  reg [31:0] fifo_addr_3; // @[lib.scala 374:16]
  reg [31:0] fifo_addr_2; // @[lib.scala 374:16]
  reg [31:0] fifo_addr_1; // @[lib.scala 374:16]
  reg [31:0] fifo_addr_0; // @[lib.scala 374:16]
  wire [31:0] _GEN_60 = 3'h1 == RdPtr ? fifo_addr_1 : fifo_addr_0; // @[dma_ctrl.scala 355:20]
  wire [31:0] _GEN_61 = 3'h2 == RdPtr ? fifo_addr_2 : _GEN_60; // @[dma_ctrl.scala 355:20]
  wire [31:0] _GEN_62 = 3'h3 == RdPtr ? fifo_addr_3 : _GEN_61; // @[dma_ctrl.scala 355:20]
  wire [31:0] dma_mem_addr_int = 3'h4 == RdPtr ? fifo_addr_4 : _GEN_62; // @[dma_ctrl.scala 355:20]
  wire  dma_mem_addr_in_dccm = dma_mem_addr_int[31:16] == 16'hf004; // @[lib.scala 361:39]
  wire  dma_mem_addr_in_pic = dma_mem_addr_int[31:15] == 17'h1e018; // @[lib.scala 361:39]
  wire  dma_mem_addr_in_iccm = dma_mem_addr_int[31:16] == 16'hee00; // @[lib.scala 361:39]
  wire  dma_bus_clk = dma_bus_cgc_io_l1clk; // @[dma_ctrl.scala 170:25 dma_ctrl.scala 405:28]
  wire [2:0] _GEN_90 = {{2'd0}, io_dbg_dma_dbg_ib_dbg_cmd_addr[2]}; // @[dma_ctrl.scala 195:91]
  wire [3:0] _T_17 = 3'h4 * _GEN_90; // @[dma_ctrl.scala 195:91]
  wire [18:0] _T_18 = 19'hf << _T_17; // @[dma_ctrl.scala 195:83]
  wire [18:0] _T_20 = io_dbg_dma_dbg_ib_dbg_cmd_valid ? _T_18 : 19'h0; // @[dma_ctrl.scala 195:34]
  wire [2:0] _T_23 = {1'h0,io_dbg_cmd_size}; // @[Cat.scala 29:58]
  wire [2:0] fifo_sz_in = io_dbg_dma_dbg_ib_dbg_cmd_valid ? _T_23 : 3'h0; // @[dma_ctrl.scala 197:33]
  wire  fifo_write_in = io_dbg_dma_dbg_ib_dbg_cmd_valid & io_dbg_dma_dbg_ib_dbg_cmd_write; // @[dma_ctrl.scala 199:33]
  reg  dbg_dma_bubble_bus; // @[dma_ctrl.scala 377:12]
  wire  _T_31 = io_dbg_dma_dbg_ib_dbg_cmd_valid & io_dbg_dma_dbg_ib_dbg_cmd_type[1]; // @[dma_ctrl.scala 206:136]
  reg [2:0] WrPtr; // @[Reg.scala 27:20]
  wire  _T_33 = 3'h0 == WrPtr; // @[dma_ctrl.scala 206:188]
  wire  _T_34 = _T_31 & _T_33; // @[dma_ctrl.scala 206:181]
  wire  _T_41 = 3'h1 == WrPtr; // @[dma_ctrl.scala 206:188]
  wire  _T_42 = _T_31 & _T_41; // @[dma_ctrl.scala 206:181]
  wire  _T_49 = 3'h2 == WrPtr; // @[dma_ctrl.scala 206:188]
  wire  _T_50 = _T_31 & _T_49; // @[dma_ctrl.scala 206:181]
  wire  _T_57 = 3'h3 == WrPtr; // @[dma_ctrl.scala 206:188]
  wire  _T_58 = _T_31 & _T_57; // @[dma_ctrl.scala 206:181]
  wire  _T_65 = 3'h4 == WrPtr; // @[dma_ctrl.scala 206:188]
  wire  _T_66 = _T_31 & _T_65; // @[dma_ctrl.scala 206:181]
  wire [4:0] fifo_cmd_en = {_T_66,_T_58,_T_50,_T_42,_T_34}; // @[Cat.scala 29:58]
  wire  _T_75 = _T_31 & io_dbg_dma_dbg_ib_dbg_cmd_write; // @[dma_ctrl.scala 208:181]
  wire  _T_78 = _T_75 & _T_33; // @[dma_ctrl.scala 208:217]
  reg  _T_598; // @[dma_ctrl.scala 226:82]
  reg  _T_591; // @[dma_ctrl.scala 226:82]
  reg  _T_584; // @[dma_ctrl.scala 226:82]
  reg  _T_577; // @[dma_ctrl.scala 226:82]
  reg  _T_570; // @[dma_ctrl.scala 226:82]
  wire [4:0] fifo_valid = {_T_598,_T_591,_T_584,_T_577,_T_570}; // @[Cat.scala 29:58]
  wire [4:0] _T_990 = fifo_valid >> RdPtr; // @[dma_ctrl.scala 303:38]
  reg  _T_760; // @[dma_ctrl.scala 234:89]
  reg  _T_753; // @[dma_ctrl.scala 234:89]
  reg  _T_746; // @[dma_ctrl.scala 234:89]
  reg  _T_739; // @[dma_ctrl.scala 234:89]
  reg  _T_732; // @[dma_ctrl.scala 234:89]
  wire [4:0] fifo_done = {_T_760,_T_753,_T_746,_T_739,_T_732}; // @[Cat.scala 29:58]
  wire [4:0] _T_992 = fifo_done >> RdPtr; // @[dma_ctrl.scala 303:58]
  wire  _T_994 = ~_T_992[0]; // @[dma_ctrl.scala 303:48]
  wire  _T_995 = _T_990[0] & _T_994; // @[dma_ctrl.scala 303:46]
  wire  dma_buffer_c1_clk = dma_buffer_c1cgc_io_l1clk; // @[dma_ctrl.scala 172:31 dma_ctrl.scala 393:33]
  reg  _T_886; // @[Reg.scala 27:20]
  reg  _T_884; // @[Reg.scala 27:20]
  reg  _T_882; // @[Reg.scala 27:20]
  reg  _T_880; // @[Reg.scala 27:20]
  reg  _T_878; // @[Reg.scala 27:20]
  wire [4:0] fifo_dbg = {_T_886,_T_884,_T_882,_T_880,_T_878}; // @[Cat.scala 29:58]
  wire [4:0] _T_996 = fifo_dbg >> RdPtr; // @[dma_ctrl.scala 303:77]
  wire  _T_998 = ~_T_996[0]; // @[dma_ctrl.scala 303:68]
  wire  _T_999 = _T_995 & _T_998; // @[dma_ctrl.scala 303:66]
  wire  _T_1000 = dma_mem_addr_in_dccm | dma_mem_addr_in_iccm; // @[dma_ctrl.scala 303:111]
  wire  _T_1001 = ~_T_1000; // @[dma_ctrl.scala 303:88]
  wire  dma_address_error = _T_999 & _T_1001; // @[dma_ctrl.scala 303:85]
  wire  _T_1009 = ~dma_address_error; // @[dma_ctrl.scala 304:68]
  wire  _T_1010 = _T_995 & _T_1009; // @[dma_ctrl.scala 304:66]
  reg [2:0] fifo_sz_4; // @[Reg.scala 27:20]
  reg [2:0] fifo_sz_3; // @[Reg.scala 27:20]
  reg [2:0] fifo_sz_2; // @[Reg.scala 27:20]
  reg [2:0] fifo_sz_1; // @[Reg.scala 27:20]
  reg [2:0] fifo_sz_0; // @[Reg.scala 27:20]
  wire [2:0] _GEN_65 = 3'h1 == RdPtr ? fifo_sz_1 : fifo_sz_0; // @[dma_ctrl.scala 356:20]
  wire [2:0] _GEN_66 = 3'h2 == RdPtr ? fifo_sz_2 : _GEN_65; // @[dma_ctrl.scala 356:20]
  wire [2:0] _GEN_67 = 3'h3 == RdPtr ? fifo_sz_3 : _GEN_66; // @[dma_ctrl.scala 356:20]
  wire [2:0] dma_mem_sz_int = 3'h4 == RdPtr ? fifo_sz_4 : _GEN_67; // @[dma_ctrl.scala 356:20]
  wire  _T_1012 = dma_mem_sz_int == 3'h1; // @[dma_ctrl.scala 305:28]
  wire  _T_1014 = _T_1012 & dma_mem_addr_int[0]; // @[dma_ctrl.scala 305:37]
  wire  _T_1016 = dma_mem_sz_int == 3'h2; // @[dma_ctrl.scala 306:29]
  wire  _T_1018 = |dma_mem_addr_int[1:0]; // @[dma_ctrl.scala 306:64]
  wire  _T_1019 = _T_1016 & _T_1018; // @[dma_ctrl.scala 306:38]
  wire  _T_1020 = _T_1014 | _T_1019; // @[dma_ctrl.scala 305:60]
  wire  _T_1022 = dma_mem_sz_int == 3'h3; // @[dma_ctrl.scala 307:29]
  wire  _T_1024 = |dma_mem_addr_int[2:0]; // @[dma_ctrl.scala 307:64]
  wire  _T_1025 = _T_1022 & _T_1024; // @[dma_ctrl.scala 307:38]
  wire  _T_1026 = _T_1020 | _T_1025; // @[dma_ctrl.scala 306:70]
  wire  _T_1028 = dma_mem_sz_int[1:0] == 2'h2; // @[dma_ctrl.scala 308:55]
  wire  _T_1030 = dma_mem_sz_int[1:0] == 2'h3; // @[dma_ctrl.scala 308:88]
  wire  _T_1031 = _T_1028 | _T_1030; // @[dma_ctrl.scala 308:64]
  wire  _T_1032 = ~_T_1031; // @[dma_ctrl.scala 308:31]
  wire  _T_1033 = dma_mem_addr_in_iccm & _T_1032; // @[dma_ctrl.scala 308:29]
  wire  _T_1034 = _T_1026 | _T_1033; // @[dma_ctrl.scala 307:70]
  wire  _T_1035 = dma_mem_addr_in_dccm & io_lsu_dma_dma_lsc_ctl_dma_mem_write; // @[dma_ctrl.scala 309:29]
  wire  _T_1042 = _T_1035 & _T_1032; // @[dma_ctrl.scala 309:68]
  wire  _T_1043 = _T_1034 | _T_1042; // @[dma_ctrl.scala 308:108]
  wire  _T_1046 = io_lsu_dma_dma_lsc_ctl_dma_mem_write & _T_1016; // @[dma_ctrl.scala 310:45]
  wire  _T_1048 = dma_mem_addr_int[2:0] == 3'h0; // @[dma_ctrl.scala 310:114]
  reg [7:0] fifo_byteen_4; // @[Reg.scala 27:20]
  reg [7:0] fifo_byteen_3; // @[Reg.scala 27:20]
  reg [7:0] fifo_byteen_2; // @[Reg.scala 27:20]
  reg [7:0] fifo_byteen_1; // @[Reg.scala 27:20]
  reg [7:0] fifo_byteen_0; // @[Reg.scala 27:20]
  wire [7:0] _GEN_70 = 3'h1 == RdPtr ? fifo_byteen_1 : fifo_byteen_0; // @[dma_ctrl.scala 359:20]
  wire [7:0] _GEN_71 = 3'h2 == RdPtr ? fifo_byteen_2 : _GEN_70; // @[dma_ctrl.scala 359:20]
  wire [7:0] _GEN_72 = 3'h3 == RdPtr ? fifo_byteen_3 : _GEN_71; // @[dma_ctrl.scala 359:20]
  wire [7:0] dma_mem_byteen = 3'h4 == RdPtr ? fifo_byteen_4 : _GEN_72; // @[dma_ctrl.scala 359:20]
  wire [3:0] _T_1071 = _T_1048 ? dma_mem_byteen[3:0] : 4'h0; // @[Mux.scala 27:72]
  wire  _T_1051 = dma_mem_addr_int[2:0] == 3'h1; // @[dma_ctrl.scala 311:32]
  wire [3:0] _T_1072 = _T_1051 ? dma_mem_byteen[4:1] : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_1079 = _T_1071 | _T_1072; // @[Mux.scala 27:72]
  wire  _T_1054 = dma_mem_addr_int[2:0] == 3'h2; // @[dma_ctrl.scala 312:32]
  wire [3:0] _T_1073 = _T_1054 ? dma_mem_byteen[5:2] : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_1080 = _T_1079 | _T_1073; // @[Mux.scala 27:72]
  wire  _T_1057 = dma_mem_addr_int[2:0] == 3'h3; // @[dma_ctrl.scala 313:32]
  wire [3:0] _T_1074 = _T_1057 ? dma_mem_byteen[6:3] : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_1081 = _T_1080 | _T_1074; // @[Mux.scala 27:72]
  wire  _T_1060 = dma_mem_addr_int[2:0] == 3'h4; // @[dma_ctrl.scala 314:32]
  wire [3:0] _T_1075 = _T_1060 ? dma_mem_byteen[7:4] : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_1082 = _T_1081 | _T_1075; // @[Mux.scala 27:72]
  wire  _T_1063 = dma_mem_addr_int[2:0] == 3'h5; // @[dma_ctrl.scala 315:32]
  wire [2:0] _T_1076 = _T_1063 ? dma_mem_byteen[7:5] : 3'h0; // @[Mux.scala 27:72]
  wire [3:0] _GEN_91 = {{1'd0}, _T_1076}; // @[Mux.scala 27:72]
  wire [3:0] _T_1083 = _T_1082 | _GEN_91; // @[Mux.scala 27:72]
  wire  _T_1066 = dma_mem_addr_int[2:0] == 3'h6; // @[dma_ctrl.scala 316:32]
  wire [1:0] _T_1077 = _T_1066 ? dma_mem_byteen[7:6] : 2'h0; // @[Mux.scala 27:72]
  wire [3:0] _GEN_92 = {{2'd0}, _T_1077}; // @[Mux.scala 27:72]
  wire [3:0] _T_1084 = _T_1083 | _GEN_92; // @[Mux.scala 27:72]
  wire  _T_1069 = dma_mem_addr_int[2:0] == 3'h7; // @[dma_ctrl.scala 317:32]
  wire  _T_1078 = _T_1069 & dma_mem_byteen[7]; // @[Mux.scala 27:72]
  wire [3:0] _GEN_93 = {{3'd0}, _T_1078}; // @[Mux.scala 27:72]
  wire [3:0] _T_1085 = _T_1084 | _GEN_93; // @[Mux.scala 27:72]
  wire  _T_1087 = _T_1085 != 4'hf; // @[dma_ctrl.scala 317:66]
  wire  _T_1088 = _T_1046 & _T_1087; // @[dma_ctrl.scala 310:78]
  wire  _T_1089 = _T_1043 | _T_1088; // @[dma_ctrl.scala 309:145]
  wire  _T_1092 = io_lsu_dma_dma_lsc_ctl_dma_mem_write & _T_1022; // @[dma_ctrl.scala 318:45]
  wire  _T_1094 = dma_mem_byteen == 8'hf; // @[dma_ctrl.scala 318:103]
  wire  _T_1096 = dma_mem_byteen == 8'hf0; // @[dma_ctrl.scala 318:139]
  wire  _T_1097 = _T_1094 | _T_1096; // @[dma_ctrl.scala 318:116]
  wire  _T_1099 = dma_mem_byteen == 8'hff; // @[dma_ctrl.scala 318:175]
  wire  _T_1100 = _T_1097 | _T_1099; // @[dma_ctrl.scala 318:152]
  wire  _T_1101 = ~_T_1100; // @[dma_ctrl.scala 318:80]
  wire  _T_1102 = _T_1092 & _T_1101; // @[dma_ctrl.scala 318:78]
  wire  _T_1103 = _T_1089 | _T_1102; // @[dma_ctrl.scala 317:79]
  wire  dma_alignment_error = _T_1010 & _T_1103; // @[dma_ctrl.scala 304:87]
  wire  _T_79 = dma_address_error | dma_alignment_error; // @[dma_ctrl.scala 208:258]
  wire  _T_80 = 3'h0 == RdPtr; // @[dma_ctrl.scala 208:288]
  wire  _T_81 = _T_79 & _T_80; // @[dma_ctrl.scala 208:281]
  wire  _T_82 = _T_78 | _T_81; // @[dma_ctrl.scala 208:236]
  wire  _T_83 = 3'h0 == io_lsu_dma_dma_dccm_ctl_dccm_dma_rtag; // @[dma_ctrl.scala 208:350]
  wire  _T_84 = io_lsu_dma_dma_dccm_ctl_dccm_dma_rvalid & _T_83; // @[dma_ctrl.scala 208:343]
  wire  _T_85 = _T_82 | _T_84; // @[dma_ctrl.scala 208:300]
  wire  _T_86 = 3'h0 == io_iccm_dma_rtag; // @[dma_ctrl.scala 208:423]
  wire  _T_87 = io_iccm_dma_rvalid & _T_86; // @[dma_ctrl.scala 208:416]
  wire  _T_88 = _T_85 | _T_87; // @[dma_ctrl.scala 208:394]
  wire  _T_96 = _T_75 & _T_41; // @[dma_ctrl.scala 208:217]
  wire  _T_98 = 3'h1 == RdPtr; // @[dma_ctrl.scala 208:288]
  wire  _T_99 = _T_79 & _T_98; // @[dma_ctrl.scala 208:281]
  wire  _T_100 = _T_96 | _T_99; // @[dma_ctrl.scala 208:236]
  wire  _T_101 = 3'h1 == io_lsu_dma_dma_dccm_ctl_dccm_dma_rtag; // @[dma_ctrl.scala 208:350]
  wire  _T_102 = io_lsu_dma_dma_dccm_ctl_dccm_dma_rvalid & _T_101; // @[dma_ctrl.scala 208:343]
  wire  _T_103 = _T_100 | _T_102; // @[dma_ctrl.scala 208:300]
  wire  _T_104 = 3'h1 == io_iccm_dma_rtag; // @[dma_ctrl.scala 208:423]
  wire  _T_105 = io_iccm_dma_rvalid & _T_104; // @[dma_ctrl.scala 208:416]
  wire  _T_106 = _T_103 | _T_105; // @[dma_ctrl.scala 208:394]
  wire  _T_114 = _T_75 & _T_49; // @[dma_ctrl.scala 208:217]
  wire  _T_116 = 3'h2 == RdPtr; // @[dma_ctrl.scala 208:288]
  wire  _T_117 = _T_79 & _T_116; // @[dma_ctrl.scala 208:281]
  wire  _T_118 = _T_114 | _T_117; // @[dma_ctrl.scala 208:236]
  wire  _T_119 = 3'h2 == io_lsu_dma_dma_dccm_ctl_dccm_dma_rtag; // @[dma_ctrl.scala 208:350]
  wire  _T_120 = io_lsu_dma_dma_dccm_ctl_dccm_dma_rvalid & _T_119; // @[dma_ctrl.scala 208:343]
  wire  _T_121 = _T_118 | _T_120; // @[dma_ctrl.scala 208:300]
  wire  _T_122 = 3'h2 == io_iccm_dma_rtag; // @[dma_ctrl.scala 208:423]
  wire  _T_123 = io_iccm_dma_rvalid & _T_122; // @[dma_ctrl.scala 208:416]
  wire  _T_124 = _T_121 | _T_123; // @[dma_ctrl.scala 208:394]
  wire  _T_132 = _T_75 & _T_57; // @[dma_ctrl.scala 208:217]
  wire  _T_134 = 3'h3 == RdPtr; // @[dma_ctrl.scala 208:288]
  wire  _T_135 = _T_79 & _T_134; // @[dma_ctrl.scala 208:281]
  wire  _T_136 = _T_132 | _T_135; // @[dma_ctrl.scala 208:236]
  wire  _T_137 = 3'h3 == io_lsu_dma_dma_dccm_ctl_dccm_dma_rtag; // @[dma_ctrl.scala 208:350]
  wire  _T_138 = io_lsu_dma_dma_dccm_ctl_dccm_dma_rvalid & _T_137; // @[dma_ctrl.scala 208:343]
  wire  _T_139 = _T_136 | _T_138; // @[dma_ctrl.scala 208:300]
  wire  _T_140 = 3'h3 == io_iccm_dma_rtag; // @[dma_ctrl.scala 208:423]
  wire  _T_141 = io_iccm_dma_rvalid & _T_140; // @[dma_ctrl.scala 208:416]
  wire  _T_142 = _T_139 | _T_141; // @[dma_ctrl.scala 208:394]
  wire  _T_150 = _T_75 & _T_65; // @[dma_ctrl.scala 208:217]
  wire  _T_152 = 3'h4 == RdPtr; // @[dma_ctrl.scala 208:288]
  wire  _T_153 = _T_79 & _T_152; // @[dma_ctrl.scala 208:281]
  wire  _T_154 = _T_150 | _T_153; // @[dma_ctrl.scala 208:236]
  wire  _T_155 = 3'h4 == io_lsu_dma_dma_dccm_ctl_dccm_dma_rtag; // @[dma_ctrl.scala 208:350]
  wire  _T_156 = io_lsu_dma_dma_dccm_ctl_dccm_dma_rvalid & _T_155; // @[dma_ctrl.scala 208:343]
  wire  _T_157 = _T_154 | _T_156; // @[dma_ctrl.scala 208:300]
  wire  _T_158 = 3'h4 == io_iccm_dma_rtag; // @[dma_ctrl.scala 208:423]
  wire  _T_159 = io_iccm_dma_rvalid & _T_158; // @[dma_ctrl.scala 208:416]
  wire  _T_160 = _T_157 | _T_159; // @[dma_ctrl.scala 208:394]
  wire [4:0] fifo_data_en = {_T_160,_T_142,_T_124,_T_106,_T_88}; // @[Cat.scala 29:58]
  wire  _T_165 = io_lsu_dma_dma_lsc_ctl_dma_dccm_req | io_ifu_dma_dma_mem_ctl_dma_iccm_req; // @[dma_ctrl.scala 210:95]
  wire  _T_166 = ~io_lsu_dma_dma_lsc_ctl_dma_mem_write; // @[dma_ctrl.scala 210:136]
  wire  _T_167 = _T_165 & _T_166; // @[dma_ctrl.scala 210:134]
  wire  _T_169 = _T_167 & _T_80; // @[dma_ctrl.scala 210:174]
  wire  _T_174 = _T_167 & _T_98; // @[dma_ctrl.scala 210:174]
  wire  _T_179 = _T_167 & _T_116; // @[dma_ctrl.scala 210:174]
  wire  _T_184 = _T_167 & _T_134; // @[dma_ctrl.scala 210:174]
  wire  _T_189 = _T_167 & _T_152; // @[dma_ctrl.scala 210:174]
  wire [4:0] fifo_pend_en = {_T_189,_T_184,_T_179,_T_174,_T_169}; // @[Cat.scala 29:58]
  wire  _T_1127 = _T_995 & _T_996[0]; // @[dma_ctrl.scala 328:66]
  wire  _T_1129 = _T_1000 | dma_mem_addr_in_pic; // @[dma_ctrl.scala 328:134]
  wire  _T_1130 = ~_T_1129; // @[dma_ctrl.scala 328:88]
  wire  _T_1133 = dma_mem_sz_int[1:0] != 2'h2; // @[dma_ctrl.scala 328:191]
  wire  _T_1134 = _T_1130 | _T_1133; // @[dma_ctrl.scala 328:167]
  wire  dma_dbg_cmd_error = _T_1127 & _T_1134; // @[dma_ctrl.scala 328:84]
  wire  _T_197 = _T_79 | dma_dbg_cmd_error; // @[dma_ctrl.scala 212:114]
  wire  _T_199 = _T_197 & _T_80; // @[dma_ctrl.scala 212:135]
  wire  _T_200 = io_lsu_dma_dma_dccm_ctl_dccm_dma_rvalid & io_lsu_dma_dma_dccm_ctl_dccm_dma_ecc_error; // @[dma_ctrl.scala 212:198]
  wire  _T_202 = _T_200 & _T_83; // @[dma_ctrl.scala 212:244]
  wire  _T_203 = _T_199 | _T_202; // @[dma_ctrl.scala 212:154]
  wire  _T_204 = io_iccm_dma_rvalid & io_iccm_dma_ecc_error; // @[dma_ctrl.scala 212:318]
  wire  _T_206 = _T_204 & _T_86; // @[dma_ctrl.scala 212:343]
  wire  _T_207 = _T_203 | _T_206; // @[dma_ctrl.scala 212:295]
  wire  _T_213 = _T_197 & _T_98; // @[dma_ctrl.scala 212:135]
  wire  _T_216 = _T_200 & _T_101; // @[dma_ctrl.scala 212:244]
  wire  _T_217 = _T_213 | _T_216; // @[dma_ctrl.scala 212:154]
  wire  _T_220 = _T_204 & _T_104; // @[dma_ctrl.scala 212:343]
  wire  _T_221 = _T_217 | _T_220; // @[dma_ctrl.scala 212:295]
  wire  _T_227 = _T_197 & _T_116; // @[dma_ctrl.scala 212:135]
  wire  _T_230 = _T_200 & _T_119; // @[dma_ctrl.scala 212:244]
  wire  _T_231 = _T_227 | _T_230; // @[dma_ctrl.scala 212:154]
  wire  _T_234 = _T_204 & _T_122; // @[dma_ctrl.scala 212:343]
  wire  _T_235 = _T_231 | _T_234; // @[dma_ctrl.scala 212:295]
  wire  _T_241 = _T_197 & _T_134; // @[dma_ctrl.scala 212:135]
  wire  _T_244 = _T_200 & _T_137; // @[dma_ctrl.scala 212:244]
  wire  _T_245 = _T_241 | _T_244; // @[dma_ctrl.scala 212:154]
  wire  _T_248 = _T_204 & _T_140; // @[dma_ctrl.scala 212:343]
  wire  _T_249 = _T_245 | _T_248; // @[dma_ctrl.scala 212:295]
  wire  _T_255 = _T_197 & _T_152; // @[dma_ctrl.scala 212:135]
  wire  _T_258 = _T_200 & _T_155; // @[dma_ctrl.scala 212:244]
  wire  _T_259 = _T_255 | _T_258; // @[dma_ctrl.scala 212:154]
  wire  _T_262 = _T_204 & _T_158; // @[dma_ctrl.scala 212:343]
  wire  _T_263 = _T_259 | _T_262; // @[dma_ctrl.scala 212:295]
  wire [4:0] fifo_error_en = {_T_263,_T_249,_T_235,_T_221,_T_207}; // @[Cat.scala 29:58]
  wire [1:0] _T_436 = {1'h0,io_lsu_dma_dma_dccm_ctl_dccm_dma_ecc_error}; // @[Cat.scala 29:58]
  wire [1:0] _T_439 = {1'h0,io_iccm_dma_ecc_error}; // @[Cat.scala 29:58]
  wire [1:0] _T_442 = {_T_197,dma_alignment_error}; // @[Cat.scala 29:58]
  wire [1:0] _T_443 = _T_87 ? _T_439 : _T_442; // @[dma_ctrl.scala 222:209]
  wire [1:0] fifo_error_in_0 = _T_84 ? _T_436 : _T_443; // @[dma_ctrl.scala 222:60]
  wire  _T_269 = |fifo_error_in_0; // @[dma_ctrl.scala 214:83]
  reg [1:0] fifo_error_0; // @[dma_ctrl.scala 228:85]
  wire  _T_272 = |fifo_error_0; // @[dma_ctrl.scala 214:125]
  wire [1:0] _T_454 = _T_105 ? _T_439 : _T_442; // @[dma_ctrl.scala 222:209]
  wire [1:0] fifo_error_in_1 = _T_102 ? _T_436 : _T_454; // @[dma_ctrl.scala 222:60]
  wire  _T_276 = |fifo_error_in_1; // @[dma_ctrl.scala 214:83]
  reg [1:0] fifo_error_1; // @[dma_ctrl.scala 228:85]
  wire  _T_279 = |fifo_error_1; // @[dma_ctrl.scala 214:125]
  wire [1:0] _T_465 = _T_123 ? _T_439 : _T_442; // @[dma_ctrl.scala 222:209]
  wire [1:0] fifo_error_in_2 = _T_120 ? _T_436 : _T_465; // @[dma_ctrl.scala 222:60]
  wire  _T_283 = |fifo_error_in_2; // @[dma_ctrl.scala 214:83]
  reg [1:0] fifo_error_2; // @[dma_ctrl.scala 228:85]
  wire  _T_286 = |fifo_error_2; // @[dma_ctrl.scala 214:125]
  wire [1:0] _T_476 = _T_141 ? _T_439 : _T_442; // @[dma_ctrl.scala 222:209]
  wire [1:0] fifo_error_in_3 = _T_138 ? _T_436 : _T_476; // @[dma_ctrl.scala 222:60]
  wire  _T_290 = |fifo_error_in_3; // @[dma_ctrl.scala 214:83]
  reg [1:0] fifo_error_3; // @[dma_ctrl.scala 228:85]
  wire  _T_293 = |fifo_error_3; // @[dma_ctrl.scala 214:125]
  wire [1:0] _T_487 = _T_159 ? _T_439 : _T_442; // @[dma_ctrl.scala 222:209]
  wire [1:0] fifo_error_in_4 = _T_156 ? _T_436 : _T_487; // @[dma_ctrl.scala 222:60]
  wire  _T_297 = |fifo_error_in_4; // @[dma_ctrl.scala 214:83]
  reg [1:0] fifo_error_4; // @[dma_ctrl.scala 228:85]
  wire  _T_300 = |fifo_error_4; // @[dma_ctrl.scala 214:125]
  wire  _T_309 = _T_272 | fifo_error_en[0]; // @[dma_ctrl.scala 216:78]
  wire  _T_311 = _T_165 & io_lsu_dma_dma_lsc_ctl_dma_mem_write; // @[dma_ctrl.scala 216:176]
  wire  _T_312 = _T_309 | _T_311; // @[dma_ctrl.scala 216:97]
  wire  _T_314 = _T_312 & _T_80; // @[dma_ctrl.scala 216:217]
  wire  _T_317 = _T_314 | _T_84; // @[dma_ctrl.scala 216:236]
  wire  _T_320 = _T_317 | _T_87; // @[dma_ctrl.scala 216:330]
  wire  _T_323 = _T_279 | fifo_error_en[1]; // @[dma_ctrl.scala 216:78]
  wire  _T_326 = _T_323 | _T_311; // @[dma_ctrl.scala 216:97]
  wire  _T_328 = _T_326 & _T_98; // @[dma_ctrl.scala 216:217]
  wire  _T_331 = _T_328 | _T_102; // @[dma_ctrl.scala 216:236]
  wire  _T_334 = _T_331 | _T_105; // @[dma_ctrl.scala 216:330]
  wire  _T_337 = _T_286 | fifo_error_en[2]; // @[dma_ctrl.scala 216:78]
  wire  _T_340 = _T_337 | _T_311; // @[dma_ctrl.scala 216:97]
  wire  _T_342 = _T_340 & _T_116; // @[dma_ctrl.scala 216:217]
  wire  _T_345 = _T_342 | _T_120; // @[dma_ctrl.scala 216:236]
  wire  _T_348 = _T_345 | _T_123; // @[dma_ctrl.scala 216:330]
  wire  _T_351 = _T_293 | fifo_error_en[3]; // @[dma_ctrl.scala 216:78]
  wire  _T_354 = _T_351 | _T_311; // @[dma_ctrl.scala 216:97]
  wire  _T_356 = _T_354 & _T_134; // @[dma_ctrl.scala 216:217]
  wire  _T_359 = _T_356 | _T_138; // @[dma_ctrl.scala 216:236]
  wire  _T_362 = _T_359 | _T_141; // @[dma_ctrl.scala 216:330]
  wire  _T_365 = _T_300 | fifo_error_en[4]; // @[dma_ctrl.scala 216:78]
  wire  _T_368 = _T_365 | _T_311; // @[dma_ctrl.scala 216:97]
  wire  _T_370 = _T_368 & _T_152; // @[dma_ctrl.scala 216:217]
  wire  _T_373 = _T_370 | _T_156; // @[dma_ctrl.scala 216:236]
  wire  _T_376 = _T_373 | _T_159; // @[dma_ctrl.scala 216:330]
  wire [4:0] fifo_done_en = {_T_376,_T_362,_T_348,_T_334,_T_320}; // @[Cat.scala 29:58]
  wire  _T_383 = fifo_done_en[0] | fifo_done[0]; // @[dma_ctrl.scala 218:75]
  wire  _T_384 = _T_383 & io_dma_bus_clk_en; // @[dma_ctrl.scala 218:91]
  wire  _T_387 = fifo_done_en[1] | fifo_done[1]; // @[dma_ctrl.scala 218:75]
  wire  _T_388 = _T_387 & io_dma_bus_clk_en; // @[dma_ctrl.scala 218:91]
  wire  _T_391 = fifo_done_en[2] | fifo_done[2]; // @[dma_ctrl.scala 218:75]
  wire  _T_392 = _T_391 & io_dma_bus_clk_en; // @[dma_ctrl.scala 218:91]
  wire  _T_395 = fifo_done_en[3] | fifo_done[3]; // @[dma_ctrl.scala 218:75]
  wire  _T_396 = _T_395 & io_dma_bus_clk_en; // @[dma_ctrl.scala 218:91]
  wire  _T_399 = fifo_done_en[4] | fifo_done[4]; // @[dma_ctrl.scala 218:75]
  wire  _T_400 = _T_399 & io_dma_bus_clk_en; // @[dma_ctrl.scala 218:91]
  wire [4:0] fifo_done_bus_en = {_T_400,_T_396,_T_392,_T_388,_T_384}; // @[Cat.scala 29:58]
  reg [2:0] RspPtr; // @[Reg.scala 27:20]
  wire  _T_408 = 3'h0 == RspPtr; // @[dma_ctrl.scala 220:150]
  wire  _T_409 = io_dma_dbg_cmd_done & _T_408; // @[dma_ctrl.scala 220:143]
  wire  _T_413 = 3'h1 == RspPtr; // @[dma_ctrl.scala 220:150]
  wire  _T_414 = io_dma_dbg_cmd_done & _T_413; // @[dma_ctrl.scala 220:143]
  wire  _T_418 = 3'h2 == RspPtr; // @[dma_ctrl.scala 220:150]
  wire  _T_419 = io_dma_dbg_cmd_done & _T_418; // @[dma_ctrl.scala 220:143]
  wire  _T_423 = 3'h3 == RspPtr; // @[dma_ctrl.scala 220:150]
  wire  _T_424 = io_dma_dbg_cmd_done & _T_423; // @[dma_ctrl.scala 220:143]
  wire  _T_428 = 3'h4 == RspPtr; // @[dma_ctrl.scala 220:150]
  wire  _T_429 = io_dma_dbg_cmd_done & _T_428; // @[dma_ctrl.scala 220:143]
  wire [4:0] fifo_reset = {_T_429,_T_424,_T_419,_T_414,_T_409}; // @[Cat.scala 29:58]
  wire  _T_491 = fifo_error_en[0] & _T_269; // @[dma_ctrl.scala 224:77]
  wire [63:0] _T_493 = {32'h0,fifo_addr_0}; // @[Cat.scala 29:58]
  wire [63:0] _T_498 = {io_dbg_dma_dbg_dctl_dbg_cmd_wrdata,io_dbg_dma_dbg_dctl_dbg_cmd_wrdata}; // @[Cat.scala 29:58]
  wire [63:0] _T_500 = io_dbg_dma_dbg_ib_dbg_cmd_valid ? _T_498 : 64'h0; // @[dma_ctrl.scala 224:347]
  wire  _T_506 = fifo_error_en[1] & _T_276; // @[dma_ctrl.scala 224:77]
  wire [63:0] _T_508 = {32'h0,fifo_addr_1}; // @[Cat.scala 29:58]
  wire  _T_521 = fifo_error_en[2] & _T_283; // @[dma_ctrl.scala 224:77]
  wire [63:0] _T_523 = {32'h0,fifo_addr_2}; // @[Cat.scala 29:58]
  wire  _T_536 = fifo_error_en[3] & _T_290; // @[dma_ctrl.scala 224:77]
  wire [63:0] _T_538 = {32'h0,fifo_addr_3}; // @[Cat.scala 29:58]
  wire  _T_551 = fifo_error_en[4] & _T_297; // @[dma_ctrl.scala 224:77]
  wire [63:0] _T_553 = {32'h0,fifo_addr_4}; // @[Cat.scala 29:58]
  wire  _T_566 = fifo_cmd_en[0] | fifo_valid[0]; // @[dma_ctrl.scala 226:86]
  wire  _T_568 = ~fifo_reset[0]; // @[dma_ctrl.scala 226:125]
  wire  _T_573 = fifo_cmd_en[1] | fifo_valid[1]; // @[dma_ctrl.scala 226:86]
  wire  _T_575 = ~fifo_reset[1]; // @[dma_ctrl.scala 226:125]
  wire  _T_580 = fifo_cmd_en[2] | fifo_valid[2]; // @[dma_ctrl.scala 226:86]
  wire  _T_582 = ~fifo_reset[2]; // @[dma_ctrl.scala 226:125]
  wire  _T_587 = fifo_cmd_en[3] | fifo_valid[3]; // @[dma_ctrl.scala 226:86]
  wire  _T_589 = ~fifo_reset[3]; // @[dma_ctrl.scala 226:125]
  wire  _T_594 = fifo_cmd_en[4] | fifo_valid[4]; // @[dma_ctrl.scala 226:86]
  wire  _T_596 = ~fifo_reset[4]; // @[dma_ctrl.scala 226:125]
  wire [1:0] _T_605 = fifo_error_en[0] ? fifo_error_in_0 : fifo_error_0; // @[dma_ctrl.scala 228:89]
  wire [1:0] _T_609 = _T_568 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [1:0] _T_614 = fifo_error_en[1] ? fifo_error_in_1 : fifo_error_1; // @[dma_ctrl.scala 228:89]
  wire [1:0] _T_618 = _T_575 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [1:0] _T_623 = fifo_error_en[2] ? fifo_error_in_2 : fifo_error_2; // @[dma_ctrl.scala 228:89]
  wire [1:0] _T_627 = _T_582 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [1:0] _T_632 = fifo_error_en[3] ? fifo_error_in_3 : fifo_error_3; // @[dma_ctrl.scala 228:89]
  wire [1:0] _T_636 = _T_589 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [1:0] _T_641 = fifo_error_en[4] ? fifo_error_in_4 : fifo_error_4; // @[dma_ctrl.scala 228:89]
  wire [1:0] _T_645 = _T_596 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  reg  _T_721; // @[dma_ctrl.scala 232:89]
  reg  _T_714; // @[dma_ctrl.scala 232:89]
  reg  _T_707; // @[dma_ctrl.scala 232:89]
  reg  _T_700; // @[dma_ctrl.scala 232:89]
  reg  _T_693; // @[dma_ctrl.scala 232:89]
  wire [4:0] fifo_rpend = {_T_721,_T_714,_T_707,_T_700,_T_693}; // @[Cat.scala 29:58]
  wire  _T_689 = fifo_pend_en[0] | fifo_rpend[0]; // @[dma_ctrl.scala 232:93]
  wire  _T_696 = fifo_pend_en[1] | fifo_rpend[1]; // @[dma_ctrl.scala 232:93]
  wire  _T_703 = fifo_pend_en[2] | fifo_rpend[2]; // @[dma_ctrl.scala 232:93]
  wire  _T_710 = fifo_pend_en[3] | fifo_rpend[3]; // @[dma_ctrl.scala 232:93]
  wire  _T_717 = fifo_pend_en[4] | fifo_rpend[4]; // @[dma_ctrl.scala 232:93]
  reg  _T_799; // @[dma_ctrl.scala 236:89]
  reg  _T_792; // @[dma_ctrl.scala 236:89]
  reg  _T_785; // @[dma_ctrl.scala 236:89]
  reg  _T_778; // @[dma_ctrl.scala 236:89]
  reg  _T_771; // @[dma_ctrl.scala 236:89]
  wire [4:0] fifo_done_bus = {_T_799,_T_792,_T_785,_T_778,_T_771}; // @[Cat.scala 29:58]
  wire  _T_767 = fifo_done_bus_en[0] | fifo_done_bus[0]; // @[dma_ctrl.scala 236:93]
  wire  _T_774 = fifo_done_bus_en[1] | fifo_done_bus[1]; // @[dma_ctrl.scala 236:93]
  wire  _T_781 = fifo_done_bus_en[2] | fifo_done_bus[2]; // @[dma_ctrl.scala 236:93]
  wire  _T_788 = fifo_done_bus_en[3] | fifo_done_bus[3]; // @[dma_ctrl.scala 236:93]
  wire  _T_795 = fifo_done_bus_en[4] | fifo_done_bus[4]; // @[dma_ctrl.scala 236:93]
  wire [7:0] fifo_byteen_in = _T_20[7:0]; // @[dma_ctrl.scala 195:28]
  reg  _T_850; // @[Reg.scala 27:20]
  reg  _T_852; // @[Reg.scala 27:20]
  reg  _T_854; // @[Reg.scala 27:20]
  reg  _T_856; // @[Reg.scala 27:20]
  reg  _T_858; // @[Reg.scala 27:20]
  wire [4:0] fifo_write = {_T_858,_T_856,_T_854,_T_852,_T_850}; // @[Cat.scala 29:58]
  reg [63:0] fifo_data_0; // @[lib.scala 374:16]
  reg [63:0] fifo_data_1; // @[lib.scala 374:16]
  reg [63:0] fifo_data_2; // @[lib.scala 374:16]
  reg [63:0] fifo_data_3; // @[lib.scala 374:16]
  reg [63:0] fifo_data_4; // @[lib.scala 374:16]
  wire  _T_931 = WrPtr == 3'h4; // @[dma_ctrl.scala 260:30]
  wire [2:0] _T_934 = WrPtr + 3'h1; // @[dma_ctrl.scala 260:76]
  wire  _T_936 = RdPtr == 3'h4; // @[dma_ctrl.scala 262:30]
  wire [2:0] _T_939 = RdPtr + 3'h1; // @[dma_ctrl.scala 262:76]
  wire  _T_941 = RspPtr == 3'h4; // @[dma_ctrl.scala 264:31]
  wire [2:0] _T_944 = RspPtr + 3'h1; // @[dma_ctrl.scala 264:78]
  wire  WrPtrEn = |fifo_cmd_en; // @[dma_ctrl.scala 266:30]
  wire  RdPtrEn = _T_165 | _T_197; // @[dma_ctrl.scala 268:93]
  wire  _T_1143 = |fifo_valid; // @[dma_ctrl.scala 338:30]
  wire  fifo_empty = ~_T_1143; // @[dma_ctrl.scala 338:17]
  wire [4:0] _T_1106 = fifo_valid >> RspPtr; // @[dma_ctrl.scala 324:39]
  wire [4:0] _T_1108 = fifo_dbg >> RspPtr; // @[dma_ctrl.scala 324:58]
  wire  _T_1110 = _T_1106[0] & _T_1108[0]; // @[dma_ctrl.scala 324:48]
  wire [4:0] _T_1111 = fifo_done >> RspPtr; // @[dma_ctrl.scala 324:78]
  wire [31:0] _GEN_44 = 3'h1 == RspPtr ? fifo_addr_1 : fifo_addr_0; // @[dma_ctrl.scala 325:49]
  wire [31:0] _GEN_45 = 3'h2 == RspPtr ? fifo_addr_2 : _GEN_44; // @[dma_ctrl.scala 325:49]
  wire [31:0] _GEN_46 = 3'h3 == RspPtr ? fifo_addr_3 : _GEN_45; // @[dma_ctrl.scala 325:49]
  wire [31:0] _GEN_47 = 3'h4 == RspPtr ? fifo_addr_4 : _GEN_46; // @[dma_ctrl.scala 325:49]
  wire [63:0] _GEN_49 = 3'h1 == RspPtr ? fifo_data_1 : fifo_data_0; // @[dma_ctrl.scala 325:71]
  wire [63:0] _GEN_50 = 3'h2 == RspPtr ? fifo_data_2 : _GEN_49; // @[dma_ctrl.scala 325:71]
  wire [63:0] _GEN_51 = 3'h3 == RspPtr ? fifo_data_3 : _GEN_50; // @[dma_ctrl.scala 325:71]
  wire [63:0] _GEN_52 = 3'h4 == RspPtr ? fifo_data_4 : _GEN_51; // @[dma_ctrl.scala 325:71]
  wire [1:0] _GEN_54 = 3'h1 == RspPtr ? fifo_error_1 : fifo_error_0; // @[dma_ctrl.scala 326:47]
  wire [1:0] _GEN_55 = 3'h2 == RspPtr ? fifo_error_2 : _GEN_54; // @[dma_ctrl.scala 326:47]
  wire [1:0] _GEN_56 = 3'h3 == RspPtr ? fifo_error_3 : _GEN_55; // @[dma_ctrl.scala 326:47]
  wire [1:0] _GEN_57 = 3'h4 == RspPtr ? fifo_error_4 : _GEN_56; // @[dma_ctrl.scala 326:47]
  wire  _T_1136 = dma_mem_addr_in_dccm | dma_mem_addr_in_pic; // @[dma_ctrl.scala 332:80]
  wire [4:0] _T_1165 = fifo_rpend >> RdPtr; // @[dma_ctrl.scala 351:54]
  wire  _T_1167 = ~_T_1165[0]; // @[dma_ctrl.scala 351:43]
  wire  _T_1168 = _T_990[0] & _T_1167; // @[dma_ctrl.scala 351:41]
  wire  _T_1172 = _T_1168 & _T_994; // @[dma_ctrl.scala 351:62]
  wire  _T_1175 = ~_T_197; // @[dma_ctrl.scala 351:84]
  wire  dma_mem_req = _T_1172 & _T_1175; // @[dma_ctrl.scala 351:82]
  wire  _T_1137 = dma_mem_req & _T_1136; // @[dma_ctrl.scala 332:56]
  reg [2:0] dma_nack_count; // @[Reg.scala 27:20]
  wire  _T_1138 = dma_nack_count >= io_dec_dma_tlu_dma_dec_tlu_dma_qos_prty; // @[dma_ctrl.scala 332:121]
  wire  _T_1140 = dma_mem_req & dma_mem_addr_in_iccm; // @[dma_ctrl.scala 333:56]
  wire  _T_1147 = ~_T_165; // @[dma_ctrl.scala 343:77]
  wire [2:0] _T_1149 = _T_1147 ? 3'h7 : 3'h0; // @[Bitwise.scala 72:12]
  wire [2:0] _T_1151 = _T_1149 & dma_nack_count; // @[dma_ctrl.scala 343:155]
  wire  _T_1155 = dma_mem_req & _T_1147; // @[dma_ctrl.scala 343:203]
  wire [2:0] _T_1158 = dma_nack_count + 3'h1; // @[dma_ctrl.scala 343:304]
  wire  _T_1184 = io_lsu_dma_dma_lsc_ctl_dma_mem_write & _T_1096; // @[dma_ctrl.scala 357:84]
  wire [31:0] _T_1188 = {dma_mem_addr_int[31:3],1'h1,dma_mem_addr_int[1:0]}; // @[Cat.scala 29:58]
  wire  _T_1196 = io_lsu_dma_dma_lsc_ctl_dma_mem_write & _T_1097; // @[dma_ctrl.scala 358:84]
  wire [4:0] _T_1199 = fifo_write >> RdPtr; // @[dma_ctrl.scala 360:53]
  wire [63:0] _GEN_75 = 3'h1 == RdPtr ? fifo_data_1 : fifo_data_0; // @[dma_ctrl.scala 361:40]
  wire [63:0] _GEN_76 = 3'h2 == RdPtr ? fifo_data_2 : _GEN_75; // @[dma_ctrl.scala 361:40]
  wire [63:0] _GEN_77 = 3'h3 == RdPtr ? fifo_data_3 : _GEN_76; // @[dma_ctrl.scala 361:40]
  reg  dma_dbg_cmd_done_q; // @[dma_ctrl.scala 381:12]
  wire  bus_rsp_valid = io_dma_axi_b_valid | io_dma_axi_r_valid; // @[dma_ctrl.scala 501:60]
  wire  _T_1215 = bus_rsp_valid | io_dbg_dma_dbg_ib_dbg_cmd_valid; // @[dma_ctrl.scala 387:60]
  wire  _T_1216 = _T_1215 | io_dma_dbg_cmd_done; // @[dma_ctrl.scala 387:94]
  wire  _T_1217 = _T_1216 | dma_dbg_cmd_done_q; // @[dma_ctrl.scala 387:116]
  wire  _T_1219 = _T_1217 | _T_1143; // @[dma_ctrl.scala 387:137]
  wire  _T_1271 = ~_T_1108[0]; // @[dma_ctrl.scala 481:50]
  wire  _T_1272 = _T_1106[0] & _T_1271; // @[dma_ctrl.scala 481:48]
  wire [4:0] _T_1273 = fifo_done_bus >> RspPtr; // @[dma_ctrl.scala 481:83]
  wire  axi_rsp_valid = _T_1272 & _T_1273[0]; // @[dma_ctrl.scala 481:68]
  wire [4:0] _T_1275 = fifo_write >> RspPtr; // @[dma_ctrl.scala 483:39]
  wire  axi_rsp_write = _T_1275[0]; // @[dma_ctrl.scala 483:39]
  wire [1:0] _T_1278 = _GEN_57[1] ? 2'h3 : 2'h0; // @[dma_ctrl.scala 484:64]
  wire  _T_1281 = ~axi_rsp_write; // @[dma_ctrl.scala 494:46]
  rvclkhdr rvclkhdr ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_io_l1clk),
    .io_clk(rvclkhdr_io_clk),
    .io_en(rvclkhdr_io_en),
    .io_scan_mode(rvclkhdr_io_scan_mode)
  );
  rvclkhdr rvclkhdr_1 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_1_io_l1clk),
    .io_clk(rvclkhdr_1_io_clk),
    .io_en(rvclkhdr_1_io_en),
    .io_scan_mode(rvclkhdr_1_io_scan_mode)
  );
  rvclkhdr rvclkhdr_2 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_2_io_l1clk),
    .io_clk(rvclkhdr_2_io_clk),
    .io_en(rvclkhdr_2_io_en),
    .io_scan_mode(rvclkhdr_2_io_scan_mode)
  );
  rvclkhdr rvclkhdr_3 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_3_io_l1clk),
    .io_clk(rvclkhdr_3_io_clk),
    .io_en(rvclkhdr_3_io_en),
    .io_scan_mode(rvclkhdr_3_io_scan_mode)
  );
  rvclkhdr rvclkhdr_4 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_4_io_l1clk),
    .io_clk(rvclkhdr_4_io_clk),
    .io_en(rvclkhdr_4_io_en),
    .io_scan_mode(rvclkhdr_4_io_scan_mode)
  );
  rvclkhdr rvclkhdr_5 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_5_io_l1clk),
    .io_clk(rvclkhdr_5_io_clk),
    .io_en(rvclkhdr_5_io_en),
    .io_scan_mode(rvclkhdr_5_io_scan_mode)
  );
  rvclkhdr rvclkhdr_6 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_6_io_l1clk),
    .io_clk(rvclkhdr_6_io_clk),
    .io_en(rvclkhdr_6_io_en),
    .io_scan_mode(rvclkhdr_6_io_scan_mode)
  );
  rvclkhdr rvclkhdr_7 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_7_io_l1clk),
    .io_clk(rvclkhdr_7_io_clk),
    .io_en(rvclkhdr_7_io_en),
    .io_scan_mode(rvclkhdr_7_io_scan_mode)
  );
  rvclkhdr rvclkhdr_8 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_8_io_l1clk),
    .io_clk(rvclkhdr_8_io_clk),
    .io_en(rvclkhdr_8_io_en),
    .io_scan_mode(rvclkhdr_8_io_scan_mode)
  );
  rvclkhdr rvclkhdr_9 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_9_io_l1clk),
    .io_clk(rvclkhdr_9_io_clk),
    .io_en(rvclkhdr_9_io_en),
    .io_scan_mode(rvclkhdr_9_io_scan_mode)
  );
  rvclkhdr dma_buffer_c1cgc ( // @[dma_ctrl.scala 389:32]
    .io_l1clk(dma_buffer_c1cgc_io_l1clk),
    .io_clk(dma_buffer_c1cgc_io_clk),
    .io_en(dma_buffer_c1cgc_io_en),
    .io_scan_mode(dma_buffer_c1cgc_io_scan_mode)
  );
  rvclkhdr dma_free_cgc ( // @[dma_ctrl.scala 395:28]
    .io_l1clk(dma_free_cgc_io_l1clk),
    .io_clk(dma_free_cgc_io_clk),
    .io_en(dma_free_cgc_io_en),
    .io_scan_mode(dma_free_cgc_io_scan_mode)
  );
  rvclkhdr dma_bus_cgc ( // @[dma_ctrl.scala 401:27]
    .io_l1clk(dma_bus_cgc_io_l1clk),
    .io_clk(dma_bus_cgc_io_clk),
    .io_en(dma_bus_cgc_io_en),
    .io_scan_mode(dma_bus_cgc_io_scan_mode)
  );
  rvclkhdr rvclkhdr_10 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_10_io_l1clk),
    .io_clk(rvclkhdr_10_io_clk),
    .io_en(rvclkhdr_10_io_en),
    .io_scan_mode(rvclkhdr_10_io_scan_mode)
  );
  rvclkhdr rvclkhdr_11 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_11_io_l1clk),
    .io_clk(rvclkhdr_11_io_clk),
    .io_en(rvclkhdr_11_io_en),
    .io_scan_mode(rvclkhdr_11_io_scan_mode)
  );
  rvclkhdr rvclkhdr_12 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_12_io_l1clk),
    .io_clk(rvclkhdr_12_io_clk),
    .io_en(rvclkhdr_12_io_en),
    .io_scan_mode(rvclkhdr_12_io_scan_mode)
  );
  assign io_dma_dbg_rddata = _GEN_47[2] ? _GEN_52[63:32] : _GEN_52[31:0]; // @[dma_ctrl.scala 325:25]
  assign io_dma_dbg_cmd_done = _T_1110 & _T_1111[0]; // @[dma_ctrl.scala 324:25]
  assign io_dma_dbg_cmd_fail = |_GEN_57; // @[dma_ctrl.scala 326:25]
  assign io_dbg_dma_io_dma_dbg_ready = fifo_empty & dbg_dma_bubble_bus; // @[dma_ctrl.scala 323:36]
  assign io_dec_dma_dctl_dma_dma_dccm_stall_any = io_dec_dma_tlu_dma_dma_dccm_stall_any; // @[dma_ctrl.scala 335:42]
  assign io_dec_dma_tlu_dma_dma_pmu_dccm_read = io_lsu_dma_dma_lsc_ctl_dma_dccm_req & _T_166; // @[dma_ctrl.scala 365:42]
  assign io_dec_dma_tlu_dma_dma_pmu_dccm_write = io_lsu_dma_dma_lsc_ctl_dma_dccm_req & io_lsu_dma_dma_lsc_ctl_dma_mem_write; // @[dma_ctrl.scala 366:42]
  assign io_dec_dma_tlu_dma_dma_pmu_any_read = _T_165 & _T_166; // @[dma_ctrl.scala 367:42]
  assign io_dec_dma_tlu_dma_dma_pmu_any_write = _T_165 & io_lsu_dma_dma_lsc_ctl_dma_mem_write; // @[dma_ctrl.scala 368:42]
  assign io_dec_dma_tlu_dma_dma_dccm_stall_any = _T_1137 & _T_1138; // @[dma_ctrl.scala 332:41]
  assign io_dec_dma_tlu_dma_dma_iccm_stall_any = io_ifu_dma_dma_ifc_dma_iccm_stall_any; // @[dma_ctrl.scala 334:41]
  assign io_dma_axi_b_valid = axi_rsp_valid & axi_rsp_write; // @[dma_ctrl.scala 490:27]
  assign io_dma_axi_r_valid = axi_rsp_valid & _T_1281; // @[dma_ctrl.scala 494:27]
  assign io_dma_axi_r_bits_resp = _GEN_57[0] ? 2'h2 : _T_1278; // @[dma_ctrl.scala 495:41]
  assign io_lsu_dma_dma_lsc_ctl_dma_dccm_req = _T_1137 & io_lsu_dma_dccm_ready; // @[dma_ctrl.scala 352:40]
  assign io_lsu_dma_dma_lsc_ctl_dma_mem_addr = _T_1184 ? _T_1188 : dma_mem_addr_int; // @[dma_ctrl.scala 357:40]
  assign io_lsu_dma_dma_lsc_ctl_dma_mem_sz = _T_1196 ? 3'h2 : dma_mem_sz_int; // @[dma_ctrl.scala 358:40]
  assign io_lsu_dma_dma_lsc_ctl_dma_mem_write = _T_1199[0]; // @[dma_ctrl.scala 360:40]
  assign io_lsu_dma_dma_lsc_ctl_dma_mem_wdata = 3'h4 == RdPtr ? fifo_data_4 : _GEN_77; // @[dma_ctrl.scala 361:40]
  assign io_lsu_dma_dma_dccm_ctl_dma_mem_addr = io_lsu_dma_dma_lsc_ctl_dma_mem_addr; // @[dma_ctrl.scala 503:40]
  assign io_lsu_dma_dma_dccm_ctl_dma_mem_wdata = io_lsu_dma_dma_lsc_ctl_dma_mem_wdata; // @[dma_ctrl.scala 504:41]
  assign io_lsu_dma_dma_mem_tag = RdPtr; // @[dma_ctrl.scala 354:28]
  assign io_ifu_dma_dma_ifc_dma_iccm_stall_any = _T_1140 & _T_1138; // @[dma_ctrl.scala 333:41]
  assign io_ifu_dma_dma_mem_ctl_dma_iccm_req = _T_1140 & io_iccm_ready; // @[dma_ctrl.scala 353:40]
  assign io_ifu_dma_dma_mem_ctl_dma_mem_addr = io_lsu_dma_dma_lsc_ctl_dma_mem_addr; // @[dma_ctrl.scala 506:39]
  assign io_ifu_dma_dma_mem_ctl_dma_mem_sz = io_lsu_dma_dma_lsc_ctl_dma_mem_sz; // @[dma_ctrl.scala 505:37]
  assign io_ifu_dma_dma_mem_ctl_dma_mem_write = io_lsu_dma_dma_lsc_ctl_dma_mem_write; // @[dma_ctrl.scala 508:40]
  assign io_ifu_dma_dma_mem_ctl_dma_mem_wdata = io_lsu_dma_dma_lsc_ctl_dma_mem_wdata; // @[dma_ctrl.scala 507:40]
  assign io_ifu_dma_dma_mem_ctl_dma_mem_tag = io_lsu_dma_dma_mem_tag; // @[dma_ctrl.scala 509:38]
  assign rvclkhdr_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_io_en = fifo_cmd_en[0]; // @[lib.scala 371:17]
  assign rvclkhdr_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_1_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_1_io_en = fifo_cmd_en[1]; // @[lib.scala 371:17]
  assign rvclkhdr_1_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_2_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_2_io_en = fifo_cmd_en[2]; // @[lib.scala 371:17]
  assign rvclkhdr_2_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_3_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_3_io_en = fifo_cmd_en[3]; // @[lib.scala 371:17]
  assign rvclkhdr_3_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_4_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_4_io_en = fifo_cmd_en[4]; // @[lib.scala 371:17]
  assign rvclkhdr_4_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_5_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_5_io_en = fifo_data_en[0]; // @[lib.scala 371:17]
  assign rvclkhdr_5_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_6_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_6_io_en = fifo_data_en[1]; // @[lib.scala 371:17]
  assign rvclkhdr_6_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_7_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_7_io_en = fifo_data_en[2]; // @[lib.scala 371:17]
  assign rvclkhdr_7_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_8_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_8_io_en = fifo_data_en[3]; // @[lib.scala 371:17]
  assign rvclkhdr_8_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_9_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_9_io_en = fifo_data_en[4]; // @[lib.scala 371:17]
  assign rvclkhdr_9_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign dma_buffer_c1cgc_io_clk = clock; // @[dma_ctrl.scala 392:33]
  assign dma_buffer_c1cgc_io_en = io_dbg_dma_dbg_ib_dbg_cmd_valid | io_clk_override; // @[dma_ctrl.scala 390:33]
  assign dma_buffer_c1cgc_io_scan_mode = io_scan_mode; // @[dma_ctrl.scala 391:33]
  assign dma_free_cgc_io_clk = clock; // @[dma_ctrl.scala 398:29]
  assign dma_free_cgc_io_en = _T_1219 | io_clk_override; // @[dma_ctrl.scala 396:29]
  assign dma_free_cgc_io_scan_mode = io_scan_mode; // @[dma_ctrl.scala 397:29]
  assign dma_bus_cgc_io_clk = clock; // @[dma_ctrl.scala 404:28]
  assign dma_bus_cgc_io_en = io_dma_bus_clk_en; // @[dma_ctrl.scala 402:28]
  assign dma_bus_cgc_io_scan_mode = io_scan_mode; // @[dma_ctrl.scala 403:28]
  assign rvclkhdr_10_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_10_io_en = 1'h0; // @[lib.scala 371:17]
  assign rvclkhdr_10_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_11_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_11_io_en = 1'h0; // @[lib.scala 371:17]
  assign rvclkhdr_11_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_12_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_12_io_en = 1'h0; // @[lib.scala 371:17]
  assign rvclkhdr_12_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  RdPtr = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  fifo_addr_4 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  fifo_addr_3 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  fifo_addr_2 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  fifo_addr_1 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  fifo_addr_0 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  dbg_dma_bubble_bus = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  WrPtr = _RAND_7[2:0];
  _RAND_8 = {1{`RANDOM}};
  _T_598 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  _T_591 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  _T_584 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  _T_577 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  _T_570 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  _T_760 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  _T_753 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  _T_746 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  _T_739 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  _T_732 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  _T_886 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  _T_884 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  _T_882 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  _T_880 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  _T_878 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  fifo_sz_4 = _RAND_23[2:0];
  _RAND_24 = {1{`RANDOM}};
  fifo_sz_3 = _RAND_24[2:0];
  _RAND_25 = {1{`RANDOM}};
  fifo_sz_2 = _RAND_25[2:0];
  _RAND_26 = {1{`RANDOM}};
  fifo_sz_1 = _RAND_26[2:0];
  _RAND_27 = {1{`RANDOM}};
  fifo_sz_0 = _RAND_27[2:0];
  _RAND_28 = {1{`RANDOM}};
  fifo_byteen_4 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  fifo_byteen_3 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  fifo_byteen_2 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  fifo_byteen_1 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  fifo_byteen_0 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  fifo_error_0 = _RAND_33[1:0];
  _RAND_34 = {1{`RANDOM}};
  fifo_error_1 = _RAND_34[1:0];
  _RAND_35 = {1{`RANDOM}};
  fifo_error_2 = _RAND_35[1:0];
  _RAND_36 = {1{`RANDOM}};
  fifo_error_3 = _RAND_36[1:0];
  _RAND_37 = {1{`RANDOM}};
  fifo_error_4 = _RAND_37[1:0];
  _RAND_38 = {1{`RANDOM}};
  RspPtr = _RAND_38[2:0];
  _RAND_39 = {1{`RANDOM}};
  _T_721 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  _T_714 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  _T_707 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  _T_700 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  _T_693 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  _T_799 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  _T_792 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  _T_785 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  _T_778 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  _T_771 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  _T_850 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  _T_852 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  _T_854 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  _T_856 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  _T_858 = _RAND_53[0:0];
  _RAND_54 = {2{`RANDOM}};
  fifo_data_0 = _RAND_54[63:0];
  _RAND_55 = {2{`RANDOM}};
  fifo_data_1 = _RAND_55[63:0];
  _RAND_56 = {2{`RANDOM}};
  fifo_data_2 = _RAND_56[63:0];
  _RAND_57 = {2{`RANDOM}};
  fifo_data_3 = _RAND_57[63:0];
  _RAND_58 = {2{`RANDOM}};
  fifo_data_4 = _RAND_58[63:0];
  _RAND_59 = {1{`RANDOM}};
  dma_nack_count = _RAND_59[2:0];
  _RAND_60 = {1{`RANDOM}};
  dma_dbg_cmd_done_q = _RAND_60[0:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    RdPtr = 3'h0;
  end
  if (reset) begin
    fifo_addr_4 = 32'h0;
  end
  if (reset) begin
    fifo_addr_3 = 32'h0;
  end
  if (reset) begin
    fifo_addr_2 = 32'h0;
  end
  if (reset) begin
    fifo_addr_1 = 32'h0;
  end
  if (reset) begin
    fifo_addr_0 = 32'h0;
  end
  if (reset) begin
    dbg_dma_bubble_bus = 1'h0;
  end
  if (reset) begin
    WrPtr = 3'h0;
  end
  if (reset) begin
    _T_598 = 1'h0;
  end
  if (reset) begin
    _T_591 = 1'h0;
  end
  if (reset) begin
    _T_584 = 1'h0;
  end
  if (reset) begin
    _T_577 = 1'h0;
  end
  if (reset) begin
    _T_570 = 1'h0;
  end
  if (reset) begin
    _T_760 = 1'h0;
  end
  if (reset) begin
    _T_753 = 1'h0;
  end
  if (reset) begin
    _T_746 = 1'h0;
  end
  if (reset) begin
    _T_739 = 1'h0;
  end
  if (reset) begin
    _T_732 = 1'h0;
  end
  if (reset) begin
    _T_886 = 1'h0;
  end
  if (reset) begin
    _T_884 = 1'h0;
  end
  if (reset) begin
    _T_882 = 1'h0;
  end
  if (reset) begin
    _T_880 = 1'h0;
  end
  if (reset) begin
    _T_878 = 1'h0;
  end
  if (reset) begin
    fifo_sz_4 = 3'h0;
  end
  if (reset) begin
    fifo_sz_3 = 3'h0;
  end
  if (reset) begin
    fifo_sz_2 = 3'h0;
  end
  if (reset) begin
    fifo_sz_1 = 3'h0;
  end
  if (reset) begin
    fifo_sz_0 = 3'h0;
  end
  if (reset) begin
    fifo_byteen_4 = 8'h0;
  end
  if (reset) begin
    fifo_byteen_3 = 8'h0;
  end
  if (reset) begin
    fifo_byteen_2 = 8'h0;
  end
  if (reset) begin
    fifo_byteen_1 = 8'h0;
  end
  if (reset) begin
    fifo_byteen_0 = 8'h0;
  end
  if (reset) begin
    fifo_error_0 = 2'h0;
  end
  if (reset) begin
    fifo_error_1 = 2'h0;
  end
  if (reset) begin
    fifo_error_2 = 2'h0;
  end
  if (reset) begin
    fifo_error_3 = 2'h0;
  end
  if (reset) begin
    fifo_error_4 = 2'h0;
  end
  if (reset) begin
    RspPtr = 3'h0;
  end
  if (reset) begin
    _T_721 = 1'h0;
  end
  if (reset) begin
    _T_714 = 1'h0;
  end
  if (reset) begin
    _T_707 = 1'h0;
  end
  if (reset) begin
    _T_700 = 1'h0;
  end
  if (reset) begin
    _T_693 = 1'h0;
  end
  if (reset) begin
    _T_799 = 1'h0;
  end
  if (reset) begin
    _T_792 = 1'h0;
  end
  if (reset) begin
    _T_785 = 1'h0;
  end
  if (reset) begin
    _T_778 = 1'h0;
  end
  if (reset) begin
    _T_771 = 1'h0;
  end
  if (reset) begin
    _T_850 = 1'h0;
  end
  if (reset) begin
    _T_852 = 1'h0;
  end
  if (reset) begin
    _T_854 = 1'h0;
  end
  if (reset) begin
    _T_856 = 1'h0;
  end
  if (reset) begin
    _T_858 = 1'h0;
  end
  if (reset) begin
    fifo_data_0 = 64'h0;
  end
  if (reset) begin
    fifo_data_1 = 64'h0;
  end
  if (reset) begin
    fifo_data_2 = 64'h0;
  end
  if (reset) begin
    fifo_data_3 = 64'h0;
  end
  if (reset) begin
    fifo_data_4 = 64'h0;
  end
  if (reset) begin
    dma_nack_count = 3'h0;
  end
  if (reset) begin
    dma_dbg_cmd_done_q = 1'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge dma_free_clk or posedge reset) begin
    if (reset) begin
      RdPtr <= 3'h0;
    end else if (RdPtrEn) begin
      if (_T_936) begin
        RdPtr <= 3'h0;
      end else begin
        RdPtr <= _T_939;
      end
    end
  end
  always @(posedge rvclkhdr_4_io_l1clk or posedge reset) begin
    if (reset) begin
      fifo_addr_4 <= 32'h0;
    end else if (io_dbg_dma_dbg_ib_dbg_cmd_valid) begin
      fifo_addr_4 <= io_dbg_dma_dbg_ib_dbg_cmd_addr;
    end else begin
      fifo_addr_4 <= 32'h0;
    end
  end
  always @(posedge rvclkhdr_3_io_l1clk or posedge reset) begin
    if (reset) begin
      fifo_addr_3 <= 32'h0;
    end else if (io_dbg_dma_dbg_ib_dbg_cmd_valid) begin
      fifo_addr_3 <= io_dbg_dma_dbg_ib_dbg_cmd_addr;
    end else begin
      fifo_addr_3 <= 32'h0;
    end
  end
  always @(posedge rvclkhdr_2_io_l1clk or posedge reset) begin
    if (reset) begin
      fifo_addr_2 <= 32'h0;
    end else if (io_dbg_dma_dbg_ib_dbg_cmd_valid) begin
      fifo_addr_2 <= io_dbg_dma_dbg_ib_dbg_cmd_addr;
    end else begin
      fifo_addr_2 <= 32'h0;
    end
  end
  always @(posedge rvclkhdr_1_io_l1clk or posedge reset) begin
    if (reset) begin
      fifo_addr_1 <= 32'h0;
    end else if (io_dbg_dma_dbg_ib_dbg_cmd_valid) begin
      fifo_addr_1 <= io_dbg_dma_dbg_ib_dbg_cmd_addr;
    end else begin
      fifo_addr_1 <= 32'h0;
    end
  end
  always @(posedge rvclkhdr_io_l1clk or posedge reset) begin
    if (reset) begin
      fifo_addr_0 <= 32'h0;
    end else if (io_dbg_dma_dbg_ib_dbg_cmd_valid) begin
      fifo_addr_0 <= io_dbg_dma_dbg_ib_dbg_cmd_addr;
    end else begin
      fifo_addr_0 <= 32'h0;
    end
  end
  always @(posedge dma_bus_clk or posedge reset) begin
    if (reset) begin
      dbg_dma_bubble_bus <= 1'h0;
    end else begin
      dbg_dma_bubble_bus <= io_dbg_dma_io_dbg_dma_bubble;
    end
  end
  always @(posedge dma_free_clk or posedge reset) begin
    if (reset) begin
      WrPtr <= 3'h0;
    end else if (WrPtrEn) begin
      if (_T_931) begin
        WrPtr <= 3'h0;
      end else begin
        WrPtr <= _T_934;
      end
    end
  end
  always @(posedge dma_free_clk or posedge reset) begin
    if (reset) begin
      _T_598 <= 1'h0;
    end else begin
      _T_598 <= _T_594 & _T_596;
    end
  end
  always @(posedge dma_free_clk or posedge reset) begin
    if (reset) begin
      _T_591 <= 1'h0;
    end else begin
      _T_591 <= _T_587 & _T_589;
    end
  end
  always @(posedge dma_free_clk or posedge reset) begin
    if (reset) begin
      _T_584 <= 1'h0;
    end else begin
      _T_584 <= _T_580 & _T_582;
    end
  end
  always @(posedge dma_free_clk or posedge reset) begin
    if (reset) begin
      _T_577 <= 1'h0;
    end else begin
      _T_577 <= _T_573 & _T_575;
    end
  end
  always @(posedge dma_free_clk or posedge reset) begin
    if (reset) begin
      _T_570 <= 1'h0;
    end else begin
      _T_570 <= _T_566 & _T_568;
    end
  end
  always @(posedge dma_free_clk or posedge reset) begin
    if (reset) begin
      _T_760 <= 1'h0;
    end else begin
      _T_760 <= _T_399 & _T_596;
    end
  end
  always @(posedge dma_free_clk or posedge reset) begin
    if (reset) begin
      _T_753 <= 1'h0;
    end else begin
      _T_753 <= _T_395 & _T_589;
    end
  end
  always @(posedge dma_free_clk or posedge reset) begin
    if (reset) begin
      _T_746 <= 1'h0;
    end else begin
      _T_746 <= _T_391 & _T_582;
    end
  end
  always @(posedge dma_free_clk or posedge reset) begin
    if (reset) begin
      _T_739 <= 1'h0;
    end else begin
      _T_739 <= _T_387 & _T_575;
    end
  end
  always @(posedge dma_free_clk or posedge reset) begin
    if (reset) begin
      _T_732 <= 1'h0;
    end else begin
      _T_732 <= _T_383 & _T_568;
    end
  end
  always @(posedge dma_buffer_c1_clk or posedge reset) begin
    if (reset) begin
      _T_886 <= 1'h0;
    end else if (fifo_cmd_en[4]) begin
      _T_886 <= io_dbg_dma_dbg_ib_dbg_cmd_valid;
    end
  end
  always @(posedge dma_buffer_c1_clk or posedge reset) begin
    if (reset) begin
      _T_884 <= 1'h0;
    end else if (fifo_cmd_en[3]) begin
      _T_884 <= io_dbg_dma_dbg_ib_dbg_cmd_valid;
    end
  end
  always @(posedge dma_buffer_c1_clk or posedge reset) begin
    if (reset) begin
      _T_882 <= 1'h0;
    end else if (fifo_cmd_en[2]) begin
      _T_882 <= io_dbg_dma_dbg_ib_dbg_cmd_valid;
    end
  end
  always @(posedge dma_buffer_c1_clk or posedge reset) begin
    if (reset) begin
      _T_880 <= 1'h0;
    end else if (fifo_cmd_en[1]) begin
      _T_880 <= io_dbg_dma_dbg_ib_dbg_cmd_valid;
    end
  end
  always @(posedge dma_buffer_c1_clk or posedge reset) begin
    if (reset) begin
      _T_878 <= 1'h0;
    end else if (fifo_cmd_en[0]) begin
      _T_878 <= io_dbg_dma_dbg_ib_dbg_cmd_valid;
    end
  end
  always @(posedge dma_buffer_c1_clk or posedge reset) begin
    if (reset) begin
      fifo_sz_4 <= 3'h0;
    end else if (fifo_cmd_en[4]) begin
      if (io_dbg_dma_dbg_ib_dbg_cmd_valid) begin
        fifo_sz_4 <= _T_23;
      end else begin
        fifo_sz_4 <= 3'h0;
      end
    end
  end
  always @(posedge dma_buffer_c1_clk or posedge reset) begin
    if (reset) begin
      fifo_sz_3 <= 3'h0;
    end else if (fifo_cmd_en[3]) begin
      if (io_dbg_dma_dbg_ib_dbg_cmd_valid) begin
        fifo_sz_3 <= _T_23;
      end else begin
        fifo_sz_3 <= 3'h0;
      end
    end
  end
  always @(posedge dma_buffer_c1_clk or posedge reset) begin
    if (reset) begin
      fifo_sz_2 <= 3'h0;
    end else if (fifo_cmd_en[2]) begin
      if (io_dbg_dma_dbg_ib_dbg_cmd_valid) begin
        fifo_sz_2 <= _T_23;
      end else begin
        fifo_sz_2 <= 3'h0;
      end
    end
  end
  always @(posedge dma_buffer_c1_clk or posedge reset) begin
    if (reset) begin
      fifo_sz_1 <= 3'h0;
    end else if (fifo_cmd_en[1]) begin
      if (io_dbg_dma_dbg_ib_dbg_cmd_valid) begin
        fifo_sz_1 <= _T_23;
      end else begin
        fifo_sz_1 <= 3'h0;
      end
    end
  end
  always @(posedge dma_buffer_c1_clk or posedge reset) begin
    if (reset) begin
      fifo_sz_0 <= 3'h0;
    end else if (fifo_cmd_en[0]) begin
      fifo_sz_0 <= fifo_sz_in;
    end
  end
  always @(posedge dma_buffer_c1_clk or posedge reset) begin
    if (reset) begin
      fifo_byteen_4 <= 8'h0;
    end else if (fifo_cmd_en[4]) begin
      fifo_byteen_4 <= fifo_byteen_in;
    end
  end
  always @(posedge dma_buffer_c1_clk or posedge reset) begin
    if (reset) begin
      fifo_byteen_3 <= 8'h0;
    end else if (fifo_cmd_en[3]) begin
      fifo_byteen_3 <= fifo_byteen_in;
    end
  end
  always @(posedge dma_buffer_c1_clk or posedge reset) begin
    if (reset) begin
      fifo_byteen_2 <= 8'h0;
    end else if (fifo_cmd_en[2]) begin
      fifo_byteen_2 <= fifo_byteen_in;
    end
  end
  always @(posedge dma_buffer_c1_clk or posedge reset) begin
    if (reset) begin
      fifo_byteen_1 <= 8'h0;
    end else if (fifo_cmd_en[1]) begin
      fifo_byteen_1 <= fifo_byteen_in;
    end
  end
  always @(posedge dma_buffer_c1_clk or posedge reset) begin
    if (reset) begin
      fifo_byteen_0 <= 8'h0;
    end else if (fifo_cmd_en[0]) begin
      fifo_byteen_0 <= fifo_byteen_in;
    end
  end
  always @(posedge dma_free_clk or posedge reset) begin
    if (reset) begin
      fifo_error_0 <= 2'h0;
    end else begin
      fifo_error_0 <= _T_605 & _T_609;
    end
  end
  always @(posedge dma_free_clk or posedge reset) begin
    if (reset) begin
      fifo_error_1 <= 2'h0;
    end else begin
      fifo_error_1 <= _T_614 & _T_618;
    end
  end
  always @(posedge dma_free_clk or posedge reset) begin
    if (reset) begin
      fifo_error_2 <= 2'h0;
    end else begin
      fifo_error_2 <= _T_623 & _T_627;
    end
  end
  always @(posedge dma_free_clk or posedge reset) begin
    if (reset) begin
      fifo_error_3 <= 2'h0;
    end else begin
      fifo_error_3 <= _T_632 & _T_636;
    end
  end
  always @(posedge dma_free_clk or posedge reset) begin
    if (reset) begin
      fifo_error_4 <= 2'h0;
    end else begin
      fifo_error_4 <= _T_641 & _T_645;
    end
  end
  always @(posedge dma_free_clk or posedge reset) begin
    if (reset) begin
      RspPtr <= 3'h0;
    end else if (io_dma_dbg_cmd_done) begin
      if (_T_941) begin
        RspPtr <= 3'h0;
      end else begin
        RspPtr <= _T_944;
      end
    end
  end
  always @(posedge dma_free_clk or posedge reset) begin
    if (reset) begin
      _T_721 <= 1'h0;
    end else begin
      _T_721 <= _T_717 & _T_596;
    end
  end
  always @(posedge dma_free_clk or posedge reset) begin
    if (reset) begin
      _T_714 <= 1'h0;
    end else begin
      _T_714 <= _T_710 & _T_589;
    end
  end
  always @(posedge dma_free_clk or posedge reset) begin
    if (reset) begin
      _T_707 <= 1'h0;
    end else begin
      _T_707 <= _T_703 & _T_582;
    end
  end
  always @(posedge dma_free_clk or posedge reset) begin
    if (reset) begin
      _T_700 <= 1'h0;
    end else begin
      _T_700 <= _T_696 & _T_575;
    end
  end
  always @(posedge dma_free_clk or posedge reset) begin
    if (reset) begin
      _T_693 <= 1'h0;
    end else begin
      _T_693 <= _T_689 & _T_568;
    end
  end
  always @(posedge dma_free_clk or posedge reset) begin
    if (reset) begin
      _T_799 <= 1'h0;
    end else begin
      _T_799 <= _T_795 & _T_596;
    end
  end
  always @(posedge dma_free_clk or posedge reset) begin
    if (reset) begin
      _T_792 <= 1'h0;
    end else begin
      _T_792 <= _T_788 & _T_589;
    end
  end
  always @(posedge dma_free_clk or posedge reset) begin
    if (reset) begin
      _T_785 <= 1'h0;
    end else begin
      _T_785 <= _T_781 & _T_582;
    end
  end
  always @(posedge dma_free_clk or posedge reset) begin
    if (reset) begin
      _T_778 <= 1'h0;
    end else begin
      _T_778 <= _T_774 & _T_575;
    end
  end
  always @(posedge dma_free_clk or posedge reset) begin
    if (reset) begin
      _T_771 <= 1'h0;
    end else begin
      _T_771 <= _T_767 & _T_568;
    end
  end
  always @(posedge dma_buffer_c1_clk or posedge reset) begin
    if (reset) begin
      _T_850 <= 1'h0;
    end else if (fifo_cmd_en[0]) begin
      _T_850 <= fifo_write_in;
    end
  end
  always @(posedge dma_buffer_c1_clk or posedge reset) begin
    if (reset) begin
      _T_852 <= 1'h0;
    end else if (fifo_cmd_en[1]) begin
      _T_852 <= fifo_write_in;
    end
  end
  always @(posedge dma_buffer_c1_clk or posedge reset) begin
    if (reset) begin
      _T_854 <= 1'h0;
    end else if (fifo_cmd_en[2]) begin
      _T_854 <= fifo_write_in;
    end
  end
  always @(posedge dma_buffer_c1_clk or posedge reset) begin
    if (reset) begin
      _T_856 <= 1'h0;
    end else if (fifo_cmd_en[3]) begin
      _T_856 <= fifo_write_in;
    end
  end
  always @(posedge dma_buffer_c1_clk or posedge reset) begin
    if (reset) begin
      _T_858 <= 1'h0;
    end else if (fifo_cmd_en[4]) begin
      _T_858 <= fifo_write_in;
    end
  end
  always @(posedge rvclkhdr_5_io_l1clk or posedge reset) begin
    if (reset) begin
      fifo_data_0 <= 64'h0;
    end else if (_T_491) begin
      fifo_data_0 <= _T_493;
    end else if (_T_84) begin
      fifo_data_0 <= io_lsu_dma_dma_dccm_ctl_dccm_dma_rdata;
    end else if (_T_87) begin
      fifo_data_0 <= io_iccm_dma_rdata;
    end else if (io_dbg_dma_dbg_ib_dbg_cmd_valid) begin
      fifo_data_0 <= _T_498;
    end else begin
      fifo_data_0 <= 64'h0;
    end
  end
  always @(posedge rvclkhdr_6_io_l1clk or posedge reset) begin
    if (reset) begin
      fifo_data_1 <= 64'h0;
    end else if (_T_506) begin
      fifo_data_1 <= _T_508;
    end else if (_T_102) begin
      fifo_data_1 <= io_lsu_dma_dma_dccm_ctl_dccm_dma_rdata;
    end else if (_T_105) begin
      fifo_data_1 <= io_iccm_dma_rdata;
    end else if (io_dbg_dma_dbg_ib_dbg_cmd_valid) begin
      fifo_data_1 <= _T_498;
    end else begin
      fifo_data_1 <= 64'h0;
    end
  end
  always @(posedge rvclkhdr_7_io_l1clk or posedge reset) begin
    if (reset) begin
      fifo_data_2 <= 64'h0;
    end else if (_T_521) begin
      fifo_data_2 <= _T_523;
    end else if (_T_120) begin
      fifo_data_2 <= io_lsu_dma_dma_dccm_ctl_dccm_dma_rdata;
    end else if (_T_123) begin
      fifo_data_2 <= io_iccm_dma_rdata;
    end else if (io_dbg_dma_dbg_ib_dbg_cmd_valid) begin
      fifo_data_2 <= _T_498;
    end else begin
      fifo_data_2 <= 64'h0;
    end
  end
  always @(posedge rvclkhdr_8_io_l1clk or posedge reset) begin
    if (reset) begin
      fifo_data_3 <= 64'h0;
    end else if (_T_536) begin
      fifo_data_3 <= _T_538;
    end else if (_T_138) begin
      fifo_data_3 <= io_lsu_dma_dma_dccm_ctl_dccm_dma_rdata;
    end else if (_T_141) begin
      fifo_data_3 <= io_iccm_dma_rdata;
    end else if (io_dbg_dma_dbg_ib_dbg_cmd_valid) begin
      fifo_data_3 <= _T_498;
    end else begin
      fifo_data_3 <= 64'h0;
    end
  end
  always @(posedge rvclkhdr_9_io_l1clk or posedge reset) begin
    if (reset) begin
      fifo_data_4 <= 64'h0;
    end else if (_T_551) begin
      fifo_data_4 <= _T_553;
    end else if (_T_156) begin
      fifo_data_4 <= io_lsu_dma_dma_dccm_ctl_dccm_dma_rdata;
    end else if (_T_159) begin
      fifo_data_4 <= io_iccm_dma_rdata;
    end else begin
      fifo_data_4 <= _T_500;
    end
  end
  always @(posedge dma_free_clk or posedge reset) begin
    if (reset) begin
      dma_nack_count <= 3'h0;
    end else if (dma_mem_req) begin
      if (_T_1138) begin
        dma_nack_count <= _T_1151;
      end else if (_T_1155) begin
        dma_nack_count <= _T_1158;
      end else begin
        dma_nack_count <= 3'h0;
      end
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      dma_dbg_cmd_done_q <= 1'h0;
    end else begin
      dma_dbg_cmd_done_q <= io_dma_dbg_cmd_done;
    end
  end
endmodule
module axi4_to_ahb(
  input         clock,
  input         reset,
  input         io_scan_mode,
  input         io_bus_clk_en,
  input         io_clk_override,
  output        io_axi_aw_ready,
  input         io_axi_aw_valid,
  input  [31:0] io_axi_aw_bits_addr,
  input  [2:0]  io_axi_aw_bits_size,
  output        io_axi_w_ready,
  input         io_axi_w_valid,
  input  [7:0]  io_axi_w_bits_strb,
  input         io_axi_b_ready,
  input         io_axi_ar_valid,
  input  [31:0] io_axi_ar_bits_addr,
  input  [2:0]  io_axi_ar_bits_size,
  input         io_ahb_in_hready,
  input         io_ahb_in_hresp,
  output [1:0]  io_ahb_out_htrans,
  output        io_ahb_out_hwrite
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
`endif // RANDOMIZE_REG_INIT
  wire  rvclkhdr_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_1_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_1_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_1_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_1_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_2_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_2_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_2_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_2_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_3_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_3_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_3_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_3_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_4_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_4_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_4_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_4_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_5_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_5_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_5_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_5_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_6_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_6_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_6_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_6_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_7_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_7_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_7_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_7_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_8_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_8_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_8_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_8_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_9_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_9_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_9_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_9_io_scan_mode; // @[lib.scala 343:22]
  wire  ahbm_clk = rvclkhdr_7_io_l1clk; // @[axi4_to_ahb.scala 31:22 axi4_to_ahb.scala 340:12]
  reg [2:0] buf_state; // @[axi4_to_ahb.scala 37:45]
  wire  _T_49 = 3'h0 == buf_state; // @[Conditional.scala 37:30]
  wire  bus_clk = rvclkhdr_io_l1clk; // @[axi4_to_ahb.scala 57:21 axi4_to_ahb.scala 169:11]
  reg  wrbuf_vld; // @[axi4_to_ahb.scala 308:51]
  reg  wrbuf_data_vld; // @[axi4_to_ahb.scala 309:51]
  wire  wr_cmd_vld = wrbuf_vld & wrbuf_data_vld; // @[axi4_to_ahb.scala 146:27]
  wire  master_valid = wr_cmd_vld | io_axi_ar_valid; // @[axi4_to_ahb.scala 147:30]
  wire  _T_101 = 3'h1 == buf_state; // @[Conditional.scala 37:30]
  reg  ahb_hready_q; // @[axi4_to_ahb.scala 328:52]
  reg [1:0] ahb_htrans_q; // @[axi4_to_ahb.scala 329:52]
  wire  _T_108 = ahb_htrans_q != 2'h0; // @[axi4_to_ahb.scala 190:58]
  wire  _T_109 = ahb_hready_q & _T_108; // @[axi4_to_ahb.scala 190:36]
  wire  ahbm_addr_clk = rvclkhdr_8_io_l1clk; // @[axi4_to_ahb.scala 32:27 axi4_to_ahb.scala 341:17]
  reg  ahb_hwrite_q; // @[axi4_to_ahb.scala 330:57]
  wire  _T_110 = ~ahb_hwrite_q; // @[axi4_to_ahb.scala 190:72]
  wire  _T_111 = _T_109 & _T_110; // @[axi4_to_ahb.scala 190:70]
  wire  _T_136 = 3'h6 == buf_state; // @[Conditional.scala 37:30]
  reg  ahb_hresp_q; // @[axi4_to_ahb.scala 331:52]
  wire  _T_156 = ahb_hready_q | ahb_hresp_q; // @[axi4_to_ahb.scala 204:37]
  wire  _T_175 = 3'h7 == buf_state; // @[Conditional.scala 37:30]
  wire  _T_186 = 3'h3 == buf_state; // @[Conditional.scala 37:30]
  wire  _T_188 = 3'h2 == buf_state; // @[Conditional.scala 37:30]
  wire  _T_189 = ahb_hready_q & ahb_hwrite_q; // @[axi4_to_ahb.scala 236:33]
  wire  _T_192 = _T_189 & _T_108; // @[axi4_to_ahb.scala 236:48]
  wire  _T_281 = 3'h4 == buf_state; // @[Conditional.scala 37:30]
  wire  _GEN_15 = _T_281 & _T_192; // @[Conditional.scala 39:67]
  wire  _GEN_19 = _T_188 ? _T_192 : _GEN_15; // @[Conditional.scala 39:67]
  wire  _GEN_40 = _T_186 ? 1'h0 : _GEN_19; // @[Conditional.scala 39:67]
  wire  _GEN_59 = _T_175 ? 1'h0 : _GEN_40; // @[Conditional.scala 39:67]
  wire  _GEN_79 = _T_136 ? 1'h0 : _GEN_59; // @[Conditional.scala 39:67]
  wire  _GEN_95 = _T_101 ? 1'h0 : _GEN_79; // @[Conditional.scala 39:67]
  wire  trxn_done = _T_49 ? 1'h0 : _GEN_95; // @[Conditional.scala 40:58]
  reg  cmd_doneQ; // @[axi4_to_ahb.scala 326:52]
  wire  _T_282 = cmd_doneQ & ahb_hready_q; // @[axi4_to_ahb.scala 246:34]
  wire  _T_283 = _T_282 | ahb_hresp_q; // @[axi4_to_ahb.scala 246:50]
  wire  _T_440 = 3'h5 == buf_state; // @[Conditional.scala 37:30]
  wire  _GEN_1 = _T_440 & io_axi_b_ready; // @[Conditional.scala 39:67]
  wire  _GEN_3 = _T_281 ? _T_283 : _GEN_1; // @[Conditional.scala 39:67]
  wire  _GEN_20 = _T_188 ? trxn_done : _GEN_3; // @[Conditional.scala 39:67]
  wire  _GEN_35 = _T_186 ? _T_156 : _GEN_20; // @[Conditional.scala 39:67]
  wire  _GEN_51 = _T_175 ? _T_111 : _GEN_35; // @[Conditional.scala 39:67]
  wire  _GEN_69 = _T_136 ? _T_156 : _GEN_51; // @[Conditional.scala 39:67]
  wire  _GEN_83 = _T_101 ? _T_111 : _GEN_69; // @[Conditional.scala 39:67]
  wire  buf_state_en = _T_49 ? master_valid : _GEN_83; // @[Conditional.scala 40:58]
  wire [1:0] _T_14 = wr_cmd_vld ? 2'h3 : 2'h0; // @[axi4_to_ahb.scala 149:20]
  wire [2:0] master_opc = {{1'd0}, _T_14}; // @[axi4_to_ahb.scala 149:14]
  wire  _T_51 = master_opc[2:1] == 2'h1; // @[axi4_to_ahb.scala 175:41]
  wire  _GEN_8 = _T_281 & _T_51; // @[Conditional.scala 39:67]
  wire  _GEN_29 = _T_188 ? 1'h0 : _GEN_8; // @[Conditional.scala 39:67]
  wire  _GEN_46 = _T_186 ? 1'h0 : _GEN_29; // @[Conditional.scala 39:67]
  wire  _GEN_63 = _T_175 ? 1'h0 : _GEN_46; // @[Conditional.scala 39:67]
  wire  _GEN_81 = _T_136 ? 1'h0 : _GEN_63; // @[Conditional.scala 39:67]
  wire  _GEN_97 = _T_101 ? 1'h0 : _GEN_81; // @[Conditional.scala 39:67]
  wire  buf_write_in = _T_49 ? _T_51 : _GEN_97; // @[Conditional.scala 40:58]
  wire [2:0] _T_53 = buf_write_in ? 3'h2 : 3'h1; // @[axi4_to_ahb.scala 176:26]
  wire  _T_103 = master_opc == 3'h0; // @[axi4_to_ahb.scala 189:61]
  wire  _T_104 = master_valid & _T_103; // @[axi4_to_ahb.scala 189:41]
  wire [2:0] _T_106 = _T_104 ? 3'h6 : 3'h3; // @[axi4_to_ahb.scala 189:26]
  wire  _T_124 = _T_106 == 3'h6; // @[axi4_to_ahb.scala 193:174]
  wire  _T_125 = _T_111 & _T_124; // @[axi4_to_ahb.scala 193:88]
  wire  _T_137 = ~ahb_hresp_q; // @[axi4_to_ahb.scala 201:39]
  wire  _T_138 = ahb_hready_q & _T_137; // @[axi4_to_ahb.scala 201:37]
  wire  _T_141 = master_valid & _T_51; // @[axi4_to_ahb.scala 201:70]
  wire  _T_142 = ~_T_141; // @[axi4_to_ahb.scala 201:55]
  wire  _T_143 = _T_138 & _T_142; // @[axi4_to_ahb.scala 201:53]
  wire  _T_285 = buf_state_en & _T_137; // @[axi4_to_ahb.scala 247:36]
  wire  _T_286 = _T_285 & io_axi_b_ready; // @[axi4_to_ahb.scala 247:51]
  wire  _GEN_4 = _T_281 & _T_286; // @[Conditional.scala 39:67]
  wire  _GEN_26 = _T_188 ? 1'h0 : _GEN_4; // @[Conditional.scala 39:67]
  wire  _GEN_45 = _T_186 ? 1'h0 : _GEN_26; // @[Conditional.scala 39:67]
  wire  _GEN_62 = _T_175 ? 1'h0 : _GEN_45; // @[Conditional.scala 39:67]
  wire  _GEN_66 = _T_136 ? _T_143 : _GEN_62; // @[Conditional.scala 39:67]
  wire  _GEN_86 = _T_101 ? _T_125 : _GEN_66; // @[Conditional.scala 39:67]
  wire  master_ready = _T_49 | _GEN_86; // @[Conditional.scala 40:58]
  wire  _T_149 = master_valid & master_ready; // @[axi4_to_ahb.scala 203:82]
  wire  _T_152 = _T_149 & _T_103; // @[axi4_to_ahb.scala 203:97]
  wire [2:0] _T_154 = _T_152 ? 3'h6 : 3'h3; // @[axi4_to_ahb.scala 203:67]
  wire [2:0] _T_155 = ahb_hresp_q ? 3'h7 : _T_154; // @[axi4_to_ahb.scala 203:26]
  wire  _T_287 = ~io_axi_b_ready; // @[axi4_to_ahb.scala 248:42]
  wire  _T_288 = ahb_hresp_q | _T_287; // @[axi4_to_ahb.scala 248:40]
  wire [2:0] _T_293 = _T_51 ? 3'h2 : 3'h1; // @[axi4_to_ahb.scala 248:99]
  wire [2:0] _T_294 = master_valid ? _T_293 : 3'h0; // @[axi4_to_ahb.scala 248:65]
  wire [2:0] _T_295 = _T_288 ? 3'h5 : _T_294; // @[axi4_to_ahb.scala 248:26]
  wire [2:0] _GEN_5 = _T_281 ? _T_295 : 3'h0; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_18 = _T_188 ? 3'h4 : _GEN_5; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_34 = _T_186 ? 3'h5 : _GEN_18; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_50 = _T_175 ? 3'h3 : _GEN_34; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_68 = _T_136 ? _T_155 : _GEN_50; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_82 = _T_101 ? _T_106 : _GEN_68; // @[Conditional.scala 39:67]
  wire [2:0] buf_nxtstate = _T_49 ? _T_53 : _GEN_82; // @[Conditional.scala 40:58]
  reg [31:0] wrbuf_addr; // @[lib.scala 374:16]
  wire [31:0] master_addr = wr_cmd_vld ? wrbuf_addr : io_axi_ar_bits_addr; // @[axi4_to_ahb.scala 150:21]
  reg [2:0] wrbuf_size; // @[Reg.scala 27:20]
  wire [2:0] master_size = wr_cmd_vld ? wrbuf_size : io_axi_ar_bits_size; // @[axi4_to_ahb.scala 151:21]
  reg [7:0] wrbuf_byteen; // @[Reg.scala 27:20]
  wire  _T_358 = buf_nxtstate != 3'h5; // @[axi4_to_ahb.scala 258:55]
  wire  _T_359 = buf_state_en & _T_358; // @[axi4_to_ahb.scala 258:39]
  wire  _GEN_14 = _T_281 ? _T_359 : _T_440; // @[Conditional.scala 39:67]
  wire  _GEN_33 = _T_188 ? 1'h0 : _GEN_14; // @[Conditional.scala 39:67]
  wire  _GEN_49 = _T_186 ? 1'h0 : _GEN_33; // @[Conditional.scala 39:67]
  wire  _GEN_52 = _T_175 ? buf_state_en : _GEN_49; // @[Conditional.scala 39:67]
  wire  _GEN_73 = _T_136 ? _T_285 : _GEN_52; // @[Conditional.scala 39:67]
  wire  _GEN_94 = _T_101 ? 1'h0 : _GEN_73; // @[Conditional.scala 39:67]
  wire  slave_valid_pre = _T_49 ? 1'h0 : _GEN_94; // @[Conditional.scala 40:58]
  wire  buf_clk = rvclkhdr_6_io_l1clk; // @[axi4_to_ahb.scala 125:21 axi4_to_ahb.scala 339:12]
  wire  _T_44 = io_axi_aw_valid & io_axi_aw_ready; // @[axi4_to_ahb.scala 167:57]
  wire  _T_45 = io_axi_w_valid & io_axi_w_ready; // @[axi4_to_ahb.scala 167:94]
  wire  _T_46 = _T_44 | _T_45; // @[axi4_to_ahb.scala 167:76]
  wire  _T_55 = buf_nxtstate == 3'h2; // @[axi4_to_ahb.scala 179:54]
  wire  _T_56 = buf_state_en & _T_55; // @[axi4_to_ahb.scala 179:38]
  wire  _T_96 = buf_nxtstate == 3'h1; // @[axi4_to_ahb.scala 184:51]
  wire  _T_126 = master_ready & master_valid; // @[axi4_to_ahb.scala 195:33]
  wire  _T_162 = buf_nxtstate == 3'h6; // @[axi4_to_ahb.scala 210:64]
  wire  _T_163 = _T_126 & _T_162; // @[axi4_to_ahb.scala 210:48]
  wire  _T_164 = _T_163 & buf_state_en; // @[axi4_to_ahb.scala 210:79]
  wire  _T_349 = buf_state_en & buf_write_in; // @[axi4_to_ahb.scala 256:33]
  wire  _T_351 = _T_349 & _T_55; // @[axi4_to_ahb.scala 256:48]
  wire  _GEN_12 = _T_281 & _T_351; // @[Conditional.scala 39:67]
  wire  _GEN_32 = _T_188 ? 1'h0 : _GEN_12; // @[Conditional.scala 39:67]
  wire  _GEN_48 = _T_186 ? 1'h0 : _GEN_32; // @[Conditional.scala 39:67]
  wire  _GEN_65 = _T_175 ? 1'h0 : _GEN_48; // @[Conditional.scala 39:67]
  wire  _GEN_75 = _T_136 ? _T_164 : _GEN_65; // @[Conditional.scala 39:67]
  wire  _GEN_88 = _T_101 ? _T_126 : _GEN_75; // @[Conditional.scala 39:67]
  wire  bypass_en = _T_49 ? buf_state_en : _GEN_88; // @[Conditional.scala 40:58]
  wire [1:0] _T_99 = bypass_en ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [1:0] _T_100 = _T_99 & 2'h2; // @[axi4_to_ahb.scala 185:49]
  wire  _T_112 = ~master_valid; // @[axi4_to_ahb.scala 191:34]
  wire  _T_113 = buf_state_en & _T_112; // @[axi4_to_ahb.scala 191:32]
  reg [31:0] buf_addr; // @[lib.scala 374:16]
  wire  _T_131 = ~buf_state_en; // @[axi4_to_ahb.scala 197:48]
  wire  _T_132 = _T_131 | bypass_en; // @[axi4_to_ahb.scala 197:62]
  wire [1:0] _T_134 = _T_132 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [1:0] _T_135 = 2'h2 & _T_134; // @[axi4_to_ahb.scala 197:36]
  wire  _T_169 = buf_nxtstate != 3'h6; // @[axi4_to_ahb.scala 212:63]
  wire  _T_170 = _T_169 & buf_state_en; // @[axi4_to_ahb.scala 212:78]
  wire  _T_171 = ~_T_170; // @[axi4_to_ahb.scala 212:47]
  wire [1:0] _T_173 = _T_171 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [1:0] _T_174 = 2'h2 & _T_173; // @[axi4_to_ahb.scala 212:36]
  wire [1:0] _T_184 = _T_131 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [1:0] _T_185 = 2'h2 & _T_184; // @[axi4_to_ahb.scala 222:41]
  reg [2:0] buf_cmd_byte_ptrQ; // @[Reg.scala 27:20]
  reg [7:0] buf_byteen; // @[Reg.scala 27:20]
  wire [2:0] _T_197 = buf_cmd_byte_ptrQ + 3'h1; // @[axi4_to_ahb.scala 142:52]
  wire  _T_200 = 3'h0 >= _T_197; // @[axi4_to_ahb.scala 143:62]
  wire  _T_201 = buf_byteen[0] & _T_200; // @[axi4_to_ahb.scala 143:48]
  wire  _T_203 = 3'h1 >= _T_197; // @[axi4_to_ahb.scala 143:62]
  wire  _T_204 = buf_byteen[1] & _T_203; // @[axi4_to_ahb.scala 143:48]
  wire  _T_206 = 3'h2 >= _T_197; // @[axi4_to_ahb.scala 143:62]
  wire  _T_207 = buf_byteen[2] & _T_206; // @[axi4_to_ahb.scala 143:48]
  wire  _T_209 = 3'h3 >= _T_197; // @[axi4_to_ahb.scala 143:62]
  wire  _T_210 = buf_byteen[3] & _T_209; // @[axi4_to_ahb.scala 143:48]
  wire  _T_212 = 3'h4 >= _T_197; // @[axi4_to_ahb.scala 143:62]
  wire  _T_213 = buf_byteen[4] & _T_212; // @[axi4_to_ahb.scala 143:48]
  wire  _T_215 = 3'h5 >= _T_197; // @[axi4_to_ahb.scala 143:62]
  wire  _T_216 = buf_byteen[5] & _T_215; // @[axi4_to_ahb.scala 143:48]
  wire  _T_218 = 3'h6 >= _T_197; // @[axi4_to_ahb.scala 143:62]
  wire  _T_219 = buf_byteen[6] & _T_218; // @[axi4_to_ahb.scala 143:48]
  wire [2:0] _T_224 = _T_219 ? 3'h6 : 3'h7; // @[Mux.scala 98:16]
  wire [2:0] _T_225 = _T_216 ? 3'h5 : _T_224; // @[Mux.scala 98:16]
  wire [2:0] _T_226 = _T_213 ? 3'h4 : _T_225; // @[Mux.scala 98:16]
  wire [2:0] _T_227 = _T_210 ? 3'h3 : _T_226; // @[Mux.scala 98:16]
  wire [2:0] _T_228 = _T_207 ? 3'h2 : _T_227; // @[Mux.scala 98:16]
  wire [2:0] _T_229 = _T_204 ? 3'h1 : _T_228; // @[Mux.scala 98:16]
  wire [2:0] _T_230 = _T_201 ? 3'h0 : _T_229; // @[Mux.scala 98:16]
  wire  _T_232 = buf_cmd_byte_ptrQ == 3'h7; // @[axi4_to_ahb.scala 241:65]
  reg  buf_aligned; // @[Reg.scala 27:20]
  wire  _T_233 = buf_aligned | _T_232; // @[axi4_to_ahb.scala 241:44]
  wire [7:0] _T_271 = buf_byteen >> _T_230; // @[axi4_to_ahb.scala 241:92]
  wire  _T_273 = ~_T_271[0]; // @[axi4_to_ahb.scala 241:163]
  wire  _T_274 = _T_233 | _T_273; // @[axi4_to_ahb.scala 241:79]
  wire  _T_275 = trxn_done & _T_274; // @[axi4_to_ahb.scala 241:29]
  wire  _T_346 = _T_232 | _T_273; // @[axi4_to_ahb.scala 255:38]
  wire  _T_347 = _T_109 & _T_346; // @[axi4_to_ahb.scala 254:80]
  wire  _T_348 = ahb_hresp_q | _T_347; // @[axi4_to_ahb.scala 254:34]
  wire  _GEN_11 = _T_281 & _T_348; // @[Conditional.scala 39:67]
  wire  _GEN_24 = _T_188 ? _T_275 : _GEN_11; // @[Conditional.scala 39:67]
  wire  _GEN_43 = _T_186 ? 1'h0 : _GEN_24; // @[Conditional.scala 39:67]
  wire  _GEN_61 = _T_175 ? 1'h0 : _GEN_43; // @[Conditional.scala 39:67]
  wire  _GEN_74 = _T_136 ? _T_113 : _GEN_61; // @[Conditional.scala 39:67]
  wire  _GEN_84 = _T_101 ? _T_113 : _GEN_74; // @[Conditional.scala 39:67]
  wire  cmd_done = _T_49 ? 1'h0 : _GEN_84; // @[Conditional.scala 40:58]
  wire  _T_276 = cmd_done | cmd_doneQ; // @[axi4_to_ahb.scala 242:47]
  wire  _T_277 = ~_T_276; // @[axi4_to_ahb.scala 242:36]
  wire [1:0] _T_279 = _T_277 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [1:0] _T_280 = _T_279 & 2'h2; // @[axi4_to_ahb.scala 242:61]
  wire  _T_300 = _T_55 | _T_96; // @[axi4_to_ahb.scala 252:62]
  wire  _T_301 = buf_state_en & _T_300; // @[axi4_to_ahb.scala 252:33]
  wire  _T_354 = _T_277 | bypass_en; // @[axi4_to_ahb.scala 257:61]
  wire [1:0] _T_356 = _T_354 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [1:0] _T_357 = _T_356 & 2'h2; // @[axi4_to_ahb.scala 257:75]
  wire  _T_364 = trxn_done | bypass_en; // @[axi4_to_ahb.scala 260:40]
  wire  _GEN_9 = _T_281 & _T_301; // @[Conditional.scala 39:67]
  wire  _GEN_30 = _T_188 ? 1'h0 : _GEN_9; // @[Conditional.scala 39:67]
  wire  _GEN_47 = _T_186 ? 1'h0 : _GEN_30; // @[Conditional.scala 39:67]
  wire  _GEN_64 = _T_175 ? 1'h0 : _GEN_47; // @[Conditional.scala 39:67]
  wire  _GEN_67 = _T_136 ? _T_152 : _GEN_64; // @[Conditional.scala 39:67]
  wire  _GEN_87 = _T_101 ? master_ready : _GEN_67; // @[Conditional.scala 39:67]
  wire  buf_wr_en = _T_49 ? buf_state_en : _GEN_87; // @[Conditional.scala 40:58]
  wire  _GEN_10 = _T_281 & buf_wr_en; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_13 = _T_281 ? _T_357 : 2'h0; // @[Conditional.scala 39:67]
  wire  _GEN_16 = _T_281 & _T_364; // @[Conditional.scala 39:67]
  wire  _GEN_21 = _T_188 ? buf_state_en : _GEN_16; // @[Conditional.scala 39:67]
  wire  _GEN_22 = _T_188 & buf_state_en; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_25 = _T_188 ? _T_280 : _GEN_13; // @[Conditional.scala 39:67]
  wire  _GEN_31 = _T_188 ? 1'h0 : _GEN_10; // @[Conditional.scala 39:67]
  wire  _GEN_36 = _T_186 ? buf_state_en : _GEN_31; // @[Conditional.scala 39:67]
  wire  _GEN_39 = _T_186 ? buf_state_en : _GEN_22; // @[Conditional.scala 39:67]
  wire  _GEN_41 = _T_186 ? 1'h0 : _GEN_21; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_44 = _T_186 ? 2'h0 : _GEN_25; // @[Conditional.scala 39:67]
  wire  _GEN_53 = _T_175 ? buf_state_en : _GEN_39; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_55 = _T_175 ? _T_185 : _GEN_44; // @[Conditional.scala 39:67]
  wire  _GEN_56 = _T_175 ? 1'h0 : _GEN_36; // @[Conditional.scala 39:67]
  wire  _GEN_60 = _T_175 ? 1'h0 : _GEN_41; // @[Conditional.scala 39:67]
  wire  _GEN_70 = _T_136 ? buf_state_en : _GEN_56; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_77 = _T_136 ? _T_174 : _GEN_55; // @[Conditional.scala 39:67]
  wire  _GEN_78 = _T_136 ? buf_wr_en : _GEN_53; // @[Conditional.scala 39:67]
  wire  _GEN_80 = _T_136 ? 1'h0 : _GEN_60; // @[Conditional.scala 39:67]
  wire  _GEN_85 = _T_101 ? buf_state_en : _GEN_78; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_90 = _T_101 ? _T_135 : _GEN_77; // @[Conditional.scala 39:67]
  wire  _GEN_91 = _T_101 ? 1'h0 : _GEN_70; // @[Conditional.scala 39:67]
  wire  _GEN_96 = _T_101 ? 1'h0 : _GEN_80; // @[Conditional.scala 39:67]
  wire  buf_data_wr_en = _T_49 ? _T_56 : _GEN_91; // @[Conditional.scala 40:58]
  wire  buf_cmd_byte_ptr_en = _T_49 ? buf_state_en : _GEN_96; // @[Conditional.scala 40:58]
  wire  slvbuf_wr_en = _T_49 ? 1'h0 : _GEN_85; // @[Conditional.scala 40:58]
  wire  _T_535 = master_size[1:0] == 2'h0; // @[axi4_to_ahb.scala 278:24]
  wire  _T_536 = _T_103 | _T_535; // @[axi4_to_ahb.scala 277:48]
  wire  _T_538 = master_size[1:0] == 2'h1; // @[axi4_to_ahb.scala 278:54]
  wire  _T_539 = _T_536 | _T_538; // @[axi4_to_ahb.scala 278:33]
  wire  _T_541 = master_size[1:0] == 2'h2; // @[axi4_to_ahb.scala 278:93]
  wire  _T_542 = _T_539 | _T_541; // @[axi4_to_ahb.scala 278:72]
  wire  _T_544 = master_size[1:0] == 2'h3; // @[axi4_to_ahb.scala 279:25]
  wire  _T_546 = wrbuf_byteen == 8'h3; // @[axi4_to_ahb.scala 279:62]
  wire  _T_548 = wrbuf_byteen == 8'hc; // @[axi4_to_ahb.scala 279:97]
  wire  _T_549 = _T_546 | _T_548; // @[axi4_to_ahb.scala 279:74]
  wire  _T_551 = wrbuf_byteen == 8'h30; // @[axi4_to_ahb.scala 279:132]
  wire  _T_552 = _T_549 | _T_551; // @[axi4_to_ahb.scala 279:109]
  wire  _T_554 = wrbuf_byteen == 8'hc0; // @[axi4_to_ahb.scala 279:168]
  wire  _T_555 = _T_552 | _T_554; // @[axi4_to_ahb.scala 279:145]
  wire  _T_557 = wrbuf_byteen == 8'hf; // @[axi4_to_ahb.scala 280:28]
  wire  _T_558 = _T_555 | _T_557; // @[axi4_to_ahb.scala 279:181]
  wire  _T_560 = wrbuf_byteen == 8'hf0; // @[axi4_to_ahb.scala 280:63]
  wire  _T_561 = _T_558 | _T_560; // @[axi4_to_ahb.scala 280:40]
  wire  _T_563 = wrbuf_byteen == 8'hff; // @[axi4_to_ahb.scala 280:99]
  wire  _T_564 = _T_561 | _T_563; // @[axi4_to_ahb.scala 280:76]
  wire  _T_565 = _T_544 & _T_564; // @[axi4_to_ahb.scala 279:38]
  wire  buf_aligned_in = _T_542 | _T_565; // @[axi4_to_ahb.scala 278:106]
  wire  _T_444 = buf_aligned_in & _T_51; // @[axi4_to_ahb.scala 272:60]
  wire [2:0] _T_461 = _T_548 ? 3'h7 : 3'h0; // @[Bitwise.scala 72:12]
  wire [2:0] _T_462 = 3'h2 & _T_461; // @[axi4_to_ahb.scala 135:15]
  wire  _T_468 = _T_560 | _T_546; // @[axi4_to_ahb.scala 136:56]
  wire [2:0] _T_470 = _T_468 ? 3'h7 : 3'h0; // @[Bitwise.scala 72:12]
  wire [2:0] _T_471 = 3'h4 & _T_470; // @[axi4_to_ahb.scala 136:15]
  wire [2:0] _T_472 = _T_462 | _T_471; // @[axi4_to_ahb.scala 135:63]
  wire [2:0] _T_476 = _T_554 ? 3'h7 : 3'h0; // @[Bitwise.scala 72:12]
  wire [2:0] _T_477 = 3'h6 & _T_476; // @[axi4_to_ahb.scala 137:15]
  wire [2:0] _T_478 = _T_472 | _T_477; // @[axi4_to_ahb.scala 136:96]
  wire [2:0] _T_485 = _T_444 ? _T_478 : master_addr[2:0]; // @[axi4_to_ahb.scala 272:43]
  reg  buf_write; // @[Reg.scala 27:20]
  wire  wrbuf_en = _T_44 & master_ready; // @[axi4_to_ahb.scala 298:49]
  wire  wrbuf_data_en = _T_45 & master_ready; // @[axi4_to_ahb.scala 299:52]
  wire  wrbuf_cmd_sent = _T_149 & _T_51; // @[axi4_to_ahb.scala 300:49]
  wire  _T_622 = ~wrbuf_en; // @[axi4_to_ahb.scala 301:33]
  wire  wrbuf_rst = wrbuf_cmd_sent & _T_622; // @[axi4_to_ahb.scala 301:31]
  wire  _T_624 = ~wrbuf_cmd_sent; // @[axi4_to_ahb.scala 303:36]
  wire  _T_625 = wrbuf_vld & _T_624; // @[axi4_to_ahb.scala 303:34]
  wire  _T_626 = ~_T_625; // @[axi4_to_ahb.scala 303:22]
  wire  _T_629 = wrbuf_data_vld & _T_624; // @[axi4_to_ahb.scala 304:38]
  wire  _T_630 = ~_T_629; // @[axi4_to_ahb.scala 304:21]
  wire  _T_636 = wrbuf_en | wrbuf_vld; // @[axi4_to_ahb.scala 308:55]
  wire  _T_637 = ~wrbuf_rst; // @[axi4_to_ahb.scala 308:91]
  wire  _T_641 = wrbuf_data_en | wrbuf_data_vld; // @[axi4_to_ahb.scala 309:55]
  wire  _T_691 = ~slave_valid_pre; // @[axi4_to_ahb.scala 326:92]
  wire  _T_704 = buf_wr_en | slvbuf_wr_en; // @[axi4_to_ahb.scala 334:43]
  wire  _T_705 = _T_704 | io_clk_override; // @[axi4_to_ahb.scala 334:58]
  wire  _T_708 = io_ahb_in_hready & io_ahb_out_htrans[1]; // @[axi4_to_ahb.scala 335:57]
  wire  _T_709 = _T_708 | io_clk_override; // @[axi4_to_ahb.scala 335:81]
  wire  _T_711 = buf_state != 3'h0; // @[axi4_to_ahb.scala 336:50]
  wire  _T_712 = _T_711 | io_clk_override; // @[axi4_to_ahb.scala 336:60]
  rvclkhdr rvclkhdr ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_io_l1clk),
    .io_clk(rvclkhdr_io_clk),
    .io_en(rvclkhdr_io_en),
    .io_scan_mode(rvclkhdr_io_scan_mode)
  );
  rvclkhdr rvclkhdr_1 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_1_io_l1clk),
    .io_clk(rvclkhdr_1_io_clk),
    .io_en(rvclkhdr_1_io_en),
    .io_scan_mode(rvclkhdr_1_io_scan_mode)
  );
  rvclkhdr rvclkhdr_2 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_2_io_l1clk),
    .io_clk(rvclkhdr_2_io_clk),
    .io_en(rvclkhdr_2_io_en),
    .io_scan_mode(rvclkhdr_2_io_scan_mode)
  );
  rvclkhdr rvclkhdr_3 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_3_io_l1clk),
    .io_clk(rvclkhdr_3_io_clk),
    .io_en(rvclkhdr_3_io_en),
    .io_scan_mode(rvclkhdr_3_io_scan_mode)
  );
  rvclkhdr rvclkhdr_4 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_4_io_l1clk),
    .io_clk(rvclkhdr_4_io_clk),
    .io_en(rvclkhdr_4_io_en),
    .io_scan_mode(rvclkhdr_4_io_scan_mode)
  );
  rvclkhdr rvclkhdr_5 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_5_io_l1clk),
    .io_clk(rvclkhdr_5_io_clk),
    .io_en(rvclkhdr_5_io_en),
    .io_scan_mode(rvclkhdr_5_io_scan_mode)
  );
  rvclkhdr rvclkhdr_6 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_6_io_l1clk),
    .io_clk(rvclkhdr_6_io_clk),
    .io_en(rvclkhdr_6_io_en),
    .io_scan_mode(rvclkhdr_6_io_scan_mode)
  );
  rvclkhdr rvclkhdr_7 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_7_io_l1clk),
    .io_clk(rvclkhdr_7_io_clk),
    .io_en(rvclkhdr_7_io_en),
    .io_scan_mode(rvclkhdr_7_io_scan_mode)
  );
  rvclkhdr rvclkhdr_8 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_8_io_l1clk),
    .io_clk(rvclkhdr_8_io_clk),
    .io_en(rvclkhdr_8_io_en),
    .io_scan_mode(rvclkhdr_8_io_scan_mode)
  );
  rvclkhdr rvclkhdr_9 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_9_io_l1clk),
    .io_clk(rvclkhdr_9_io_clk),
    .io_en(rvclkhdr_9_io_en),
    .io_scan_mode(rvclkhdr_9_io_scan_mode)
  );
  assign io_axi_aw_ready = _T_626 & master_ready; // @[axi4_to_ahb.scala 303:19]
  assign io_axi_w_ready = _T_630 & master_ready; // @[axi4_to_ahb.scala 304:18]
  assign io_ahb_out_htrans = _T_49 ? _T_100 : _GEN_90; // @[axi4_to_ahb.scala 29:21 axi4_to_ahb.scala 185:25 axi4_to_ahb.scala 197:25 axi4_to_ahb.scala 212:25 axi4_to_ahb.scala 222:25 axi4_to_ahb.scala 242:25 axi4_to_ahb.scala 257:25]
  assign io_ahb_out_hwrite = bypass_en ? _T_51 : buf_write; // @[axi4_to_ahb.scala 288:21]
  assign rvclkhdr_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_io_en = io_bus_clk_en; // @[lib.scala 345:16]
  assign rvclkhdr_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_1_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_1_io_en = io_bus_clk_en & _T_46; // @[lib.scala 345:16]
  assign rvclkhdr_1_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_2_io_clk = rvclkhdr_io_l1clk; // @[lib.scala 370:18]
  assign rvclkhdr_2_io_en = _T_44 & master_ready; // @[lib.scala 371:17]
  assign rvclkhdr_2_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_3_io_clk = rvclkhdr_io_l1clk; // @[lib.scala 370:18]
  assign rvclkhdr_3_io_en = _T_45 & master_ready; // @[lib.scala 371:17]
  assign rvclkhdr_3_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_4_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_4_io_en = buf_wr_en & io_bus_clk_en; // @[lib.scala 371:17]
  assign rvclkhdr_4_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_5_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_5_io_en = buf_data_wr_en & io_bus_clk_en; // @[lib.scala 371:17]
  assign rvclkhdr_5_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_6_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_6_io_en = io_bus_clk_en & _T_705; // @[lib.scala 345:16]
  assign rvclkhdr_6_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_7_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_7_io_en = io_bus_clk_en; // @[lib.scala 345:16]
  assign rvclkhdr_7_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_8_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_8_io_en = io_bus_clk_en & _T_709; // @[lib.scala 345:16]
  assign rvclkhdr_8_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_9_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_9_io_en = io_bus_clk_en & _T_712; // @[lib.scala 345:16]
  assign rvclkhdr_9_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  buf_state = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  wrbuf_vld = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  wrbuf_data_vld = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  ahb_hready_q = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  ahb_htrans_q = _RAND_4[1:0];
  _RAND_5 = {1{`RANDOM}};
  ahb_hwrite_q = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  ahb_hresp_q = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  cmd_doneQ = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  wrbuf_addr = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  wrbuf_size = _RAND_9[2:0];
  _RAND_10 = {1{`RANDOM}};
  wrbuf_byteen = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  buf_addr = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  buf_cmd_byte_ptrQ = _RAND_12[2:0];
  _RAND_13 = {1{`RANDOM}};
  buf_byteen = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  buf_aligned = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  buf_write = _RAND_15[0:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    buf_state = 3'h0;
  end
  if (reset) begin
    wrbuf_vld = 1'h0;
  end
  if (reset) begin
    wrbuf_data_vld = 1'h0;
  end
  if (reset) begin
    ahb_hready_q = 1'h0;
  end
  if (reset) begin
    ahb_htrans_q = 2'h0;
  end
  if (reset) begin
    ahb_hwrite_q = 1'h0;
  end
  if (reset) begin
    ahb_hresp_q = 1'h0;
  end
  if (reset) begin
    cmd_doneQ = 1'h0;
  end
  if (reset) begin
    wrbuf_addr = 32'h0;
  end
  if (reset) begin
    wrbuf_size = 3'h0;
  end
  if (reset) begin
    wrbuf_byteen = 8'h0;
  end
  if (reset) begin
    buf_addr = 32'h0;
  end
  if (reset) begin
    buf_cmd_byte_ptrQ = 3'h0;
  end
  if (reset) begin
    buf_byteen = 8'h0;
  end
  if (reset) begin
    buf_aligned = 1'h0;
  end
  if (reset) begin
    buf_write = 1'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge ahbm_clk or posedge reset) begin
    if (reset) begin
      buf_state <= 3'h0;
    end else if (buf_state_en) begin
      if (_T_49) begin
        if (buf_write_in) begin
          buf_state <= 3'h2;
        end else begin
          buf_state <= 3'h1;
        end
      end else if (_T_101) begin
        if (_T_104) begin
          buf_state <= 3'h6;
        end else begin
          buf_state <= 3'h3;
        end
      end else if (_T_136) begin
        if (ahb_hresp_q) begin
          buf_state <= 3'h7;
        end else if (_T_152) begin
          buf_state <= 3'h6;
        end else begin
          buf_state <= 3'h3;
        end
      end else if (_T_175) begin
        buf_state <= 3'h3;
      end else if (_T_186) begin
        buf_state <= 3'h5;
      end else if (_T_188) begin
        buf_state <= 3'h4;
      end else if (_T_281) begin
        if (_T_288) begin
          buf_state <= 3'h5;
        end else if (master_valid) begin
          if (_T_51) begin
            buf_state <= 3'h2;
          end else begin
            buf_state <= 3'h1;
          end
        end else begin
          buf_state <= 3'h0;
        end
      end else begin
        buf_state <= 3'h0;
      end
    end
  end
  always @(posedge bus_clk or posedge reset) begin
    if (reset) begin
      wrbuf_vld <= 1'h0;
    end else begin
      wrbuf_vld <= _T_636 & _T_637;
    end
  end
  always @(posedge bus_clk or posedge reset) begin
    if (reset) begin
      wrbuf_data_vld <= 1'h0;
    end else begin
      wrbuf_data_vld <= _T_641 & _T_637;
    end
  end
  always @(posedge ahbm_clk or posedge reset) begin
    if (reset) begin
      ahb_hready_q <= 1'h0;
    end else begin
      ahb_hready_q <= io_ahb_in_hready;
    end
  end
  always @(posedge ahbm_clk or posedge reset) begin
    if (reset) begin
      ahb_htrans_q <= 2'h0;
    end else begin
      ahb_htrans_q <= io_ahb_out_htrans;
    end
  end
  always @(posedge ahbm_addr_clk or posedge reset) begin
    if (reset) begin
      ahb_hwrite_q <= 1'h0;
    end else begin
      ahb_hwrite_q <= io_ahb_out_hwrite;
    end
  end
  always @(posedge ahbm_clk or posedge reset) begin
    if (reset) begin
      ahb_hresp_q <= 1'h0;
    end else begin
      ahb_hresp_q <= io_ahb_in_hresp;
    end
  end
  always @(posedge ahbm_clk or posedge reset) begin
    if (reset) begin
      cmd_doneQ <= 1'h0;
    end else begin
      cmd_doneQ <= _T_276 & _T_691;
    end
  end
  always @(posedge rvclkhdr_2_io_l1clk or posedge reset) begin
    if (reset) begin
      wrbuf_addr <= 32'h0;
    end else begin
      wrbuf_addr <= io_axi_aw_bits_addr;
    end
  end
  always @(posedge bus_clk or posedge reset) begin
    if (reset) begin
      wrbuf_size <= 3'h0;
    end else if (wrbuf_en) begin
      wrbuf_size <= io_axi_aw_bits_size;
    end
  end
  always @(posedge bus_clk or posedge reset) begin
    if (reset) begin
      wrbuf_byteen <= 8'h0;
    end else if (wrbuf_data_en) begin
      wrbuf_byteen <= io_axi_w_bits_strb;
    end
  end
  always @(posedge rvclkhdr_4_io_l1clk or posedge reset) begin
    if (reset) begin
      buf_addr <= 32'h0;
    end else begin
      buf_addr <= {master_addr[31:3],_T_485};
    end
  end
  always @(posedge ahbm_clk or posedge reset) begin
    if (reset) begin
      buf_cmd_byte_ptrQ <= 3'h0;
    end else if (buf_cmd_byte_ptr_en) begin
      if (_T_49) begin
        if (buf_write_in) begin
          if (wrbuf_byteen[0]) begin
            buf_cmd_byte_ptrQ <= 3'h0;
          end else if (wrbuf_byteen[1]) begin
            buf_cmd_byte_ptrQ <= 3'h1;
          end else if (wrbuf_byteen[2]) begin
            buf_cmd_byte_ptrQ <= 3'h2;
          end else if (wrbuf_byteen[3]) begin
            buf_cmd_byte_ptrQ <= 3'h3;
          end else if (wrbuf_byteen[4]) begin
            buf_cmd_byte_ptrQ <= 3'h4;
          end else if (wrbuf_byteen[5]) begin
            buf_cmd_byte_ptrQ <= 3'h5;
          end else if (wrbuf_byteen[6]) begin
            buf_cmd_byte_ptrQ <= 3'h6;
          end else begin
            buf_cmd_byte_ptrQ <= 3'h7;
          end
        end else begin
          buf_cmd_byte_ptrQ <= master_addr[2:0];
        end
      end else if (_T_101) begin
        if (bypass_en) begin
          buf_cmd_byte_ptrQ <= master_addr[2:0];
        end else begin
          buf_cmd_byte_ptrQ <= buf_addr[2:0];
        end
      end else if (_T_136) begin
        if (bypass_en) begin
          buf_cmd_byte_ptrQ <= master_addr[2:0];
        end else begin
          buf_cmd_byte_ptrQ <= buf_addr[2:0];
        end
      end else if (_T_175) begin
        buf_cmd_byte_ptrQ <= buf_addr[2:0];
      end else if (_T_186) begin
        buf_cmd_byte_ptrQ <= 3'h0;
      end else if (_T_188) begin
        if (trxn_done) begin
          if (_T_201) begin
            buf_cmd_byte_ptrQ <= 3'h0;
          end else if (_T_204) begin
            buf_cmd_byte_ptrQ <= 3'h1;
          end else if (_T_207) begin
            buf_cmd_byte_ptrQ <= 3'h2;
          end else if (_T_210) begin
            buf_cmd_byte_ptrQ <= 3'h3;
          end else if (_T_213) begin
            buf_cmd_byte_ptrQ <= 3'h4;
          end else if (_T_216) begin
            buf_cmd_byte_ptrQ <= 3'h5;
          end else if (_T_219) begin
            buf_cmd_byte_ptrQ <= 3'h6;
          end else begin
            buf_cmd_byte_ptrQ <= 3'h7;
          end
        end
      end else if (_T_281) begin
        if (bypass_en) begin
          if (wrbuf_byteen[0]) begin
            buf_cmd_byte_ptrQ <= 3'h0;
          end else if (wrbuf_byteen[1]) begin
            buf_cmd_byte_ptrQ <= 3'h1;
          end else if (wrbuf_byteen[2]) begin
            buf_cmd_byte_ptrQ <= 3'h2;
          end else if (wrbuf_byteen[3]) begin
            buf_cmd_byte_ptrQ <= 3'h3;
          end else if (wrbuf_byteen[4]) begin
            buf_cmd_byte_ptrQ <= 3'h4;
          end else if (wrbuf_byteen[5]) begin
            buf_cmd_byte_ptrQ <= 3'h5;
          end else if (wrbuf_byteen[6]) begin
            buf_cmd_byte_ptrQ <= 3'h6;
          end else begin
            buf_cmd_byte_ptrQ <= 3'h7;
          end
        end else if (trxn_done) begin
          if (_T_201) begin
            buf_cmd_byte_ptrQ <= 3'h0;
          end else if (_T_204) begin
            buf_cmd_byte_ptrQ <= 3'h1;
          end else if (_T_207) begin
            buf_cmd_byte_ptrQ <= 3'h2;
          end else if (_T_210) begin
            buf_cmd_byte_ptrQ <= 3'h3;
          end else if (_T_213) begin
            buf_cmd_byte_ptrQ <= 3'h4;
          end else if (_T_216) begin
            buf_cmd_byte_ptrQ <= 3'h5;
          end else if (_T_219) begin
            buf_cmd_byte_ptrQ <= 3'h6;
          end else begin
            buf_cmd_byte_ptrQ <= 3'h7;
          end
        end
      end else begin
        buf_cmd_byte_ptrQ <= 3'h0;
      end
    end
  end
  always @(posedge buf_clk or posedge reset) begin
    if (reset) begin
      buf_byteen <= 8'h0;
    end else if (buf_wr_en) begin
      buf_byteen <= wrbuf_byteen;
    end
  end
  always @(posedge buf_clk or posedge reset) begin
    if (reset) begin
      buf_aligned <= 1'h0;
    end else if (buf_wr_en) begin
      buf_aligned <= buf_aligned_in;
    end
  end
  always @(posedge buf_clk or posedge reset) begin
    if (reset) begin
      buf_write <= 1'h0;
    end else if (buf_wr_en) begin
      if (_T_49) begin
        buf_write <= _T_51;
      end else if (_T_101) begin
        buf_write <= 1'h0;
      end else if (_T_136) begin
        buf_write <= 1'h0;
      end else if (_T_175) begin
        buf_write <= 1'h0;
      end else if (_T_186) begin
        buf_write <= 1'h0;
      end else if (_T_188) begin
        buf_write <= 1'h0;
      end else begin
        buf_write <= _GEN_8;
      end
    end
  end
endmodule
module ahb_to_axi4(
  input         clock,
  input         reset,
  input         io_scan_mode,
  input         io_bus_clk_en,
  output        io_axi_aw_valid,
  output        io_axi_ar_valid,
  input         io_axi_r_valid,
  input  [1:0]  io_axi_r_bits_resp,
  output        io_ahb_sig_in_hready,
  output        io_ahb_sig_in_hresp,
  input  [31:0] io_ahb_sig_out_haddr,
  input  [2:0]  io_ahb_sig_out_hsize,
  input  [1:0]  io_ahb_sig_out_htrans,
  input         io_ahb_sig_out_hwrite,
  input         io_ahb_hsel,
  input         io_ahb_hreadyin
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
`endif // RANDOMIZE_REG_INIT
  wire  rvclkhdr_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_1_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_1_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_1_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_1_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_2_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_2_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_2_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_2_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_3_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_3_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_3_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_3_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_4_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_4_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_4_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_4_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_5_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_5_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_5_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_5_io_scan_mode; // @[lib.scala 343:22]
  wire  ahb_addr_clk = rvclkhdr_1_io_l1clk; // @[ahb_to_axi4.scala 45:33 ahb_to_axi4.scala 134:31]
  reg [31:0] ahb_haddr_q; // @[ahb_to_axi4.scala 127:65]
  wire  ahb_addr_in_dccm = ahb_haddr_q[31:16] == 16'hf004; // @[lib.scala 87:29]
  wire  ahb_addr_in_iccm = ahb_haddr_q[31:16] == 16'hee00; // @[lib.scala 87:29]
  wire  ahb_clk = rvclkhdr_io_l1clk; // @[ahb_to_axi4.scala 44:33 ahb_to_axi4.scala 133:31]
  reg [1:0] buf_state; // @[Reg.scala 27:20]
  wire  _T_7 = 2'h0 == buf_state; // @[Conditional.scala 37:30]
  wire  ahb_hready = io_ahb_sig_in_hready & io_ahb_hreadyin; // @[ahb_to_axi4.scala 105:55]
  wire  _T_10 = ahb_hready & io_ahb_sig_out_htrans[1]; // @[ahb_to_axi4.scala 77:34]
  wire  _T_11 = _T_10 & io_ahb_hsel; // @[ahb_to_axi4.scala 77:61]
  wire  _T_12 = 2'h1 == buf_state; // @[Conditional.scala 37:30]
  wire  _T_14 = io_ahb_sig_out_htrans == 2'h0; // @[ahb_to_axi4.scala 80:79]
  wire  _T_15 = io_ahb_sig_in_hresp | _T_14; // @[ahb_to_axi4.scala 80:48]
  wire  _T_16 = ~io_ahb_hsel; // @[ahb_to_axi4.scala 80:93]
  wire  _T_17 = _T_15 | _T_16; // @[ahb_to_axi4.scala 80:91]
  wire  bus_clk = rvclkhdr_5_io_l1clk; // @[ahb_to_axi4.scala 58:33 ahb_to_axi4.scala 181:27]
  reg  cmdbuf_vld; // @[ahb_to_axi4.scala 140:61]
  wire  _T_153 = io_axi_aw_valid | io_axi_ar_valid; // @[ahb_to_axi4.scala 138:86]
  wire  _T_154 = ~_T_153; // @[ahb_to_axi4.scala 138:48]
  wire  cmdbuf_full = cmdbuf_vld & _T_154; // @[ahb_to_axi4.scala 138:46]
  wire  _T_21 = ~cmdbuf_full; // @[ahb_to_axi4.scala 81:24]
  wire  _T_22 = _T_21 | io_ahb_sig_in_hresp; // @[ahb_to_axi4.scala 81:37]
  wire  _T_25 = io_ahb_sig_out_htrans == 2'h1; // @[ahb_to_axi4.scala 82:92]
  wire  _T_26 = _T_25 & io_ahb_hsel; // @[ahb_to_axi4.scala 82:110]
  wire  _T_27 = io_ahb_sig_in_hresp | _T_26; // @[ahb_to_axi4.scala 82:60]
  wire  _T_28 = ~_T_27; // @[ahb_to_axi4.scala 82:38]
  wire  _T_29 = _T_21 & _T_28; // @[ahb_to_axi4.scala 82:36]
  wire  _T_30 = 2'h2 == buf_state; // @[Conditional.scala 37:30]
  wire  _T_34 = ~io_ahb_sig_in_hresp; // @[ahb_to_axi4.scala 87:23]
  wire  _T_36 = _T_34 & _T_21; // @[ahb_to_axi4.scala 87:44]
  wire  _T_37 = 2'h3 == buf_state; // @[Conditional.scala 37:30]
  reg  cmdbuf_write; // @[Reg.scala 27:20]
  wire  _T_38 = ~cmdbuf_write; // @[ahb_to_axi4.scala 91:40]
  wire  _T_39 = io_axi_r_valid & _T_38; // @[ahb_to_axi4.scala 91:38]
  wire  _T_41 = |io_axi_r_bits_resp; // @[ahb_to_axi4.scala 93:68]
  wire  _GEN_1 = _T_37 & _T_39; // @[Conditional.scala 39:67]
  wire  _GEN_5 = _T_30 ? _T_22 : _GEN_1; // @[Conditional.scala 39:67]
  wire  _GEN_10 = _T_12 ? _T_22 : _GEN_5; // @[Conditional.scala 39:67]
  wire  buf_state_en = _T_7 ? _T_11 : _GEN_10; // @[Conditional.scala 40:58]
  wire  _T_42 = buf_state_en & _T_41; // @[ahb_to_axi4.scala 93:41]
  wire  _GEN_2 = _T_37 & buf_state_en; // @[Conditional.scala 39:67]
  wire  _GEN_3 = _T_37 & _T_42; // @[Conditional.scala 39:67]
  wire  _GEN_6 = _T_30 & _T_36; // @[Conditional.scala 39:67]
  wire  _GEN_7 = _T_30 ? 1'h0 : _GEN_2; // @[Conditional.scala 39:67]
  wire  _GEN_11 = _T_12 ? _T_29 : _GEN_6; // @[Conditional.scala 39:67]
  wire  _GEN_12 = _T_12 ? 1'h0 : _GEN_7; // @[Conditional.scala 39:67]
  wire  cmdbuf_wr_en = _T_7 ? 1'h0 : _GEN_11; // @[Conditional.scala 40:58]
  wire  buf_rdata_en = _T_7 ? 1'h0 : _GEN_12; // @[Conditional.scala 40:58]
  reg [2:0] ahb_hsize_q; // @[ahb_to_axi4.scala 125:65]
  wire  _T_53 = ahb_hsize_q == 3'h1; // @[ahb_to_axi4.scala 99:30]
  wire  _T_61 = ahb_hsize_q == 3'h2; // @[ahb_to_axi4.scala 100:30]
  wire  _T_69 = ahb_hsize_q == 3'h3; // @[ahb_to_axi4.scala 101:30]
  reg  ahb_hready_q; // @[ahb_to_axi4.scala 123:60]
  wire  _T_74 = ~ahb_hready_q; // @[ahb_to_axi4.scala 104:80]
  reg  ahb_hresp_q; // @[ahb_to_axi4.scala 122:60]
  wire  _T_75 = ahb_hresp_q & _T_74; // @[ahb_to_axi4.scala 104:78]
  wire  _T_77 = buf_state == 2'h0; // @[ahb_to_axi4.scala 104:124]
  wire  _T_78 = _T_21 | _T_77; // @[ahb_to_axi4.scala 104:111]
  wire  _T_79 = buf_state == 2'h2; // @[ahb_to_axi4.scala 104:149]
  wire  _T_80 = buf_state == 2'h3; // @[ahb_to_axi4.scala 104:168]
  wire  _T_81 = _T_79 | _T_80; // @[ahb_to_axi4.scala 104:156]
  wire  _T_82 = ~_T_81; // @[ahb_to_axi4.scala 104:137]
  wire  _T_83 = _T_78 & _T_82; // @[ahb_to_axi4.scala 104:135]
  reg  buf_read_error; // @[ahb_to_axi4.scala 119:60]
  wire  _T_84 = ~buf_read_error; // @[ahb_to_axi4.scala 104:181]
  wire  _T_85 = _T_83 & _T_84; // @[ahb_to_axi4.scala 104:179]
  wire [1:0] _T_89 = io_ahb_hsel ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  reg [1:0] ahb_htrans_q; // @[ahb_to_axi4.scala 124:60]
  wire  _T_94 = ahb_htrans_q != 2'h0; // @[ahb_to_axi4.scala 108:61]
  wire  _T_95 = buf_state != 2'h0; // @[ahb_to_axi4.scala 108:83]
  wire  _T_96 = _T_94 & _T_95; // @[ahb_to_axi4.scala 108:70]
  wire  _T_97 = ahb_addr_in_dccm | ahb_addr_in_iccm; // @[ahb_to_axi4.scala 109:26]
  wire  _T_98 = ~_T_97; // @[ahb_to_axi4.scala 109:7]
  reg  ahb_hwrite_q; // @[ahb_to_axi4.scala 126:65]
  wire  _T_99 = ahb_addr_in_dccm & ahb_hwrite_q; // @[ahb_to_axi4.scala 110:46]
  wire  _T_100 = ahb_addr_in_iccm | _T_99; // @[ahb_to_axi4.scala 110:26]
  wire  _T_102 = ahb_hsize_q[1:0] == 2'h2; // @[ahb_to_axi4.scala 110:86]
  wire  _T_104 = ahb_hsize_q[1:0] == 2'h3; // @[ahb_to_axi4.scala 110:115]
  wire  _T_105 = _T_102 | _T_104; // @[ahb_to_axi4.scala 110:95]
  wire  _T_106 = ~_T_105; // @[ahb_to_axi4.scala 110:66]
  wire  _T_107 = _T_100 & _T_106; // @[ahb_to_axi4.scala 110:64]
  wire  _T_108 = _T_98 | _T_107; // @[ahb_to_axi4.scala 109:47]
  wire  _T_112 = _T_53 & ahb_haddr_q[0]; // @[ahb_to_axi4.scala 111:35]
  wire  _T_113 = _T_108 | _T_112; // @[ahb_to_axi4.scala 110:126]
  wire  _T_117 = |ahb_haddr_q[1:0]; // @[ahb_to_axi4.scala 112:56]
  wire  _T_118 = _T_61 & _T_117; // @[ahb_to_axi4.scala 112:35]
  wire  _T_119 = _T_113 | _T_118; // @[ahb_to_axi4.scala 111:55]
  wire  _T_123 = |ahb_haddr_q[2:0]; // @[ahb_to_axi4.scala 113:56]
  wire  _T_124 = _T_69 & _T_123; // @[ahb_to_axi4.scala 113:35]
  wire  _T_125 = _T_119 | _T_124; // @[ahb_to_axi4.scala 112:61]
  wire  _T_126 = _T_96 & _T_125; // @[ahb_to_axi4.scala 108:94]
  wire  _T_127 = _T_126 | buf_read_error; // @[ahb_to_axi4.scala 113:63]
  wire  _T_146 = ~cmdbuf_wr_en; // @[ahb_to_axi4.scala 137:113]
  wire  _T_147 = _T_153 & _T_146; // @[ahb_to_axi4.scala 137:111]
  wire  _T_149 = io_ahb_sig_in_hresp & _T_38; // @[ahb_to_axi4.scala 137:151]
  wire  cmdbuf_rst = _T_147 | _T_149; // @[ahb_to_axi4.scala 137:128]
  wire  _T_157 = cmdbuf_wr_en | cmdbuf_vld; // @[ahb_to_axi4.scala 140:66]
  wire  _T_158 = ~cmdbuf_rst; // @[ahb_to_axi4.scala 140:110]
  rvclkhdr rvclkhdr ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_io_l1clk),
    .io_clk(rvclkhdr_io_clk),
    .io_en(rvclkhdr_io_en),
    .io_scan_mode(rvclkhdr_io_scan_mode)
  );
  rvclkhdr rvclkhdr_1 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_1_io_l1clk),
    .io_clk(rvclkhdr_1_io_clk),
    .io_en(rvclkhdr_1_io_en),
    .io_scan_mode(rvclkhdr_1_io_scan_mode)
  );
  rvclkhdr rvclkhdr_2 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_2_io_l1clk),
    .io_clk(rvclkhdr_2_io_clk),
    .io_en(rvclkhdr_2_io_en),
    .io_scan_mode(rvclkhdr_2_io_scan_mode)
  );
  rvclkhdr rvclkhdr_3 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_3_io_l1clk),
    .io_clk(rvclkhdr_3_io_clk),
    .io_en(rvclkhdr_3_io_en),
    .io_scan_mode(rvclkhdr_3_io_scan_mode)
  );
  rvclkhdr rvclkhdr_4 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_4_io_l1clk),
    .io_clk(rvclkhdr_4_io_clk),
    .io_en(rvclkhdr_4_io_en),
    .io_scan_mode(rvclkhdr_4_io_scan_mode)
  );
  rvclkhdr rvclkhdr_5 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_5_io_l1clk),
    .io_clk(rvclkhdr_5_io_clk),
    .io_en(rvclkhdr_5_io_en),
    .io_scan_mode(rvclkhdr_5_io_scan_mode)
  );
  assign io_axi_aw_valid = cmdbuf_vld & cmdbuf_write; // @[ahb_to_axi4.scala 20:10 ahb_to_axi4.scala 157:28]
  assign io_axi_ar_valid = cmdbuf_vld & _T_38; // @[ahb_to_axi4.scala 20:10 ahb_to_axi4.scala 172:28]
  assign io_ahb_sig_in_hready = io_ahb_sig_in_hresp ? _T_75 : _T_85; // @[ahb_to_axi4.scala 104:38]
  assign io_ahb_sig_in_hresp = _T_127 | _T_75; // @[ahb_to_axi4.scala 108:38]
  assign rvclkhdr_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_io_en = io_bus_clk_en; // @[lib.scala 345:16]
  assign rvclkhdr_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_1_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_1_io_en = io_bus_clk_en & _T_10; // @[lib.scala 345:16]
  assign rvclkhdr_1_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_2_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_2_io_en = io_bus_clk_en & buf_rdata_en; // @[lib.scala 345:16]
  assign rvclkhdr_2_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_3_io_clk = rvclkhdr_5_io_l1clk; // @[lib.scala 370:18]
  assign rvclkhdr_3_io_en = _T_7 ? 1'h0 : _GEN_11; // @[lib.scala 371:17]
  assign rvclkhdr_3_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_4_io_clk = rvclkhdr_5_io_l1clk; // @[lib.scala 370:18]
  assign rvclkhdr_4_io_en = _T_7 ? 1'h0 : _GEN_11; // @[lib.scala 371:17]
  assign rvclkhdr_4_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_5_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_5_io_en = io_bus_clk_en; // @[lib.scala 345:16]
  assign rvclkhdr_5_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ahb_haddr_q = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  buf_state = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  cmdbuf_vld = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  cmdbuf_write = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  ahb_hsize_q = _RAND_4[2:0];
  _RAND_5 = {1{`RANDOM}};
  ahb_hready_q = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  ahb_hresp_q = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  buf_read_error = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  ahb_htrans_q = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  ahb_hwrite_q = _RAND_9[0:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    ahb_haddr_q = 32'h0;
  end
  if (reset) begin
    buf_state = 2'h0;
  end
  if (reset) begin
    cmdbuf_vld = 1'h0;
  end
  if (reset) begin
    cmdbuf_write = 1'h0;
  end
  if (reset) begin
    ahb_hsize_q = 3'h0;
  end
  if (reset) begin
    ahb_hready_q = 1'h0;
  end
  if (reset) begin
    ahb_hresp_q = 1'h0;
  end
  if (reset) begin
    buf_read_error = 1'h0;
  end
  if (reset) begin
    ahb_htrans_q = 2'h0;
  end
  if (reset) begin
    ahb_hwrite_q = 1'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge ahb_addr_clk or posedge reset) begin
    if (reset) begin
      ahb_haddr_q <= 32'h0;
    end else begin
      ahb_haddr_q <= io_ahb_sig_out_haddr;
    end
  end
  always @(posedge ahb_clk or posedge reset) begin
    if (reset) begin
      buf_state <= 2'h0;
    end else if (buf_state_en) begin
      if (_T_7) begin
        if (io_ahb_sig_out_hwrite) begin
          buf_state <= 2'h1;
        end else begin
          buf_state <= 2'h2;
        end
      end else if (_T_12) begin
        if (_T_17) begin
          buf_state <= 2'h0;
        end else if (io_ahb_sig_out_hwrite) begin
          buf_state <= 2'h1;
        end else begin
          buf_state <= 2'h2;
        end
      end else if (_T_30) begin
        if (io_ahb_sig_in_hresp) begin
          buf_state <= 2'h0;
        end else begin
          buf_state <= 2'h3;
        end
      end else begin
        buf_state <= 2'h0;
      end
    end
  end
  always @(posedge bus_clk or posedge reset) begin
    if (reset) begin
      cmdbuf_vld <= 1'h0;
    end else begin
      cmdbuf_vld <= _T_157 & _T_158;
    end
  end
  always @(posedge bus_clk or posedge reset) begin
    if (reset) begin
      cmdbuf_write <= 1'h0;
    end else if (cmdbuf_wr_en) begin
      cmdbuf_write <= ahb_hwrite_q;
    end
  end
  always @(posedge ahb_addr_clk or posedge reset) begin
    if (reset) begin
      ahb_hsize_q <= 3'h0;
    end else begin
      ahb_hsize_q <= io_ahb_sig_out_hsize;
    end
  end
  always @(posedge ahb_clk or posedge reset) begin
    if (reset) begin
      ahb_hready_q <= 1'h0;
    end else begin
      ahb_hready_q <= io_ahb_sig_in_hready & io_ahb_hreadyin;
    end
  end
  always @(posedge ahb_clk or posedge reset) begin
    if (reset) begin
      ahb_hresp_q <= 1'h0;
    end else begin
      ahb_hresp_q <= io_ahb_sig_in_hresp;
    end
  end
  always @(posedge ahb_clk or posedge reset) begin
    if (reset) begin
      buf_read_error <= 1'h0;
    end else if (_T_7) begin
      buf_read_error <= 1'h0;
    end else if (_T_12) begin
      buf_read_error <= 1'h0;
    end else if (_T_30) begin
      buf_read_error <= 1'h0;
    end else begin
      buf_read_error <= _GEN_3;
    end
  end
  always @(posedge ahb_clk or posedge reset) begin
    if (reset) begin
      ahb_htrans_q <= 2'h0;
    end else begin
      ahb_htrans_q <= _T_89 & io_ahb_sig_out_htrans;
    end
  end
  always @(posedge ahb_addr_clk or posedge reset) begin
    if (reset) begin
      ahb_hwrite_q <= 1'h0;
    end else begin
      ahb_hwrite_q <= io_ahb_sig_out_hwrite;
    end
  end
endmodule
module quasar(
  input         clock,
  input         reset,
  input         io_lsu_ahb_in_hready,
  input         io_lsu_ahb_in_hresp,
  input         io_ifu_ahb_in_hready,
  input         io_ifu_ahb_in_hresp,
  input         io_sb_ahb_in_hready,
  input         io_sb_ahb_in_hresp,
  input  [31:0] io_dma_ahb_sig_out_haddr,
  input  [2:0]  io_dma_ahb_sig_out_hsize,
  input  [1:0]  io_dma_ahb_sig_out_htrans,
  input         io_dma_ahb_sig_out_hwrite,
  input         io_dma_ahb_hsel,
  input         io_dma_ahb_hreadyin,
  input         io_dbg_rst_l,
  input  [30:0] io_rst_vec,
  input         io_nmi_int,
  input  [30:0] io_nmi_vec,
  output        io_core_rst_l,
  output [1:0]  io_rv_trace_pkt_rv_i_valid_ip,
  output [31:0] io_rv_trace_pkt_rv_i_insn_ip,
  output [31:0] io_rv_trace_pkt_rv_i_address_ip,
  output [1:0]  io_rv_trace_pkt_rv_i_exception_ip,
  output [4:0]  io_rv_trace_pkt_rv_i_ecause_ip,
  output [1:0]  io_rv_trace_pkt_rv_i_interrupt_ip,
  output [31:0] io_rv_trace_pkt_rv_i_tval_ip,
  output        io_dccm_clk_override,
  output        io_icm_clk_override,
  output        io_dec_tlu_core_ecc_disable,
  input         io_i_cpu_halt_req,
  input         io_i_cpu_run_req,
  output        io_o_cpu_halt_ack,
  output        io_o_cpu_halt_status,
  output        io_o_cpu_run_ack,
  output        io_o_debug_mode_status,
  input  [27:0] io_core_id,
  input         io_mpc_debug_halt_req,
  input         io_mpc_debug_run_req,
  input         io_mpc_reset_run_req,
  output        io_mpc_debug_halt_ack,
  output        io_mpc_debug_run_ack,
  output        io_debug_brkpt_status,
  output        io_dec_tlu_perfcnt0,
  output        io_dec_tlu_perfcnt1,
  output        io_dec_tlu_perfcnt2,
  output        io_dec_tlu_perfcnt3,
  output        io_dccm_wren,
  output        io_dccm_rden,
  output [15:0] io_dccm_wr_addr_lo,
  output [15:0] io_dccm_wr_addr_hi,
  output [15:0] io_dccm_rd_addr_lo,
  output [15:0] io_dccm_rd_addr_hi,
  output [38:0] io_dccm_wr_data_lo,
  output [38:0] io_dccm_wr_data_hi,
  input  [38:0] io_dccm_rd_data_lo,
  input  [38:0] io_dccm_rd_data_hi,
  output [30:0] io_ic_rw_addr,
  output [1:0]  io_ic_tag_valid,
  output        io_ic_rd_en,
  output [70:0] io_ic_debug_wr_data,
  output [9:0]  io_ic_debug_addr,
  input  [63:0] io_ic_rd_data,
  input  [70:0] io_ic_debug_rd_data,
  input  [25:0] io_ic_tag_debug_rd_data,
  input  [1:0]  io_ic_eccerr,
  input  [1:0]  io_ic_rd_hit,
  input         io_ic_tag_perr,
  output        io_ic_debug_rd_en,
  output        io_ic_debug_wr_en,
  output        io_ic_debug_tag_array,
  output [1:0]  io_ic_debug_way,
  output [63:0] io_ic_premux_data,
  output        io_ic_sel_premux_data,
  output [14:0] io_iccm_rw_addr,
  output        io_iccm_buf_correct_ecc,
  output        io_iccm_correction_state,
  output        io_iccm_wren,
  output        io_iccm_rden,
  output [2:0]  io_iccm_wr_size,
  output [77:0] io_iccm_wr_data,
  input  [63:0] io_iccm_rd_data,
  input  [77:0] io_iccm_rd_data_ecc,
  input         io_lsu_bus_clk_en,
  input         io_ifu_bus_clk_en,
  input         io_dbg_bus_clk_en,
  input         io_dma_bus_clk_en,
  input         io_dmi_reg_en,
  input  [6:0]  io_dmi_reg_addr,
  input         io_dmi_reg_wr_en,
  input  [31:0] io_dmi_reg_wdata,
  input  [30:0] io_extintsrc_req,
  input         io_timer_int,
  input         io_soft_int,
  input         io_scan_mode
);
  wire  ifu_clock; // @[quasar.scala 72:19]
  wire  ifu_reset; // @[quasar.scala 72:19]
  wire  ifu_io_exu_flush_final; // @[quasar.scala 72:19]
  wire [30:0] ifu_io_exu_flush_path_final; // @[quasar.scala 72:19]
  wire  ifu_io_free_clk; // @[quasar.scala 72:19]
  wire  ifu_io_active_clk; // @[quasar.scala 72:19]
  wire  ifu_io_ifu_dec_dec_aln_aln_dec_dec_i0_decode_d; // @[quasar.scala 72:19]
  wire [15:0] ifu_io_ifu_dec_dec_aln_aln_dec_ifu_i0_cinst; // @[quasar.scala 72:19]
  wire  ifu_io_ifu_dec_dec_aln_aln_ib_ifu_i0_icaf; // @[quasar.scala 72:19]
  wire [1:0] ifu_io_ifu_dec_dec_aln_aln_ib_ifu_i0_icaf_type; // @[quasar.scala 72:19]
  wire  ifu_io_ifu_dec_dec_aln_aln_ib_ifu_i0_icaf_f1; // @[quasar.scala 72:19]
  wire  ifu_io_ifu_dec_dec_aln_aln_ib_ifu_i0_dbecc; // @[quasar.scala 72:19]
  wire [7:0] ifu_io_ifu_dec_dec_aln_aln_ib_ifu_i0_bp_index; // @[quasar.scala 72:19]
  wire [7:0] ifu_io_ifu_dec_dec_aln_aln_ib_ifu_i0_bp_fghr; // @[quasar.scala 72:19]
  wire [4:0] ifu_io_ifu_dec_dec_aln_aln_ib_ifu_i0_bp_btag; // @[quasar.scala 72:19]
  wire  ifu_io_ifu_dec_dec_aln_aln_ib_ifu_i0_valid; // @[quasar.scala 72:19]
  wire [31:0] ifu_io_ifu_dec_dec_aln_aln_ib_ifu_i0_instr; // @[quasar.scala 72:19]
  wire [30:0] ifu_io_ifu_dec_dec_aln_aln_ib_ifu_i0_pc; // @[quasar.scala 72:19]
  wire  ifu_io_ifu_dec_dec_aln_aln_ib_ifu_i0_pc4; // @[quasar.scala 72:19]
  wire  ifu_io_ifu_dec_dec_aln_aln_ib_i0_brp_valid; // @[quasar.scala 72:19]
  wire [11:0] ifu_io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_toffset; // @[quasar.scala 72:19]
  wire [1:0] ifu_io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_hist; // @[quasar.scala 72:19]
  wire  ifu_io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_br_error; // @[quasar.scala 72:19]
  wire  ifu_io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_br_start_error; // @[quasar.scala 72:19]
  wire [30:0] ifu_io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_prett; // @[quasar.scala 72:19]
  wire  ifu_io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_way; // @[quasar.scala 72:19]
  wire  ifu_io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_ret; // @[quasar.scala 72:19]
  wire  ifu_io_ifu_dec_dec_aln_ifu_pmu_instr_aligned; // @[quasar.scala 72:19]
  wire  ifu_io_ifu_dec_dec_mem_ctrl_dec_tlu_flush_err_wb; // @[quasar.scala 72:19]
  wire  ifu_io_ifu_dec_dec_mem_ctrl_dec_tlu_i0_commit_cmt; // @[quasar.scala 72:19]
  wire  ifu_io_ifu_dec_dec_mem_ctrl_dec_tlu_force_halt; // @[quasar.scala 72:19]
  wire  ifu_io_ifu_dec_dec_mem_ctrl_dec_tlu_fence_i_wb; // @[quasar.scala 72:19]
  wire [70:0] ifu_io_ifu_dec_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_wrdata; // @[quasar.scala 72:19]
  wire [16:0] ifu_io_ifu_dec_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_dicawics; // @[quasar.scala 72:19]
  wire  ifu_io_ifu_dec_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_rd_valid; // @[quasar.scala 72:19]
  wire  ifu_io_ifu_dec_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_wr_valid; // @[quasar.scala 72:19]
  wire  ifu_io_ifu_dec_dec_mem_ctrl_dec_tlu_core_ecc_disable; // @[quasar.scala 72:19]
  wire  ifu_io_ifu_dec_dec_mem_ctrl_ifu_pmu_ic_miss; // @[quasar.scala 72:19]
  wire  ifu_io_ifu_dec_dec_mem_ctrl_ifu_pmu_ic_hit; // @[quasar.scala 72:19]
  wire  ifu_io_ifu_dec_dec_mem_ctrl_ifu_pmu_bus_error; // @[quasar.scala 72:19]
  wire  ifu_io_ifu_dec_dec_mem_ctrl_ifu_pmu_bus_busy; // @[quasar.scala 72:19]
  wire  ifu_io_ifu_dec_dec_mem_ctrl_ifu_ic_error_start; // @[quasar.scala 72:19]
  wire  ifu_io_ifu_dec_dec_mem_ctrl_ifu_iccm_rd_ecc_single_err; // @[quasar.scala 72:19]
  wire [70:0] ifu_io_ifu_dec_dec_mem_ctrl_ifu_ic_debug_rd_data; // @[quasar.scala 72:19]
  wire  ifu_io_ifu_dec_dec_mem_ctrl_ifu_ic_debug_rd_data_valid; // @[quasar.scala 72:19]
  wire  ifu_io_ifu_dec_dec_mem_ctrl_ifu_miss_state_idle; // @[quasar.scala 72:19]
  wire  ifu_io_ifu_dec_dec_ifc_dec_tlu_flush_noredir_wb; // @[quasar.scala 72:19]
  wire [31:0] ifu_io_ifu_dec_dec_ifc_dec_tlu_mrac_ff; // @[quasar.scala 72:19]
  wire  ifu_io_ifu_dec_dec_ifc_ifu_pmu_fetch_stall; // @[quasar.scala 72:19]
  wire  ifu_io_ifu_dec_dec_bp_dec_tlu_br0_r_pkt_valid; // @[quasar.scala 72:19]
  wire [1:0] ifu_io_ifu_dec_dec_bp_dec_tlu_br0_r_pkt_bits_hist; // @[quasar.scala 72:19]
  wire  ifu_io_ifu_dec_dec_bp_dec_tlu_br0_r_pkt_bits_br_error; // @[quasar.scala 72:19]
  wire  ifu_io_ifu_dec_dec_bp_dec_tlu_br0_r_pkt_bits_br_start_error; // @[quasar.scala 72:19]
  wire  ifu_io_ifu_dec_dec_bp_dec_tlu_br0_r_pkt_bits_way; // @[quasar.scala 72:19]
  wire  ifu_io_ifu_dec_dec_bp_dec_tlu_br0_r_pkt_bits_middle; // @[quasar.scala 72:19]
  wire  ifu_io_ifu_dec_dec_bp_dec_tlu_flush_leak_one_wb; // @[quasar.scala 72:19]
  wire  ifu_io_ifu_dec_dec_bp_dec_tlu_bpred_disable; // @[quasar.scala 72:19]
  wire [7:0] ifu_io_exu_ifu_exu_bp_exu_i0_br_index_r; // @[quasar.scala 72:19]
  wire [7:0] ifu_io_exu_ifu_exu_bp_exu_i0_br_fghr_r; // @[quasar.scala 72:19]
  wire  ifu_io_exu_ifu_exu_bp_exu_mp_pkt_bits_misp; // @[quasar.scala 72:19]
  wire  ifu_io_exu_ifu_exu_bp_exu_mp_pkt_bits_ataken; // @[quasar.scala 72:19]
  wire  ifu_io_exu_ifu_exu_bp_exu_mp_pkt_bits_boffset; // @[quasar.scala 72:19]
  wire  ifu_io_exu_ifu_exu_bp_exu_mp_pkt_bits_pc4; // @[quasar.scala 72:19]
  wire [1:0] ifu_io_exu_ifu_exu_bp_exu_mp_pkt_bits_hist; // @[quasar.scala 72:19]
  wire [11:0] ifu_io_exu_ifu_exu_bp_exu_mp_pkt_bits_toffset; // @[quasar.scala 72:19]
  wire  ifu_io_exu_ifu_exu_bp_exu_mp_pkt_bits_pcall; // @[quasar.scala 72:19]
  wire  ifu_io_exu_ifu_exu_bp_exu_mp_pkt_bits_pret; // @[quasar.scala 72:19]
  wire  ifu_io_exu_ifu_exu_bp_exu_mp_pkt_bits_pja; // @[quasar.scala 72:19]
  wire  ifu_io_exu_ifu_exu_bp_exu_mp_pkt_bits_way; // @[quasar.scala 72:19]
  wire [7:0] ifu_io_exu_ifu_exu_bp_exu_mp_eghr; // @[quasar.scala 72:19]
  wire [7:0] ifu_io_exu_ifu_exu_bp_exu_mp_fghr; // @[quasar.scala 72:19]
  wire [7:0] ifu_io_exu_ifu_exu_bp_exu_mp_index; // @[quasar.scala 72:19]
  wire [4:0] ifu_io_exu_ifu_exu_bp_exu_mp_btag; // @[quasar.scala 72:19]
  wire [14:0] ifu_io_iccm_rw_addr; // @[quasar.scala 72:19]
  wire  ifu_io_iccm_buf_correct_ecc; // @[quasar.scala 72:19]
  wire  ifu_io_iccm_correction_state; // @[quasar.scala 72:19]
  wire  ifu_io_iccm_wren; // @[quasar.scala 72:19]
  wire  ifu_io_iccm_rden; // @[quasar.scala 72:19]
  wire [2:0] ifu_io_iccm_wr_size; // @[quasar.scala 72:19]
  wire [77:0] ifu_io_iccm_wr_data; // @[quasar.scala 72:19]
  wire [63:0] ifu_io_iccm_rd_data; // @[quasar.scala 72:19]
  wire [77:0] ifu_io_iccm_rd_data_ecc; // @[quasar.scala 72:19]
  wire [30:0] ifu_io_ic_rw_addr; // @[quasar.scala 72:19]
  wire [1:0] ifu_io_ic_tag_valid; // @[quasar.scala 72:19]
  wire  ifu_io_ic_rd_en; // @[quasar.scala 72:19]
  wire [70:0] ifu_io_ic_debug_wr_data; // @[quasar.scala 72:19]
  wire [9:0] ifu_io_ic_debug_addr; // @[quasar.scala 72:19]
  wire [63:0] ifu_io_ic_rd_data; // @[quasar.scala 72:19]
  wire [70:0] ifu_io_ic_debug_rd_data; // @[quasar.scala 72:19]
  wire [25:0] ifu_io_ic_tag_debug_rd_data; // @[quasar.scala 72:19]
  wire [1:0] ifu_io_ic_eccerr; // @[quasar.scala 72:19]
  wire [1:0] ifu_io_ic_rd_hit; // @[quasar.scala 72:19]
  wire  ifu_io_ic_tag_perr; // @[quasar.scala 72:19]
  wire  ifu_io_ic_debug_rd_en; // @[quasar.scala 72:19]
  wire  ifu_io_ic_debug_wr_en; // @[quasar.scala 72:19]
  wire  ifu_io_ic_debug_tag_array; // @[quasar.scala 72:19]
  wire [1:0] ifu_io_ic_debug_way; // @[quasar.scala 72:19]
  wire [63:0] ifu_io_ic_premux_data; // @[quasar.scala 72:19]
  wire  ifu_io_ic_sel_premux_data; // @[quasar.scala 72:19]
  wire  ifu_io_ifu_ar_valid; // @[quasar.scala 72:19]
  wire [31:0] ifu_io_ifu_ar_bits_addr; // @[quasar.scala 72:19]
  wire  ifu_io_ifu_bus_clk_en; // @[quasar.scala 72:19]
  wire  ifu_io_ifu_dma_dma_ifc_dma_iccm_stall_any; // @[quasar.scala 72:19]
  wire  ifu_io_ifu_dma_dma_mem_ctl_dma_iccm_req; // @[quasar.scala 72:19]
  wire [31:0] ifu_io_ifu_dma_dma_mem_ctl_dma_mem_addr; // @[quasar.scala 72:19]
  wire [2:0] ifu_io_ifu_dma_dma_mem_ctl_dma_mem_sz; // @[quasar.scala 72:19]
  wire  ifu_io_ifu_dma_dma_mem_ctl_dma_mem_write; // @[quasar.scala 72:19]
  wire [63:0] ifu_io_ifu_dma_dma_mem_ctl_dma_mem_wdata; // @[quasar.scala 72:19]
  wire [2:0] ifu_io_ifu_dma_dma_mem_ctl_dma_mem_tag; // @[quasar.scala 72:19]
  wire  ifu_io_iccm_dma_ecc_error; // @[quasar.scala 72:19]
  wire  ifu_io_iccm_dma_rvalid; // @[quasar.scala 72:19]
  wire [63:0] ifu_io_iccm_dma_rdata; // @[quasar.scala 72:19]
  wire [2:0] ifu_io_iccm_dma_rtag; // @[quasar.scala 72:19]
  wire  ifu_io_iccm_ready; // @[quasar.scala 72:19]
  wire  ifu_io_iccm_dma_sb_error; // @[quasar.scala 72:19]
  wire  ifu_io_dec_tlu_flush_lower_wb; // @[quasar.scala 72:19]
  wire  ifu_io_scan_mode; // @[quasar.scala 72:19]
  wire  dec_clock; // @[quasar.scala 73:19]
  wire  dec_reset; // @[quasar.scala 73:19]
  wire  dec_io_free_clk; // @[quasar.scala 73:19]
  wire  dec_io_active_clk; // @[quasar.scala 73:19]
  wire  dec_io_lsu_fastint_stall_any; // @[quasar.scala 73:19]
  wire  dec_io_dec_pause_state_cg; // @[quasar.scala 73:19]
  wire [30:0] dec_io_rst_vec; // @[quasar.scala 73:19]
  wire  dec_io_nmi_int; // @[quasar.scala 73:19]
  wire [30:0] dec_io_nmi_vec; // @[quasar.scala 73:19]
  wire  dec_io_i_cpu_halt_req; // @[quasar.scala 73:19]
  wire  dec_io_i_cpu_run_req; // @[quasar.scala 73:19]
  wire  dec_io_o_cpu_halt_status; // @[quasar.scala 73:19]
  wire  dec_io_o_cpu_halt_ack; // @[quasar.scala 73:19]
  wire  dec_io_o_cpu_run_ack; // @[quasar.scala 73:19]
  wire  dec_io_o_debug_mode_status; // @[quasar.scala 73:19]
  wire [27:0] dec_io_core_id; // @[quasar.scala 73:19]
  wire  dec_io_mpc_debug_halt_req; // @[quasar.scala 73:19]
  wire  dec_io_mpc_debug_run_req; // @[quasar.scala 73:19]
  wire  dec_io_mpc_reset_run_req; // @[quasar.scala 73:19]
  wire  dec_io_mpc_debug_halt_ack; // @[quasar.scala 73:19]
  wire  dec_io_mpc_debug_run_ack; // @[quasar.scala 73:19]
  wire  dec_io_debug_brkpt_status; // @[quasar.scala 73:19]
  wire  dec_io_lsu_pmu_misaligned_m; // @[quasar.scala 73:19]
  wire [30:0] dec_io_lsu_fir_addr; // @[quasar.scala 73:19]
  wire [1:0] dec_io_lsu_fir_error; // @[quasar.scala 73:19]
  wire [3:0] dec_io_lsu_trigger_match_m; // @[quasar.scala 73:19]
  wire  dec_io_lsu_idle_any; // @[quasar.scala 73:19]
  wire  dec_io_lsu_error_pkt_r_valid; // @[quasar.scala 73:19]
  wire  dec_io_lsu_error_pkt_r_bits_single_ecc_error; // @[quasar.scala 73:19]
  wire  dec_io_lsu_error_pkt_r_bits_inst_type; // @[quasar.scala 73:19]
  wire  dec_io_lsu_error_pkt_r_bits_exc_type; // @[quasar.scala 73:19]
  wire [3:0] dec_io_lsu_error_pkt_r_bits_mscause; // @[quasar.scala 73:19]
  wire [31:0] dec_io_lsu_error_pkt_r_bits_addr; // @[quasar.scala 73:19]
  wire  dec_io_lsu_single_ecc_error_incr; // @[quasar.scala 73:19]
  wire [31:0] dec_io_exu_div_result; // @[quasar.scala 73:19]
  wire  dec_io_exu_div_wren; // @[quasar.scala 73:19]
  wire [31:0] dec_io_lsu_result_m; // @[quasar.scala 73:19]
  wire [31:0] dec_io_lsu_result_corr_r; // @[quasar.scala 73:19]
  wire  dec_io_lsu_load_stall_any; // @[quasar.scala 73:19]
  wire  dec_io_lsu_store_stall_any; // @[quasar.scala 73:19]
  wire  dec_io_iccm_dma_sb_error; // @[quasar.scala 73:19]
  wire  dec_io_exu_flush_final; // @[quasar.scala 73:19]
  wire  dec_io_timer_int; // @[quasar.scala 73:19]
  wire  dec_io_soft_int; // @[quasar.scala 73:19]
  wire  dec_io_dbg_halt_req; // @[quasar.scala 73:19]
  wire  dec_io_dbg_resume_req; // @[quasar.scala 73:19]
  wire  dec_io_dec_tlu_dbg_halted; // @[quasar.scala 73:19]
  wire  dec_io_dec_tlu_debug_mode; // @[quasar.scala 73:19]
  wire  dec_io_dec_tlu_resume_ack; // @[quasar.scala 73:19]
  wire  dec_io_dec_tlu_mpc_halted_only; // @[quasar.scala 73:19]
  wire [31:0] dec_io_dec_dbg_rddata; // @[quasar.scala 73:19]
  wire  dec_io_dec_dbg_cmd_done; // @[quasar.scala 73:19]
  wire  dec_io_dec_dbg_cmd_fail; // @[quasar.scala 73:19]
  wire  dec_io_trigger_pkt_any_0_select; // @[quasar.scala 73:19]
  wire  dec_io_trigger_pkt_any_0_match_pkt; // @[quasar.scala 73:19]
  wire  dec_io_trigger_pkt_any_0_store; // @[quasar.scala 73:19]
  wire  dec_io_trigger_pkt_any_0_load; // @[quasar.scala 73:19]
  wire [31:0] dec_io_trigger_pkt_any_0_tdata2; // @[quasar.scala 73:19]
  wire  dec_io_trigger_pkt_any_1_select; // @[quasar.scala 73:19]
  wire  dec_io_trigger_pkt_any_1_match_pkt; // @[quasar.scala 73:19]
  wire  dec_io_trigger_pkt_any_1_store; // @[quasar.scala 73:19]
  wire  dec_io_trigger_pkt_any_1_load; // @[quasar.scala 73:19]
  wire [31:0] dec_io_trigger_pkt_any_1_tdata2; // @[quasar.scala 73:19]
  wire  dec_io_trigger_pkt_any_2_select; // @[quasar.scala 73:19]
  wire  dec_io_trigger_pkt_any_2_match_pkt; // @[quasar.scala 73:19]
  wire  dec_io_trigger_pkt_any_2_store; // @[quasar.scala 73:19]
  wire  dec_io_trigger_pkt_any_2_load; // @[quasar.scala 73:19]
  wire [31:0] dec_io_trigger_pkt_any_2_tdata2; // @[quasar.scala 73:19]
  wire  dec_io_trigger_pkt_any_3_select; // @[quasar.scala 73:19]
  wire  dec_io_trigger_pkt_any_3_match_pkt; // @[quasar.scala 73:19]
  wire  dec_io_trigger_pkt_any_3_store; // @[quasar.scala 73:19]
  wire  dec_io_trigger_pkt_any_3_load; // @[quasar.scala 73:19]
  wire [31:0] dec_io_trigger_pkt_any_3_tdata2; // @[quasar.scala 73:19]
  wire  dec_io_exu_i0_br_way_r; // @[quasar.scala 73:19]
  wire  dec_io_lsu_p_valid; // @[quasar.scala 73:19]
  wire  dec_io_lsu_p_bits_fast_int; // @[quasar.scala 73:19]
  wire  dec_io_lsu_p_bits_by; // @[quasar.scala 73:19]
  wire  dec_io_lsu_p_bits_half; // @[quasar.scala 73:19]
  wire  dec_io_lsu_p_bits_word; // @[quasar.scala 73:19]
  wire  dec_io_lsu_p_bits_load; // @[quasar.scala 73:19]
  wire  dec_io_lsu_p_bits_store; // @[quasar.scala 73:19]
  wire  dec_io_lsu_p_bits_unsign; // @[quasar.scala 73:19]
  wire  dec_io_lsu_p_bits_store_data_bypass_d; // @[quasar.scala 73:19]
  wire  dec_io_lsu_p_bits_load_ldst_bypass_d; // @[quasar.scala 73:19]
  wire [11:0] dec_io_dec_lsu_offset_d; // @[quasar.scala 73:19]
  wire  dec_io_dec_tlu_i0_kill_writeb_r; // @[quasar.scala 73:19]
  wire  dec_io_dec_tlu_perfcnt0; // @[quasar.scala 73:19]
  wire  dec_io_dec_tlu_perfcnt1; // @[quasar.scala 73:19]
  wire  dec_io_dec_tlu_perfcnt2; // @[quasar.scala 73:19]
  wire  dec_io_dec_tlu_perfcnt3; // @[quasar.scala 73:19]
  wire  dec_io_dec_lsu_valid_raw_d; // @[quasar.scala 73:19]
  wire [1:0] dec_io_rv_trace_pkt_rv_i_valid_ip; // @[quasar.scala 73:19]
  wire [31:0] dec_io_rv_trace_pkt_rv_i_insn_ip; // @[quasar.scala 73:19]
  wire [31:0] dec_io_rv_trace_pkt_rv_i_address_ip; // @[quasar.scala 73:19]
  wire [1:0] dec_io_rv_trace_pkt_rv_i_exception_ip; // @[quasar.scala 73:19]
  wire [4:0] dec_io_rv_trace_pkt_rv_i_ecause_ip; // @[quasar.scala 73:19]
  wire [1:0] dec_io_rv_trace_pkt_rv_i_interrupt_ip; // @[quasar.scala 73:19]
  wire [31:0] dec_io_rv_trace_pkt_rv_i_tval_ip; // @[quasar.scala 73:19]
  wire  dec_io_dec_tlu_misc_clk_override; // @[quasar.scala 73:19]
  wire  dec_io_dec_tlu_lsu_clk_override; // @[quasar.scala 73:19]
  wire  dec_io_dec_tlu_bus_clk_override; // @[quasar.scala 73:19]
  wire  dec_io_dec_tlu_pic_clk_override; // @[quasar.scala 73:19]
  wire  dec_io_dec_tlu_dccm_clk_override; // @[quasar.scala 73:19]
  wire  dec_io_dec_tlu_icm_clk_override; // @[quasar.scala 73:19]
  wire  dec_io_scan_mode; // @[quasar.scala 73:19]
  wire  dec_io_ifu_dec_dec_aln_aln_dec_dec_i0_decode_d; // @[quasar.scala 73:19]
  wire [15:0] dec_io_ifu_dec_dec_aln_aln_dec_ifu_i0_cinst; // @[quasar.scala 73:19]
  wire  dec_io_ifu_dec_dec_aln_aln_ib_ifu_i0_icaf; // @[quasar.scala 73:19]
  wire [1:0] dec_io_ifu_dec_dec_aln_aln_ib_ifu_i0_icaf_type; // @[quasar.scala 73:19]
  wire  dec_io_ifu_dec_dec_aln_aln_ib_ifu_i0_icaf_f1; // @[quasar.scala 73:19]
  wire  dec_io_ifu_dec_dec_aln_aln_ib_ifu_i0_dbecc; // @[quasar.scala 73:19]
  wire [7:0] dec_io_ifu_dec_dec_aln_aln_ib_ifu_i0_bp_index; // @[quasar.scala 73:19]
  wire [7:0] dec_io_ifu_dec_dec_aln_aln_ib_ifu_i0_bp_fghr; // @[quasar.scala 73:19]
  wire [4:0] dec_io_ifu_dec_dec_aln_aln_ib_ifu_i0_bp_btag; // @[quasar.scala 73:19]
  wire  dec_io_ifu_dec_dec_aln_aln_ib_ifu_i0_valid; // @[quasar.scala 73:19]
  wire [31:0] dec_io_ifu_dec_dec_aln_aln_ib_ifu_i0_instr; // @[quasar.scala 73:19]
  wire [30:0] dec_io_ifu_dec_dec_aln_aln_ib_ifu_i0_pc; // @[quasar.scala 73:19]
  wire  dec_io_ifu_dec_dec_aln_aln_ib_ifu_i0_pc4; // @[quasar.scala 73:19]
  wire  dec_io_ifu_dec_dec_aln_aln_ib_i0_brp_valid; // @[quasar.scala 73:19]
  wire [11:0] dec_io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_toffset; // @[quasar.scala 73:19]
  wire [1:0] dec_io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_hist; // @[quasar.scala 73:19]
  wire  dec_io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_br_error; // @[quasar.scala 73:19]
  wire  dec_io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_br_start_error; // @[quasar.scala 73:19]
  wire [30:0] dec_io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_prett; // @[quasar.scala 73:19]
  wire  dec_io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_way; // @[quasar.scala 73:19]
  wire  dec_io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_ret; // @[quasar.scala 73:19]
  wire  dec_io_ifu_dec_dec_aln_ifu_pmu_instr_aligned; // @[quasar.scala 73:19]
  wire  dec_io_ifu_dec_dec_mem_ctrl_dec_tlu_flush_err_wb; // @[quasar.scala 73:19]
  wire  dec_io_ifu_dec_dec_mem_ctrl_dec_tlu_i0_commit_cmt; // @[quasar.scala 73:19]
  wire  dec_io_ifu_dec_dec_mem_ctrl_dec_tlu_force_halt; // @[quasar.scala 73:19]
  wire  dec_io_ifu_dec_dec_mem_ctrl_dec_tlu_fence_i_wb; // @[quasar.scala 73:19]
  wire [70:0] dec_io_ifu_dec_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_wrdata; // @[quasar.scala 73:19]
  wire [16:0] dec_io_ifu_dec_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_dicawics; // @[quasar.scala 73:19]
  wire  dec_io_ifu_dec_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_rd_valid; // @[quasar.scala 73:19]
  wire  dec_io_ifu_dec_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_wr_valid; // @[quasar.scala 73:19]
  wire  dec_io_ifu_dec_dec_mem_ctrl_dec_tlu_core_ecc_disable; // @[quasar.scala 73:19]
  wire  dec_io_ifu_dec_dec_mem_ctrl_ifu_pmu_ic_miss; // @[quasar.scala 73:19]
  wire  dec_io_ifu_dec_dec_mem_ctrl_ifu_pmu_ic_hit; // @[quasar.scala 73:19]
  wire  dec_io_ifu_dec_dec_mem_ctrl_ifu_pmu_bus_error; // @[quasar.scala 73:19]
  wire  dec_io_ifu_dec_dec_mem_ctrl_ifu_pmu_bus_busy; // @[quasar.scala 73:19]
  wire  dec_io_ifu_dec_dec_mem_ctrl_ifu_ic_error_start; // @[quasar.scala 73:19]
  wire  dec_io_ifu_dec_dec_mem_ctrl_ifu_iccm_rd_ecc_single_err; // @[quasar.scala 73:19]
  wire [70:0] dec_io_ifu_dec_dec_mem_ctrl_ifu_ic_debug_rd_data; // @[quasar.scala 73:19]
  wire  dec_io_ifu_dec_dec_mem_ctrl_ifu_ic_debug_rd_data_valid; // @[quasar.scala 73:19]
  wire  dec_io_ifu_dec_dec_mem_ctrl_ifu_miss_state_idle; // @[quasar.scala 73:19]
  wire  dec_io_ifu_dec_dec_ifc_dec_tlu_flush_noredir_wb; // @[quasar.scala 73:19]
  wire [31:0] dec_io_ifu_dec_dec_ifc_dec_tlu_mrac_ff; // @[quasar.scala 73:19]
  wire  dec_io_ifu_dec_dec_ifc_ifu_pmu_fetch_stall; // @[quasar.scala 73:19]
  wire  dec_io_ifu_dec_dec_bp_dec_tlu_br0_r_pkt_valid; // @[quasar.scala 73:19]
  wire [1:0] dec_io_ifu_dec_dec_bp_dec_tlu_br0_r_pkt_bits_hist; // @[quasar.scala 73:19]
  wire  dec_io_ifu_dec_dec_bp_dec_tlu_br0_r_pkt_bits_br_error; // @[quasar.scala 73:19]
  wire  dec_io_ifu_dec_dec_bp_dec_tlu_br0_r_pkt_bits_br_start_error; // @[quasar.scala 73:19]
  wire  dec_io_ifu_dec_dec_bp_dec_tlu_br0_r_pkt_bits_way; // @[quasar.scala 73:19]
  wire  dec_io_ifu_dec_dec_bp_dec_tlu_br0_r_pkt_bits_middle; // @[quasar.scala 73:19]
  wire  dec_io_ifu_dec_dec_bp_dec_tlu_flush_leak_one_wb; // @[quasar.scala 73:19]
  wire  dec_io_ifu_dec_dec_bp_dec_tlu_bpred_disable; // @[quasar.scala 73:19]
  wire  dec_io_dec_exu_dec_alu_dec_i0_alu_decode_d; // @[quasar.scala 73:19]
  wire  dec_io_dec_exu_dec_alu_dec_csr_ren_d; // @[quasar.scala 73:19]
  wire [11:0] dec_io_dec_exu_dec_alu_dec_i0_br_immed_d; // @[quasar.scala 73:19]
  wire [30:0] dec_io_dec_exu_dec_alu_exu_i0_pc_x; // @[quasar.scala 73:19]
  wire  dec_io_dec_exu_dec_div_div_p_valid; // @[quasar.scala 73:19]
  wire  dec_io_dec_exu_dec_div_div_p_bits_unsign; // @[quasar.scala 73:19]
  wire  dec_io_dec_exu_dec_div_div_p_bits_rem; // @[quasar.scala 73:19]
  wire  dec_io_dec_exu_dec_div_dec_div_cancel; // @[quasar.scala 73:19]
  wire [1:0] dec_io_dec_exu_decode_exu_dec_data_en; // @[quasar.scala 73:19]
  wire [1:0] dec_io_dec_exu_decode_exu_dec_ctl_en; // @[quasar.scala 73:19]
  wire  dec_io_dec_exu_decode_exu_i0_ap_land; // @[quasar.scala 73:19]
  wire  dec_io_dec_exu_decode_exu_i0_ap_lor; // @[quasar.scala 73:19]
  wire  dec_io_dec_exu_decode_exu_i0_ap_lxor; // @[quasar.scala 73:19]
  wire  dec_io_dec_exu_decode_exu_i0_ap_sll; // @[quasar.scala 73:19]
  wire  dec_io_dec_exu_decode_exu_i0_ap_srl; // @[quasar.scala 73:19]
  wire  dec_io_dec_exu_decode_exu_i0_ap_sra; // @[quasar.scala 73:19]
  wire  dec_io_dec_exu_decode_exu_i0_ap_beq; // @[quasar.scala 73:19]
  wire  dec_io_dec_exu_decode_exu_i0_ap_bne; // @[quasar.scala 73:19]
  wire  dec_io_dec_exu_decode_exu_i0_ap_blt; // @[quasar.scala 73:19]
  wire  dec_io_dec_exu_decode_exu_i0_ap_bge; // @[quasar.scala 73:19]
  wire  dec_io_dec_exu_decode_exu_i0_ap_add; // @[quasar.scala 73:19]
  wire  dec_io_dec_exu_decode_exu_i0_ap_sub; // @[quasar.scala 73:19]
  wire  dec_io_dec_exu_decode_exu_i0_ap_slt; // @[quasar.scala 73:19]
  wire  dec_io_dec_exu_decode_exu_i0_ap_unsign; // @[quasar.scala 73:19]
  wire  dec_io_dec_exu_decode_exu_i0_ap_jal; // @[quasar.scala 73:19]
  wire  dec_io_dec_exu_decode_exu_i0_ap_predict_t; // @[quasar.scala 73:19]
  wire  dec_io_dec_exu_decode_exu_i0_ap_predict_nt; // @[quasar.scala 73:19]
  wire  dec_io_dec_exu_decode_exu_i0_ap_csr_write; // @[quasar.scala 73:19]
  wire  dec_io_dec_exu_decode_exu_i0_ap_csr_imm; // @[quasar.scala 73:19]
  wire  dec_io_dec_exu_decode_exu_dec_i0_predict_p_d_valid; // @[quasar.scala 73:19]
  wire  dec_io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_pc4; // @[quasar.scala 73:19]
  wire [1:0] dec_io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_hist; // @[quasar.scala 73:19]
  wire [11:0] dec_io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_toffset; // @[quasar.scala 73:19]
  wire  dec_io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_br_error; // @[quasar.scala 73:19]
  wire  dec_io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_br_start_error; // @[quasar.scala 73:19]
  wire [30:0] dec_io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_prett; // @[quasar.scala 73:19]
  wire  dec_io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_pcall; // @[quasar.scala 73:19]
  wire  dec_io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_pret; // @[quasar.scala 73:19]
  wire  dec_io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_pja; // @[quasar.scala 73:19]
  wire  dec_io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_way; // @[quasar.scala 73:19]
  wire [7:0] dec_io_dec_exu_decode_exu_i0_predict_fghr_d; // @[quasar.scala 73:19]
  wire [7:0] dec_io_dec_exu_decode_exu_i0_predict_index_d; // @[quasar.scala 73:19]
  wire [4:0] dec_io_dec_exu_decode_exu_i0_predict_btag_d; // @[quasar.scala 73:19]
  wire  dec_io_dec_exu_decode_exu_dec_i0_rs1_en_d; // @[quasar.scala 73:19]
  wire  dec_io_dec_exu_decode_exu_dec_i0_rs2_en_d; // @[quasar.scala 73:19]
  wire [31:0] dec_io_dec_exu_decode_exu_dec_i0_immed_d; // @[quasar.scala 73:19]
  wire [31:0] dec_io_dec_exu_decode_exu_dec_i0_rs1_bypass_data_d; // @[quasar.scala 73:19]
  wire [31:0] dec_io_dec_exu_decode_exu_dec_i0_rs2_bypass_data_d; // @[quasar.scala 73:19]
  wire  dec_io_dec_exu_decode_exu_dec_i0_select_pc_d; // @[quasar.scala 73:19]
  wire [1:0] dec_io_dec_exu_decode_exu_dec_i0_rs1_bypass_en_d; // @[quasar.scala 73:19]
  wire [1:0] dec_io_dec_exu_decode_exu_dec_i0_rs2_bypass_en_d; // @[quasar.scala 73:19]
  wire  dec_io_dec_exu_decode_exu_mul_p_valid; // @[quasar.scala 73:19]
  wire  dec_io_dec_exu_decode_exu_mul_p_bits_rs1_sign; // @[quasar.scala 73:19]
  wire  dec_io_dec_exu_decode_exu_mul_p_bits_rs2_sign; // @[quasar.scala 73:19]
  wire  dec_io_dec_exu_decode_exu_mul_p_bits_low; // @[quasar.scala 73:19]
  wire [30:0] dec_io_dec_exu_decode_exu_pred_correct_npc_x; // @[quasar.scala 73:19]
  wire  dec_io_dec_exu_decode_exu_dec_extint_stall; // @[quasar.scala 73:19]
  wire [31:0] dec_io_dec_exu_decode_exu_exu_i0_result_x; // @[quasar.scala 73:19]
  wire [31:0] dec_io_dec_exu_decode_exu_exu_csr_rs1_x; // @[quasar.scala 73:19]
  wire [29:0] dec_io_dec_exu_tlu_exu_dec_tlu_meihap; // @[quasar.scala 73:19]
  wire  dec_io_dec_exu_tlu_exu_dec_tlu_flush_lower_r; // @[quasar.scala 73:19]
  wire [30:0] dec_io_dec_exu_tlu_exu_dec_tlu_flush_path_r; // @[quasar.scala 73:19]
  wire [1:0] dec_io_dec_exu_tlu_exu_exu_i0_br_hist_r; // @[quasar.scala 73:19]
  wire  dec_io_dec_exu_tlu_exu_exu_i0_br_error_r; // @[quasar.scala 73:19]
  wire  dec_io_dec_exu_tlu_exu_exu_i0_br_start_error_r; // @[quasar.scala 73:19]
  wire  dec_io_dec_exu_tlu_exu_exu_i0_br_valid_r; // @[quasar.scala 73:19]
  wire  dec_io_dec_exu_tlu_exu_exu_i0_br_mp_r; // @[quasar.scala 73:19]
  wire  dec_io_dec_exu_tlu_exu_exu_i0_br_middle_r; // @[quasar.scala 73:19]
  wire  dec_io_dec_exu_tlu_exu_exu_pmu_i0_br_misp; // @[quasar.scala 73:19]
  wire  dec_io_dec_exu_tlu_exu_exu_pmu_i0_br_ataken; // @[quasar.scala 73:19]
  wire  dec_io_dec_exu_tlu_exu_exu_pmu_i0_pc4; // @[quasar.scala 73:19]
  wire [30:0] dec_io_dec_exu_tlu_exu_exu_npc_r; // @[quasar.scala 73:19]
  wire [30:0] dec_io_dec_exu_ib_exu_dec_i0_pc_d; // @[quasar.scala 73:19]
  wire  dec_io_dec_exu_ib_exu_dec_debug_wdata_rs1_d; // @[quasar.scala 73:19]
  wire [31:0] dec_io_dec_exu_gpr_exu_gpr_i0_rs1_d; // @[quasar.scala 73:19]
  wire [31:0] dec_io_dec_exu_gpr_exu_gpr_i0_rs2_d; // @[quasar.scala 73:19]
  wire  dec_io_lsu_dec_tlu_busbuff_lsu_pmu_bus_misaligned; // @[quasar.scala 73:19]
  wire  dec_io_lsu_dec_tlu_busbuff_lsu_pmu_bus_error; // @[quasar.scala 73:19]
  wire  dec_io_lsu_dec_tlu_busbuff_lsu_pmu_bus_busy; // @[quasar.scala 73:19]
  wire  dec_io_lsu_dec_tlu_busbuff_dec_tlu_external_ldfwd_disable; // @[quasar.scala 73:19]
  wire  dec_io_lsu_dec_tlu_busbuff_dec_tlu_wb_coalescing_disable; // @[quasar.scala 73:19]
  wire  dec_io_lsu_dec_tlu_busbuff_dec_tlu_sideeffect_posted_disable; // @[quasar.scala 73:19]
  wire  dec_io_lsu_dec_tlu_busbuff_lsu_imprecise_error_load_any; // @[quasar.scala 73:19]
  wire  dec_io_lsu_dec_tlu_busbuff_lsu_imprecise_error_store_any; // @[quasar.scala 73:19]
  wire [31:0] dec_io_lsu_dec_tlu_busbuff_lsu_imprecise_error_addr_any; // @[quasar.scala 73:19]
  wire  dec_io_lsu_dec_dctl_busbuff_lsu_nonblock_load_valid_m; // @[quasar.scala 73:19]
  wire [1:0] dec_io_lsu_dec_dctl_busbuff_lsu_nonblock_load_tag_m; // @[quasar.scala 73:19]
  wire  dec_io_lsu_dec_dctl_busbuff_lsu_nonblock_load_inv_r; // @[quasar.scala 73:19]
  wire [1:0] dec_io_lsu_dec_dctl_busbuff_lsu_nonblock_load_inv_tag_r; // @[quasar.scala 73:19]
  wire  dec_io_lsu_dec_dctl_busbuff_lsu_nonblock_load_data_valid; // @[quasar.scala 73:19]
  wire  dec_io_lsu_dec_dctl_busbuff_lsu_nonblock_load_data_error; // @[quasar.scala 73:19]
  wire [1:0] dec_io_lsu_dec_dctl_busbuff_lsu_nonblock_load_data_tag; // @[quasar.scala 73:19]
  wire [31:0] dec_io_lsu_dec_dctl_busbuff_lsu_nonblock_load_data; // @[quasar.scala 73:19]
  wire  dec_io_lsu_tlu_lsu_pmu_load_external_m; // @[quasar.scala 73:19]
  wire  dec_io_lsu_tlu_lsu_pmu_store_external_m; // @[quasar.scala 73:19]
  wire  dec_io_dec_dbg_dbg_ib_dbg_cmd_valid; // @[quasar.scala 73:19]
  wire  dec_io_dec_dbg_dbg_ib_dbg_cmd_write; // @[quasar.scala 73:19]
  wire [1:0] dec_io_dec_dbg_dbg_ib_dbg_cmd_type; // @[quasar.scala 73:19]
  wire [31:0] dec_io_dec_dbg_dbg_ib_dbg_cmd_addr; // @[quasar.scala 73:19]
  wire [31:0] dec_io_dec_dbg_dbg_dctl_dbg_cmd_wrdata; // @[quasar.scala 73:19]
  wire  dec_io_dec_dma_dctl_dma_dma_dccm_stall_any; // @[quasar.scala 73:19]
  wire  dec_io_dec_dma_tlu_dma_dma_pmu_dccm_read; // @[quasar.scala 73:19]
  wire  dec_io_dec_dma_tlu_dma_dma_pmu_dccm_write; // @[quasar.scala 73:19]
  wire  dec_io_dec_dma_tlu_dma_dma_pmu_any_read; // @[quasar.scala 73:19]
  wire  dec_io_dec_dma_tlu_dma_dma_pmu_any_write; // @[quasar.scala 73:19]
  wire [2:0] dec_io_dec_dma_tlu_dma_dec_tlu_dma_qos_prty; // @[quasar.scala 73:19]
  wire  dec_io_dec_dma_tlu_dma_dma_dccm_stall_any; // @[quasar.scala 73:19]
  wire  dec_io_dec_dma_tlu_dma_dma_iccm_stall_any; // @[quasar.scala 73:19]
  wire [7:0] dec_io_dec_pic_pic_claimid; // @[quasar.scala 73:19]
  wire [3:0] dec_io_dec_pic_pic_pl; // @[quasar.scala 73:19]
  wire  dec_io_dec_pic_mhwakeup; // @[quasar.scala 73:19]
  wire [3:0] dec_io_dec_pic_dec_tlu_meicurpl; // @[quasar.scala 73:19]
  wire [3:0] dec_io_dec_pic_dec_tlu_meipt; // @[quasar.scala 73:19]
  wire  dec_io_dec_pic_mexintpend; // @[quasar.scala 73:19]
  wire  dbg_clock; // @[quasar.scala 74:19]
  wire  dbg_reset; // @[quasar.scala 74:19]
  wire [1:0] dbg_io_dbg_cmd_size; // @[quasar.scala 74:19]
  wire  dbg_io_dbg_core_rst_l; // @[quasar.scala 74:19]
  wire [31:0] dbg_io_core_dbg_rddata; // @[quasar.scala 74:19]
  wire  dbg_io_core_dbg_cmd_done; // @[quasar.scala 74:19]
  wire  dbg_io_core_dbg_cmd_fail; // @[quasar.scala 74:19]
  wire  dbg_io_dbg_halt_req; // @[quasar.scala 74:19]
  wire  dbg_io_dbg_resume_req; // @[quasar.scala 74:19]
  wire  dbg_io_dec_tlu_debug_mode; // @[quasar.scala 74:19]
  wire  dbg_io_dec_tlu_dbg_halted; // @[quasar.scala 74:19]
  wire  dbg_io_dec_tlu_mpc_halted_only; // @[quasar.scala 74:19]
  wire  dbg_io_dec_tlu_resume_ack; // @[quasar.scala 74:19]
  wire  dbg_io_dmi_reg_en; // @[quasar.scala 74:19]
  wire [6:0] dbg_io_dmi_reg_addr; // @[quasar.scala 74:19]
  wire  dbg_io_dmi_reg_wr_en; // @[quasar.scala 74:19]
  wire [31:0] dbg_io_dmi_reg_wdata; // @[quasar.scala 74:19]
  wire  dbg_io_sb_axi_aw_valid; // @[quasar.scala 74:19]
  wire [31:0] dbg_io_sb_axi_aw_bits_addr; // @[quasar.scala 74:19]
  wire [2:0] dbg_io_sb_axi_aw_bits_size; // @[quasar.scala 74:19]
  wire  dbg_io_sb_axi_w_valid; // @[quasar.scala 74:19]
  wire [7:0] dbg_io_sb_axi_w_bits_strb; // @[quasar.scala 74:19]
  wire  dbg_io_sb_axi_ar_valid; // @[quasar.scala 74:19]
  wire [31:0] dbg_io_sb_axi_ar_bits_addr; // @[quasar.scala 74:19]
  wire [2:0] dbg_io_sb_axi_ar_bits_size; // @[quasar.scala 74:19]
  wire  dbg_io_dbg_dec_dbg_ib_dbg_cmd_valid; // @[quasar.scala 74:19]
  wire  dbg_io_dbg_dec_dbg_ib_dbg_cmd_write; // @[quasar.scala 74:19]
  wire [1:0] dbg_io_dbg_dec_dbg_ib_dbg_cmd_type; // @[quasar.scala 74:19]
  wire [31:0] dbg_io_dbg_dec_dbg_ib_dbg_cmd_addr; // @[quasar.scala 74:19]
  wire [31:0] dbg_io_dbg_dec_dbg_dctl_dbg_cmd_wrdata; // @[quasar.scala 74:19]
  wire  dbg_io_dbg_dma_dbg_ib_dbg_cmd_valid; // @[quasar.scala 74:19]
  wire  dbg_io_dbg_dma_dbg_ib_dbg_cmd_write; // @[quasar.scala 74:19]
  wire [1:0] dbg_io_dbg_dma_dbg_ib_dbg_cmd_type; // @[quasar.scala 74:19]
  wire [31:0] dbg_io_dbg_dma_dbg_ib_dbg_cmd_addr; // @[quasar.scala 74:19]
  wire [31:0] dbg_io_dbg_dma_dbg_dctl_dbg_cmd_wrdata; // @[quasar.scala 74:19]
  wire  dbg_io_dbg_dma_io_dbg_dma_bubble; // @[quasar.scala 74:19]
  wire  dbg_io_dbg_dma_io_dma_dbg_ready; // @[quasar.scala 74:19]
  wire  dbg_io_dbg_bus_clk_en; // @[quasar.scala 74:19]
  wire  dbg_io_dbg_rst_l; // @[quasar.scala 74:19]
  wire  dbg_io_clk_override; // @[quasar.scala 74:19]
  wire  dbg_io_scan_mode; // @[quasar.scala 74:19]
  wire  exu_clock; // @[quasar.scala 75:19]
  wire  exu_reset; // @[quasar.scala 75:19]
  wire  exu_io_scan_mode; // @[quasar.scala 75:19]
  wire  exu_io_dec_exu_dec_alu_dec_i0_alu_decode_d; // @[quasar.scala 75:19]
  wire  exu_io_dec_exu_dec_alu_dec_csr_ren_d; // @[quasar.scala 75:19]
  wire [11:0] exu_io_dec_exu_dec_alu_dec_i0_br_immed_d; // @[quasar.scala 75:19]
  wire [30:0] exu_io_dec_exu_dec_alu_exu_i0_pc_x; // @[quasar.scala 75:19]
  wire  exu_io_dec_exu_dec_div_div_p_valid; // @[quasar.scala 75:19]
  wire  exu_io_dec_exu_dec_div_div_p_bits_unsign; // @[quasar.scala 75:19]
  wire  exu_io_dec_exu_dec_div_div_p_bits_rem; // @[quasar.scala 75:19]
  wire  exu_io_dec_exu_dec_div_dec_div_cancel; // @[quasar.scala 75:19]
  wire [1:0] exu_io_dec_exu_decode_exu_dec_data_en; // @[quasar.scala 75:19]
  wire [1:0] exu_io_dec_exu_decode_exu_dec_ctl_en; // @[quasar.scala 75:19]
  wire  exu_io_dec_exu_decode_exu_i0_ap_land; // @[quasar.scala 75:19]
  wire  exu_io_dec_exu_decode_exu_i0_ap_lor; // @[quasar.scala 75:19]
  wire  exu_io_dec_exu_decode_exu_i0_ap_lxor; // @[quasar.scala 75:19]
  wire  exu_io_dec_exu_decode_exu_i0_ap_sll; // @[quasar.scala 75:19]
  wire  exu_io_dec_exu_decode_exu_i0_ap_srl; // @[quasar.scala 75:19]
  wire  exu_io_dec_exu_decode_exu_i0_ap_sra; // @[quasar.scala 75:19]
  wire  exu_io_dec_exu_decode_exu_i0_ap_beq; // @[quasar.scala 75:19]
  wire  exu_io_dec_exu_decode_exu_i0_ap_bne; // @[quasar.scala 75:19]
  wire  exu_io_dec_exu_decode_exu_i0_ap_blt; // @[quasar.scala 75:19]
  wire  exu_io_dec_exu_decode_exu_i0_ap_bge; // @[quasar.scala 75:19]
  wire  exu_io_dec_exu_decode_exu_i0_ap_add; // @[quasar.scala 75:19]
  wire  exu_io_dec_exu_decode_exu_i0_ap_sub; // @[quasar.scala 75:19]
  wire  exu_io_dec_exu_decode_exu_i0_ap_slt; // @[quasar.scala 75:19]
  wire  exu_io_dec_exu_decode_exu_i0_ap_unsign; // @[quasar.scala 75:19]
  wire  exu_io_dec_exu_decode_exu_i0_ap_jal; // @[quasar.scala 75:19]
  wire  exu_io_dec_exu_decode_exu_i0_ap_predict_t; // @[quasar.scala 75:19]
  wire  exu_io_dec_exu_decode_exu_i0_ap_predict_nt; // @[quasar.scala 75:19]
  wire  exu_io_dec_exu_decode_exu_i0_ap_csr_write; // @[quasar.scala 75:19]
  wire  exu_io_dec_exu_decode_exu_i0_ap_csr_imm; // @[quasar.scala 75:19]
  wire  exu_io_dec_exu_decode_exu_dec_i0_predict_p_d_valid; // @[quasar.scala 75:19]
  wire  exu_io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_pc4; // @[quasar.scala 75:19]
  wire [1:0] exu_io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_hist; // @[quasar.scala 75:19]
  wire [11:0] exu_io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_toffset; // @[quasar.scala 75:19]
  wire  exu_io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_br_error; // @[quasar.scala 75:19]
  wire  exu_io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_br_start_error; // @[quasar.scala 75:19]
  wire [30:0] exu_io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_prett; // @[quasar.scala 75:19]
  wire  exu_io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_pcall; // @[quasar.scala 75:19]
  wire  exu_io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_pret; // @[quasar.scala 75:19]
  wire  exu_io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_pja; // @[quasar.scala 75:19]
  wire  exu_io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_way; // @[quasar.scala 75:19]
  wire [7:0] exu_io_dec_exu_decode_exu_i0_predict_fghr_d; // @[quasar.scala 75:19]
  wire [7:0] exu_io_dec_exu_decode_exu_i0_predict_index_d; // @[quasar.scala 75:19]
  wire [4:0] exu_io_dec_exu_decode_exu_i0_predict_btag_d; // @[quasar.scala 75:19]
  wire  exu_io_dec_exu_decode_exu_dec_i0_rs1_en_d; // @[quasar.scala 75:19]
  wire  exu_io_dec_exu_decode_exu_dec_i0_rs2_en_d; // @[quasar.scala 75:19]
  wire [31:0] exu_io_dec_exu_decode_exu_dec_i0_immed_d; // @[quasar.scala 75:19]
  wire [31:0] exu_io_dec_exu_decode_exu_dec_i0_rs1_bypass_data_d; // @[quasar.scala 75:19]
  wire [31:0] exu_io_dec_exu_decode_exu_dec_i0_rs2_bypass_data_d; // @[quasar.scala 75:19]
  wire  exu_io_dec_exu_decode_exu_dec_i0_select_pc_d; // @[quasar.scala 75:19]
  wire [1:0] exu_io_dec_exu_decode_exu_dec_i0_rs1_bypass_en_d; // @[quasar.scala 75:19]
  wire [1:0] exu_io_dec_exu_decode_exu_dec_i0_rs2_bypass_en_d; // @[quasar.scala 75:19]
  wire  exu_io_dec_exu_decode_exu_mul_p_valid; // @[quasar.scala 75:19]
  wire  exu_io_dec_exu_decode_exu_mul_p_bits_rs1_sign; // @[quasar.scala 75:19]
  wire  exu_io_dec_exu_decode_exu_mul_p_bits_rs2_sign; // @[quasar.scala 75:19]
  wire  exu_io_dec_exu_decode_exu_mul_p_bits_low; // @[quasar.scala 75:19]
  wire [30:0] exu_io_dec_exu_decode_exu_pred_correct_npc_x; // @[quasar.scala 75:19]
  wire  exu_io_dec_exu_decode_exu_dec_extint_stall; // @[quasar.scala 75:19]
  wire [31:0] exu_io_dec_exu_decode_exu_exu_i0_result_x; // @[quasar.scala 75:19]
  wire [31:0] exu_io_dec_exu_decode_exu_exu_csr_rs1_x; // @[quasar.scala 75:19]
  wire [29:0] exu_io_dec_exu_tlu_exu_dec_tlu_meihap; // @[quasar.scala 75:19]
  wire  exu_io_dec_exu_tlu_exu_dec_tlu_flush_lower_r; // @[quasar.scala 75:19]
  wire [30:0] exu_io_dec_exu_tlu_exu_dec_tlu_flush_path_r; // @[quasar.scala 75:19]
  wire [1:0] exu_io_dec_exu_tlu_exu_exu_i0_br_hist_r; // @[quasar.scala 75:19]
  wire  exu_io_dec_exu_tlu_exu_exu_i0_br_error_r; // @[quasar.scala 75:19]
  wire  exu_io_dec_exu_tlu_exu_exu_i0_br_start_error_r; // @[quasar.scala 75:19]
  wire [7:0] exu_io_dec_exu_tlu_exu_exu_i0_br_index_r; // @[quasar.scala 75:19]
  wire  exu_io_dec_exu_tlu_exu_exu_i0_br_valid_r; // @[quasar.scala 75:19]
  wire  exu_io_dec_exu_tlu_exu_exu_i0_br_mp_r; // @[quasar.scala 75:19]
  wire  exu_io_dec_exu_tlu_exu_exu_i0_br_middle_r; // @[quasar.scala 75:19]
  wire  exu_io_dec_exu_tlu_exu_exu_pmu_i0_br_misp; // @[quasar.scala 75:19]
  wire  exu_io_dec_exu_tlu_exu_exu_pmu_i0_br_ataken; // @[quasar.scala 75:19]
  wire  exu_io_dec_exu_tlu_exu_exu_pmu_i0_pc4; // @[quasar.scala 75:19]
  wire [30:0] exu_io_dec_exu_tlu_exu_exu_npc_r; // @[quasar.scala 75:19]
  wire [30:0] exu_io_dec_exu_ib_exu_dec_i0_pc_d; // @[quasar.scala 75:19]
  wire  exu_io_dec_exu_ib_exu_dec_debug_wdata_rs1_d; // @[quasar.scala 75:19]
  wire [31:0] exu_io_dec_exu_gpr_exu_gpr_i0_rs1_d; // @[quasar.scala 75:19]
  wire [31:0] exu_io_dec_exu_gpr_exu_gpr_i0_rs2_d; // @[quasar.scala 75:19]
  wire [7:0] exu_io_exu_bp_exu_i0_br_fghr_r; // @[quasar.scala 75:19]
  wire  exu_io_exu_bp_exu_i0_br_way_r; // @[quasar.scala 75:19]
  wire  exu_io_exu_bp_exu_mp_pkt_bits_misp; // @[quasar.scala 75:19]
  wire  exu_io_exu_bp_exu_mp_pkt_bits_ataken; // @[quasar.scala 75:19]
  wire  exu_io_exu_bp_exu_mp_pkt_bits_boffset; // @[quasar.scala 75:19]
  wire  exu_io_exu_bp_exu_mp_pkt_bits_pc4; // @[quasar.scala 75:19]
  wire [1:0] exu_io_exu_bp_exu_mp_pkt_bits_hist; // @[quasar.scala 75:19]
  wire [11:0] exu_io_exu_bp_exu_mp_pkt_bits_toffset; // @[quasar.scala 75:19]
  wire  exu_io_exu_bp_exu_mp_pkt_bits_pcall; // @[quasar.scala 75:19]
  wire  exu_io_exu_bp_exu_mp_pkt_bits_pret; // @[quasar.scala 75:19]
  wire  exu_io_exu_bp_exu_mp_pkt_bits_pja; // @[quasar.scala 75:19]
  wire  exu_io_exu_bp_exu_mp_pkt_bits_way; // @[quasar.scala 75:19]
  wire [7:0] exu_io_exu_bp_exu_mp_eghr; // @[quasar.scala 75:19]
  wire [7:0] exu_io_exu_bp_exu_mp_fghr; // @[quasar.scala 75:19]
  wire [7:0] exu_io_exu_bp_exu_mp_index; // @[quasar.scala 75:19]
  wire [4:0] exu_io_exu_bp_exu_mp_btag; // @[quasar.scala 75:19]
  wire  exu_io_exu_flush_final; // @[quasar.scala 75:19]
  wire [31:0] exu_io_exu_div_result; // @[quasar.scala 75:19]
  wire  exu_io_exu_div_wren; // @[quasar.scala 75:19]
  wire [31:0] exu_io_dbg_cmd_wrdata; // @[quasar.scala 75:19]
  wire [31:0] exu_io_lsu_exu_exu_lsu_rs1_d; // @[quasar.scala 75:19]
  wire [31:0] exu_io_lsu_exu_exu_lsu_rs2_d; // @[quasar.scala 75:19]
  wire [30:0] exu_io_exu_flush_path_final; // @[quasar.scala 75:19]
  wire  lsu_clock; // @[quasar.scala 76:19]
  wire  lsu_reset; // @[quasar.scala 76:19]
  wire  lsu_io_clk_override; // @[quasar.scala 76:19]
  wire  lsu_io_lsu_dma_dma_lsc_ctl_dma_dccm_req; // @[quasar.scala 76:19]
  wire [31:0] lsu_io_lsu_dma_dma_lsc_ctl_dma_mem_addr; // @[quasar.scala 76:19]
  wire [2:0] lsu_io_lsu_dma_dma_lsc_ctl_dma_mem_sz; // @[quasar.scala 76:19]
  wire  lsu_io_lsu_dma_dma_lsc_ctl_dma_mem_write; // @[quasar.scala 76:19]
  wire [63:0] lsu_io_lsu_dma_dma_lsc_ctl_dma_mem_wdata; // @[quasar.scala 76:19]
  wire [31:0] lsu_io_lsu_dma_dma_dccm_ctl_dma_mem_addr; // @[quasar.scala 76:19]
  wire [63:0] lsu_io_lsu_dma_dma_dccm_ctl_dma_mem_wdata; // @[quasar.scala 76:19]
  wire  lsu_io_lsu_dma_dma_dccm_ctl_dccm_dma_rvalid; // @[quasar.scala 76:19]
  wire  lsu_io_lsu_dma_dma_dccm_ctl_dccm_dma_ecc_error; // @[quasar.scala 76:19]
  wire [2:0] lsu_io_lsu_dma_dma_dccm_ctl_dccm_dma_rtag; // @[quasar.scala 76:19]
  wire [63:0] lsu_io_lsu_dma_dma_dccm_ctl_dccm_dma_rdata; // @[quasar.scala 76:19]
  wire  lsu_io_lsu_dma_dccm_ready; // @[quasar.scala 76:19]
  wire [2:0] lsu_io_lsu_dma_dma_mem_tag; // @[quasar.scala 76:19]
  wire  lsu_io_lsu_pic_picm_wren; // @[quasar.scala 76:19]
  wire  lsu_io_lsu_pic_picm_rden; // @[quasar.scala 76:19]
  wire  lsu_io_lsu_pic_picm_mken; // @[quasar.scala 76:19]
  wire [31:0] lsu_io_lsu_pic_picm_rdaddr; // @[quasar.scala 76:19]
  wire [31:0] lsu_io_lsu_pic_picm_wraddr; // @[quasar.scala 76:19]
  wire [31:0] lsu_io_lsu_pic_picm_wr_data; // @[quasar.scala 76:19]
  wire [31:0] lsu_io_lsu_pic_picm_rd_data; // @[quasar.scala 76:19]
  wire [31:0] lsu_io_lsu_exu_exu_lsu_rs1_d; // @[quasar.scala 76:19]
  wire [31:0] lsu_io_lsu_exu_exu_lsu_rs2_d; // @[quasar.scala 76:19]
  wire  lsu_io_lsu_dec_tlu_busbuff_lsu_pmu_bus_misaligned; // @[quasar.scala 76:19]
  wire  lsu_io_lsu_dec_tlu_busbuff_lsu_pmu_bus_error; // @[quasar.scala 76:19]
  wire  lsu_io_lsu_dec_tlu_busbuff_lsu_pmu_bus_busy; // @[quasar.scala 76:19]
  wire  lsu_io_lsu_dec_tlu_busbuff_dec_tlu_external_ldfwd_disable; // @[quasar.scala 76:19]
  wire  lsu_io_lsu_dec_tlu_busbuff_dec_tlu_wb_coalescing_disable; // @[quasar.scala 76:19]
  wire  lsu_io_lsu_dec_tlu_busbuff_dec_tlu_sideeffect_posted_disable; // @[quasar.scala 76:19]
  wire  lsu_io_lsu_dec_tlu_busbuff_lsu_imprecise_error_load_any; // @[quasar.scala 76:19]
  wire  lsu_io_lsu_dec_tlu_busbuff_lsu_imprecise_error_store_any; // @[quasar.scala 76:19]
  wire [31:0] lsu_io_lsu_dec_tlu_busbuff_lsu_imprecise_error_addr_any; // @[quasar.scala 76:19]
  wire  lsu_io_lsu_dec_dctl_busbuff_lsu_nonblock_load_valid_m; // @[quasar.scala 76:19]
  wire [1:0] lsu_io_lsu_dec_dctl_busbuff_lsu_nonblock_load_tag_m; // @[quasar.scala 76:19]
  wire  lsu_io_lsu_dec_dctl_busbuff_lsu_nonblock_load_inv_r; // @[quasar.scala 76:19]
  wire [1:0] lsu_io_lsu_dec_dctl_busbuff_lsu_nonblock_load_inv_tag_r; // @[quasar.scala 76:19]
  wire  lsu_io_lsu_dec_dctl_busbuff_lsu_nonblock_load_data_valid; // @[quasar.scala 76:19]
  wire  lsu_io_lsu_dec_dctl_busbuff_lsu_nonblock_load_data_error; // @[quasar.scala 76:19]
  wire [1:0] lsu_io_lsu_dec_dctl_busbuff_lsu_nonblock_load_data_tag; // @[quasar.scala 76:19]
  wire [31:0] lsu_io_lsu_dec_dctl_busbuff_lsu_nonblock_load_data; // @[quasar.scala 76:19]
  wire  lsu_io_dccm_wren; // @[quasar.scala 76:19]
  wire  lsu_io_dccm_rden; // @[quasar.scala 76:19]
  wire [15:0] lsu_io_dccm_wr_addr_lo; // @[quasar.scala 76:19]
  wire [15:0] lsu_io_dccm_wr_addr_hi; // @[quasar.scala 76:19]
  wire [15:0] lsu_io_dccm_rd_addr_lo; // @[quasar.scala 76:19]
  wire [15:0] lsu_io_dccm_rd_addr_hi; // @[quasar.scala 76:19]
  wire [38:0] lsu_io_dccm_wr_data_lo; // @[quasar.scala 76:19]
  wire [38:0] lsu_io_dccm_wr_data_hi; // @[quasar.scala 76:19]
  wire [38:0] lsu_io_dccm_rd_data_lo; // @[quasar.scala 76:19]
  wire [38:0] lsu_io_dccm_rd_data_hi; // @[quasar.scala 76:19]
  wire  lsu_io_lsu_tlu_lsu_pmu_load_external_m; // @[quasar.scala 76:19]
  wire  lsu_io_lsu_tlu_lsu_pmu_store_external_m; // @[quasar.scala 76:19]
  wire  lsu_io_axi_aw_valid; // @[quasar.scala 76:19]
  wire [31:0] lsu_io_axi_aw_bits_addr; // @[quasar.scala 76:19]
  wire [2:0] lsu_io_axi_aw_bits_size; // @[quasar.scala 76:19]
  wire  lsu_io_axi_w_valid; // @[quasar.scala 76:19]
  wire [7:0] lsu_io_axi_w_bits_strb; // @[quasar.scala 76:19]
  wire  lsu_io_axi_ar_valid; // @[quasar.scala 76:19]
  wire [31:0] lsu_io_axi_ar_bits_addr; // @[quasar.scala 76:19]
  wire [2:0] lsu_io_axi_ar_bits_size; // @[quasar.scala 76:19]
  wire  lsu_io_dec_tlu_flush_lower_r; // @[quasar.scala 76:19]
  wire  lsu_io_dec_tlu_i0_kill_writeb_r; // @[quasar.scala 76:19]
  wire  lsu_io_dec_tlu_force_halt; // @[quasar.scala 76:19]
  wire  lsu_io_dec_tlu_core_ecc_disable; // @[quasar.scala 76:19]
  wire [11:0] lsu_io_dec_lsu_offset_d; // @[quasar.scala 76:19]
  wire  lsu_io_lsu_p_valid; // @[quasar.scala 76:19]
  wire  lsu_io_lsu_p_bits_fast_int; // @[quasar.scala 76:19]
  wire  lsu_io_lsu_p_bits_by; // @[quasar.scala 76:19]
  wire  lsu_io_lsu_p_bits_half; // @[quasar.scala 76:19]
  wire  lsu_io_lsu_p_bits_word; // @[quasar.scala 76:19]
  wire  lsu_io_lsu_p_bits_load; // @[quasar.scala 76:19]
  wire  lsu_io_lsu_p_bits_store; // @[quasar.scala 76:19]
  wire  lsu_io_lsu_p_bits_unsign; // @[quasar.scala 76:19]
  wire  lsu_io_lsu_p_bits_store_data_bypass_d; // @[quasar.scala 76:19]
  wire  lsu_io_lsu_p_bits_load_ldst_bypass_d; // @[quasar.scala 76:19]
  wire  lsu_io_trigger_pkt_any_0_select; // @[quasar.scala 76:19]
  wire  lsu_io_trigger_pkt_any_0_match_pkt; // @[quasar.scala 76:19]
  wire  lsu_io_trigger_pkt_any_0_store; // @[quasar.scala 76:19]
  wire  lsu_io_trigger_pkt_any_0_load; // @[quasar.scala 76:19]
  wire [31:0] lsu_io_trigger_pkt_any_0_tdata2; // @[quasar.scala 76:19]
  wire  lsu_io_trigger_pkt_any_1_select; // @[quasar.scala 76:19]
  wire  lsu_io_trigger_pkt_any_1_match_pkt; // @[quasar.scala 76:19]
  wire  lsu_io_trigger_pkt_any_1_store; // @[quasar.scala 76:19]
  wire  lsu_io_trigger_pkt_any_1_load; // @[quasar.scala 76:19]
  wire [31:0] lsu_io_trigger_pkt_any_1_tdata2; // @[quasar.scala 76:19]
  wire  lsu_io_trigger_pkt_any_2_select; // @[quasar.scala 76:19]
  wire  lsu_io_trigger_pkt_any_2_match_pkt; // @[quasar.scala 76:19]
  wire  lsu_io_trigger_pkt_any_2_store; // @[quasar.scala 76:19]
  wire  lsu_io_trigger_pkt_any_2_load; // @[quasar.scala 76:19]
  wire [31:0] lsu_io_trigger_pkt_any_2_tdata2; // @[quasar.scala 76:19]
  wire  lsu_io_trigger_pkt_any_3_select; // @[quasar.scala 76:19]
  wire  lsu_io_trigger_pkt_any_3_match_pkt; // @[quasar.scala 76:19]
  wire  lsu_io_trigger_pkt_any_3_store; // @[quasar.scala 76:19]
  wire  lsu_io_trigger_pkt_any_3_load; // @[quasar.scala 76:19]
  wire [31:0] lsu_io_trigger_pkt_any_3_tdata2; // @[quasar.scala 76:19]
  wire  lsu_io_dec_lsu_valid_raw_d; // @[quasar.scala 76:19]
  wire [31:0] lsu_io_dec_tlu_mrac_ff; // @[quasar.scala 76:19]
  wire [31:0] lsu_io_lsu_result_m; // @[quasar.scala 76:19]
  wire [31:0] lsu_io_lsu_result_corr_r; // @[quasar.scala 76:19]
  wire  lsu_io_lsu_load_stall_any; // @[quasar.scala 76:19]
  wire  lsu_io_lsu_store_stall_any; // @[quasar.scala 76:19]
  wire  lsu_io_lsu_fastint_stall_any; // @[quasar.scala 76:19]
  wire  lsu_io_lsu_idle_any; // @[quasar.scala 76:19]
  wire [30:0] lsu_io_lsu_fir_addr; // @[quasar.scala 76:19]
  wire [1:0] lsu_io_lsu_fir_error; // @[quasar.scala 76:19]
  wire  lsu_io_lsu_single_ecc_error_incr; // @[quasar.scala 76:19]
  wire  lsu_io_lsu_error_pkt_r_valid; // @[quasar.scala 76:19]
  wire  lsu_io_lsu_error_pkt_r_bits_single_ecc_error; // @[quasar.scala 76:19]
  wire  lsu_io_lsu_error_pkt_r_bits_inst_type; // @[quasar.scala 76:19]
  wire  lsu_io_lsu_error_pkt_r_bits_exc_type; // @[quasar.scala 76:19]
  wire [3:0] lsu_io_lsu_error_pkt_r_bits_mscause; // @[quasar.scala 76:19]
  wire [31:0] lsu_io_lsu_error_pkt_r_bits_addr; // @[quasar.scala 76:19]
  wire  lsu_io_lsu_pmu_misaligned_m; // @[quasar.scala 76:19]
  wire [3:0] lsu_io_lsu_trigger_match_m; // @[quasar.scala 76:19]
  wire  lsu_io_lsu_bus_clk_en; // @[quasar.scala 76:19]
  wire  lsu_io_scan_mode; // @[quasar.scala 76:19]
  wire  lsu_io_free_clk; // @[quasar.scala 76:19]
  wire  pic_ctrl_inst_clock; // @[quasar.scala 77:29]
  wire  pic_ctrl_inst_reset; // @[quasar.scala 77:29]
  wire  pic_ctrl_inst_io_scan_mode; // @[quasar.scala 77:29]
  wire  pic_ctrl_inst_io_free_clk; // @[quasar.scala 77:29]
  wire  pic_ctrl_inst_io_active_clk; // @[quasar.scala 77:29]
  wire  pic_ctrl_inst_io_clk_override; // @[quasar.scala 77:29]
  wire [31:0] pic_ctrl_inst_io_extintsrc_req; // @[quasar.scala 77:29]
  wire  pic_ctrl_inst_io_lsu_pic_picm_wren; // @[quasar.scala 77:29]
  wire  pic_ctrl_inst_io_lsu_pic_picm_rden; // @[quasar.scala 77:29]
  wire  pic_ctrl_inst_io_lsu_pic_picm_mken; // @[quasar.scala 77:29]
  wire [31:0] pic_ctrl_inst_io_lsu_pic_picm_rdaddr; // @[quasar.scala 77:29]
  wire [31:0] pic_ctrl_inst_io_lsu_pic_picm_wraddr; // @[quasar.scala 77:29]
  wire [31:0] pic_ctrl_inst_io_lsu_pic_picm_wr_data; // @[quasar.scala 77:29]
  wire [31:0] pic_ctrl_inst_io_lsu_pic_picm_rd_data; // @[quasar.scala 77:29]
  wire [7:0] pic_ctrl_inst_io_dec_pic_pic_claimid; // @[quasar.scala 77:29]
  wire [3:0] pic_ctrl_inst_io_dec_pic_pic_pl; // @[quasar.scala 77:29]
  wire  pic_ctrl_inst_io_dec_pic_mhwakeup; // @[quasar.scala 77:29]
  wire [3:0] pic_ctrl_inst_io_dec_pic_dec_tlu_meicurpl; // @[quasar.scala 77:29]
  wire [3:0] pic_ctrl_inst_io_dec_pic_dec_tlu_meipt; // @[quasar.scala 77:29]
  wire  pic_ctrl_inst_io_dec_pic_mexintpend; // @[quasar.scala 77:29]
  wire  dma_ctrl_clock; // @[quasar.scala 78:24]
  wire  dma_ctrl_reset; // @[quasar.scala 78:24]
  wire  dma_ctrl_io_free_clk; // @[quasar.scala 78:24]
  wire  dma_ctrl_io_dma_bus_clk_en; // @[quasar.scala 78:24]
  wire  dma_ctrl_io_clk_override; // @[quasar.scala 78:24]
  wire  dma_ctrl_io_scan_mode; // @[quasar.scala 78:24]
  wire [1:0] dma_ctrl_io_dbg_cmd_size; // @[quasar.scala 78:24]
  wire [31:0] dma_ctrl_io_dma_dbg_rddata; // @[quasar.scala 78:24]
  wire  dma_ctrl_io_dma_dbg_cmd_done; // @[quasar.scala 78:24]
  wire  dma_ctrl_io_dma_dbg_cmd_fail; // @[quasar.scala 78:24]
  wire  dma_ctrl_io_dbg_dma_dbg_ib_dbg_cmd_valid; // @[quasar.scala 78:24]
  wire  dma_ctrl_io_dbg_dma_dbg_ib_dbg_cmd_write; // @[quasar.scala 78:24]
  wire [1:0] dma_ctrl_io_dbg_dma_dbg_ib_dbg_cmd_type; // @[quasar.scala 78:24]
  wire [31:0] dma_ctrl_io_dbg_dma_dbg_ib_dbg_cmd_addr; // @[quasar.scala 78:24]
  wire [31:0] dma_ctrl_io_dbg_dma_dbg_dctl_dbg_cmd_wrdata; // @[quasar.scala 78:24]
  wire  dma_ctrl_io_dbg_dma_io_dbg_dma_bubble; // @[quasar.scala 78:24]
  wire  dma_ctrl_io_dbg_dma_io_dma_dbg_ready; // @[quasar.scala 78:24]
  wire  dma_ctrl_io_dec_dma_dctl_dma_dma_dccm_stall_any; // @[quasar.scala 78:24]
  wire  dma_ctrl_io_dec_dma_tlu_dma_dma_pmu_dccm_read; // @[quasar.scala 78:24]
  wire  dma_ctrl_io_dec_dma_tlu_dma_dma_pmu_dccm_write; // @[quasar.scala 78:24]
  wire  dma_ctrl_io_dec_dma_tlu_dma_dma_pmu_any_read; // @[quasar.scala 78:24]
  wire  dma_ctrl_io_dec_dma_tlu_dma_dma_pmu_any_write; // @[quasar.scala 78:24]
  wire [2:0] dma_ctrl_io_dec_dma_tlu_dma_dec_tlu_dma_qos_prty; // @[quasar.scala 78:24]
  wire  dma_ctrl_io_dec_dma_tlu_dma_dma_dccm_stall_any; // @[quasar.scala 78:24]
  wire  dma_ctrl_io_dec_dma_tlu_dma_dma_iccm_stall_any; // @[quasar.scala 78:24]
  wire  dma_ctrl_io_iccm_dma_rvalid; // @[quasar.scala 78:24]
  wire  dma_ctrl_io_iccm_dma_ecc_error; // @[quasar.scala 78:24]
  wire [2:0] dma_ctrl_io_iccm_dma_rtag; // @[quasar.scala 78:24]
  wire [63:0] dma_ctrl_io_iccm_dma_rdata; // @[quasar.scala 78:24]
  wire  dma_ctrl_io_iccm_ready; // @[quasar.scala 78:24]
  wire  dma_ctrl_io_dma_axi_b_valid; // @[quasar.scala 78:24]
  wire  dma_ctrl_io_dma_axi_r_valid; // @[quasar.scala 78:24]
  wire [1:0] dma_ctrl_io_dma_axi_r_bits_resp; // @[quasar.scala 78:24]
  wire  dma_ctrl_io_lsu_dma_dma_lsc_ctl_dma_dccm_req; // @[quasar.scala 78:24]
  wire [31:0] dma_ctrl_io_lsu_dma_dma_lsc_ctl_dma_mem_addr; // @[quasar.scala 78:24]
  wire [2:0] dma_ctrl_io_lsu_dma_dma_lsc_ctl_dma_mem_sz; // @[quasar.scala 78:24]
  wire  dma_ctrl_io_lsu_dma_dma_lsc_ctl_dma_mem_write; // @[quasar.scala 78:24]
  wire [63:0] dma_ctrl_io_lsu_dma_dma_lsc_ctl_dma_mem_wdata; // @[quasar.scala 78:24]
  wire [31:0] dma_ctrl_io_lsu_dma_dma_dccm_ctl_dma_mem_addr; // @[quasar.scala 78:24]
  wire [63:0] dma_ctrl_io_lsu_dma_dma_dccm_ctl_dma_mem_wdata; // @[quasar.scala 78:24]
  wire  dma_ctrl_io_lsu_dma_dma_dccm_ctl_dccm_dma_rvalid; // @[quasar.scala 78:24]
  wire  dma_ctrl_io_lsu_dma_dma_dccm_ctl_dccm_dma_ecc_error; // @[quasar.scala 78:24]
  wire [2:0] dma_ctrl_io_lsu_dma_dma_dccm_ctl_dccm_dma_rtag; // @[quasar.scala 78:24]
  wire [63:0] dma_ctrl_io_lsu_dma_dma_dccm_ctl_dccm_dma_rdata; // @[quasar.scala 78:24]
  wire  dma_ctrl_io_lsu_dma_dccm_ready; // @[quasar.scala 78:24]
  wire [2:0] dma_ctrl_io_lsu_dma_dma_mem_tag; // @[quasar.scala 78:24]
  wire  dma_ctrl_io_ifu_dma_dma_ifc_dma_iccm_stall_any; // @[quasar.scala 78:24]
  wire  dma_ctrl_io_ifu_dma_dma_mem_ctl_dma_iccm_req; // @[quasar.scala 78:24]
  wire [31:0] dma_ctrl_io_ifu_dma_dma_mem_ctl_dma_mem_addr; // @[quasar.scala 78:24]
  wire [2:0] dma_ctrl_io_ifu_dma_dma_mem_ctl_dma_mem_sz; // @[quasar.scala 78:24]
  wire  dma_ctrl_io_ifu_dma_dma_mem_ctl_dma_mem_write; // @[quasar.scala 78:24]
  wire [63:0] dma_ctrl_io_ifu_dma_dma_mem_ctl_dma_mem_wdata; // @[quasar.scala 78:24]
  wire [2:0] dma_ctrl_io_ifu_dma_dma_mem_ctl_dma_mem_tag; // @[quasar.scala 78:24]
  wire  rvclkhdr_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_1_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_1_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_1_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_1_io_scan_mode; // @[lib.scala 343:22]
  wire  axi4_to_ahb_clock; // @[quasar.scala 242:32]
  wire  axi4_to_ahb_reset; // @[quasar.scala 242:32]
  wire  axi4_to_ahb_io_scan_mode; // @[quasar.scala 242:32]
  wire  axi4_to_ahb_io_bus_clk_en; // @[quasar.scala 242:32]
  wire  axi4_to_ahb_io_clk_override; // @[quasar.scala 242:32]
  wire  axi4_to_ahb_io_axi_aw_ready; // @[quasar.scala 242:32]
  wire  axi4_to_ahb_io_axi_aw_valid; // @[quasar.scala 242:32]
  wire [31:0] axi4_to_ahb_io_axi_aw_bits_addr; // @[quasar.scala 242:32]
  wire [2:0] axi4_to_ahb_io_axi_aw_bits_size; // @[quasar.scala 242:32]
  wire  axi4_to_ahb_io_axi_w_ready; // @[quasar.scala 242:32]
  wire  axi4_to_ahb_io_axi_w_valid; // @[quasar.scala 242:32]
  wire [7:0] axi4_to_ahb_io_axi_w_bits_strb; // @[quasar.scala 242:32]
  wire  axi4_to_ahb_io_axi_b_ready; // @[quasar.scala 242:32]
  wire  axi4_to_ahb_io_axi_ar_valid; // @[quasar.scala 242:32]
  wire [31:0] axi4_to_ahb_io_axi_ar_bits_addr; // @[quasar.scala 242:32]
  wire [2:0] axi4_to_ahb_io_axi_ar_bits_size; // @[quasar.scala 242:32]
  wire  axi4_to_ahb_io_ahb_in_hready; // @[quasar.scala 242:32]
  wire  axi4_to_ahb_io_ahb_in_hresp; // @[quasar.scala 242:32]
  wire [1:0] axi4_to_ahb_io_ahb_out_htrans; // @[quasar.scala 242:32]
  wire  axi4_to_ahb_io_ahb_out_hwrite; // @[quasar.scala 242:32]
  wire  axi4_to_ahb_1_clock; // @[quasar.scala 243:33]
  wire  axi4_to_ahb_1_reset; // @[quasar.scala 243:33]
  wire  axi4_to_ahb_1_io_scan_mode; // @[quasar.scala 243:33]
  wire  axi4_to_ahb_1_io_bus_clk_en; // @[quasar.scala 243:33]
  wire  axi4_to_ahb_1_io_clk_override; // @[quasar.scala 243:33]
  wire  axi4_to_ahb_1_io_axi_aw_ready; // @[quasar.scala 243:33]
  wire  axi4_to_ahb_1_io_axi_aw_valid; // @[quasar.scala 243:33]
  wire [31:0] axi4_to_ahb_1_io_axi_aw_bits_addr; // @[quasar.scala 243:33]
  wire [2:0] axi4_to_ahb_1_io_axi_aw_bits_size; // @[quasar.scala 243:33]
  wire  axi4_to_ahb_1_io_axi_w_ready; // @[quasar.scala 243:33]
  wire  axi4_to_ahb_1_io_axi_w_valid; // @[quasar.scala 243:33]
  wire [7:0] axi4_to_ahb_1_io_axi_w_bits_strb; // @[quasar.scala 243:33]
  wire  axi4_to_ahb_1_io_axi_b_ready; // @[quasar.scala 243:33]
  wire  axi4_to_ahb_1_io_axi_ar_valid; // @[quasar.scala 243:33]
  wire [31:0] axi4_to_ahb_1_io_axi_ar_bits_addr; // @[quasar.scala 243:33]
  wire [2:0] axi4_to_ahb_1_io_axi_ar_bits_size; // @[quasar.scala 243:33]
  wire  axi4_to_ahb_1_io_ahb_in_hready; // @[quasar.scala 243:33]
  wire  axi4_to_ahb_1_io_ahb_in_hresp; // @[quasar.scala 243:33]
  wire [1:0] axi4_to_ahb_1_io_ahb_out_htrans; // @[quasar.scala 243:33]
  wire  axi4_to_ahb_1_io_ahb_out_hwrite; // @[quasar.scala 243:33]
  wire  axi4_to_ahb_2_clock; // @[quasar.scala 244:33]
  wire  axi4_to_ahb_2_reset; // @[quasar.scala 244:33]
  wire  axi4_to_ahb_2_io_scan_mode; // @[quasar.scala 244:33]
  wire  axi4_to_ahb_2_io_bus_clk_en; // @[quasar.scala 244:33]
  wire  axi4_to_ahb_2_io_clk_override; // @[quasar.scala 244:33]
  wire  axi4_to_ahb_2_io_axi_aw_ready; // @[quasar.scala 244:33]
  wire  axi4_to_ahb_2_io_axi_aw_valid; // @[quasar.scala 244:33]
  wire [31:0] axi4_to_ahb_2_io_axi_aw_bits_addr; // @[quasar.scala 244:33]
  wire [2:0] axi4_to_ahb_2_io_axi_aw_bits_size; // @[quasar.scala 244:33]
  wire  axi4_to_ahb_2_io_axi_w_ready; // @[quasar.scala 244:33]
  wire  axi4_to_ahb_2_io_axi_w_valid; // @[quasar.scala 244:33]
  wire [7:0] axi4_to_ahb_2_io_axi_w_bits_strb; // @[quasar.scala 244:33]
  wire  axi4_to_ahb_2_io_axi_b_ready; // @[quasar.scala 244:33]
  wire  axi4_to_ahb_2_io_axi_ar_valid; // @[quasar.scala 244:33]
  wire [31:0] axi4_to_ahb_2_io_axi_ar_bits_addr; // @[quasar.scala 244:33]
  wire [2:0] axi4_to_ahb_2_io_axi_ar_bits_size; // @[quasar.scala 244:33]
  wire  axi4_to_ahb_2_io_ahb_in_hready; // @[quasar.scala 244:33]
  wire  axi4_to_ahb_2_io_ahb_in_hresp; // @[quasar.scala 244:33]
  wire [1:0] axi4_to_ahb_2_io_ahb_out_htrans; // @[quasar.scala 244:33]
  wire  axi4_to_ahb_2_io_ahb_out_hwrite; // @[quasar.scala 244:33]
  wire  ahb_to_axi4_clock; // @[quasar.scala 245:33]
  wire  ahb_to_axi4_reset; // @[quasar.scala 245:33]
  wire  ahb_to_axi4_io_scan_mode; // @[quasar.scala 245:33]
  wire  ahb_to_axi4_io_bus_clk_en; // @[quasar.scala 245:33]
  wire  ahb_to_axi4_io_axi_aw_valid; // @[quasar.scala 245:33]
  wire  ahb_to_axi4_io_axi_ar_valid; // @[quasar.scala 245:33]
  wire  ahb_to_axi4_io_axi_r_valid; // @[quasar.scala 245:33]
  wire [1:0] ahb_to_axi4_io_axi_r_bits_resp; // @[quasar.scala 245:33]
  wire  ahb_to_axi4_io_ahb_sig_in_hready; // @[quasar.scala 245:33]
  wire  ahb_to_axi4_io_ahb_sig_in_hresp; // @[quasar.scala 245:33]
  wire [31:0] ahb_to_axi4_io_ahb_sig_out_haddr; // @[quasar.scala 245:33]
  wire [2:0] ahb_to_axi4_io_ahb_sig_out_hsize; // @[quasar.scala 245:33]
  wire [1:0] ahb_to_axi4_io_ahb_sig_out_htrans; // @[quasar.scala 245:33]
  wire  ahb_to_axi4_io_ahb_sig_out_hwrite; // @[quasar.scala 245:33]
  wire  ahb_to_axi4_io_ahb_hsel; // @[quasar.scala 245:33]
  wire  ahb_to_axi4_io_ahb_hreadyin; // @[quasar.scala 245:33]
  wire  _T_1 = dbg_io_dbg_core_rst_l; // @[quasar.scala 80:67]
  wire  _T_2 = _T_1 | io_scan_mode; // @[quasar.scala 80:70]
  wire  _T_5 = ~dec_io_dec_pause_state_cg; // @[quasar.scala 81:23]
  wire  _T_6 = _T_5 | dec_io_dec_exu_tlu_exu_dec_tlu_flush_lower_r; // @[quasar.scala 81:50]
  ifu ifu ( // @[quasar.scala 72:19]
    .clock(ifu_clock),
    .reset(ifu_reset),
    .io_exu_flush_final(ifu_io_exu_flush_final),
    .io_exu_flush_path_final(ifu_io_exu_flush_path_final),
    .io_free_clk(ifu_io_free_clk),
    .io_active_clk(ifu_io_active_clk),
    .io_ifu_dec_dec_aln_aln_dec_dec_i0_decode_d(ifu_io_ifu_dec_dec_aln_aln_dec_dec_i0_decode_d),
    .io_ifu_dec_dec_aln_aln_dec_ifu_i0_cinst(ifu_io_ifu_dec_dec_aln_aln_dec_ifu_i0_cinst),
    .io_ifu_dec_dec_aln_aln_ib_ifu_i0_icaf(ifu_io_ifu_dec_dec_aln_aln_ib_ifu_i0_icaf),
    .io_ifu_dec_dec_aln_aln_ib_ifu_i0_icaf_type(ifu_io_ifu_dec_dec_aln_aln_ib_ifu_i0_icaf_type),
    .io_ifu_dec_dec_aln_aln_ib_ifu_i0_icaf_f1(ifu_io_ifu_dec_dec_aln_aln_ib_ifu_i0_icaf_f1),
    .io_ifu_dec_dec_aln_aln_ib_ifu_i0_dbecc(ifu_io_ifu_dec_dec_aln_aln_ib_ifu_i0_dbecc),
    .io_ifu_dec_dec_aln_aln_ib_ifu_i0_bp_index(ifu_io_ifu_dec_dec_aln_aln_ib_ifu_i0_bp_index),
    .io_ifu_dec_dec_aln_aln_ib_ifu_i0_bp_fghr(ifu_io_ifu_dec_dec_aln_aln_ib_ifu_i0_bp_fghr),
    .io_ifu_dec_dec_aln_aln_ib_ifu_i0_bp_btag(ifu_io_ifu_dec_dec_aln_aln_ib_ifu_i0_bp_btag),
    .io_ifu_dec_dec_aln_aln_ib_ifu_i0_valid(ifu_io_ifu_dec_dec_aln_aln_ib_ifu_i0_valid),
    .io_ifu_dec_dec_aln_aln_ib_ifu_i0_instr(ifu_io_ifu_dec_dec_aln_aln_ib_ifu_i0_instr),
    .io_ifu_dec_dec_aln_aln_ib_ifu_i0_pc(ifu_io_ifu_dec_dec_aln_aln_ib_ifu_i0_pc),
    .io_ifu_dec_dec_aln_aln_ib_ifu_i0_pc4(ifu_io_ifu_dec_dec_aln_aln_ib_ifu_i0_pc4),
    .io_ifu_dec_dec_aln_aln_ib_i0_brp_valid(ifu_io_ifu_dec_dec_aln_aln_ib_i0_brp_valid),
    .io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_toffset(ifu_io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_toffset),
    .io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_hist(ifu_io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_hist),
    .io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_br_error(ifu_io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_br_error),
    .io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_br_start_error(ifu_io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_br_start_error),
    .io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_prett(ifu_io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_prett),
    .io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_way(ifu_io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_way),
    .io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_ret(ifu_io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_ret),
    .io_ifu_dec_dec_aln_ifu_pmu_instr_aligned(ifu_io_ifu_dec_dec_aln_ifu_pmu_instr_aligned),
    .io_ifu_dec_dec_mem_ctrl_dec_tlu_flush_err_wb(ifu_io_ifu_dec_dec_mem_ctrl_dec_tlu_flush_err_wb),
    .io_ifu_dec_dec_mem_ctrl_dec_tlu_i0_commit_cmt(ifu_io_ifu_dec_dec_mem_ctrl_dec_tlu_i0_commit_cmt),
    .io_ifu_dec_dec_mem_ctrl_dec_tlu_force_halt(ifu_io_ifu_dec_dec_mem_ctrl_dec_tlu_force_halt),
    .io_ifu_dec_dec_mem_ctrl_dec_tlu_fence_i_wb(ifu_io_ifu_dec_dec_mem_ctrl_dec_tlu_fence_i_wb),
    .io_ifu_dec_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_wrdata(ifu_io_ifu_dec_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_wrdata),
    .io_ifu_dec_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_dicawics(ifu_io_ifu_dec_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_dicawics),
    .io_ifu_dec_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_rd_valid(ifu_io_ifu_dec_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_rd_valid),
    .io_ifu_dec_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_wr_valid(ifu_io_ifu_dec_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_wr_valid),
    .io_ifu_dec_dec_mem_ctrl_dec_tlu_core_ecc_disable(ifu_io_ifu_dec_dec_mem_ctrl_dec_tlu_core_ecc_disable),
    .io_ifu_dec_dec_mem_ctrl_ifu_pmu_ic_miss(ifu_io_ifu_dec_dec_mem_ctrl_ifu_pmu_ic_miss),
    .io_ifu_dec_dec_mem_ctrl_ifu_pmu_ic_hit(ifu_io_ifu_dec_dec_mem_ctrl_ifu_pmu_ic_hit),
    .io_ifu_dec_dec_mem_ctrl_ifu_pmu_bus_error(ifu_io_ifu_dec_dec_mem_ctrl_ifu_pmu_bus_error),
    .io_ifu_dec_dec_mem_ctrl_ifu_pmu_bus_busy(ifu_io_ifu_dec_dec_mem_ctrl_ifu_pmu_bus_busy),
    .io_ifu_dec_dec_mem_ctrl_ifu_ic_error_start(ifu_io_ifu_dec_dec_mem_ctrl_ifu_ic_error_start),
    .io_ifu_dec_dec_mem_ctrl_ifu_iccm_rd_ecc_single_err(ifu_io_ifu_dec_dec_mem_ctrl_ifu_iccm_rd_ecc_single_err),
    .io_ifu_dec_dec_mem_ctrl_ifu_ic_debug_rd_data(ifu_io_ifu_dec_dec_mem_ctrl_ifu_ic_debug_rd_data),
    .io_ifu_dec_dec_mem_ctrl_ifu_ic_debug_rd_data_valid(ifu_io_ifu_dec_dec_mem_ctrl_ifu_ic_debug_rd_data_valid),
    .io_ifu_dec_dec_mem_ctrl_ifu_miss_state_idle(ifu_io_ifu_dec_dec_mem_ctrl_ifu_miss_state_idle),
    .io_ifu_dec_dec_ifc_dec_tlu_flush_noredir_wb(ifu_io_ifu_dec_dec_ifc_dec_tlu_flush_noredir_wb),
    .io_ifu_dec_dec_ifc_dec_tlu_mrac_ff(ifu_io_ifu_dec_dec_ifc_dec_tlu_mrac_ff),
    .io_ifu_dec_dec_ifc_ifu_pmu_fetch_stall(ifu_io_ifu_dec_dec_ifc_ifu_pmu_fetch_stall),
    .io_ifu_dec_dec_bp_dec_tlu_br0_r_pkt_valid(ifu_io_ifu_dec_dec_bp_dec_tlu_br0_r_pkt_valid),
    .io_ifu_dec_dec_bp_dec_tlu_br0_r_pkt_bits_hist(ifu_io_ifu_dec_dec_bp_dec_tlu_br0_r_pkt_bits_hist),
    .io_ifu_dec_dec_bp_dec_tlu_br0_r_pkt_bits_br_error(ifu_io_ifu_dec_dec_bp_dec_tlu_br0_r_pkt_bits_br_error),
    .io_ifu_dec_dec_bp_dec_tlu_br0_r_pkt_bits_br_start_error(ifu_io_ifu_dec_dec_bp_dec_tlu_br0_r_pkt_bits_br_start_error),
    .io_ifu_dec_dec_bp_dec_tlu_br0_r_pkt_bits_way(ifu_io_ifu_dec_dec_bp_dec_tlu_br0_r_pkt_bits_way),
    .io_ifu_dec_dec_bp_dec_tlu_br0_r_pkt_bits_middle(ifu_io_ifu_dec_dec_bp_dec_tlu_br0_r_pkt_bits_middle),
    .io_ifu_dec_dec_bp_dec_tlu_flush_leak_one_wb(ifu_io_ifu_dec_dec_bp_dec_tlu_flush_leak_one_wb),
    .io_ifu_dec_dec_bp_dec_tlu_bpred_disable(ifu_io_ifu_dec_dec_bp_dec_tlu_bpred_disable),
    .io_exu_ifu_exu_bp_exu_i0_br_index_r(ifu_io_exu_ifu_exu_bp_exu_i0_br_index_r),
    .io_exu_ifu_exu_bp_exu_i0_br_fghr_r(ifu_io_exu_ifu_exu_bp_exu_i0_br_fghr_r),
    .io_exu_ifu_exu_bp_exu_mp_pkt_bits_misp(ifu_io_exu_ifu_exu_bp_exu_mp_pkt_bits_misp),
    .io_exu_ifu_exu_bp_exu_mp_pkt_bits_ataken(ifu_io_exu_ifu_exu_bp_exu_mp_pkt_bits_ataken),
    .io_exu_ifu_exu_bp_exu_mp_pkt_bits_boffset(ifu_io_exu_ifu_exu_bp_exu_mp_pkt_bits_boffset),
    .io_exu_ifu_exu_bp_exu_mp_pkt_bits_pc4(ifu_io_exu_ifu_exu_bp_exu_mp_pkt_bits_pc4),
    .io_exu_ifu_exu_bp_exu_mp_pkt_bits_hist(ifu_io_exu_ifu_exu_bp_exu_mp_pkt_bits_hist),
    .io_exu_ifu_exu_bp_exu_mp_pkt_bits_toffset(ifu_io_exu_ifu_exu_bp_exu_mp_pkt_bits_toffset),
    .io_exu_ifu_exu_bp_exu_mp_pkt_bits_pcall(ifu_io_exu_ifu_exu_bp_exu_mp_pkt_bits_pcall),
    .io_exu_ifu_exu_bp_exu_mp_pkt_bits_pret(ifu_io_exu_ifu_exu_bp_exu_mp_pkt_bits_pret),
    .io_exu_ifu_exu_bp_exu_mp_pkt_bits_pja(ifu_io_exu_ifu_exu_bp_exu_mp_pkt_bits_pja),
    .io_exu_ifu_exu_bp_exu_mp_pkt_bits_way(ifu_io_exu_ifu_exu_bp_exu_mp_pkt_bits_way),
    .io_exu_ifu_exu_bp_exu_mp_eghr(ifu_io_exu_ifu_exu_bp_exu_mp_eghr),
    .io_exu_ifu_exu_bp_exu_mp_fghr(ifu_io_exu_ifu_exu_bp_exu_mp_fghr),
    .io_exu_ifu_exu_bp_exu_mp_index(ifu_io_exu_ifu_exu_bp_exu_mp_index),
    .io_exu_ifu_exu_bp_exu_mp_btag(ifu_io_exu_ifu_exu_bp_exu_mp_btag),
    .io_iccm_rw_addr(ifu_io_iccm_rw_addr),
    .io_iccm_buf_correct_ecc(ifu_io_iccm_buf_correct_ecc),
    .io_iccm_correction_state(ifu_io_iccm_correction_state),
    .io_iccm_wren(ifu_io_iccm_wren),
    .io_iccm_rden(ifu_io_iccm_rden),
    .io_iccm_wr_size(ifu_io_iccm_wr_size),
    .io_iccm_wr_data(ifu_io_iccm_wr_data),
    .io_iccm_rd_data(ifu_io_iccm_rd_data),
    .io_iccm_rd_data_ecc(ifu_io_iccm_rd_data_ecc),
    .io_ic_rw_addr(ifu_io_ic_rw_addr),
    .io_ic_tag_valid(ifu_io_ic_tag_valid),
    .io_ic_rd_en(ifu_io_ic_rd_en),
    .io_ic_debug_wr_data(ifu_io_ic_debug_wr_data),
    .io_ic_debug_addr(ifu_io_ic_debug_addr),
    .io_ic_rd_data(ifu_io_ic_rd_data),
    .io_ic_debug_rd_data(ifu_io_ic_debug_rd_data),
    .io_ic_tag_debug_rd_data(ifu_io_ic_tag_debug_rd_data),
    .io_ic_eccerr(ifu_io_ic_eccerr),
    .io_ic_rd_hit(ifu_io_ic_rd_hit),
    .io_ic_tag_perr(ifu_io_ic_tag_perr),
    .io_ic_debug_rd_en(ifu_io_ic_debug_rd_en),
    .io_ic_debug_wr_en(ifu_io_ic_debug_wr_en),
    .io_ic_debug_tag_array(ifu_io_ic_debug_tag_array),
    .io_ic_debug_way(ifu_io_ic_debug_way),
    .io_ic_premux_data(ifu_io_ic_premux_data),
    .io_ic_sel_premux_data(ifu_io_ic_sel_premux_data),
    .io_ifu_ar_valid(ifu_io_ifu_ar_valid),
    .io_ifu_ar_bits_addr(ifu_io_ifu_ar_bits_addr),
    .io_ifu_bus_clk_en(ifu_io_ifu_bus_clk_en),
    .io_ifu_dma_dma_ifc_dma_iccm_stall_any(ifu_io_ifu_dma_dma_ifc_dma_iccm_stall_any),
    .io_ifu_dma_dma_mem_ctl_dma_iccm_req(ifu_io_ifu_dma_dma_mem_ctl_dma_iccm_req),
    .io_ifu_dma_dma_mem_ctl_dma_mem_addr(ifu_io_ifu_dma_dma_mem_ctl_dma_mem_addr),
    .io_ifu_dma_dma_mem_ctl_dma_mem_sz(ifu_io_ifu_dma_dma_mem_ctl_dma_mem_sz),
    .io_ifu_dma_dma_mem_ctl_dma_mem_write(ifu_io_ifu_dma_dma_mem_ctl_dma_mem_write),
    .io_ifu_dma_dma_mem_ctl_dma_mem_wdata(ifu_io_ifu_dma_dma_mem_ctl_dma_mem_wdata),
    .io_ifu_dma_dma_mem_ctl_dma_mem_tag(ifu_io_ifu_dma_dma_mem_ctl_dma_mem_tag),
    .io_iccm_dma_ecc_error(ifu_io_iccm_dma_ecc_error),
    .io_iccm_dma_rvalid(ifu_io_iccm_dma_rvalid),
    .io_iccm_dma_rdata(ifu_io_iccm_dma_rdata),
    .io_iccm_dma_rtag(ifu_io_iccm_dma_rtag),
    .io_iccm_ready(ifu_io_iccm_ready),
    .io_iccm_dma_sb_error(ifu_io_iccm_dma_sb_error),
    .io_dec_tlu_flush_lower_wb(ifu_io_dec_tlu_flush_lower_wb),
    .io_scan_mode(ifu_io_scan_mode)
  );
  dec dec ( // @[quasar.scala 73:19]
    .clock(dec_clock),
    .reset(dec_reset),
    .io_free_clk(dec_io_free_clk),
    .io_active_clk(dec_io_active_clk),
    .io_lsu_fastint_stall_any(dec_io_lsu_fastint_stall_any),
    .io_dec_pause_state_cg(dec_io_dec_pause_state_cg),
    .io_rst_vec(dec_io_rst_vec),
    .io_nmi_int(dec_io_nmi_int),
    .io_nmi_vec(dec_io_nmi_vec),
    .io_i_cpu_halt_req(dec_io_i_cpu_halt_req),
    .io_i_cpu_run_req(dec_io_i_cpu_run_req),
    .io_o_cpu_halt_status(dec_io_o_cpu_halt_status),
    .io_o_cpu_halt_ack(dec_io_o_cpu_halt_ack),
    .io_o_cpu_run_ack(dec_io_o_cpu_run_ack),
    .io_o_debug_mode_status(dec_io_o_debug_mode_status),
    .io_core_id(dec_io_core_id),
    .io_mpc_debug_halt_req(dec_io_mpc_debug_halt_req),
    .io_mpc_debug_run_req(dec_io_mpc_debug_run_req),
    .io_mpc_reset_run_req(dec_io_mpc_reset_run_req),
    .io_mpc_debug_halt_ack(dec_io_mpc_debug_halt_ack),
    .io_mpc_debug_run_ack(dec_io_mpc_debug_run_ack),
    .io_debug_brkpt_status(dec_io_debug_brkpt_status),
    .io_lsu_pmu_misaligned_m(dec_io_lsu_pmu_misaligned_m),
    .io_lsu_fir_addr(dec_io_lsu_fir_addr),
    .io_lsu_fir_error(dec_io_lsu_fir_error),
    .io_lsu_trigger_match_m(dec_io_lsu_trigger_match_m),
    .io_lsu_idle_any(dec_io_lsu_idle_any),
    .io_lsu_error_pkt_r_valid(dec_io_lsu_error_pkt_r_valid),
    .io_lsu_error_pkt_r_bits_single_ecc_error(dec_io_lsu_error_pkt_r_bits_single_ecc_error),
    .io_lsu_error_pkt_r_bits_inst_type(dec_io_lsu_error_pkt_r_bits_inst_type),
    .io_lsu_error_pkt_r_bits_exc_type(dec_io_lsu_error_pkt_r_bits_exc_type),
    .io_lsu_error_pkt_r_bits_mscause(dec_io_lsu_error_pkt_r_bits_mscause),
    .io_lsu_error_pkt_r_bits_addr(dec_io_lsu_error_pkt_r_bits_addr),
    .io_lsu_single_ecc_error_incr(dec_io_lsu_single_ecc_error_incr),
    .io_exu_div_result(dec_io_exu_div_result),
    .io_exu_div_wren(dec_io_exu_div_wren),
    .io_lsu_result_m(dec_io_lsu_result_m),
    .io_lsu_result_corr_r(dec_io_lsu_result_corr_r),
    .io_lsu_load_stall_any(dec_io_lsu_load_stall_any),
    .io_lsu_store_stall_any(dec_io_lsu_store_stall_any),
    .io_iccm_dma_sb_error(dec_io_iccm_dma_sb_error),
    .io_exu_flush_final(dec_io_exu_flush_final),
    .io_timer_int(dec_io_timer_int),
    .io_soft_int(dec_io_soft_int),
    .io_dbg_halt_req(dec_io_dbg_halt_req),
    .io_dbg_resume_req(dec_io_dbg_resume_req),
    .io_dec_tlu_dbg_halted(dec_io_dec_tlu_dbg_halted),
    .io_dec_tlu_debug_mode(dec_io_dec_tlu_debug_mode),
    .io_dec_tlu_resume_ack(dec_io_dec_tlu_resume_ack),
    .io_dec_tlu_mpc_halted_only(dec_io_dec_tlu_mpc_halted_only),
    .io_dec_dbg_rddata(dec_io_dec_dbg_rddata),
    .io_dec_dbg_cmd_done(dec_io_dec_dbg_cmd_done),
    .io_dec_dbg_cmd_fail(dec_io_dec_dbg_cmd_fail),
    .io_trigger_pkt_any_0_select(dec_io_trigger_pkt_any_0_select),
    .io_trigger_pkt_any_0_match_pkt(dec_io_trigger_pkt_any_0_match_pkt),
    .io_trigger_pkt_any_0_store(dec_io_trigger_pkt_any_0_store),
    .io_trigger_pkt_any_0_load(dec_io_trigger_pkt_any_0_load),
    .io_trigger_pkt_any_0_tdata2(dec_io_trigger_pkt_any_0_tdata2),
    .io_trigger_pkt_any_1_select(dec_io_trigger_pkt_any_1_select),
    .io_trigger_pkt_any_1_match_pkt(dec_io_trigger_pkt_any_1_match_pkt),
    .io_trigger_pkt_any_1_store(dec_io_trigger_pkt_any_1_store),
    .io_trigger_pkt_any_1_load(dec_io_trigger_pkt_any_1_load),
    .io_trigger_pkt_any_1_tdata2(dec_io_trigger_pkt_any_1_tdata2),
    .io_trigger_pkt_any_2_select(dec_io_trigger_pkt_any_2_select),
    .io_trigger_pkt_any_2_match_pkt(dec_io_trigger_pkt_any_2_match_pkt),
    .io_trigger_pkt_any_2_store(dec_io_trigger_pkt_any_2_store),
    .io_trigger_pkt_any_2_load(dec_io_trigger_pkt_any_2_load),
    .io_trigger_pkt_any_2_tdata2(dec_io_trigger_pkt_any_2_tdata2),
    .io_trigger_pkt_any_3_select(dec_io_trigger_pkt_any_3_select),
    .io_trigger_pkt_any_3_match_pkt(dec_io_trigger_pkt_any_3_match_pkt),
    .io_trigger_pkt_any_3_store(dec_io_trigger_pkt_any_3_store),
    .io_trigger_pkt_any_3_load(dec_io_trigger_pkt_any_3_load),
    .io_trigger_pkt_any_3_tdata2(dec_io_trigger_pkt_any_3_tdata2),
    .io_exu_i0_br_way_r(dec_io_exu_i0_br_way_r),
    .io_lsu_p_valid(dec_io_lsu_p_valid),
    .io_lsu_p_bits_fast_int(dec_io_lsu_p_bits_fast_int),
    .io_lsu_p_bits_by(dec_io_lsu_p_bits_by),
    .io_lsu_p_bits_half(dec_io_lsu_p_bits_half),
    .io_lsu_p_bits_word(dec_io_lsu_p_bits_word),
    .io_lsu_p_bits_load(dec_io_lsu_p_bits_load),
    .io_lsu_p_bits_store(dec_io_lsu_p_bits_store),
    .io_lsu_p_bits_unsign(dec_io_lsu_p_bits_unsign),
    .io_lsu_p_bits_store_data_bypass_d(dec_io_lsu_p_bits_store_data_bypass_d),
    .io_lsu_p_bits_load_ldst_bypass_d(dec_io_lsu_p_bits_load_ldst_bypass_d),
    .io_dec_lsu_offset_d(dec_io_dec_lsu_offset_d),
    .io_dec_tlu_i0_kill_writeb_r(dec_io_dec_tlu_i0_kill_writeb_r),
    .io_dec_tlu_perfcnt0(dec_io_dec_tlu_perfcnt0),
    .io_dec_tlu_perfcnt1(dec_io_dec_tlu_perfcnt1),
    .io_dec_tlu_perfcnt2(dec_io_dec_tlu_perfcnt2),
    .io_dec_tlu_perfcnt3(dec_io_dec_tlu_perfcnt3),
    .io_dec_lsu_valid_raw_d(dec_io_dec_lsu_valid_raw_d),
    .io_rv_trace_pkt_rv_i_valid_ip(dec_io_rv_trace_pkt_rv_i_valid_ip),
    .io_rv_trace_pkt_rv_i_insn_ip(dec_io_rv_trace_pkt_rv_i_insn_ip),
    .io_rv_trace_pkt_rv_i_address_ip(dec_io_rv_trace_pkt_rv_i_address_ip),
    .io_rv_trace_pkt_rv_i_exception_ip(dec_io_rv_trace_pkt_rv_i_exception_ip),
    .io_rv_trace_pkt_rv_i_ecause_ip(dec_io_rv_trace_pkt_rv_i_ecause_ip),
    .io_rv_trace_pkt_rv_i_interrupt_ip(dec_io_rv_trace_pkt_rv_i_interrupt_ip),
    .io_rv_trace_pkt_rv_i_tval_ip(dec_io_rv_trace_pkt_rv_i_tval_ip),
    .io_dec_tlu_misc_clk_override(dec_io_dec_tlu_misc_clk_override),
    .io_dec_tlu_lsu_clk_override(dec_io_dec_tlu_lsu_clk_override),
    .io_dec_tlu_bus_clk_override(dec_io_dec_tlu_bus_clk_override),
    .io_dec_tlu_pic_clk_override(dec_io_dec_tlu_pic_clk_override),
    .io_dec_tlu_dccm_clk_override(dec_io_dec_tlu_dccm_clk_override),
    .io_dec_tlu_icm_clk_override(dec_io_dec_tlu_icm_clk_override),
    .io_scan_mode(dec_io_scan_mode),
    .io_ifu_dec_dec_aln_aln_dec_dec_i0_decode_d(dec_io_ifu_dec_dec_aln_aln_dec_dec_i0_decode_d),
    .io_ifu_dec_dec_aln_aln_dec_ifu_i0_cinst(dec_io_ifu_dec_dec_aln_aln_dec_ifu_i0_cinst),
    .io_ifu_dec_dec_aln_aln_ib_ifu_i0_icaf(dec_io_ifu_dec_dec_aln_aln_ib_ifu_i0_icaf),
    .io_ifu_dec_dec_aln_aln_ib_ifu_i0_icaf_type(dec_io_ifu_dec_dec_aln_aln_ib_ifu_i0_icaf_type),
    .io_ifu_dec_dec_aln_aln_ib_ifu_i0_icaf_f1(dec_io_ifu_dec_dec_aln_aln_ib_ifu_i0_icaf_f1),
    .io_ifu_dec_dec_aln_aln_ib_ifu_i0_dbecc(dec_io_ifu_dec_dec_aln_aln_ib_ifu_i0_dbecc),
    .io_ifu_dec_dec_aln_aln_ib_ifu_i0_bp_index(dec_io_ifu_dec_dec_aln_aln_ib_ifu_i0_bp_index),
    .io_ifu_dec_dec_aln_aln_ib_ifu_i0_bp_fghr(dec_io_ifu_dec_dec_aln_aln_ib_ifu_i0_bp_fghr),
    .io_ifu_dec_dec_aln_aln_ib_ifu_i0_bp_btag(dec_io_ifu_dec_dec_aln_aln_ib_ifu_i0_bp_btag),
    .io_ifu_dec_dec_aln_aln_ib_ifu_i0_valid(dec_io_ifu_dec_dec_aln_aln_ib_ifu_i0_valid),
    .io_ifu_dec_dec_aln_aln_ib_ifu_i0_instr(dec_io_ifu_dec_dec_aln_aln_ib_ifu_i0_instr),
    .io_ifu_dec_dec_aln_aln_ib_ifu_i0_pc(dec_io_ifu_dec_dec_aln_aln_ib_ifu_i0_pc),
    .io_ifu_dec_dec_aln_aln_ib_ifu_i0_pc4(dec_io_ifu_dec_dec_aln_aln_ib_ifu_i0_pc4),
    .io_ifu_dec_dec_aln_aln_ib_i0_brp_valid(dec_io_ifu_dec_dec_aln_aln_ib_i0_brp_valid),
    .io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_toffset(dec_io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_toffset),
    .io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_hist(dec_io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_hist),
    .io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_br_error(dec_io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_br_error),
    .io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_br_start_error(dec_io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_br_start_error),
    .io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_prett(dec_io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_prett),
    .io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_way(dec_io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_way),
    .io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_ret(dec_io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_ret),
    .io_ifu_dec_dec_aln_ifu_pmu_instr_aligned(dec_io_ifu_dec_dec_aln_ifu_pmu_instr_aligned),
    .io_ifu_dec_dec_mem_ctrl_dec_tlu_flush_err_wb(dec_io_ifu_dec_dec_mem_ctrl_dec_tlu_flush_err_wb),
    .io_ifu_dec_dec_mem_ctrl_dec_tlu_i0_commit_cmt(dec_io_ifu_dec_dec_mem_ctrl_dec_tlu_i0_commit_cmt),
    .io_ifu_dec_dec_mem_ctrl_dec_tlu_force_halt(dec_io_ifu_dec_dec_mem_ctrl_dec_tlu_force_halt),
    .io_ifu_dec_dec_mem_ctrl_dec_tlu_fence_i_wb(dec_io_ifu_dec_dec_mem_ctrl_dec_tlu_fence_i_wb),
    .io_ifu_dec_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_wrdata(dec_io_ifu_dec_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_wrdata),
    .io_ifu_dec_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_dicawics(dec_io_ifu_dec_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_dicawics),
    .io_ifu_dec_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_rd_valid(dec_io_ifu_dec_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_rd_valid),
    .io_ifu_dec_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_wr_valid(dec_io_ifu_dec_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_wr_valid),
    .io_ifu_dec_dec_mem_ctrl_dec_tlu_core_ecc_disable(dec_io_ifu_dec_dec_mem_ctrl_dec_tlu_core_ecc_disable),
    .io_ifu_dec_dec_mem_ctrl_ifu_pmu_ic_miss(dec_io_ifu_dec_dec_mem_ctrl_ifu_pmu_ic_miss),
    .io_ifu_dec_dec_mem_ctrl_ifu_pmu_ic_hit(dec_io_ifu_dec_dec_mem_ctrl_ifu_pmu_ic_hit),
    .io_ifu_dec_dec_mem_ctrl_ifu_pmu_bus_error(dec_io_ifu_dec_dec_mem_ctrl_ifu_pmu_bus_error),
    .io_ifu_dec_dec_mem_ctrl_ifu_pmu_bus_busy(dec_io_ifu_dec_dec_mem_ctrl_ifu_pmu_bus_busy),
    .io_ifu_dec_dec_mem_ctrl_ifu_ic_error_start(dec_io_ifu_dec_dec_mem_ctrl_ifu_ic_error_start),
    .io_ifu_dec_dec_mem_ctrl_ifu_iccm_rd_ecc_single_err(dec_io_ifu_dec_dec_mem_ctrl_ifu_iccm_rd_ecc_single_err),
    .io_ifu_dec_dec_mem_ctrl_ifu_ic_debug_rd_data(dec_io_ifu_dec_dec_mem_ctrl_ifu_ic_debug_rd_data),
    .io_ifu_dec_dec_mem_ctrl_ifu_ic_debug_rd_data_valid(dec_io_ifu_dec_dec_mem_ctrl_ifu_ic_debug_rd_data_valid),
    .io_ifu_dec_dec_mem_ctrl_ifu_miss_state_idle(dec_io_ifu_dec_dec_mem_ctrl_ifu_miss_state_idle),
    .io_ifu_dec_dec_ifc_dec_tlu_flush_noredir_wb(dec_io_ifu_dec_dec_ifc_dec_tlu_flush_noredir_wb),
    .io_ifu_dec_dec_ifc_dec_tlu_mrac_ff(dec_io_ifu_dec_dec_ifc_dec_tlu_mrac_ff),
    .io_ifu_dec_dec_ifc_ifu_pmu_fetch_stall(dec_io_ifu_dec_dec_ifc_ifu_pmu_fetch_stall),
    .io_ifu_dec_dec_bp_dec_tlu_br0_r_pkt_valid(dec_io_ifu_dec_dec_bp_dec_tlu_br0_r_pkt_valid),
    .io_ifu_dec_dec_bp_dec_tlu_br0_r_pkt_bits_hist(dec_io_ifu_dec_dec_bp_dec_tlu_br0_r_pkt_bits_hist),
    .io_ifu_dec_dec_bp_dec_tlu_br0_r_pkt_bits_br_error(dec_io_ifu_dec_dec_bp_dec_tlu_br0_r_pkt_bits_br_error),
    .io_ifu_dec_dec_bp_dec_tlu_br0_r_pkt_bits_br_start_error(dec_io_ifu_dec_dec_bp_dec_tlu_br0_r_pkt_bits_br_start_error),
    .io_ifu_dec_dec_bp_dec_tlu_br0_r_pkt_bits_way(dec_io_ifu_dec_dec_bp_dec_tlu_br0_r_pkt_bits_way),
    .io_ifu_dec_dec_bp_dec_tlu_br0_r_pkt_bits_middle(dec_io_ifu_dec_dec_bp_dec_tlu_br0_r_pkt_bits_middle),
    .io_ifu_dec_dec_bp_dec_tlu_flush_leak_one_wb(dec_io_ifu_dec_dec_bp_dec_tlu_flush_leak_one_wb),
    .io_ifu_dec_dec_bp_dec_tlu_bpred_disable(dec_io_ifu_dec_dec_bp_dec_tlu_bpred_disable),
    .io_dec_exu_dec_alu_dec_i0_alu_decode_d(dec_io_dec_exu_dec_alu_dec_i0_alu_decode_d),
    .io_dec_exu_dec_alu_dec_csr_ren_d(dec_io_dec_exu_dec_alu_dec_csr_ren_d),
    .io_dec_exu_dec_alu_dec_i0_br_immed_d(dec_io_dec_exu_dec_alu_dec_i0_br_immed_d),
    .io_dec_exu_dec_alu_exu_i0_pc_x(dec_io_dec_exu_dec_alu_exu_i0_pc_x),
    .io_dec_exu_dec_div_div_p_valid(dec_io_dec_exu_dec_div_div_p_valid),
    .io_dec_exu_dec_div_div_p_bits_unsign(dec_io_dec_exu_dec_div_div_p_bits_unsign),
    .io_dec_exu_dec_div_div_p_bits_rem(dec_io_dec_exu_dec_div_div_p_bits_rem),
    .io_dec_exu_dec_div_dec_div_cancel(dec_io_dec_exu_dec_div_dec_div_cancel),
    .io_dec_exu_decode_exu_dec_data_en(dec_io_dec_exu_decode_exu_dec_data_en),
    .io_dec_exu_decode_exu_dec_ctl_en(dec_io_dec_exu_decode_exu_dec_ctl_en),
    .io_dec_exu_decode_exu_i0_ap_land(dec_io_dec_exu_decode_exu_i0_ap_land),
    .io_dec_exu_decode_exu_i0_ap_lor(dec_io_dec_exu_decode_exu_i0_ap_lor),
    .io_dec_exu_decode_exu_i0_ap_lxor(dec_io_dec_exu_decode_exu_i0_ap_lxor),
    .io_dec_exu_decode_exu_i0_ap_sll(dec_io_dec_exu_decode_exu_i0_ap_sll),
    .io_dec_exu_decode_exu_i0_ap_srl(dec_io_dec_exu_decode_exu_i0_ap_srl),
    .io_dec_exu_decode_exu_i0_ap_sra(dec_io_dec_exu_decode_exu_i0_ap_sra),
    .io_dec_exu_decode_exu_i0_ap_beq(dec_io_dec_exu_decode_exu_i0_ap_beq),
    .io_dec_exu_decode_exu_i0_ap_bne(dec_io_dec_exu_decode_exu_i0_ap_bne),
    .io_dec_exu_decode_exu_i0_ap_blt(dec_io_dec_exu_decode_exu_i0_ap_blt),
    .io_dec_exu_decode_exu_i0_ap_bge(dec_io_dec_exu_decode_exu_i0_ap_bge),
    .io_dec_exu_decode_exu_i0_ap_add(dec_io_dec_exu_decode_exu_i0_ap_add),
    .io_dec_exu_decode_exu_i0_ap_sub(dec_io_dec_exu_decode_exu_i0_ap_sub),
    .io_dec_exu_decode_exu_i0_ap_slt(dec_io_dec_exu_decode_exu_i0_ap_slt),
    .io_dec_exu_decode_exu_i0_ap_unsign(dec_io_dec_exu_decode_exu_i0_ap_unsign),
    .io_dec_exu_decode_exu_i0_ap_jal(dec_io_dec_exu_decode_exu_i0_ap_jal),
    .io_dec_exu_decode_exu_i0_ap_predict_t(dec_io_dec_exu_decode_exu_i0_ap_predict_t),
    .io_dec_exu_decode_exu_i0_ap_predict_nt(dec_io_dec_exu_decode_exu_i0_ap_predict_nt),
    .io_dec_exu_decode_exu_i0_ap_csr_write(dec_io_dec_exu_decode_exu_i0_ap_csr_write),
    .io_dec_exu_decode_exu_i0_ap_csr_imm(dec_io_dec_exu_decode_exu_i0_ap_csr_imm),
    .io_dec_exu_decode_exu_dec_i0_predict_p_d_valid(dec_io_dec_exu_decode_exu_dec_i0_predict_p_d_valid),
    .io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_pc4(dec_io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_pc4),
    .io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_hist(dec_io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_hist),
    .io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_toffset(dec_io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_toffset),
    .io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_br_error(dec_io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_br_error),
    .io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_br_start_error(dec_io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_br_start_error),
    .io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_prett(dec_io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_prett),
    .io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_pcall(dec_io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_pcall),
    .io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_pret(dec_io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_pret),
    .io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_pja(dec_io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_pja),
    .io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_way(dec_io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_way),
    .io_dec_exu_decode_exu_i0_predict_fghr_d(dec_io_dec_exu_decode_exu_i0_predict_fghr_d),
    .io_dec_exu_decode_exu_i0_predict_index_d(dec_io_dec_exu_decode_exu_i0_predict_index_d),
    .io_dec_exu_decode_exu_i0_predict_btag_d(dec_io_dec_exu_decode_exu_i0_predict_btag_d),
    .io_dec_exu_decode_exu_dec_i0_rs1_en_d(dec_io_dec_exu_decode_exu_dec_i0_rs1_en_d),
    .io_dec_exu_decode_exu_dec_i0_rs2_en_d(dec_io_dec_exu_decode_exu_dec_i0_rs2_en_d),
    .io_dec_exu_decode_exu_dec_i0_immed_d(dec_io_dec_exu_decode_exu_dec_i0_immed_d),
    .io_dec_exu_decode_exu_dec_i0_rs1_bypass_data_d(dec_io_dec_exu_decode_exu_dec_i0_rs1_bypass_data_d),
    .io_dec_exu_decode_exu_dec_i0_rs2_bypass_data_d(dec_io_dec_exu_decode_exu_dec_i0_rs2_bypass_data_d),
    .io_dec_exu_decode_exu_dec_i0_select_pc_d(dec_io_dec_exu_decode_exu_dec_i0_select_pc_d),
    .io_dec_exu_decode_exu_dec_i0_rs1_bypass_en_d(dec_io_dec_exu_decode_exu_dec_i0_rs1_bypass_en_d),
    .io_dec_exu_decode_exu_dec_i0_rs2_bypass_en_d(dec_io_dec_exu_decode_exu_dec_i0_rs2_bypass_en_d),
    .io_dec_exu_decode_exu_mul_p_valid(dec_io_dec_exu_decode_exu_mul_p_valid),
    .io_dec_exu_decode_exu_mul_p_bits_rs1_sign(dec_io_dec_exu_decode_exu_mul_p_bits_rs1_sign),
    .io_dec_exu_decode_exu_mul_p_bits_rs2_sign(dec_io_dec_exu_decode_exu_mul_p_bits_rs2_sign),
    .io_dec_exu_decode_exu_mul_p_bits_low(dec_io_dec_exu_decode_exu_mul_p_bits_low),
    .io_dec_exu_decode_exu_pred_correct_npc_x(dec_io_dec_exu_decode_exu_pred_correct_npc_x),
    .io_dec_exu_decode_exu_dec_extint_stall(dec_io_dec_exu_decode_exu_dec_extint_stall),
    .io_dec_exu_decode_exu_exu_i0_result_x(dec_io_dec_exu_decode_exu_exu_i0_result_x),
    .io_dec_exu_decode_exu_exu_csr_rs1_x(dec_io_dec_exu_decode_exu_exu_csr_rs1_x),
    .io_dec_exu_tlu_exu_dec_tlu_meihap(dec_io_dec_exu_tlu_exu_dec_tlu_meihap),
    .io_dec_exu_tlu_exu_dec_tlu_flush_lower_r(dec_io_dec_exu_tlu_exu_dec_tlu_flush_lower_r),
    .io_dec_exu_tlu_exu_dec_tlu_flush_path_r(dec_io_dec_exu_tlu_exu_dec_tlu_flush_path_r),
    .io_dec_exu_tlu_exu_exu_i0_br_hist_r(dec_io_dec_exu_tlu_exu_exu_i0_br_hist_r),
    .io_dec_exu_tlu_exu_exu_i0_br_error_r(dec_io_dec_exu_tlu_exu_exu_i0_br_error_r),
    .io_dec_exu_tlu_exu_exu_i0_br_start_error_r(dec_io_dec_exu_tlu_exu_exu_i0_br_start_error_r),
    .io_dec_exu_tlu_exu_exu_i0_br_valid_r(dec_io_dec_exu_tlu_exu_exu_i0_br_valid_r),
    .io_dec_exu_tlu_exu_exu_i0_br_mp_r(dec_io_dec_exu_tlu_exu_exu_i0_br_mp_r),
    .io_dec_exu_tlu_exu_exu_i0_br_middle_r(dec_io_dec_exu_tlu_exu_exu_i0_br_middle_r),
    .io_dec_exu_tlu_exu_exu_pmu_i0_br_misp(dec_io_dec_exu_tlu_exu_exu_pmu_i0_br_misp),
    .io_dec_exu_tlu_exu_exu_pmu_i0_br_ataken(dec_io_dec_exu_tlu_exu_exu_pmu_i0_br_ataken),
    .io_dec_exu_tlu_exu_exu_pmu_i0_pc4(dec_io_dec_exu_tlu_exu_exu_pmu_i0_pc4),
    .io_dec_exu_tlu_exu_exu_npc_r(dec_io_dec_exu_tlu_exu_exu_npc_r),
    .io_dec_exu_ib_exu_dec_i0_pc_d(dec_io_dec_exu_ib_exu_dec_i0_pc_d),
    .io_dec_exu_ib_exu_dec_debug_wdata_rs1_d(dec_io_dec_exu_ib_exu_dec_debug_wdata_rs1_d),
    .io_dec_exu_gpr_exu_gpr_i0_rs1_d(dec_io_dec_exu_gpr_exu_gpr_i0_rs1_d),
    .io_dec_exu_gpr_exu_gpr_i0_rs2_d(dec_io_dec_exu_gpr_exu_gpr_i0_rs2_d),
    .io_lsu_dec_tlu_busbuff_lsu_pmu_bus_misaligned(dec_io_lsu_dec_tlu_busbuff_lsu_pmu_bus_misaligned),
    .io_lsu_dec_tlu_busbuff_lsu_pmu_bus_error(dec_io_lsu_dec_tlu_busbuff_lsu_pmu_bus_error),
    .io_lsu_dec_tlu_busbuff_lsu_pmu_bus_busy(dec_io_lsu_dec_tlu_busbuff_lsu_pmu_bus_busy),
    .io_lsu_dec_tlu_busbuff_dec_tlu_external_ldfwd_disable(dec_io_lsu_dec_tlu_busbuff_dec_tlu_external_ldfwd_disable),
    .io_lsu_dec_tlu_busbuff_dec_tlu_wb_coalescing_disable(dec_io_lsu_dec_tlu_busbuff_dec_tlu_wb_coalescing_disable),
    .io_lsu_dec_tlu_busbuff_dec_tlu_sideeffect_posted_disable(dec_io_lsu_dec_tlu_busbuff_dec_tlu_sideeffect_posted_disable),
    .io_lsu_dec_tlu_busbuff_lsu_imprecise_error_load_any(dec_io_lsu_dec_tlu_busbuff_lsu_imprecise_error_load_any),
    .io_lsu_dec_tlu_busbuff_lsu_imprecise_error_store_any(dec_io_lsu_dec_tlu_busbuff_lsu_imprecise_error_store_any),
    .io_lsu_dec_tlu_busbuff_lsu_imprecise_error_addr_any(dec_io_lsu_dec_tlu_busbuff_lsu_imprecise_error_addr_any),
    .io_lsu_dec_dctl_busbuff_lsu_nonblock_load_valid_m(dec_io_lsu_dec_dctl_busbuff_lsu_nonblock_load_valid_m),
    .io_lsu_dec_dctl_busbuff_lsu_nonblock_load_tag_m(dec_io_lsu_dec_dctl_busbuff_lsu_nonblock_load_tag_m),
    .io_lsu_dec_dctl_busbuff_lsu_nonblock_load_inv_r(dec_io_lsu_dec_dctl_busbuff_lsu_nonblock_load_inv_r),
    .io_lsu_dec_dctl_busbuff_lsu_nonblock_load_inv_tag_r(dec_io_lsu_dec_dctl_busbuff_lsu_nonblock_load_inv_tag_r),
    .io_lsu_dec_dctl_busbuff_lsu_nonblock_load_data_valid(dec_io_lsu_dec_dctl_busbuff_lsu_nonblock_load_data_valid),
    .io_lsu_dec_dctl_busbuff_lsu_nonblock_load_data_error(dec_io_lsu_dec_dctl_busbuff_lsu_nonblock_load_data_error),
    .io_lsu_dec_dctl_busbuff_lsu_nonblock_load_data_tag(dec_io_lsu_dec_dctl_busbuff_lsu_nonblock_load_data_tag),
    .io_lsu_dec_dctl_busbuff_lsu_nonblock_load_data(dec_io_lsu_dec_dctl_busbuff_lsu_nonblock_load_data),
    .io_lsu_tlu_lsu_pmu_load_external_m(dec_io_lsu_tlu_lsu_pmu_load_external_m),
    .io_lsu_tlu_lsu_pmu_store_external_m(dec_io_lsu_tlu_lsu_pmu_store_external_m),
    .io_dec_dbg_dbg_ib_dbg_cmd_valid(dec_io_dec_dbg_dbg_ib_dbg_cmd_valid),
    .io_dec_dbg_dbg_ib_dbg_cmd_write(dec_io_dec_dbg_dbg_ib_dbg_cmd_write),
    .io_dec_dbg_dbg_ib_dbg_cmd_type(dec_io_dec_dbg_dbg_ib_dbg_cmd_type),
    .io_dec_dbg_dbg_ib_dbg_cmd_addr(dec_io_dec_dbg_dbg_ib_dbg_cmd_addr),
    .io_dec_dbg_dbg_dctl_dbg_cmd_wrdata(dec_io_dec_dbg_dbg_dctl_dbg_cmd_wrdata),
    .io_dec_dma_dctl_dma_dma_dccm_stall_any(dec_io_dec_dma_dctl_dma_dma_dccm_stall_any),
    .io_dec_dma_tlu_dma_dma_pmu_dccm_read(dec_io_dec_dma_tlu_dma_dma_pmu_dccm_read),
    .io_dec_dma_tlu_dma_dma_pmu_dccm_write(dec_io_dec_dma_tlu_dma_dma_pmu_dccm_write),
    .io_dec_dma_tlu_dma_dma_pmu_any_read(dec_io_dec_dma_tlu_dma_dma_pmu_any_read),
    .io_dec_dma_tlu_dma_dma_pmu_any_write(dec_io_dec_dma_tlu_dma_dma_pmu_any_write),
    .io_dec_dma_tlu_dma_dec_tlu_dma_qos_prty(dec_io_dec_dma_tlu_dma_dec_tlu_dma_qos_prty),
    .io_dec_dma_tlu_dma_dma_dccm_stall_any(dec_io_dec_dma_tlu_dma_dma_dccm_stall_any),
    .io_dec_dma_tlu_dma_dma_iccm_stall_any(dec_io_dec_dma_tlu_dma_dma_iccm_stall_any),
    .io_dec_pic_pic_claimid(dec_io_dec_pic_pic_claimid),
    .io_dec_pic_pic_pl(dec_io_dec_pic_pic_pl),
    .io_dec_pic_mhwakeup(dec_io_dec_pic_mhwakeup),
    .io_dec_pic_dec_tlu_meicurpl(dec_io_dec_pic_dec_tlu_meicurpl),
    .io_dec_pic_dec_tlu_meipt(dec_io_dec_pic_dec_tlu_meipt),
    .io_dec_pic_mexintpend(dec_io_dec_pic_mexintpend)
  );
  dbg dbg ( // @[quasar.scala 74:19]
    .clock(dbg_clock),
    .reset(dbg_reset),
    .io_dbg_cmd_size(dbg_io_dbg_cmd_size),
    .io_dbg_core_rst_l(dbg_io_dbg_core_rst_l),
    .io_core_dbg_rddata(dbg_io_core_dbg_rddata),
    .io_core_dbg_cmd_done(dbg_io_core_dbg_cmd_done),
    .io_core_dbg_cmd_fail(dbg_io_core_dbg_cmd_fail),
    .io_dbg_halt_req(dbg_io_dbg_halt_req),
    .io_dbg_resume_req(dbg_io_dbg_resume_req),
    .io_dec_tlu_debug_mode(dbg_io_dec_tlu_debug_mode),
    .io_dec_tlu_dbg_halted(dbg_io_dec_tlu_dbg_halted),
    .io_dec_tlu_mpc_halted_only(dbg_io_dec_tlu_mpc_halted_only),
    .io_dec_tlu_resume_ack(dbg_io_dec_tlu_resume_ack),
    .io_dmi_reg_en(dbg_io_dmi_reg_en),
    .io_dmi_reg_addr(dbg_io_dmi_reg_addr),
    .io_dmi_reg_wr_en(dbg_io_dmi_reg_wr_en),
    .io_dmi_reg_wdata(dbg_io_dmi_reg_wdata),
    .io_sb_axi_aw_valid(dbg_io_sb_axi_aw_valid),
    .io_sb_axi_aw_bits_addr(dbg_io_sb_axi_aw_bits_addr),
    .io_sb_axi_aw_bits_size(dbg_io_sb_axi_aw_bits_size),
    .io_sb_axi_w_valid(dbg_io_sb_axi_w_valid),
    .io_sb_axi_w_bits_strb(dbg_io_sb_axi_w_bits_strb),
    .io_sb_axi_ar_valid(dbg_io_sb_axi_ar_valid),
    .io_sb_axi_ar_bits_addr(dbg_io_sb_axi_ar_bits_addr),
    .io_sb_axi_ar_bits_size(dbg_io_sb_axi_ar_bits_size),
    .io_dbg_dec_dbg_ib_dbg_cmd_valid(dbg_io_dbg_dec_dbg_ib_dbg_cmd_valid),
    .io_dbg_dec_dbg_ib_dbg_cmd_write(dbg_io_dbg_dec_dbg_ib_dbg_cmd_write),
    .io_dbg_dec_dbg_ib_dbg_cmd_type(dbg_io_dbg_dec_dbg_ib_dbg_cmd_type),
    .io_dbg_dec_dbg_ib_dbg_cmd_addr(dbg_io_dbg_dec_dbg_ib_dbg_cmd_addr),
    .io_dbg_dec_dbg_dctl_dbg_cmd_wrdata(dbg_io_dbg_dec_dbg_dctl_dbg_cmd_wrdata),
    .io_dbg_dma_dbg_ib_dbg_cmd_valid(dbg_io_dbg_dma_dbg_ib_dbg_cmd_valid),
    .io_dbg_dma_dbg_ib_dbg_cmd_write(dbg_io_dbg_dma_dbg_ib_dbg_cmd_write),
    .io_dbg_dma_dbg_ib_dbg_cmd_type(dbg_io_dbg_dma_dbg_ib_dbg_cmd_type),
    .io_dbg_dma_dbg_ib_dbg_cmd_addr(dbg_io_dbg_dma_dbg_ib_dbg_cmd_addr),
    .io_dbg_dma_dbg_dctl_dbg_cmd_wrdata(dbg_io_dbg_dma_dbg_dctl_dbg_cmd_wrdata),
    .io_dbg_dma_io_dbg_dma_bubble(dbg_io_dbg_dma_io_dbg_dma_bubble),
    .io_dbg_dma_io_dma_dbg_ready(dbg_io_dbg_dma_io_dma_dbg_ready),
    .io_dbg_bus_clk_en(dbg_io_dbg_bus_clk_en),
    .io_dbg_rst_l(dbg_io_dbg_rst_l),
    .io_clk_override(dbg_io_clk_override),
    .io_scan_mode(dbg_io_scan_mode)
  );
  exu exu ( // @[quasar.scala 75:19]
    .clock(exu_clock),
    .reset(exu_reset),
    .io_scan_mode(exu_io_scan_mode),
    .io_dec_exu_dec_alu_dec_i0_alu_decode_d(exu_io_dec_exu_dec_alu_dec_i0_alu_decode_d),
    .io_dec_exu_dec_alu_dec_csr_ren_d(exu_io_dec_exu_dec_alu_dec_csr_ren_d),
    .io_dec_exu_dec_alu_dec_i0_br_immed_d(exu_io_dec_exu_dec_alu_dec_i0_br_immed_d),
    .io_dec_exu_dec_alu_exu_i0_pc_x(exu_io_dec_exu_dec_alu_exu_i0_pc_x),
    .io_dec_exu_dec_div_div_p_valid(exu_io_dec_exu_dec_div_div_p_valid),
    .io_dec_exu_dec_div_div_p_bits_unsign(exu_io_dec_exu_dec_div_div_p_bits_unsign),
    .io_dec_exu_dec_div_div_p_bits_rem(exu_io_dec_exu_dec_div_div_p_bits_rem),
    .io_dec_exu_dec_div_dec_div_cancel(exu_io_dec_exu_dec_div_dec_div_cancel),
    .io_dec_exu_decode_exu_dec_data_en(exu_io_dec_exu_decode_exu_dec_data_en),
    .io_dec_exu_decode_exu_dec_ctl_en(exu_io_dec_exu_decode_exu_dec_ctl_en),
    .io_dec_exu_decode_exu_i0_ap_land(exu_io_dec_exu_decode_exu_i0_ap_land),
    .io_dec_exu_decode_exu_i0_ap_lor(exu_io_dec_exu_decode_exu_i0_ap_lor),
    .io_dec_exu_decode_exu_i0_ap_lxor(exu_io_dec_exu_decode_exu_i0_ap_lxor),
    .io_dec_exu_decode_exu_i0_ap_sll(exu_io_dec_exu_decode_exu_i0_ap_sll),
    .io_dec_exu_decode_exu_i0_ap_srl(exu_io_dec_exu_decode_exu_i0_ap_srl),
    .io_dec_exu_decode_exu_i0_ap_sra(exu_io_dec_exu_decode_exu_i0_ap_sra),
    .io_dec_exu_decode_exu_i0_ap_beq(exu_io_dec_exu_decode_exu_i0_ap_beq),
    .io_dec_exu_decode_exu_i0_ap_bne(exu_io_dec_exu_decode_exu_i0_ap_bne),
    .io_dec_exu_decode_exu_i0_ap_blt(exu_io_dec_exu_decode_exu_i0_ap_blt),
    .io_dec_exu_decode_exu_i0_ap_bge(exu_io_dec_exu_decode_exu_i0_ap_bge),
    .io_dec_exu_decode_exu_i0_ap_add(exu_io_dec_exu_decode_exu_i0_ap_add),
    .io_dec_exu_decode_exu_i0_ap_sub(exu_io_dec_exu_decode_exu_i0_ap_sub),
    .io_dec_exu_decode_exu_i0_ap_slt(exu_io_dec_exu_decode_exu_i0_ap_slt),
    .io_dec_exu_decode_exu_i0_ap_unsign(exu_io_dec_exu_decode_exu_i0_ap_unsign),
    .io_dec_exu_decode_exu_i0_ap_jal(exu_io_dec_exu_decode_exu_i0_ap_jal),
    .io_dec_exu_decode_exu_i0_ap_predict_t(exu_io_dec_exu_decode_exu_i0_ap_predict_t),
    .io_dec_exu_decode_exu_i0_ap_predict_nt(exu_io_dec_exu_decode_exu_i0_ap_predict_nt),
    .io_dec_exu_decode_exu_i0_ap_csr_write(exu_io_dec_exu_decode_exu_i0_ap_csr_write),
    .io_dec_exu_decode_exu_i0_ap_csr_imm(exu_io_dec_exu_decode_exu_i0_ap_csr_imm),
    .io_dec_exu_decode_exu_dec_i0_predict_p_d_valid(exu_io_dec_exu_decode_exu_dec_i0_predict_p_d_valid),
    .io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_pc4(exu_io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_pc4),
    .io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_hist(exu_io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_hist),
    .io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_toffset(exu_io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_toffset),
    .io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_br_error(exu_io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_br_error),
    .io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_br_start_error(exu_io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_br_start_error),
    .io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_prett(exu_io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_prett),
    .io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_pcall(exu_io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_pcall),
    .io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_pret(exu_io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_pret),
    .io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_pja(exu_io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_pja),
    .io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_way(exu_io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_way),
    .io_dec_exu_decode_exu_i0_predict_fghr_d(exu_io_dec_exu_decode_exu_i0_predict_fghr_d),
    .io_dec_exu_decode_exu_i0_predict_index_d(exu_io_dec_exu_decode_exu_i0_predict_index_d),
    .io_dec_exu_decode_exu_i0_predict_btag_d(exu_io_dec_exu_decode_exu_i0_predict_btag_d),
    .io_dec_exu_decode_exu_dec_i0_rs1_en_d(exu_io_dec_exu_decode_exu_dec_i0_rs1_en_d),
    .io_dec_exu_decode_exu_dec_i0_rs2_en_d(exu_io_dec_exu_decode_exu_dec_i0_rs2_en_d),
    .io_dec_exu_decode_exu_dec_i0_immed_d(exu_io_dec_exu_decode_exu_dec_i0_immed_d),
    .io_dec_exu_decode_exu_dec_i0_rs1_bypass_data_d(exu_io_dec_exu_decode_exu_dec_i0_rs1_bypass_data_d),
    .io_dec_exu_decode_exu_dec_i0_rs2_bypass_data_d(exu_io_dec_exu_decode_exu_dec_i0_rs2_bypass_data_d),
    .io_dec_exu_decode_exu_dec_i0_select_pc_d(exu_io_dec_exu_decode_exu_dec_i0_select_pc_d),
    .io_dec_exu_decode_exu_dec_i0_rs1_bypass_en_d(exu_io_dec_exu_decode_exu_dec_i0_rs1_bypass_en_d),
    .io_dec_exu_decode_exu_dec_i0_rs2_bypass_en_d(exu_io_dec_exu_decode_exu_dec_i0_rs2_bypass_en_d),
    .io_dec_exu_decode_exu_mul_p_valid(exu_io_dec_exu_decode_exu_mul_p_valid),
    .io_dec_exu_decode_exu_mul_p_bits_rs1_sign(exu_io_dec_exu_decode_exu_mul_p_bits_rs1_sign),
    .io_dec_exu_decode_exu_mul_p_bits_rs2_sign(exu_io_dec_exu_decode_exu_mul_p_bits_rs2_sign),
    .io_dec_exu_decode_exu_mul_p_bits_low(exu_io_dec_exu_decode_exu_mul_p_bits_low),
    .io_dec_exu_decode_exu_pred_correct_npc_x(exu_io_dec_exu_decode_exu_pred_correct_npc_x),
    .io_dec_exu_decode_exu_dec_extint_stall(exu_io_dec_exu_decode_exu_dec_extint_stall),
    .io_dec_exu_decode_exu_exu_i0_result_x(exu_io_dec_exu_decode_exu_exu_i0_result_x),
    .io_dec_exu_decode_exu_exu_csr_rs1_x(exu_io_dec_exu_decode_exu_exu_csr_rs1_x),
    .io_dec_exu_tlu_exu_dec_tlu_meihap(exu_io_dec_exu_tlu_exu_dec_tlu_meihap),
    .io_dec_exu_tlu_exu_dec_tlu_flush_lower_r(exu_io_dec_exu_tlu_exu_dec_tlu_flush_lower_r),
    .io_dec_exu_tlu_exu_dec_tlu_flush_path_r(exu_io_dec_exu_tlu_exu_dec_tlu_flush_path_r),
    .io_dec_exu_tlu_exu_exu_i0_br_hist_r(exu_io_dec_exu_tlu_exu_exu_i0_br_hist_r),
    .io_dec_exu_tlu_exu_exu_i0_br_error_r(exu_io_dec_exu_tlu_exu_exu_i0_br_error_r),
    .io_dec_exu_tlu_exu_exu_i0_br_start_error_r(exu_io_dec_exu_tlu_exu_exu_i0_br_start_error_r),
    .io_dec_exu_tlu_exu_exu_i0_br_index_r(exu_io_dec_exu_tlu_exu_exu_i0_br_index_r),
    .io_dec_exu_tlu_exu_exu_i0_br_valid_r(exu_io_dec_exu_tlu_exu_exu_i0_br_valid_r),
    .io_dec_exu_tlu_exu_exu_i0_br_mp_r(exu_io_dec_exu_tlu_exu_exu_i0_br_mp_r),
    .io_dec_exu_tlu_exu_exu_i0_br_middle_r(exu_io_dec_exu_tlu_exu_exu_i0_br_middle_r),
    .io_dec_exu_tlu_exu_exu_pmu_i0_br_misp(exu_io_dec_exu_tlu_exu_exu_pmu_i0_br_misp),
    .io_dec_exu_tlu_exu_exu_pmu_i0_br_ataken(exu_io_dec_exu_tlu_exu_exu_pmu_i0_br_ataken),
    .io_dec_exu_tlu_exu_exu_pmu_i0_pc4(exu_io_dec_exu_tlu_exu_exu_pmu_i0_pc4),
    .io_dec_exu_tlu_exu_exu_npc_r(exu_io_dec_exu_tlu_exu_exu_npc_r),
    .io_dec_exu_ib_exu_dec_i0_pc_d(exu_io_dec_exu_ib_exu_dec_i0_pc_d),
    .io_dec_exu_ib_exu_dec_debug_wdata_rs1_d(exu_io_dec_exu_ib_exu_dec_debug_wdata_rs1_d),
    .io_dec_exu_gpr_exu_gpr_i0_rs1_d(exu_io_dec_exu_gpr_exu_gpr_i0_rs1_d),
    .io_dec_exu_gpr_exu_gpr_i0_rs2_d(exu_io_dec_exu_gpr_exu_gpr_i0_rs2_d),
    .io_exu_bp_exu_i0_br_fghr_r(exu_io_exu_bp_exu_i0_br_fghr_r),
    .io_exu_bp_exu_i0_br_way_r(exu_io_exu_bp_exu_i0_br_way_r),
    .io_exu_bp_exu_mp_pkt_bits_misp(exu_io_exu_bp_exu_mp_pkt_bits_misp),
    .io_exu_bp_exu_mp_pkt_bits_ataken(exu_io_exu_bp_exu_mp_pkt_bits_ataken),
    .io_exu_bp_exu_mp_pkt_bits_boffset(exu_io_exu_bp_exu_mp_pkt_bits_boffset),
    .io_exu_bp_exu_mp_pkt_bits_pc4(exu_io_exu_bp_exu_mp_pkt_bits_pc4),
    .io_exu_bp_exu_mp_pkt_bits_hist(exu_io_exu_bp_exu_mp_pkt_bits_hist),
    .io_exu_bp_exu_mp_pkt_bits_toffset(exu_io_exu_bp_exu_mp_pkt_bits_toffset),
    .io_exu_bp_exu_mp_pkt_bits_pcall(exu_io_exu_bp_exu_mp_pkt_bits_pcall),
    .io_exu_bp_exu_mp_pkt_bits_pret(exu_io_exu_bp_exu_mp_pkt_bits_pret),
    .io_exu_bp_exu_mp_pkt_bits_pja(exu_io_exu_bp_exu_mp_pkt_bits_pja),
    .io_exu_bp_exu_mp_pkt_bits_way(exu_io_exu_bp_exu_mp_pkt_bits_way),
    .io_exu_bp_exu_mp_eghr(exu_io_exu_bp_exu_mp_eghr),
    .io_exu_bp_exu_mp_fghr(exu_io_exu_bp_exu_mp_fghr),
    .io_exu_bp_exu_mp_index(exu_io_exu_bp_exu_mp_index),
    .io_exu_bp_exu_mp_btag(exu_io_exu_bp_exu_mp_btag),
    .io_exu_flush_final(exu_io_exu_flush_final),
    .io_exu_div_result(exu_io_exu_div_result),
    .io_exu_div_wren(exu_io_exu_div_wren),
    .io_dbg_cmd_wrdata(exu_io_dbg_cmd_wrdata),
    .io_lsu_exu_exu_lsu_rs1_d(exu_io_lsu_exu_exu_lsu_rs1_d),
    .io_lsu_exu_exu_lsu_rs2_d(exu_io_lsu_exu_exu_lsu_rs2_d),
    .io_exu_flush_path_final(exu_io_exu_flush_path_final)
  );
  lsu lsu ( // @[quasar.scala 76:19]
    .clock(lsu_clock),
    .reset(lsu_reset),
    .io_clk_override(lsu_io_clk_override),
    .io_lsu_dma_dma_lsc_ctl_dma_dccm_req(lsu_io_lsu_dma_dma_lsc_ctl_dma_dccm_req),
    .io_lsu_dma_dma_lsc_ctl_dma_mem_addr(lsu_io_lsu_dma_dma_lsc_ctl_dma_mem_addr),
    .io_lsu_dma_dma_lsc_ctl_dma_mem_sz(lsu_io_lsu_dma_dma_lsc_ctl_dma_mem_sz),
    .io_lsu_dma_dma_lsc_ctl_dma_mem_write(lsu_io_lsu_dma_dma_lsc_ctl_dma_mem_write),
    .io_lsu_dma_dma_lsc_ctl_dma_mem_wdata(lsu_io_lsu_dma_dma_lsc_ctl_dma_mem_wdata),
    .io_lsu_dma_dma_dccm_ctl_dma_mem_addr(lsu_io_lsu_dma_dma_dccm_ctl_dma_mem_addr),
    .io_lsu_dma_dma_dccm_ctl_dma_mem_wdata(lsu_io_lsu_dma_dma_dccm_ctl_dma_mem_wdata),
    .io_lsu_dma_dma_dccm_ctl_dccm_dma_rvalid(lsu_io_lsu_dma_dma_dccm_ctl_dccm_dma_rvalid),
    .io_lsu_dma_dma_dccm_ctl_dccm_dma_ecc_error(lsu_io_lsu_dma_dma_dccm_ctl_dccm_dma_ecc_error),
    .io_lsu_dma_dma_dccm_ctl_dccm_dma_rtag(lsu_io_lsu_dma_dma_dccm_ctl_dccm_dma_rtag),
    .io_lsu_dma_dma_dccm_ctl_dccm_dma_rdata(lsu_io_lsu_dma_dma_dccm_ctl_dccm_dma_rdata),
    .io_lsu_dma_dccm_ready(lsu_io_lsu_dma_dccm_ready),
    .io_lsu_dma_dma_mem_tag(lsu_io_lsu_dma_dma_mem_tag),
    .io_lsu_pic_picm_wren(lsu_io_lsu_pic_picm_wren),
    .io_lsu_pic_picm_rden(lsu_io_lsu_pic_picm_rden),
    .io_lsu_pic_picm_mken(lsu_io_lsu_pic_picm_mken),
    .io_lsu_pic_picm_rdaddr(lsu_io_lsu_pic_picm_rdaddr),
    .io_lsu_pic_picm_wraddr(lsu_io_lsu_pic_picm_wraddr),
    .io_lsu_pic_picm_wr_data(lsu_io_lsu_pic_picm_wr_data),
    .io_lsu_pic_picm_rd_data(lsu_io_lsu_pic_picm_rd_data),
    .io_lsu_exu_exu_lsu_rs1_d(lsu_io_lsu_exu_exu_lsu_rs1_d),
    .io_lsu_exu_exu_lsu_rs2_d(lsu_io_lsu_exu_exu_lsu_rs2_d),
    .io_lsu_dec_tlu_busbuff_lsu_pmu_bus_misaligned(lsu_io_lsu_dec_tlu_busbuff_lsu_pmu_bus_misaligned),
    .io_lsu_dec_tlu_busbuff_lsu_pmu_bus_error(lsu_io_lsu_dec_tlu_busbuff_lsu_pmu_bus_error),
    .io_lsu_dec_tlu_busbuff_lsu_pmu_bus_busy(lsu_io_lsu_dec_tlu_busbuff_lsu_pmu_bus_busy),
    .io_lsu_dec_tlu_busbuff_dec_tlu_external_ldfwd_disable(lsu_io_lsu_dec_tlu_busbuff_dec_tlu_external_ldfwd_disable),
    .io_lsu_dec_tlu_busbuff_dec_tlu_wb_coalescing_disable(lsu_io_lsu_dec_tlu_busbuff_dec_tlu_wb_coalescing_disable),
    .io_lsu_dec_tlu_busbuff_dec_tlu_sideeffect_posted_disable(lsu_io_lsu_dec_tlu_busbuff_dec_tlu_sideeffect_posted_disable),
    .io_lsu_dec_tlu_busbuff_lsu_imprecise_error_load_any(lsu_io_lsu_dec_tlu_busbuff_lsu_imprecise_error_load_any),
    .io_lsu_dec_tlu_busbuff_lsu_imprecise_error_store_any(lsu_io_lsu_dec_tlu_busbuff_lsu_imprecise_error_store_any),
    .io_lsu_dec_tlu_busbuff_lsu_imprecise_error_addr_any(lsu_io_lsu_dec_tlu_busbuff_lsu_imprecise_error_addr_any),
    .io_lsu_dec_dctl_busbuff_lsu_nonblock_load_valid_m(lsu_io_lsu_dec_dctl_busbuff_lsu_nonblock_load_valid_m),
    .io_lsu_dec_dctl_busbuff_lsu_nonblock_load_tag_m(lsu_io_lsu_dec_dctl_busbuff_lsu_nonblock_load_tag_m),
    .io_lsu_dec_dctl_busbuff_lsu_nonblock_load_inv_r(lsu_io_lsu_dec_dctl_busbuff_lsu_nonblock_load_inv_r),
    .io_lsu_dec_dctl_busbuff_lsu_nonblock_load_inv_tag_r(lsu_io_lsu_dec_dctl_busbuff_lsu_nonblock_load_inv_tag_r),
    .io_lsu_dec_dctl_busbuff_lsu_nonblock_load_data_valid(lsu_io_lsu_dec_dctl_busbuff_lsu_nonblock_load_data_valid),
    .io_lsu_dec_dctl_busbuff_lsu_nonblock_load_data_error(lsu_io_lsu_dec_dctl_busbuff_lsu_nonblock_load_data_error),
    .io_lsu_dec_dctl_busbuff_lsu_nonblock_load_data_tag(lsu_io_lsu_dec_dctl_busbuff_lsu_nonblock_load_data_tag),
    .io_lsu_dec_dctl_busbuff_lsu_nonblock_load_data(lsu_io_lsu_dec_dctl_busbuff_lsu_nonblock_load_data),
    .io_dccm_wren(lsu_io_dccm_wren),
    .io_dccm_rden(lsu_io_dccm_rden),
    .io_dccm_wr_addr_lo(lsu_io_dccm_wr_addr_lo),
    .io_dccm_wr_addr_hi(lsu_io_dccm_wr_addr_hi),
    .io_dccm_rd_addr_lo(lsu_io_dccm_rd_addr_lo),
    .io_dccm_rd_addr_hi(lsu_io_dccm_rd_addr_hi),
    .io_dccm_wr_data_lo(lsu_io_dccm_wr_data_lo),
    .io_dccm_wr_data_hi(lsu_io_dccm_wr_data_hi),
    .io_dccm_rd_data_lo(lsu_io_dccm_rd_data_lo),
    .io_dccm_rd_data_hi(lsu_io_dccm_rd_data_hi),
    .io_lsu_tlu_lsu_pmu_load_external_m(lsu_io_lsu_tlu_lsu_pmu_load_external_m),
    .io_lsu_tlu_lsu_pmu_store_external_m(lsu_io_lsu_tlu_lsu_pmu_store_external_m),
    .io_axi_aw_valid(lsu_io_axi_aw_valid),
    .io_axi_aw_bits_addr(lsu_io_axi_aw_bits_addr),
    .io_axi_aw_bits_size(lsu_io_axi_aw_bits_size),
    .io_axi_w_valid(lsu_io_axi_w_valid),
    .io_axi_w_bits_strb(lsu_io_axi_w_bits_strb),
    .io_axi_ar_valid(lsu_io_axi_ar_valid),
    .io_axi_ar_bits_addr(lsu_io_axi_ar_bits_addr),
    .io_axi_ar_bits_size(lsu_io_axi_ar_bits_size),
    .io_dec_tlu_flush_lower_r(lsu_io_dec_tlu_flush_lower_r),
    .io_dec_tlu_i0_kill_writeb_r(lsu_io_dec_tlu_i0_kill_writeb_r),
    .io_dec_tlu_force_halt(lsu_io_dec_tlu_force_halt),
    .io_dec_tlu_core_ecc_disable(lsu_io_dec_tlu_core_ecc_disable),
    .io_dec_lsu_offset_d(lsu_io_dec_lsu_offset_d),
    .io_lsu_p_valid(lsu_io_lsu_p_valid),
    .io_lsu_p_bits_fast_int(lsu_io_lsu_p_bits_fast_int),
    .io_lsu_p_bits_by(lsu_io_lsu_p_bits_by),
    .io_lsu_p_bits_half(lsu_io_lsu_p_bits_half),
    .io_lsu_p_bits_word(lsu_io_lsu_p_bits_word),
    .io_lsu_p_bits_load(lsu_io_lsu_p_bits_load),
    .io_lsu_p_bits_store(lsu_io_lsu_p_bits_store),
    .io_lsu_p_bits_unsign(lsu_io_lsu_p_bits_unsign),
    .io_lsu_p_bits_store_data_bypass_d(lsu_io_lsu_p_bits_store_data_bypass_d),
    .io_lsu_p_bits_load_ldst_bypass_d(lsu_io_lsu_p_bits_load_ldst_bypass_d),
    .io_trigger_pkt_any_0_select(lsu_io_trigger_pkt_any_0_select),
    .io_trigger_pkt_any_0_match_pkt(lsu_io_trigger_pkt_any_0_match_pkt),
    .io_trigger_pkt_any_0_store(lsu_io_trigger_pkt_any_0_store),
    .io_trigger_pkt_any_0_load(lsu_io_trigger_pkt_any_0_load),
    .io_trigger_pkt_any_0_tdata2(lsu_io_trigger_pkt_any_0_tdata2),
    .io_trigger_pkt_any_1_select(lsu_io_trigger_pkt_any_1_select),
    .io_trigger_pkt_any_1_match_pkt(lsu_io_trigger_pkt_any_1_match_pkt),
    .io_trigger_pkt_any_1_store(lsu_io_trigger_pkt_any_1_store),
    .io_trigger_pkt_any_1_load(lsu_io_trigger_pkt_any_1_load),
    .io_trigger_pkt_any_1_tdata2(lsu_io_trigger_pkt_any_1_tdata2),
    .io_trigger_pkt_any_2_select(lsu_io_trigger_pkt_any_2_select),
    .io_trigger_pkt_any_2_match_pkt(lsu_io_trigger_pkt_any_2_match_pkt),
    .io_trigger_pkt_any_2_store(lsu_io_trigger_pkt_any_2_store),
    .io_trigger_pkt_any_2_load(lsu_io_trigger_pkt_any_2_load),
    .io_trigger_pkt_any_2_tdata2(lsu_io_trigger_pkt_any_2_tdata2),
    .io_trigger_pkt_any_3_select(lsu_io_trigger_pkt_any_3_select),
    .io_trigger_pkt_any_3_match_pkt(lsu_io_trigger_pkt_any_3_match_pkt),
    .io_trigger_pkt_any_3_store(lsu_io_trigger_pkt_any_3_store),
    .io_trigger_pkt_any_3_load(lsu_io_trigger_pkt_any_3_load),
    .io_trigger_pkt_any_3_tdata2(lsu_io_trigger_pkt_any_3_tdata2),
    .io_dec_lsu_valid_raw_d(lsu_io_dec_lsu_valid_raw_d),
    .io_dec_tlu_mrac_ff(lsu_io_dec_tlu_mrac_ff),
    .io_lsu_result_m(lsu_io_lsu_result_m),
    .io_lsu_result_corr_r(lsu_io_lsu_result_corr_r),
    .io_lsu_load_stall_any(lsu_io_lsu_load_stall_any),
    .io_lsu_store_stall_any(lsu_io_lsu_store_stall_any),
    .io_lsu_fastint_stall_any(lsu_io_lsu_fastint_stall_any),
    .io_lsu_idle_any(lsu_io_lsu_idle_any),
    .io_lsu_fir_addr(lsu_io_lsu_fir_addr),
    .io_lsu_fir_error(lsu_io_lsu_fir_error),
    .io_lsu_single_ecc_error_incr(lsu_io_lsu_single_ecc_error_incr),
    .io_lsu_error_pkt_r_valid(lsu_io_lsu_error_pkt_r_valid),
    .io_lsu_error_pkt_r_bits_single_ecc_error(lsu_io_lsu_error_pkt_r_bits_single_ecc_error),
    .io_lsu_error_pkt_r_bits_inst_type(lsu_io_lsu_error_pkt_r_bits_inst_type),
    .io_lsu_error_pkt_r_bits_exc_type(lsu_io_lsu_error_pkt_r_bits_exc_type),
    .io_lsu_error_pkt_r_bits_mscause(lsu_io_lsu_error_pkt_r_bits_mscause),
    .io_lsu_error_pkt_r_bits_addr(lsu_io_lsu_error_pkt_r_bits_addr),
    .io_lsu_pmu_misaligned_m(lsu_io_lsu_pmu_misaligned_m),
    .io_lsu_trigger_match_m(lsu_io_lsu_trigger_match_m),
    .io_lsu_bus_clk_en(lsu_io_lsu_bus_clk_en),
    .io_scan_mode(lsu_io_scan_mode),
    .io_free_clk(lsu_io_free_clk)
  );
  pic_ctrl pic_ctrl_inst ( // @[quasar.scala 77:29]
    .clock(pic_ctrl_inst_clock),
    .reset(pic_ctrl_inst_reset),
    .io_scan_mode(pic_ctrl_inst_io_scan_mode),
    .io_free_clk(pic_ctrl_inst_io_free_clk),
    .io_active_clk(pic_ctrl_inst_io_active_clk),
    .io_clk_override(pic_ctrl_inst_io_clk_override),
    .io_extintsrc_req(pic_ctrl_inst_io_extintsrc_req),
    .io_lsu_pic_picm_wren(pic_ctrl_inst_io_lsu_pic_picm_wren),
    .io_lsu_pic_picm_rden(pic_ctrl_inst_io_lsu_pic_picm_rden),
    .io_lsu_pic_picm_mken(pic_ctrl_inst_io_lsu_pic_picm_mken),
    .io_lsu_pic_picm_rdaddr(pic_ctrl_inst_io_lsu_pic_picm_rdaddr),
    .io_lsu_pic_picm_wraddr(pic_ctrl_inst_io_lsu_pic_picm_wraddr),
    .io_lsu_pic_picm_wr_data(pic_ctrl_inst_io_lsu_pic_picm_wr_data),
    .io_lsu_pic_picm_rd_data(pic_ctrl_inst_io_lsu_pic_picm_rd_data),
    .io_dec_pic_pic_claimid(pic_ctrl_inst_io_dec_pic_pic_claimid),
    .io_dec_pic_pic_pl(pic_ctrl_inst_io_dec_pic_pic_pl),
    .io_dec_pic_mhwakeup(pic_ctrl_inst_io_dec_pic_mhwakeup),
    .io_dec_pic_dec_tlu_meicurpl(pic_ctrl_inst_io_dec_pic_dec_tlu_meicurpl),
    .io_dec_pic_dec_tlu_meipt(pic_ctrl_inst_io_dec_pic_dec_tlu_meipt),
    .io_dec_pic_mexintpend(pic_ctrl_inst_io_dec_pic_mexintpend)
  );
  dma_ctrl dma_ctrl ( // @[quasar.scala 78:24]
    .clock(dma_ctrl_clock),
    .reset(dma_ctrl_reset),
    .io_free_clk(dma_ctrl_io_free_clk),
    .io_dma_bus_clk_en(dma_ctrl_io_dma_bus_clk_en),
    .io_clk_override(dma_ctrl_io_clk_override),
    .io_scan_mode(dma_ctrl_io_scan_mode),
    .io_dbg_cmd_size(dma_ctrl_io_dbg_cmd_size),
    .io_dma_dbg_rddata(dma_ctrl_io_dma_dbg_rddata),
    .io_dma_dbg_cmd_done(dma_ctrl_io_dma_dbg_cmd_done),
    .io_dma_dbg_cmd_fail(dma_ctrl_io_dma_dbg_cmd_fail),
    .io_dbg_dma_dbg_ib_dbg_cmd_valid(dma_ctrl_io_dbg_dma_dbg_ib_dbg_cmd_valid),
    .io_dbg_dma_dbg_ib_dbg_cmd_write(dma_ctrl_io_dbg_dma_dbg_ib_dbg_cmd_write),
    .io_dbg_dma_dbg_ib_dbg_cmd_type(dma_ctrl_io_dbg_dma_dbg_ib_dbg_cmd_type),
    .io_dbg_dma_dbg_ib_dbg_cmd_addr(dma_ctrl_io_dbg_dma_dbg_ib_dbg_cmd_addr),
    .io_dbg_dma_dbg_dctl_dbg_cmd_wrdata(dma_ctrl_io_dbg_dma_dbg_dctl_dbg_cmd_wrdata),
    .io_dbg_dma_io_dbg_dma_bubble(dma_ctrl_io_dbg_dma_io_dbg_dma_bubble),
    .io_dbg_dma_io_dma_dbg_ready(dma_ctrl_io_dbg_dma_io_dma_dbg_ready),
    .io_dec_dma_dctl_dma_dma_dccm_stall_any(dma_ctrl_io_dec_dma_dctl_dma_dma_dccm_stall_any),
    .io_dec_dma_tlu_dma_dma_pmu_dccm_read(dma_ctrl_io_dec_dma_tlu_dma_dma_pmu_dccm_read),
    .io_dec_dma_tlu_dma_dma_pmu_dccm_write(dma_ctrl_io_dec_dma_tlu_dma_dma_pmu_dccm_write),
    .io_dec_dma_tlu_dma_dma_pmu_any_read(dma_ctrl_io_dec_dma_tlu_dma_dma_pmu_any_read),
    .io_dec_dma_tlu_dma_dma_pmu_any_write(dma_ctrl_io_dec_dma_tlu_dma_dma_pmu_any_write),
    .io_dec_dma_tlu_dma_dec_tlu_dma_qos_prty(dma_ctrl_io_dec_dma_tlu_dma_dec_tlu_dma_qos_prty),
    .io_dec_dma_tlu_dma_dma_dccm_stall_any(dma_ctrl_io_dec_dma_tlu_dma_dma_dccm_stall_any),
    .io_dec_dma_tlu_dma_dma_iccm_stall_any(dma_ctrl_io_dec_dma_tlu_dma_dma_iccm_stall_any),
    .io_iccm_dma_rvalid(dma_ctrl_io_iccm_dma_rvalid),
    .io_iccm_dma_ecc_error(dma_ctrl_io_iccm_dma_ecc_error),
    .io_iccm_dma_rtag(dma_ctrl_io_iccm_dma_rtag),
    .io_iccm_dma_rdata(dma_ctrl_io_iccm_dma_rdata),
    .io_iccm_ready(dma_ctrl_io_iccm_ready),
    .io_dma_axi_b_valid(dma_ctrl_io_dma_axi_b_valid),
    .io_dma_axi_r_valid(dma_ctrl_io_dma_axi_r_valid),
    .io_dma_axi_r_bits_resp(dma_ctrl_io_dma_axi_r_bits_resp),
    .io_lsu_dma_dma_lsc_ctl_dma_dccm_req(dma_ctrl_io_lsu_dma_dma_lsc_ctl_dma_dccm_req),
    .io_lsu_dma_dma_lsc_ctl_dma_mem_addr(dma_ctrl_io_lsu_dma_dma_lsc_ctl_dma_mem_addr),
    .io_lsu_dma_dma_lsc_ctl_dma_mem_sz(dma_ctrl_io_lsu_dma_dma_lsc_ctl_dma_mem_sz),
    .io_lsu_dma_dma_lsc_ctl_dma_mem_write(dma_ctrl_io_lsu_dma_dma_lsc_ctl_dma_mem_write),
    .io_lsu_dma_dma_lsc_ctl_dma_mem_wdata(dma_ctrl_io_lsu_dma_dma_lsc_ctl_dma_mem_wdata),
    .io_lsu_dma_dma_dccm_ctl_dma_mem_addr(dma_ctrl_io_lsu_dma_dma_dccm_ctl_dma_mem_addr),
    .io_lsu_dma_dma_dccm_ctl_dma_mem_wdata(dma_ctrl_io_lsu_dma_dma_dccm_ctl_dma_mem_wdata),
    .io_lsu_dma_dma_dccm_ctl_dccm_dma_rvalid(dma_ctrl_io_lsu_dma_dma_dccm_ctl_dccm_dma_rvalid),
    .io_lsu_dma_dma_dccm_ctl_dccm_dma_ecc_error(dma_ctrl_io_lsu_dma_dma_dccm_ctl_dccm_dma_ecc_error),
    .io_lsu_dma_dma_dccm_ctl_dccm_dma_rtag(dma_ctrl_io_lsu_dma_dma_dccm_ctl_dccm_dma_rtag),
    .io_lsu_dma_dma_dccm_ctl_dccm_dma_rdata(dma_ctrl_io_lsu_dma_dma_dccm_ctl_dccm_dma_rdata),
    .io_lsu_dma_dccm_ready(dma_ctrl_io_lsu_dma_dccm_ready),
    .io_lsu_dma_dma_mem_tag(dma_ctrl_io_lsu_dma_dma_mem_tag),
    .io_ifu_dma_dma_ifc_dma_iccm_stall_any(dma_ctrl_io_ifu_dma_dma_ifc_dma_iccm_stall_any),
    .io_ifu_dma_dma_mem_ctl_dma_iccm_req(dma_ctrl_io_ifu_dma_dma_mem_ctl_dma_iccm_req),
    .io_ifu_dma_dma_mem_ctl_dma_mem_addr(dma_ctrl_io_ifu_dma_dma_mem_ctl_dma_mem_addr),
    .io_ifu_dma_dma_mem_ctl_dma_mem_sz(dma_ctrl_io_ifu_dma_dma_mem_ctl_dma_mem_sz),
    .io_ifu_dma_dma_mem_ctl_dma_mem_write(dma_ctrl_io_ifu_dma_dma_mem_ctl_dma_mem_write),
    .io_ifu_dma_dma_mem_ctl_dma_mem_wdata(dma_ctrl_io_ifu_dma_dma_mem_ctl_dma_mem_wdata),
    .io_ifu_dma_dma_mem_ctl_dma_mem_tag(dma_ctrl_io_ifu_dma_dma_mem_ctl_dma_mem_tag)
  );
  rvclkhdr rvclkhdr ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_io_l1clk),
    .io_clk(rvclkhdr_io_clk),
    .io_en(rvclkhdr_io_en),
    .io_scan_mode(rvclkhdr_io_scan_mode)
  );
  rvclkhdr rvclkhdr_1 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_1_io_l1clk),
    .io_clk(rvclkhdr_1_io_clk),
    .io_en(rvclkhdr_1_io_en),
    .io_scan_mode(rvclkhdr_1_io_scan_mode)
  );
  axi4_to_ahb axi4_to_ahb ( // @[quasar.scala 242:32]
    .clock(axi4_to_ahb_clock),
    .reset(axi4_to_ahb_reset),
    .io_scan_mode(axi4_to_ahb_io_scan_mode),
    .io_bus_clk_en(axi4_to_ahb_io_bus_clk_en),
    .io_clk_override(axi4_to_ahb_io_clk_override),
    .io_axi_aw_ready(axi4_to_ahb_io_axi_aw_ready),
    .io_axi_aw_valid(axi4_to_ahb_io_axi_aw_valid),
    .io_axi_aw_bits_addr(axi4_to_ahb_io_axi_aw_bits_addr),
    .io_axi_aw_bits_size(axi4_to_ahb_io_axi_aw_bits_size),
    .io_axi_w_ready(axi4_to_ahb_io_axi_w_ready),
    .io_axi_w_valid(axi4_to_ahb_io_axi_w_valid),
    .io_axi_w_bits_strb(axi4_to_ahb_io_axi_w_bits_strb),
    .io_axi_b_ready(axi4_to_ahb_io_axi_b_ready),
    .io_axi_ar_valid(axi4_to_ahb_io_axi_ar_valid),
    .io_axi_ar_bits_addr(axi4_to_ahb_io_axi_ar_bits_addr),
    .io_axi_ar_bits_size(axi4_to_ahb_io_axi_ar_bits_size),
    .io_ahb_in_hready(axi4_to_ahb_io_ahb_in_hready),
    .io_ahb_in_hresp(axi4_to_ahb_io_ahb_in_hresp),
    .io_ahb_out_htrans(axi4_to_ahb_io_ahb_out_htrans),
    .io_ahb_out_hwrite(axi4_to_ahb_io_ahb_out_hwrite)
  );
  axi4_to_ahb axi4_to_ahb_1 ( // @[quasar.scala 243:33]
    .clock(axi4_to_ahb_1_clock),
    .reset(axi4_to_ahb_1_reset),
    .io_scan_mode(axi4_to_ahb_1_io_scan_mode),
    .io_bus_clk_en(axi4_to_ahb_1_io_bus_clk_en),
    .io_clk_override(axi4_to_ahb_1_io_clk_override),
    .io_axi_aw_ready(axi4_to_ahb_1_io_axi_aw_ready),
    .io_axi_aw_valid(axi4_to_ahb_1_io_axi_aw_valid),
    .io_axi_aw_bits_addr(axi4_to_ahb_1_io_axi_aw_bits_addr),
    .io_axi_aw_bits_size(axi4_to_ahb_1_io_axi_aw_bits_size),
    .io_axi_w_ready(axi4_to_ahb_1_io_axi_w_ready),
    .io_axi_w_valid(axi4_to_ahb_1_io_axi_w_valid),
    .io_axi_w_bits_strb(axi4_to_ahb_1_io_axi_w_bits_strb),
    .io_axi_b_ready(axi4_to_ahb_1_io_axi_b_ready),
    .io_axi_ar_valid(axi4_to_ahb_1_io_axi_ar_valid),
    .io_axi_ar_bits_addr(axi4_to_ahb_1_io_axi_ar_bits_addr),
    .io_axi_ar_bits_size(axi4_to_ahb_1_io_axi_ar_bits_size),
    .io_ahb_in_hready(axi4_to_ahb_1_io_ahb_in_hready),
    .io_ahb_in_hresp(axi4_to_ahb_1_io_ahb_in_hresp),
    .io_ahb_out_htrans(axi4_to_ahb_1_io_ahb_out_htrans),
    .io_ahb_out_hwrite(axi4_to_ahb_1_io_ahb_out_hwrite)
  );
  axi4_to_ahb axi4_to_ahb_2 ( // @[quasar.scala 244:33]
    .clock(axi4_to_ahb_2_clock),
    .reset(axi4_to_ahb_2_reset),
    .io_scan_mode(axi4_to_ahb_2_io_scan_mode),
    .io_bus_clk_en(axi4_to_ahb_2_io_bus_clk_en),
    .io_clk_override(axi4_to_ahb_2_io_clk_override),
    .io_axi_aw_ready(axi4_to_ahb_2_io_axi_aw_ready),
    .io_axi_aw_valid(axi4_to_ahb_2_io_axi_aw_valid),
    .io_axi_aw_bits_addr(axi4_to_ahb_2_io_axi_aw_bits_addr),
    .io_axi_aw_bits_size(axi4_to_ahb_2_io_axi_aw_bits_size),
    .io_axi_w_ready(axi4_to_ahb_2_io_axi_w_ready),
    .io_axi_w_valid(axi4_to_ahb_2_io_axi_w_valid),
    .io_axi_w_bits_strb(axi4_to_ahb_2_io_axi_w_bits_strb),
    .io_axi_b_ready(axi4_to_ahb_2_io_axi_b_ready),
    .io_axi_ar_valid(axi4_to_ahb_2_io_axi_ar_valid),
    .io_axi_ar_bits_addr(axi4_to_ahb_2_io_axi_ar_bits_addr),
    .io_axi_ar_bits_size(axi4_to_ahb_2_io_axi_ar_bits_size),
    .io_ahb_in_hready(axi4_to_ahb_2_io_ahb_in_hready),
    .io_ahb_in_hresp(axi4_to_ahb_2_io_ahb_in_hresp),
    .io_ahb_out_htrans(axi4_to_ahb_2_io_ahb_out_htrans),
    .io_ahb_out_hwrite(axi4_to_ahb_2_io_ahb_out_hwrite)
  );
  ahb_to_axi4 ahb_to_axi4 ( // @[quasar.scala 245:33]
    .clock(ahb_to_axi4_clock),
    .reset(ahb_to_axi4_reset),
    .io_scan_mode(ahb_to_axi4_io_scan_mode),
    .io_bus_clk_en(ahb_to_axi4_io_bus_clk_en),
    .io_axi_aw_valid(ahb_to_axi4_io_axi_aw_valid),
    .io_axi_ar_valid(ahb_to_axi4_io_axi_ar_valid),
    .io_axi_r_valid(ahb_to_axi4_io_axi_r_valid),
    .io_axi_r_bits_resp(ahb_to_axi4_io_axi_r_bits_resp),
    .io_ahb_sig_in_hready(ahb_to_axi4_io_ahb_sig_in_hready),
    .io_ahb_sig_in_hresp(ahb_to_axi4_io_ahb_sig_in_hresp),
    .io_ahb_sig_out_haddr(ahb_to_axi4_io_ahb_sig_out_haddr),
    .io_ahb_sig_out_hsize(ahb_to_axi4_io_ahb_sig_out_hsize),
    .io_ahb_sig_out_htrans(ahb_to_axi4_io_ahb_sig_out_htrans),
    .io_ahb_sig_out_hwrite(ahb_to_axi4_io_ahb_sig_out_hwrite),
    .io_ahb_hsel(ahb_to_axi4_io_ahb_hsel),
    .io_ahb_hreadyin(ahb_to_axi4_io_ahb_hreadyin)
  );
  assign io_core_rst_l = reset & _T_2; // @[quasar.scala 80:17]
  assign io_rv_trace_pkt_rv_i_valid_ip = dec_io_rv_trace_pkt_rv_i_valid_ip; // @[quasar.scala 220:19]
  assign io_rv_trace_pkt_rv_i_insn_ip = dec_io_rv_trace_pkt_rv_i_insn_ip; // @[quasar.scala 220:19]
  assign io_rv_trace_pkt_rv_i_address_ip = dec_io_rv_trace_pkt_rv_i_address_ip; // @[quasar.scala 220:19]
  assign io_rv_trace_pkt_rv_i_exception_ip = dec_io_rv_trace_pkt_rv_i_exception_ip; // @[quasar.scala 220:19]
  assign io_rv_trace_pkt_rv_i_ecause_ip = dec_io_rv_trace_pkt_rv_i_ecause_ip; // @[quasar.scala 220:19]
  assign io_rv_trace_pkt_rv_i_interrupt_ip = dec_io_rv_trace_pkt_rv_i_interrupt_ip; // @[quasar.scala 220:19]
  assign io_rv_trace_pkt_rv_i_tval_ip = dec_io_rv_trace_pkt_rv_i_tval_ip; // @[quasar.scala 220:19]
  assign io_dccm_clk_override = dec_io_dec_tlu_dccm_clk_override; // @[quasar.scala 223:24]
  assign io_icm_clk_override = dec_io_dec_tlu_icm_clk_override; // @[quasar.scala 224:23]
  assign io_dec_tlu_core_ecc_disable = dec_io_ifu_dec_dec_mem_ctrl_dec_tlu_core_ecc_disable; // @[quasar.scala 225:31]
  assign io_o_cpu_halt_ack = dec_io_o_cpu_halt_ack; // @[quasar.scala 226:21]
  assign io_o_cpu_halt_status = dec_io_o_cpu_halt_status; // @[quasar.scala 227:24]
  assign io_o_cpu_run_ack = dec_io_o_cpu_run_ack; // @[quasar.scala 228:20]
  assign io_o_debug_mode_status = dec_io_o_debug_mode_status; // @[quasar.scala 229:26]
  assign io_mpc_debug_halt_ack = dec_io_mpc_debug_halt_ack; // @[quasar.scala 230:25]
  assign io_mpc_debug_run_ack = dec_io_mpc_debug_run_ack; // @[quasar.scala 231:24]
  assign io_debug_brkpt_status = dec_io_debug_brkpt_status; // @[quasar.scala 232:25]
  assign io_dec_tlu_perfcnt0 = dec_io_dec_tlu_perfcnt0; // @[quasar.scala 233:23]
  assign io_dec_tlu_perfcnt1 = dec_io_dec_tlu_perfcnt1; // @[quasar.scala 234:23]
  assign io_dec_tlu_perfcnt2 = dec_io_dec_tlu_perfcnt2; // @[quasar.scala 235:23]
  assign io_dec_tlu_perfcnt3 = dec_io_dec_tlu_perfcnt3; // @[quasar.scala 236:23]
  assign io_dccm_wren = lsu_io_dccm_wren; // @[quasar.scala 238:11]
  assign io_dccm_rden = lsu_io_dccm_rden; // @[quasar.scala 238:11]
  assign io_dccm_wr_addr_lo = lsu_io_dccm_wr_addr_lo; // @[quasar.scala 238:11]
  assign io_dccm_wr_addr_hi = lsu_io_dccm_wr_addr_hi; // @[quasar.scala 238:11]
  assign io_dccm_rd_addr_lo = lsu_io_dccm_rd_addr_lo; // @[quasar.scala 238:11]
  assign io_dccm_rd_addr_hi = lsu_io_dccm_rd_addr_hi; // @[quasar.scala 238:11]
  assign io_dccm_wr_data_lo = lsu_io_dccm_wr_data_lo; // @[quasar.scala 238:11]
  assign io_dccm_wr_data_hi = lsu_io_dccm_wr_data_hi; // @[quasar.scala 238:11]
  assign io_ic_rw_addr = ifu_io_ic_rw_addr; // @[quasar.scala 101:13]
  assign io_ic_tag_valid = ifu_io_ic_tag_valid; // @[quasar.scala 101:13]
  assign io_ic_rd_en = ifu_io_ic_rd_en; // @[quasar.scala 101:13]
  assign io_ic_debug_wr_data = ifu_io_ic_debug_wr_data; // @[quasar.scala 101:13]
  assign io_ic_debug_addr = ifu_io_ic_debug_addr; // @[quasar.scala 101:13]
  assign io_ic_debug_rd_en = ifu_io_ic_debug_rd_en; // @[quasar.scala 101:13]
  assign io_ic_debug_wr_en = ifu_io_ic_debug_wr_en; // @[quasar.scala 101:13]
  assign io_ic_debug_tag_array = ifu_io_ic_debug_tag_array; // @[quasar.scala 101:13]
  assign io_ic_debug_way = ifu_io_ic_debug_way; // @[quasar.scala 101:13]
  assign io_ic_premux_data = ifu_io_ic_premux_data; // @[quasar.scala 101:13]
  assign io_ic_sel_premux_data = ifu_io_ic_sel_premux_data; // @[quasar.scala 101:13]
  assign io_iccm_rw_addr = ifu_io_iccm_rw_addr; // @[quasar.scala 102:15]
  assign io_iccm_buf_correct_ecc = ifu_io_iccm_buf_correct_ecc; // @[quasar.scala 102:15]
  assign io_iccm_correction_state = ifu_io_iccm_correction_state; // @[quasar.scala 102:15]
  assign io_iccm_wren = ifu_io_iccm_wren; // @[quasar.scala 102:15]
  assign io_iccm_rden = ifu_io_iccm_rden; // @[quasar.scala 102:15]
  assign io_iccm_wr_size = ifu_io_iccm_wr_size; // @[quasar.scala 102:15]
  assign io_iccm_wr_data = ifu_io_iccm_wr_data; // @[quasar.scala 102:15]
  assign ifu_clock = clock;
  assign ifu_reset = io_core_rst_l; // @[quasar.scala 91:13]
  assign ifu_io_exu_flush_final = dec_io_exu_flush_final; // @[quasar.scala 96:26]
  assign ifu_io_exu_flush_path_final = exu_io_exu_flush_path_final; // @[quasar.scala 97:31]
  assign ifu_io_free_clk = rvclkhdr_io_l1clk; // @[quasar.scala 93:19]
  assign ifu_io_active_clk = rvclkhdr_1_io_l1clk; // @[quasar.scala 94:21]
  assign ifu_io_ifu_dec_dec_aln_aln_dec_dec_i0_decode_d = dec_io_ifu_dec_dec_aln_aln_dec_dec_i0_decode_d; // @[quasar.scala 89:18]
  assign ifu_io_ifu_dec_dec_mem_ctrl_dec_tlu_flush_err_wb = dec_io_ifu_dec_dec_mem_ctrl_dec_tlu_flush_err_wb; // @[quasar.scala 89:18]
  assign ifu_io_ifu_dec_dec_mem_ctrl_dec_tlu_i0_commit_cmt = dec_io_ifu_dec_dec_mem_ctrl_dec_tlu_i0_commit_cmt; // @[quasar.scala 89:18]
  assign ifu_io_ifu_dec_dec_mem_ctrl_dec_tlu_force_halt = dec_io_ifu_dec_dec_mem_ctrl_dec_tlu_force_halt; // @[quasar.scala 89:18]
  assign ifu_io_ifu_dec_dec_mem_ctrl_dec_tlu_fence_i_wb = dec_io_ifu_dec_dec_mem_ctrl_dec_tlu_fence_i_wb; // @[quasar.scala 89:18]
  assign ifu_io_ifu_dec_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_wrdata = dec_io_ifu_dec_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_wrdata; // @[quasar.scala 89:18 quasar.scala 107:51]
  assign ifu_io_ifu_dec_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_dicawics = dec_io_ifu_dec_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_dicawics; // @[quasar.scala 89:18 quasar.scala 107:51]
  assign ifu_io_ifu_dec_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_rd_valid = dec_io_ifu_dec_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_rd_valid; // @[quasar.scala 89:18 quasar.scala 107:51]
  assign ifu_io_ifu_dec_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_wr_valid = dec_io_ifu_dec_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_wr_valid; // @[quasar.scala 89:18 quasar.scala 107:51]
  assign ifu_io_ifu_dec_dec_mem_ctrl_dec_tlu_core_ecc_disable = dec_io_ifu_dec_dec_mem_ctrl_dec_tlu_core_ecc_disable; // @[quasar.scala 89:18]
  assign ifu_io_ifu_dec_dec_ifc_dec_tlu_flush_noredir_wb = dec_io_ifu_dec_dec_ifc_dec_tlu_flush_noredir_wb; // @[quasar.scala 89:18]
  assign ifu_io_ifu_dec_dec_ifc_dec_tlu_mrac_ff = dec_io_ifu_dec_dec_ifc_dec_tlu_mrac_ff; // @[quasar.scala 89:18]
  assign ifu_io_ifu_dec_dec_bp_dec_tlu_br0_r_pkt_valid = dec_io_ifu_dec_dec_bp_dec_tlu_br0_r_pkt_valid; // @[quasar.scala 89:18]
  assign ifu_io_ifu_dec_dec_bp_dec_tlu_br0_r_pkt_bits_hist = dec_io_ifu_dec_dec_bp_dec_tlu_br0_r_pkt_bits_hist; // @[quasar.scala 89:18]
  assign ifu_io_ifu_dec_dec_bp_dec_tlu_br0_r_pkt_bits_br_error = dec_io_ifu_dec_dec_bp_dec_tlu_br0_r_pkt_bits_br_error; // @[quasar.scala 89:18]
  assign ifu_io_ifu_dec_dec_bp_dec_tlu_br0_r_pkt_bits_br_start_error = dec_io_ifu_dec_dec_bp_dec_tlu_br0_r_pkt_bits_br_start_error; // @[quasar.scala 89:18]
  assign ifu_io_ifu_dec_dec_bp_dec_tlu_br0_r_pkt_bits_way = dec_io_ifu_dec_dec_bp_dec_tlu_br0_r_pkt_bits_way; // @[quasar.scala 89:18]
  assign ifu_io_ifu_dec_dec_bp_dec_tlu_br0_r_pkt_bits_middle = dec_io_ifu_dec_dec_bp_dec_tlu_br0_r_pkt_bits_middle; // @[quasar.scala 89:18]
  assign ifu_io_ifu_dec_dec_bp_dec_tlu_flush_leak_one_wb = dec_io_ifu_dec_dec_bp_dec_tlu_flush_leak_one_wb; // @[quasar.scala 89:18]
  assign ifu_io_ifu_dec_dec_bp_dec_tlu_bpred_disable = dec_io_ifu_dec_dec_bp_dec_tlu_bpred_disable; // @[quasar.scala 89:18]
  assign ifu_io_exu_ifu_exu_bp_exu_i0_br_index_r = exu_io_dec_exu_tlu_exu_exu_i0_br_index_r; // @[quasar.scala 103:25 quasar.scala 105:43]
  assign ifu_io_exu_ifu_exu_bp_exu_i0_br_fghr_r = exu_io_exu_bp_exu_i0_br_fghr_r; // @[quasar.scala 103:25 quasar.scala 104:42]
  assign ifu_io_exu_ifu_exu_bp_exu_mp_pkt_bits_misp = exu_io_exu_bp_exu_mp_pkt_bits_misp; // @[quasar.scala 103:25]
  assign ifu_io_exu_ifu_exu_bp_exu_mp_pkt_bits_ataken = exu_io_exu_bp_exu_mp_pkt_bits_ataken; // @[quasar.scala 103:25]
  assign ifu_io_exu_ifu_exu_bp_exu_mp_pkt_bits_boffset = exu_io_exu_bp_exu_mp_pkt_bits_boffset; // @[quasar.scala 103:25]
  assign ifu_io_exu_ifu_exu_bp_exu_mp_pkt_bits_pc4 = exu_io_exu_bp_exu_mp_pkt_bits_pc4; // @[quasar.scala 103:25]
  assign ifu_io_exu_ifu_exu_bp_exu_mp_pkt_bits_hist = exu_io_exu_bp_exu_mp_pkt_bits_hist; // @[quasar.scala 103:25]
  assign ifu_io_exu_ifu_exu_bp_exu_mp_pkt_bits_toffset = exu_io_exu_bp_exu_mp_pkt_bits_toffset; // @[quasar.scala 103:25]
  assign ifu_io_exu_ifu_exu_bp_exu_mp_pkt_bits_pcall = exu_io_exu_bp_exu_mp_pkt_bits_pcall; // @[quasar.scala 103:25]
  assign ifu_io_exu_ifu_exu_bp_exu_mp_pkt_bits_pret = exu_io_exu_bp_exu_mp_pkt_bits_pret; // @[quasar.scala 103:25]
  assign ifu_io_exu_ifu_exu_bp_exu_mp_pkt_bits_pja = exu_io_exu_bp_exu_mp_pkt_bits_pja; // @[quasar.scala 103:25]
  assign ifu_io_exu_ifu_exu_bp_exu_mp_pkt_bits_way = exu_io_exu_bp_exu_mp_pkt_bits_way; // @[quasar.scala 103:25]
  assign ifu_io_exu_ifu_exu_bp_exu_mp_eghr = exu_io_exu_bp_exu_mp_eghr; // @[quasar.scala 103:25]
  assign ifu_io_exu_ifu_exu_bp_exu_mp_fghr = exu_io_exu_bp_exu_mp_fghr; // @[quasar.scala 103:25]
  assign ifu_io_exu_ifu_exu_bp_exu_mp_index = exu_io_exu_bp_exu_mp_index; // @[quasar.scala 103:25]
  assign ifu_io_exu_ifu_exu_bp_exu_mp_btag = exu_io_exu_bp_exu_mp_btag; // @[quasar.scala 103:25]
  assign ifu_io_iccm_rd_data = io_iccm_rd_data; // @[quasar.scala 102:15]
  assign ifu_io_iccm_rd_data_ecc = io_iccm_rd_data_ecc; // @[quasar.scala 102:15]
  assign ifu_io_ic_rd_data = io_ic_rd_data; // @[quasar.scala 101:13]
  assign ifu_io_ic_debug_rd_data = io_ic_debug_rd_data; // @[quasar.scala 101:13]
  assign ifu_io_ic_tag_debug_rd_data = io_ic_tag_debug_rd_data; // @[quasar.scala 101:13]
  assign ifu_io_ic_eccerr = io_ic_eccerr; // @[quasar.scala 101:13]
  assign ifu_io_ic_rd_hit = io_ic_rd_hit; // @[quasar.scala 101:13]
  assign ifu_io_ic_tag_perr = io_ic_tag_perr; // @[quasar.scala 101:13]
  assign ifu_io_ifu_bus_clk_en = io_ifu_bus_clk_en; // @[quasar.scala 99:25]
  assign ifu_io_ifu_dma_dma_ifc_dma_iccm_stall_any = dma_ctrl_io_ifu_dma_dma_ifc_dma_iccm_stall_any; // @[quasar.scala 100:18]
  assign ifu_io_ifu_dma_dma_mem_ctl_dma_iccm_req = dma_ctrl_io_ifu_dma_dma_mem_ctl_dma_iccm_req; // @[quasar.scala 100:18]
  assign ifu_io_ifu_dma_dma_mem_ctl_dma_mem_addr = dma_ctrl_io_ifu_dma_dma_mem_ctl_dma_mem_addr; // @[quasar.scala 100:18]
  assign ifu_io_ifu_dma_dma_mem_ctl_dma_mem_sz = dma_ctrl_io_ifu_dma_dma_mem_ctl_dma_mem_sz; // @[quasar.scala 100:18]
  assign ifu_io_ifu_dma_dma_mem_ctl_dma_mem_write = dma_ctrl_io_ifu_dma_dma_mem_ctl_dma_mem_write; // @[quasar.scala 100:18]
  assign ifu_io_ifu_dma_dma_mem_ctl_dma_mem_wdata = dma_ctrl_io_ifu_dma_dma_mem_ctl_dma_mem_wdata; // @[quasar.scala 100:18]
  assign ifu_io_ifu_dma_dma_mem_ctl_dma_mem_tag = dma_ctrl_io_ifu_dma_dma_mem_ctl_dma_mem_tag; // @[quasar.scala 100:18]
  assign ifu_io_dec_tlu_flush_lower_wb = dec_io_dec_exu_tlu_exu_dec_tlu_flush_lower_r; // @[quasar.scala 106:33]
  assign ifu_io_scan_mode = io_scan_mode; // @[quasar.scala 92:20]
  assign dec_clock = clock;
  assign dec_reset = io_core_rst_l; // @[quasar.scala 110:13]
  assign dec_io_free_clk = rvclkhdr_io_l1clk; // @[quasar.scala 111:19]
  assign dec_io_active_clk = rvclkhdr_1_io_l1clk; // @[quasar.scala 112:21]
  assign dec_io_lsu_fastint_stall_any = lsu_io_lsu_fastint_stall_any; // @[quasar.scala 113:32]
  assign dec_io_rst_vec = io_rst_vec; // @[quasar.scala 114:18]
  assign dec_io_nmi_int = io_nmi_int; // @[quasar.scala 115:18]
  assign dec_io_nmi_vec = io_nmi_vec; // @[quasar.scala 116:18]
  assign dec_io_i_cpu_halt_req = io_i_cpu_halt_req; // @[quasar.scala 117:25]
  assign dec_io_i_cpu_run_req = io_i_cpu_run_req; // @[quasar.scala 118:24]
  assign dec_io_core_id = io_core_id; // @[quasar.scala 119:18]
  assign dec_io_mpc_debug_halt_req = io_mpc_debug_halt_req; // @[quasar.scala 120:29]
  assign dec_io_mpc_debug_run_req = io_mpc_debug_run_req; // @[quasar.scala 121:28]
  assign dec_io_mpc_reset_run_req = io_mpc_reset_run_req; // @[quasar.scala 122:28]
  assign dec_io_lsu_pmu_misaligned_m = lsu_io_lsu_pmu_misaligned_m; // @[quasar.scala 125:31]
  assign dec_io_lsu_fir_addr = lsu_io_lsu_fir_addr; // @[quasar.scala 128:23]
  assign dec_io_lsu_fir_error = lsu_io_lsu_fir_error; // @[quasar.scala 129:24]
  assign dec_io_lsu_trigger_match_m = lsu_io_lsu_trigger_match_m; // @[quasar.scala 130:30]
  assign dec_io_lsu_idle_any = lsu_io_lsu_idle_any; // @[quasar.scala 132:23]
  assign dec_io_lsu_error_pkt_r_valid = lsu_io_lsu_error_pkt_r_valid; // @[quasar.scala 133:26]
  assign dec_io_lsu_error_pkt_r_bits_single_ecc_error = lsu_io_lsu_error_pkt_r_bits_single_ecc_error; // @[quasar.scala 133:26]
  assign dec_io_lsu_error_pkt_r_bits_inst_type = lsu_io_lsu_error_pkt_r_bits_inst_type; // @[quasar.scala 133:26]
  assign dec_io_lsu_error_pkt_r_bits_exc_type = lsu_io_lsu_error_pkt_r_bits_exc_type; // @[quasar.scala 133:26]
  assign dec_io_lsu_error_pkt_r_bits_mscause = lsu_io_lsu_error_pkt_r_bits_mscause; // @[quasar.scala 133:26]
  assign dec_io_lsu_error_pkt_r_bits_addr = lsu_io_lsu_error_pkt_r_bits_addr; // @[quasar.scala 133:26]
  assign dec_io_lsu_single_ecc_error_incr = lsu_io_lsu_single_ecc_error_incr; // @[quasar.scala 134:36]
  assign dec_io_exu_div_result = exu_io_exu_div_result; // @[quasar.scala 135:25]
  assign dec_io_exu_div_wren = exu_io_exu_div_wren; // @[quasar.scala 136:23]
  assign dec_io_lsu_result_m = lsu_io_lsu_result_m; // @[quasar.scala 137:23]
  assign dec_io_lsu_result_corr_r = lsu_io_lsu_result_corr_r; // @[quasar.scala 138:28]
  assign dec_io_lsu_load_stall_any = lsu_io_lsu_load_stall_any; // @[quasar.scala 139:29]
  assign dec_io_lsu_store_stall_any = lsu_io_lsu_store_stall_any; // @[quasar.scala 140:30]
  assign dec_io_iccm_dma_sb_error = ifu_io_iccm_dma_sb_error; // @[quasar.scala 141:28]
  assign dec_io_exu_flush_final = exu_io_exu_flush_final; // @[quasar.scala 142:26]
  assign dec_io_timer_int = io_timer_int; // @[quasar.scala 148:20]
  assign dec_io_soft_int = io_soft_int; // @[quasar.scala 144:19]
  assign dec_io_dbg_halt_req = dbg_io_dbg_halt_req; // @[quasar.scala 145:23]
  assign dec_io_dbg_resume_req = dbg_io_dbg_resume_req; // @[quasar.scala 146:25]
  assign dec_io_exu_i0_br_way_r = exu_io_exu_bp_exu_i0_br_way_r; // @[quasar.scala 147:26]
  assign dec_io_scan_mode = io_scan_mode; // @[quasar.scala 149:20]
  assign dec_io_ifu_dec_dec_aln_aln_dec_ifu_i0_cinst = ifu_io_ifu_dec_dec_aln_aln_dec_ifu_i0_cinst; // @[quasar.scala 89:18]
  assign dec_io_ifu_dec_dec_aln_aln_ib_ifu_i0_icaf = ifu_io_ifu_dec_dec_aln_aln_ib_ifu_i0_icaf; // @[quasar.scala 89:18]
  assign dec_io_ifu_dec_dec_aln_aln_ib_ifu_i0_icaf_type = ifu_io_ifu_dec_dec_aln_aln_ib_ifu_i0_icaf_type; // @[quasar.scala 89:18]
  assign dec_io_ifu_dec_dec_aln_aln_ib_ifu_i0_icaf_f1 = ifu_io_ifu_dec_dec_aln_aln_ib_ifu_i0_icaf_f1; // @[quasar.scala 89:18]
  assign dec_io_ifu_dec_dec_aln_aln_ib_ifu_i0_dbecc = ifu_io_ifu_dec_dec_aln_aln_ib_ifu_i0_dbecc; // @[quasar.scala 89:18]
  assign dec_io_ifu_dec_dec_aln_aln_ib_ifu_i0_bp_index = ifu_io_ifu_dec_dec_aln_aln_ib_ifu_i0_bp_index; // @[quasar.scala 89:18]
  assign dec_io_ifu_dec_dec_aln_aln_ib_ifu_i0_bp_fghr = ifu_io_ifu_dec_dec_aln_aln_ib_ifu_i0_bp_fghr; // @[quasar.scala 89:18]
  assign dec_io_ifu_dec_dec_aln_aln_ib_ifu_i0_bp_btag = ifu_io_ifu_dec_dec_aln_aln_ib_ifu_i0_bp_btag; // @[quasar.scala 89:18]
  assign dec_io_ifu_dec_dec_aln_aln_ib_ifu_i0_valid = ifu_io_ifu_dec_dec_aln_aln_ib_ifu_i0_valid; // @[quasar.scala 89:18]
  assign dec_io_ifu_dec_dec_aln_aln_ib_ifu_i0_instr = ifu_io_ifu_dec_dec_aln_aln_ib_ifu_i0_instr; // @[quasar.scala 89:18]
  assign dec_io_ifu_dec_dec_aln_aln_ib_ifu_i0_pc = ifu_io_ifu_dec_dec_aln_aln_ib_ifu_i0_pc; // @[quasar.scala 89:18]
  assign dec_io_ifu_dec_dec_aln_aln_ib_ifu_i0_pc4 = ifu_io_ifu_dec_dec_aln_aln_ib_ifu_i0_pc4; // @[quasar.scala 89:18]
  assign dec_io_ifu_dec_dec_aln_aln_ib_i0_brp_valid = ifu_io_ifu_dec_dec_aln_aln_ib_i0_brp_valid; // @[quasar.scala 89:18]
  assign dec_io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_toffset = ifu_io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_toffset; // @[quasar.scala 89:18]
  assign dec_io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_hist = ifu_io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_hist; // @[quasar.scala 89:18]
  assign dec_io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_br_error = ifu_io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_br_error; // @[quasar.scala 89:18]
  assign dec_io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_br_start_error = ifu_io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_br_start_error; // @[quasar.scala 89:18]
  assign dec_io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_prett = ifu_io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_prett; // @[quasar.scala 89:18]
  assign dec_io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_way = ifu_io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_way; // @[quasar.scala 89:18]
  assign dec_io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_ret = ifu_io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_ret; // @[quasar.scala 89:18]
  assign dec_io_ifu_dec_dec_aln_ifu_pmu_instr_aligned = ifu_io_ifu_dec_dec_aln_ifu_pmu_instr_aligned; // @[quasar.scala 89:18]
  assign dec_io_ifu_dec_dec_mem_ctrl_ifu_pmu_ic_miss = ifu_io_ifu_dec_dec_mem_ctrl_ifu_pmu_ic_miss; // @[quasar.scala 89:18]
  assign dec_io_ifu_dec_dec_mem_ctrl_ifu_pmu_ic_hit = ifu_io_ifu_dec_dec_mem_ctrl_ifu_pmu_ic_hit; // @[quasar.scala 89:18]
  assign dec_io_ifu_dec_dec_mem_ctrl_ifu_pmu_bus_error = ifu_io_ifu_dec_dec_mem_ctrl_ifu_pmu_bus_error; // @[quasar.scala 89:18]
  assign dec_io_ifu_dec_dec_mem_ctrl_ifu_pmu_bus_busy = ifu_io_ifu_dec_dec_mem_ctrl_ifu_pmu_bus_busy; // @[quasar.scala 89:18]
  assign dec_io_ifu_dec_dec_mem_ctrl_ifu_ic_error_start = ifu_io_ifu_dec_dec_mem_ctrl_ifu_ic_error_start; // @[quasar.scala 89:18]
  assign dec_io_ifu_dec_dec_mem_ctrl_ifu_iccm_rd_ecc_single_err = ifu_io_ifu_dec_dec_mem_ctrl_ifu_iccm_rd_ecc_single_err; // @[quasar.scala 89:18]
  assign dec_io_ifu_dec_dec_mem_ctrl_ifu_ic_debug_rd_data = ifu_io_ifu_dec_dec_mem_ctrl_ifu_ic_debug_rd_data; // @[quasar.scala 89:18]
  assign dec_io_ifu_dec_dec_mem_ctrl_ifu_ic_debug_rd_data_valid = ifu_io_ifu_dec_dec_mem_ctrl_ifu_ic_debug_rd_data_valid; // @[quasar.scala 89:18]
  assign dec_io_ifu_dec_dec_mem_ctrl_ifu_miss_state_idle = ifu_io_ifu_dec_dec_mem_ctrl_ifu_miss_state_idle; // @[quasar.scala 89:18]
  assign dec_io_ifu_dec_dec_ifc_ifu_pmu_fetch_stall = ifu_io_ifu_dec_dec_ifc_ifu_pmu_fetch_stall; // @[quasar.scala 89:18]
  assign dec_io_dec_exu_dec_alu_exu_i0_pc_x = exu_io_dec_exu_dec_alu_exu_i0_pc_x; // @[quasar.scala 152:18]
  assign dec_io_dec_exu_decode_exu_exu_i0_result_x = exu_io_dec_exu_decode_exu_exu_i0_result_x; // @[quasar.scala 152:18]
  assign dec_io_dec_exu_decode_exu_exu_csr_rs1_x = exu_io_dec_exu_decode_exu_exu_csr_rs1_x; // @[quasar.scala 152:18]
  assign dec_io_dec_exu_tlu_exu_exu_i0_br_hist_r = exu_io_dec_exu_tlu_exu_exu_i0_br_hist_r; // @[quasar.scala 152:18]
  assign dec_io_dec_exu_tlu_exu_exu_i0_br_error_r = exu_io_dec_exu_tlu_exu_exu_i0_br_error_r; // @[quasar.scala 152:18]
  assign dec_io_dec_exu_tlu_exu_exu_i0_br_start_error_r = exu_io_dec_exu_tlu_exu_exu_i0_br_start_error_r; // @[quasar.scala 152:18]
  assign dec_io_dec_exu_tlu_exu_exu_i0_br_valid_r = exu_io_dec_exu_tlu_exu_exu_i0_br_valid_r; // @[quasar.scala 152:18]
  assign dec_io_dec_exu_tlu_exu_exu_i0_br_mp_r = exu_io_dec_exu_tlu_exu_exu_i0_br_mp_r; // @[quasar.scala 152:18]
  assign dec_io_dec_exu_tlu_exu_exu_i0_br_middle_r = exu_io_dec_exu_tlu_exu_exu_i0_br_middle_r; // @[quasar.scala 152:18]
  assign dec_io_dec_exu_tlu_exu_exu_pmu_i0_br_misp = exu_io_dec_exu_tlu_exu_exu_pmu_i0_br_misp; // @[quasar.scala 152:18]
  assign dec_io_dec_exu_tlu_exu_exu_pmu_i0_br_ataken = exu_io_dec_exu_tlu_exu_exu_pmu_i0_br_ataken; // @[quasar.scala 152:18]
  assign dec_io_dec_exu_tlu_exu_exu_pmu_i0_pc4 = exu_io_dec_exu_tlu_exu_exu_pmu_i0_pc4; // @[quasar.scala 152:18]
  assign dec_io_dec_exu_tlu_exu_exu_npc_r = exu_io_dec_exu_tlu_exu_exu_npc_r; // @[quasar.scala 152:18]
  assign dec_io_lsu_dec_tlu_busbuff_lsu_pmu_bus_misaligned = lsu_io_lsu_dec_tlu_busbuff_lsu_pmu_bus_misaligned; // @[quasar.scala 123:18]
  assign dec_io_lsu_dec_tlu_busbuff_lsu_pmu_bus_error = lsu_io_lsu_dec_tlu_busbuff_lsu_pmu_bus_error; // @[quasar.scala 123:18]
  assign dec_io_lsu_dec_tlu_busbuff_lsu_pmu_bus_busy = lsu_io_lsu_dec_tlu_busbuff_lsu_pmu_bus_busy; // @[quasar.scala 123:18]
  assign dec_io_lsu_dec_tlu_busbuff_lsu_imprecise_error_load_any = lsu_io_lsu_dec_tlu_busbuff_lsu_imprecise_error_load_any; // @[quasar.scala 123:18]
  assign dec_io_lsu_dec_tlu_busbuff_lsu_imprecise_error_store_any = lsu_io_lsu_dec_tlu_busbuff_lsu_imprecise_error_store_any; // @[quasar.scala 123:18]
  assign dec_io_lsu_dec_tlu_busbuff_lsu_imprecise_error_addr_any = lsu_io_lsu_dec_tlu_busbuff_lsu_imprecise_error_addr_any; // @[quasar.scala 123:18]
  assign dec_io_lsu_dec_dctl_busbuff_lsu_nonblock_load_valid_m = lsu_io_lsu_dec_dctl_busbuff_lsu_nonblock_load_valid_m; // @[quasar.scala 123:18]
  assign dec_io_lsu_dec_dctl_busbuff_lsu_nonblock_load_tag_m = lsu_io_lsu_dec_dctl_busbuff_lsu_nonblock_load_tag_m; // @[quasar.scala 123:18]
  assign dec_io_lsu_dec_dctl_busbuff_lsu_nonblock_load_inv_r = lsu_io_lsu_dec_dctl_busbuff_lsu_nonblock_load_inv_r; // @[quasar.scala 123:18]
  assign dec_io_lsu_dec_dctl_busbuff_lsu_nonblock_load_inv_tag_r = lsu_io_lsu_dec_dctl_busbuff_lsu_nonblock_load_inv_tag_r; // @[quasar.scala 123:18]
  assign dec_io_lsu_dec_dctl_busbuff_lsu_nonblock_load_data_valid = lsu_io_lsu_dec_dctl_busbuff_lsu_nonblock_load_data_valid; // @[quasar.scala 123:18]
  assign dec_io_lsu_dec_dctl_busbuff_lsu_nonblock_load_data_error = lsu_io_lsu_dec_dctl_busbuff_lsu_nonblock_load_data_error; // @[quasar.scala 123:18]
  assign dec_io_lsu_dec_dctl_busbuff_lsu_nonblock_load_data_tag = lsu_io_lsu_dec_dctl_busbuff_lsu_nonblock_load_data_tag; // @[quasar.scala 123:18]
  assign dec_io_lsu_dec_dctl_busbuff_lsu_nonblock_load_data = lsu_io_lsu_dec_dctl_busbuff_lsu_nonblock_load_data; // @[quasar.scala 123:18]
  assign dec_io_lsu_tlu_lsu_pmu_load_external_m = lsu_io_lsu_tlu_lsu_pmu_load_external_m; // @[quasar.scala 124:18]
  assign dec_io_lsu_tlu_lsu_pmu_store_external_m = lsu_io_lsu_tlu_lsu_pmu_store_external_m; // @[quasar.scala 124:18]
  assign dec_io_dec_dbg_dbg_ib_dbg_cmd_valid = dbg_io_dbg_dec_dbg_ib_dbg_cmd_valid; // @[quasar.scala 131:18]
  assign dec_io_dec_dbg_dbg_ib_dbg_cmd_write = dbg_io_dbg_dec_dbg_ib_dbg_cmd_write; // @[quasar.scala 131:18]
  assign dec_io_dec_dbg_dbg_ib_dbg_cmd_type = dbg_io_dbg_dec_dbg_ib_dbg_cmd_type; // @[quasar.scala 131:18]
  assign dec_io_dec_dbg_dbg_ib_dbg_cmd_addr = dbg_io_dbg_dec_dbg_ib_dbg_cmd_addr; // @[quasar.scala 131:18]
  assign dec_io_dec_dbg_dbg_dctl_dbg_cmd_wrdata = dbg_io_dbg_dec_dbg_dctl_dbg_cmd_wrdata; // @[quasar.scala 131:18]
  assign dec_io_dec_dma_dctl_dma_dma_dccm_stall_any = dma_ctrl_io_dec_dma_dctl_dma_dma_dccm_stall_any; // @[quasar.scala 126:18]
  assign dec_io_dec_dma_tlu_dma_dma_pmu_dccm_read = dma_ctrl_io_dec_dma_tlu_dma_dma_pmu_dccm_read; // @[quasar.scala 126:18]
  assign dec_io_dec_dma_tlu_dma_dma_pmu_dccm_write = dma_ctrl_io_dec_dma_tlu_dma_dma_pmu_dccm_write; // @[quasar.scala 126:18]
  assign dec_io_dec_dma_tlu_dma_dma_pmu_any_read = dma_ctrl_io_dec_dma_tlu_dma_dma_pmu_any_read; // @[quasar.scala 126:18]
  assign dec_io_dec_dma_tlu_dma_dma_pmu_any_write = dma_ctrl_io_dec_dma_tlu_dma_dma_pmu_any_write; // @[quasar.scala 126:18]
  assign dec_io_dec_dma_tlu_dma_dma_dccm_stall_any = dma_ctrl_io_dec_dma_tlu_dma_dma_dccm_stall_any; // @[quasar.scala 126:18]
  assign dec_io_dec_dma_tlu_dma_dma_iccm_stall_any = dma_ctrl_io_dec_dma_tlu_dma_dma_iccm_stall_any; // @[quasar.scala 126:18]
  assign dec_io_dec_pic_pic_claimid = pic_ctrl_inst_io_dec_pic_pic_claimid; // @[quasar.scala 218:28]
  assign dec_io_dec_pic_pic_pl = pic_ctrl_inst_io_dec_pic_pic_pl; // @[quasar.scala 218:28]
  assign dec_io_dec_pic_mhwakeup = pic_ctrl_inst_io_dec_pic_mhwakeup; // @[quasar.scala 218:28]
  assign dec_io_dec_pic_mexintpend = pic_ctrl_inst_io_dec_pic_mexintpend; // @[quasar.scala 218:28]
  assign dbg_clock = clock;
  assign dbg_reset = io_core_rst_l; // @[quasar.scala 177:13]
  assign dbg_io_core_dbg_rddata = dma_ctrl_io_dma_dbg_cmd_done ? dma_ctrl_io_dma_dbg_rddata : dec_io_dec_dbg_rddata; // @[quasar.scala 178:26]
  assign dbg_io_core_dbg_cmd_done = dma_ctrl_io_dma_dbg_cmd_done | dec_io_dec_dbg_cmd_done; // @[quasar.scala 179:28]
  assign dbg_io_core_dbg_cmd_fail = dma_ctrl_io_dma_dbg_cmd_fail | dec_io_dec_dbg_cmd_fail; // @[quasar.scala 180:28]
  assign dbg_io_dec_tlu_debug_mode = dec_io_dec_tlu_debug_mode; // @[quasar.scala 181:29]
  assign dbg_io_dec_tlu_dbg_halted = dec_io_dec_tlu_dbg_halted; // @[quasar.scala 182:29]
  assign dbg_io_dec_tlu_mpc_halted_only = dec_io_dec_tlu_mpc_halted_only; // @[quasar.scala 183:34]
  assign dbg_io_dec_tlu_resume_ack = dec_io_dec_tlu_resume_ack; // @[quasar.scala 184:29]
  assign dbg_io_dmi_reg_en = io_dmi_reg_en; // @[quasar.scala 185:21]
  assign dbg_io_dmi_reg_addr = io_dmi_reg_addr; // @[quasar.scala 186:23]
  assign dbg_io_dmi_reg_wr_en = io_dmi_reg_wr_en; // @[quasar.scala 187:24]
  assign dbg_io_dmi_reg_wdata = io_dmi_reg_wdata; // @[quasar.scala 188:24]
  assign dbg_io_dbg_dma_io_dma_dbg_ready = dma_ctrl_io_dbg_dma_io_dma_dbg_ready; // @[quasar.scala 202:26]
  assign dbg_io_dbg_bus_clk_en = io_dbg_bus_clk_en; // @[quasar.scala 189:25]
  assign dbg_io_dbg_rst_l = io_dbg_rst_l; // @[quasar.scala 190:20]
  assign dbg_io_clk_override = dec_io_dec_tlu_misc_clk_override; // @[quasar.scala 191:23]
  assign dbg_io_scan_mode = io_scan_mode; // @[quasar.scala 192:20]
  assign exu_clock = clock;
  assign exu_reset = io_core_rst_l; // @[quasar.scala 153:13]
  assign exu_io_scan_mode = io_scan_mode; // @[quasar.scala 154:20]
  assign exu_io_dec_exu_dec_alu_dec_i0_alu_decode_d = dec_io_dec_exu_dec_alu_dec_i0_alu_decode_d; // @[quasar.scala 152:18]
  assign exu_io_dec_exu_dec_alu_dec_csr_ren_d = dec_io_dec_exu_dec_alu_dec_csr_ren_d; // @[quasar.scala 152:18]
  assign exu_io_dec_exu_dec_alu_dec_i0_br_immed_d = dec_io_dec_exu_dec_alu_dec_i0_br_immed_d; // @[quasar.scala 152:18]
  assign exu_io_dec_exu_dec_div_div_p_valid = dec_io_dec_exu_dec_div_div_p_valid; // @[quasar.scala 152:18]
  assign exu_io_dec_exu_dec_div_div_p_bits_unsign = dec_io_dec_exu_dec_div_div_p_bits_unsign; // @[quasar.scala 152:18]
  assign exu_io_dec_exu_dec_div_div_p_bits_rem = dec_io_dec_exu_dec_div_div_p_bits_rem; // @[quasar.scala 152:18]
  assign exu_io_dec_exu_dec_div_dec_div_cancel = dec_io_dec_exu_dec_div_dec_div_cancel; // @[quasar.scala 152:18]
  assign exu_io_dec_exu_decode_exu_dec_data_en = dec_io_dec_exu_decode_exu_dec_data_en; // @[quasar.scala 152:18]
  assign exu_io_dec_exu_decode_exu_dec_ctl_en = dec_io_dec_exu_decode_exu_dec_ctl_en; // @[quasar.scala 152:18]
  assign exu_io_dec_exu_decode_exu_i0_ap_land = dec_io_dec_exu_decode_exu_i0_ap_land; // @[quasar.scala 152:18]
  assign exu_io_dec_exu_decode_exu_i0_ap_lor = dec_io_dec_exu_decode_exu_i0_ap_lor; // @[quasar.scala 152:18]
  assign exu_io_dec_exu_decode_exu_i0_ap_lxor = dec_io_dec_exu_decode_exu_i0_ap_lxor; // @[quasar.scala 152:18]
  assign exu_io_dec_exu_decode_exu_i0_ap_sll = dec_io_dec_exu_decode_exu_i0_ap_sll; // @[quasar.scala 152:18]
  assign exu_io_dec_exu_decode_exu_i0_ap_srl = dec_io_dec_exu_decode_exu_i0_ap_srl; // @[quasar.scala 152:18]
  assign exu_io_dec_exu_decode_exu_i0_ap_sra = dec_io_dec_exu_decode_exu_i0_ap_sra; // @[quasar.scala 152:18]
  assign exu_io_dec_exu_decode_exu_i0_ap_beq = dec_io_dec_exu_decode_exu_i0_ap_beq; // @[quasar.scala 152:18]
  assign exu_io_dec_exu_decode_exu_i0_ap_bne = dec_io_dec_exu_decode_exu_i0_ap_bne; // @[quasar.scala 152:18]
  assign exu_io_dec_exu_decode_exu_i0_ap_blt = dec_io_dec_exu_decode_exu_i0_ap_blt; // @[quasar.scala 152:18]
  assign exu_io_dec_exu_decode_exu_i0_ap_bge = dec_io_dec_exu_decode_exu_i0_ap_bge; // @[quasar.scala 152:18]
  assign exu_io_dec_exu_decode_exu_i0_ap_add = dec_io_dec_exu_decode_exu_i0_ap_add; // @[quasar.scala 152:18]
  assign exu_io_dec_exu_decode_exu_i0_ap_sub = dec_io_dec_exu_decode_exu_i0_ap_sub; // @[quasar.scala 152:18]
  assign exu_io_dec_exu_decode_exu_i0_ap_slt = dec_io_dec_exu_decode_exu_i0_ap_slt; // @[quasar.scala 152:18]
  assign exu_io_dec_exu_decode_exu_i0_ap_unsign = dec_io_dec_exu_decode_exu_i0_ap_unsign; // @[quasar.scala 152:18]
  assign exu_io_dec_exu_decode_exu_i0_ap_jal = dec_io_dec_exu_decode_exu_i0_ap_jal; // @[quasar.scala 152:18]
  assign exu_io_dec_exu_decode_exu_i0_ap_predict_t = dec_io_dec_exu_decode_exu_i0_ap_predict_t; // @[quasar.scala 152:18]
  assign exu_io_dec_exu_decode_exu_i0_ap_predict_nt = dec_io_dec_exu_decode_exu_i0_ap_predict_nt; // @[quasar.scala 152:18]
  assign exu_io_dec_exu_decode_exu_i0_ap_csr_write = dec_io_dec_exu_decode_exu_i0_ap_csr_write; // @[quasar.scala 152:18]
  assign exu_io_dec_exu_decode_exu_i0_ap_csr_imm = dec_io_dec_exu_decode_exu_i0_ap_csr_imm; // @[quasar.scala 152:18]
  assign exu_io_dec_exu_decode_exu_dec_i0_predict_p_d_valid = dec_io_dec_exu_decode_exu_dec_i0_predict_p_d_valid; // @[quasar.scala 152:18]
  assign exu_io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_pc4 = dec_io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_pc4; // @[quasar.scala 152:18]
  assign exu_io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_hist = dec_io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_hist; // @[quasar.scala 152:18]
  assign exu_io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_toffset = dec_io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_toffset; // @[quasar.scala 152:18]
  assign exu_io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_br_error = dec_io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_br_error; // @[quasar.scala 152:18]
  assign exu_io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_br_start_error = dec_io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_br_start_error; // @[quasar.scala 152:18]
  assign exu_io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_prett = dec_io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_prett; // @[quasar.scala 152:18]
  assign exu_io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_pcall = dec_io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_pcall; // @[quasar.scala 152:18]
  assign exu_io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_pret = dec_io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_pret; // @[quasar.scala 152:18]
  assign exu_io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_pja = dec_io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_pja; // @[quasar.scala 152:18]
  assign exu_io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_way = dec_io_dec_exu_decode_exu_dec_i0_predict_p_d_bits_way; // @[quasar.scala 152:18]
  assign exu_io_dec_exu_decode_exu_i0_predict_fghr_d = dec_io_dec_exu_decode_exu_i0_predict_fghr_d; // @[quasar.scala 152:18]
  assign exu_io_dec_exu_decode_exu_i0_predict_index_d = dec_io_dec_exu_decode_exu_i0_predict_index_d; // @[quasar.scala 152:18]
  assign exu_io_dec_exu_decode_exu_i0_predict_btag_d = dec_io_dec_exu_decode_exu_i0_predict_btag_d; // @[quasar.scala 152:18]
  assign exu_io_dec_exu_decode_exu_dec_i0_rs1_en_d = dec_io_dec_exu_decode_exu_dec_i0_rs1_en_d; // @[quasar.scala 152:18]
  assign exu_io_dec_exu_decode_exu_dec_i0_rs2_en_d = dec_io_dec_exu_decode_exu_dec_i0_rs2_en_d; // @[quasar.scala 152:18]
  assign exu_io_dec_exu_decode_exu_dec_i0_immed_d = dec_io_dec_exu_decode_exu_dec_i0_immed_d; // @[quasar.scala 152:18]
  assign exu_io_dec_exu_decode_exu_dec_i0_rs1_bypass_data_d = dec_io_dec_exu_decode_exu_dec_i0_rs1_bypass_data_d; // @[quasar.scala 152:18]
  assign exu_io_dec_exu_decode_exu_dec_i0_rs2_bypass_data_d = dec_io_dec_exu_decode_exu_dec_i0_rs2_bypass_data_d; // @[quasar.scala 152:18]
  assign exu_io_dec_exu_decode_exu_dec_i0_select_pc_d = dec_io_dec_exu_decode_exu_dec_i0_select_pc_d; // @[quasar.scala 152:18]
  assign exu_io_dec_exu_decode_exu_dec_i0_rs1_bypass_en_d = dec_io_dec_exu_decode_exu_dec_i0_rs1_bypass_en_d; // @[quasar.scala 152:18]
  assign exu_io_dec_exu_decode_exu_dec_i0_rs2_bypass_en_d = dec_io_dec_exu_decode_exu_dec_i0_rs2_bypass_en_d; // @[quasar.scala 152:18]
  assign exu_io_dec_exu_decode_exu_mul_p_valid = dec_io_dec_exu_decode_exu_mul_p_valid; // @[quasar.scala 152:18]
  assign exu_io_dec_exu_decode_exu_mul_p_bits_rs1_sign = dec_io_dec_exu_decode_exu_mul_p_bits_rs1_sign; // @[quasar.scala 152:18]
  assign exu_io_dec_exu_decode_exu_mul_p_bits_rs2_sign = dec_io_dec_exu_decode_exu_mul_p_bits_rs2_sign; // @[quasar.scala 152:18]
  assign exu_io_dec_exu_decode_exu_mul_p_bits_low = dec_io_dec_exu_decode_exu_mul_p_bits_low; // @[quasar.scala 152:18]
  assign exu_io_dec_exu_decode_exu_pred_correct_npc_x = dec_io_dec_exu_decode_exu_pred_correct_npc_x; // @[quasar.scala 152:18]
  assign exu_io_dec_exu_decode_exu_dec_extint_stall = dec_io_dec_exu_decode_exu_dec_extint_stall; // @[quasar.scala 152:18]
  assign exu_io_dec_exu_tlu_exu_dec_tlu_meihap = dec_io_dec_exu_tlu_exu_dec_tlu_meihap; // @[quasar.scala 152:18]
  assign exu_io_dec_exu_tlu_exu_dec_tlu_flush_lower_r = dec_io_dec_exu_tlu_exu_dec_tlu_flush_lower_r; // @[quasar.scala 152:18]
  assign exu_io_dec_exu_tlu_exu_dec_tlu_flush_path_r = dec_io_dec_exu_tlu_exu_dec_tlu_flush_path_r; // @[quasar.scala 152:18]
  assign exu_io_dec_exu_ib_exu_dec_i0_pc_d = dec_io_dec_exu_ib_exu_dec_i0_pc_d; // @[quasar.scala 152:18]
  assign exu_io_dec_exu_ib_exu_dec_debug_wdata_rs1_d = dec_io_dec_exu_ib_exu_dec_debug_wdata_rs1_d; // @[quasar.scala 152:18]
  assign exu_io_dec_exu_gpr_exu_gpr_i0_rs1_d = dec_io_dec_exu_gpr_exu_gpr_i0_rs1_d; // @[quasar.scala 152:18]
  assign exu_io_dec_exu_gpr_exu_gpr_i0_rs2_d = dec_io_dec_exu_gpr_exu_gpr_i0_rs2_d; // @[quasar.scala 152:18]
  assign exu_io_dbg_cmd_wrdata = dbg_io_dbg_dec_dbg_dctl_dbg_cmd_wrdata; // @[quasar.scala 155:25]
  assign lsu_clock = clock;
  assign lsu_reset = io_core_rst_l; // @[quasar.scala 158:13]
  assign lsu_io_clk_override = dec_io_dec_tlu_lsu_clk_override; // @[quasar.scala 159:23]
  assign lsu_io_lsu_dma_dma_lsc_ctl_dma_dccm_req = dma_ctrl_io_lsu_dma_dma_lsc_ctl_dma_dccm_req; // @[quasar.scala 172:18]
  assign lsu_io_lsu_dma_dma_lsc_ctl_dma_mem_addr = dma_ctrl_io_lsu_dma_dma_lsc_ctl_dma_mem_addr; // @[quasar.scala 172:18]
  assign lsu_io_lsu_dma_dma_lsc_ctl_dma_mem_sz = dma_ctrl_io_lsu_dma_dma_lsc_ctl_dma_mem_sz; // @[quasar.scala 172:18]
  assign lsu_io_lsu_dma_dma_lsc_ctl_dma_mem_write = dma_ctrl_io_lsu_dma_dma_lsc_ctl_dma_mem_write; // @[quasar.scala 172:18]
  assign lsu_io_lsu_dma_dma_lsc_ctl_dma_mem_wdata = dma_ctrl_io_lsu_dma_dma_lsc_ctl_dma_mem_wdata; // @[quasar.scala 172:18]
  assign lsu_io_lsu_dma_dma_dccm_ctl_dma_mem_addr = dma_ctrl_io_lsu_dma_dma_dccm_ctl_dma_mem_addr; // @[quasar.scala 172:18]
  assign lsu_io_lsu_dma_dma_dccm_ctl_dma_mem_wdata = dma_ctrl_io_lsu_dma_dma_dccm_ctl_dma_mem_wdata; // @[quasar.scala 172:18]
  assign lsu_io_lsu_dma_dma_mem_tag = dma_ctrl_io_lsu_dma_dma_mem_tag; // @[quasar.scala 172:18]
  assign lsu_io_lsu_pic_picm_rd_data = pic_ctrl_inst_io_lsu_pic_picm_rd_data; // @[quasar.scala 217:28]
  assign lsu_io_lsu_exu_exu_lsu_rs1_d = exu_io_lsu_exu_exu_lsu_rs1_d; // @[quasar.scala 164:18]
  assign lsu_io_lsu_exu_exu_lsu_rs2_d = exu_io_lsu_exu_exu_lsu_rs2_d; // @[quasar.scala 164:18]
  assign lsu_io_lsu_dec_tlu_busbuff_dec_tlu_external_ldfwd_disable = dec_io_lsu_dec_tlu_busbuff_dec_tlu_external_ldfwd_disable; // @[quasar.scala 123:18]
  assign lsu_io_lsu_dec_tlu_busbuff_dec_tlu_wb_coalescing_disable = dec_io_lsu_dec_tlu_busbuff_dec_tlu_wb_coalescing_disable; // @[quasar.scala 123:18]
  assign lsu_io_lsu_dec_tlu_busbuff_dec_tlu_sideeffect_posted_disable = dec_io_lsu_dec_tlu_busbuff_dec_tlu_sideeffect_posted_disable; // @[quasar.scala 123:18]
  assign lsu_io_dccm_rd_data_lo = io_dccm_rd_data_lo; // @[quasar.scala 238:11]
  assign lsu_io_dccm_rd_data_hi = io_dccm_rd_data_hi; // @[quasar.scala 238:11]
  assign lsu_io_dec_tlu_flush_lower_r = dec_io_dec_exu_tlu_exu_dec_tlu_flush_lower_r; // @[quasar.scala 160:32]
  assign lsu_io_dec_tlu_i0_kill_writeb_r = dec_io_dec_tlu_i0_kill_writeb_r; // @[quasar.scala 161:35]
  assign lsu_io_dec_tlu_force_halt = dec_io_ifu_dec_dec_mem_ctrl_dec_tlu_force_halt; // @[quasar.scala 162:29]
  assign lsu_io_dec_tlu_core_ecc_disable = dec_io_ifu_dec_dec_mem_ctrl_dec_tlu_core_ecc_disable; // @[quasar.scala 163:35]
  assign lsu_io_dec_lsu_offset_d = dec_io_dec_lsu_offset_d; // @[quasar.scala 165:27]
  assign lsu_io_lsu_p_valid = dec_io_lsu_p_valid; // @[quasar.scala 166:16]
  assign lsu_io_lsu_p_bits_fast_int = dec_io_lsu_p_bits_fast_int; // @[quasar.scala 166:16]
  assign lsu_io_lsu_p_bits_by = dec_io_lsu_p_bits_by; // @[quasar.scala 166:16]
  assign lsu_io_lsu_p_bits_half = dec_io_lsu_p_bits_half; // @[quasar.scala 166:16]
  assign lsu_io_lsu_p_bits_word = dec_io_lsu_p_bits_word; // @[quasar.scala 166:16]
  assign lsu_io_lsu_p_bits_load = dec_io_lsu_p_bits_load; // @[quasar.scala 166:16]
  assign lsu_io_lsu_p_bits_store = dec_io_lsu_p_bits_store; // @[quasar.scala 166:16]
  assign lsu_io_lsu_p_bits_unsign = dec_io_lsu_p_bits_unsign; // @[quasar.scala 166:16]
  assign lsu_io_lsu_p_bits_store_data_bypass_d = dec_io_lsu_p_bits_store_data_bypass_d; // @[quasar.scala 166:16]
  assign lsu_io_lsu_p_bits_load_ldst_bypass_d = dec_io_lsu_p_bits_load_ldst_bypass_d; // @[quasar.scala 166:16]
  assign lsu_io_trigger_pkt_any_0_select = dec_io_trigger_pkt_any_0_select; // @[quasar.scala 169:26]
  assign lsu_io_trigger_pkt_any_0_match_pkt = dec_io_trigger_pkt_any_0_match_pkt; // @[quasar.scala 169:26]
  assign lsu_io_trigger_pkt_any_0_store = dec_io_trigger_pkt_any_0_store; // @[quasar.scala 169:26]
  assign lsu_io_trigger_pkt_any_0_load = dec_io_trigger_pkt_any_0_load; // @[quasar.scala 169:26]
  assign lsu_io_trigger_pkt_any_0_tdata2 = dec_io_trigger_pkt_any_0_tdata2; // @[quasar.scala 169:26]
  assign lsu_io_trigger_pkt_any_1_select = dec_io_trigger_pkt_any_1_select; // @[quasar.scala 169:26]
  assign lsu_io_trigger_pkt_any_1_match_pkt = dec_io_trigger_pkt_any_1_match_pkt; // @[quasar.scala 169:26]
  assign lsu_io_trigger_pkt_any_1_store = dec_io_trigger_pkt_any_1_store; // @[quasar.scala 169:26]
  assign lsu_io_trigger_pkt_any_1_load = dec_io_trigger_pkt_any_1_load; // @[quasar.scala 169:26]
  assign lsu_io_trigger_pkt_any_1_tdata2 = dec_io_trigger_pkt_any_1_tdata2; // @[quasar.scala 169:26]
  assign lsu_io_trigger_pkt_any_2_select = dec_io_trigger_pkt_any_2_select; // @[quasar.scala 169:26]
  assign lsu_io_trigger_pkt_any_2_match_pkt = dec_io_trigger_pkt_any_2_match_pkt; // @[quasar.scala 169:26]
  assign lsu_io_trigger_pkt_any_2_store = dec_io_trigger_pkt_any_2_store; // @[quasar.scala 169:26]
  assign lsu_io_trigger_pkt_any_2_load = dec_io_trigger_pkt_any_2_load; // @[quasar.scala 169:26]
  assign lsu_io_trigger_pkt_any_2_tdata2 = dec_io_trigger_pkt_any_2_tdata2; // @[quasar.scala 169:26]
  assign lsu_io_trigger_pkt_any_3_select = dec_io_trigger_pkt_any_3_select; // @[quasar.scala 169:26]
  assign lsu_io_trigger_pkt_any_3_match_pkt = dec_io_trigger_pkt_any_3_match_pkt; // @[quasar.scala 169:26]
  assign lsu_io_trigger_pkt_any_3_store = dec_io_trigger_pkt_any_3_store; // @[quasar.scala 169:26]
  assign lsu_io_trigger_pkt_any_3_load = dec_io_trigger_pkt_any_3_load; // @[quasar.scala 169:26]
  assign lsu_io_trigger_pkt_any_3_tdata2 = dec_io_trigger_pkt_any_3_tdata2; // @[quasar.scala 169:26]
  assign lsu_io_dec_lsu_valid_raw_d = dec_io_dec_lsu_valid_raw_d; // @[quasar.scala 167:30]
  assign lsu_io_dec_tlu_mrac_ff = dec_io_ifu_dec_dec_ifc_dec_tlu_mrac_ff; // @[quasar.scala 168:26]
  assign lsu_io_lsu_bus_clk_en = io_lsu_bus_clk_en; // @[quasar.scala 171:25]
  assign lsu_io_scan_mode = io_scan_mode; // @[quasar.scala 173:20]
  assign lsu_io_free_clk = rvclkhdr_io_l1clk; // @[quasar.scala 174:19]
  assign pic_ctrl_inst_clock = clock;
  assign pic_ctrl_inst_reset = io_core_rst_l; // @[quasar.scala 212:23]
  assign pic_ctrl_inst_io_scan_mode = io_scan_mode; // @[quasar.scala 211:30]
  assign pic_ctrl_inst_io_free_clk = rvclkhdr_io_l1clk; // @[quasar.scala 213:29]
  assign pic_ctrl_inst_io_active_clk = rvclkhdr_1_io_l1clk; // @[quasar.scala 214:31]
  assign pic_ctrl_inst_io_clk_override = dec_io_dec_tlu_pic_clk_override; // @[quasar.scala 215:33]
  assign pic_ctrl_inst_io_extintsrc_req = {{1'd0}, io_extintsrc_req}; // @[quasar.scala 216:34]
  assign pic_ctrl_inst_io_lsu_pic_picm_wren = lsu_io_lsu_pic_picm_wren; // @[quasar.scala 217:28]
  assign pic_ctrl_inst_io_lsu_pic_picm_rden = lsu_io_lsu_pic_picm_rden; // @[quasar.scala 217:28]
  assign pic_ctrl_inst_io_lsu_pic_picm_mken = lsu_io_lsu_pic_picm_mken; // @[quasar.scala 217:28]
  assign pic_ctrl_inst_io_lsu_pic_picm_rdaddr = lsu_io_lsu_pic_picm_rdaddr; // @[quasar.scala 217:28]
  assign pic_ctrl_inst_io_lsu_pic_picm_wraddr = lsu_io_lsu_pic_picm_wraddr; // @[quasar.scala 217:28]
  assign pic_ctrl_inst_io_lsu_pic_picm_wr_data = lsu_io_lsu_pic_picm_wr_data; // @[quasar.scala 217:28]
  assign pic_ctrl_inst_io_dec_pic_dec_tlu_meicurpl = dec_io_dec_pic_dec_tlu_meicurpl; // @[quasar.scala 218:28]
  assign pic_ctrl_inst_io_dec_pic_dec_tlu_meipt = dec_io_dec_pic_dec_tlu_meipt; // @[quasar.scala 218:28]
  assign dma_ctrl_clock = clock;
  assign dma_ctrl_reset = io_core_rst_l; // @[quasar.scala 196:18]
  assign dma_ctrl_io_free_clk = rvclkhdr_io_l1clk; // @[quasar.scala 197:24]
  assign dma_ctrl_io_dma_bus_clk_en = io_dma_bus_clk_en; // @[quasar.scala 198:30]
  assign dma_ctrl_io_clk_override = dec_io_dec_tlu_misc_clk_override; // @[quasar.scala 199:28]
  assign dma_ctrl_io_scan_mode = io_scan_mode; // @[quasar.scala 200:25]
  assign dma_ctrl_io_dbg_cmd_size = dbg_io_dbg_cmd_size; // @[quasar.scala 203:28]
  assign dma_ctrl_io_dbg_dma_dbg_ib_dbg_cmd_valid = dbg_io_dbg_dma_dbg_ib_dbg_cmd_valid; // @[quasar.scala 201:23]
  assign dma_ctrl_io_dbg_dma_dbg_ib_dbg_cmd_write = dbg_io_dbg_dma_dbg_ib_dbg_cmd_write; // @[quasar.scala 201:23]
  assign dma_ctrl_io_dbg_dma_dbg_ib_dbg_cmd_type = dbg_io_dbg_dma_dbg_ib_dbg_cmd_type; // @[quasar.scala 201:23]
  assign dma_ctrl_io_dbg_dma_dbg_ib_dbg_cmd_addr = dbg_io_dbg_dma_dbg_ib_dbg_cmd_addr; // @[quasar.scala 201:23]
  assign dma_ctrl_io_dbg_dma_dbg_dctl_dbg_cmd_wrdata = dbg_io_dbg_dma_dbg_dctl_dbg_cmd_wrdata; // @[quasar.scala 201:23]
  assign dma_ctrl_io_dbg_dma_io_dbg_dma_bubble = dbg_io_dbg_dma_io_dbg_dma_bubble; // @[quasar.scala 202:26]
  assign dma_ctrl_io_dec_dma_tlu_dma_dec_tlu_dma_qos_prty = dec_io_dec_dma_tlu_dma_dec_tlu_dma_qos_prty; // @[quasar.scala 126:18]
  assign dma_ctrl_io_iccm_dma_rvalid = ifu_io_iccm_dma_rvalid; // @[quasar.scala 204:31]
  assign dma_ctrl_io_iccm_dma_ecc_error = ifu_io_iccm_dma_ecc_error; // @[quasar.scala 208:34]
  assign dma_ctrl_io_iccm_dma_rtag = ifu_io_iccm_dma_rtag; // @[quasar.scala 205:29]
  assign dma_ctrl_io_iccm_dma_rdata = ifu_io_iccm_dma_rdata; // @[quasar.scala 206:30]
  assign dma_ctrl_io_iccm_ready = ifu_io_iccm_ready; // @[quasar.scala 207:26]
  assign dma_ctrl_io_lsu_dma_dma_dccm_ctl_dccm_dma_rvalid = lsu_io_lsu_dma_dma_dccm_ctl_dccm_dma_rvalid; // @[quasar.scala 172:18]
  assign dma_ctrl_io_lsu_dma_dma_dccm_ctl_dccm_dma_ecc_error = lsu_io_lsu_dma_dma_dccm_ctl_dccm_dma_ecc_error; // @[quasar.scala 172:18]
  assign dma_ctrl_io_lsu_dma_dma_dccm_ctl_dccm_dma_rtag = lsu_io_lsu_dma_dma_dccm_ctl_dccm_dma_rtag; // @[quasar.scala 172:18]
  assign dma_ctrl_io_lsu_dma_dma_dccm_ctl_dccm_dma_rdata = lsu_io_lsu_dma_dma_dccm_ctl_dccm_dma_rdata; // @[quasar.scala 172:18]
  assign dma_ctrl_io_lsu_dma_dccm_ready = lsu_io_lsu_dma_dccm_ready; // @[quasar.scala 172:18]
  assign rvclkhdr_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_io_en = 1'h1; // @[lib.scala 345:16]
  assign rvclkhdr_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_1_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_1_io_en = _T_6 | dec_io_dec_tlu_misc_clk_override; // @[lib.scala 345:16]
  assign rvclkhdr_1_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign axi4_to_ahb_clock = clock;
  assign axi4_to_ahb_reset = reset;
  assign axi4_to_ahb_io_scan_mode = io_scan_mode; // @[quasar.scala 260:33]
  assign axi4_to_ahb_io_bus_clk_en = io_dbg_bus_clk_en; // @[quasar.scala 261:34]
  assign axi4_to_ahb_io_clk_override = dec_io_dec_tlu_bus_clk_override; // @[quasar.scala 262:36]
  assign axi4_to_ahb_io_axi_aw_valid = dbg_io_sb_axi_aw_valid; // @[quasar.scala 263:27]
  assign axi4_to_ahb_io_axi_aw_bits_addr = dbg_io_sb_axi_aw_bits_addr; // @[quasar.scala 263:27]
  assign axi4_to_ahb_io_axi_aw_bits_size = dbg_io_sb_axi_aw_bits_size; // @[quasar.scala 263:27]
  assign axi4_to_ahb_io_axi_w_valid = dbg_io_sb_axi_w_valid; // @[quasar.scala 263:27]
  assign axi4_to_ahb_io_axi_w_bits_strb = dbg_io_sb_axi_w_bits_strb; // @[quasar.scala 263:27]
  assign axi4_to_ahb_io_axi_b_ready = 1'h1; // @[quasar.scala 263:27]
  assign axi4_to_ahb_io_axi_ar_valid = dbg_io_sb_axi_ar_valid; // @[quasar.scala 263:27]
  assign axi4_to_ahb_io_axi_ar_bits_addr = dbg_io_sb_axi_ar_bits_addr; // @[quasar.scala 263:27]
  assign axi4_to_ahb_io_axi_ar_bits_size = dbg_io_sb_axi_ar_bits_size; // @[quasar.scala 263:27]
  assign axi4_to_ahb_io_ahb_in_hready = io_sb_ahb_in_hready; // @[quasar.scala 264:27]
  assign axi4_to_ahb_io_ahb_in_hresp = io_sb_ahb_in_hresp; // @[quasar.scala 264:27]
  assign axi4_to_ahb_1_clock = clock;
  assign axi4_to_ahb_1_reset = reset;
  assign axi4_to_ahb_1_io_scan_mode = io_scan_mode; // @[quasar.scala 254:34]
  assign axi4_to_ahb_1_io_bus_clk_en = io_ifu_bus_clk_en; // @[quasar.scala 255:35]
  assign axi4_to_ahb_1_io_clk_override = dec_io_dec_tlu_bus_clk_override; // @[quasar.scala 256:37]
  assign axi4_to_ahb_1_io_axi_aw_valid = 1'h0; // @[quasar.scala 257:28]
  assign axi4_to_ahb_1_io_axi_aw_bits_addr = 32'h0; // @[quasar.scala 257:28]
  assign axi4_to_ahb_1_io_axi_aw_bits_size = 3'h0; // @[quasar.scala 257:28]
  assign axi4_to_ahb_1_io_axi_w_valid = 1'h0; // @[quasar.scala 257:28]
  assign axi4_to_ahb_1_io_axi_w_bits_strb = 8'h0; // @[quasar.scala 257:28]
  assign axi4_to_ahb_1_io_axi_b_ready = 1'h0; // @[quasar.scala 257:28]
  assign axi4_to_ahb_1_io_axi_ar_valid = ifu_io_ifu_ar_valid; // @[quasar.scala 257:28]
  assign axi4_to_ahb_1_io_axi_ar_bits_addr = ifu_io_ifu_ar_bits_addr; // @[quasar.scala 257:28]
  assign axi4_to_ahb_1_io_axi_ar_bits_size = 3'h3; // @[quasar.scala 257:28]
  assign axi4_to_ahb_1_io_ahb_in_hready = io_ifu_ahb_in_hready; // @[quasar.scala 258:28]
  assign axi4_to_ahb_1_io_ahb_in_hresp = io_ifu_ahb_in_hresp; // @[quasar.scala 258:28]
  assign axi4_to_ahb_2_clock = clock;
  assign axi4_to_ahb_2_reset = reset;
  assign axi4_to_ahb_2_io_scan_mode = io_scan_mode; // @[quasar.scala 247:34]
  assign axi4_to_ahb_2_io_bus_clk_en = io_lsu_bus_clk_en; // @[quasar.scala 248:35]
  assign axi4_to_ahb_2_io_clk_override = dec_io_dec_tlu_bus_clk_override; // @[quasar.scala 249:37]
  assign axi4_to_ahb_2_io_axi_aw_valid = lsu_io_axi_aw_valid; // @[quasar.scala 250:28]
  assign axi4_to_ahb_2_io_axi_aw_bits_addr = lsu_io_axi_aw_bits_addr; // @[quasar.scala 250:28]
  assign axi4_to_ahb_2_io_axi_aw_bits_size = lsu_io_axi_aw_bits_size; // @[quasar.scala 250:28]
  assign axi4_to_ahb_2_io_axi_w_valid = lsu_io_axi_w_valid; // @[quasar.scala 250:28]
  assign axi4_to_ahb_2_io_axi_w_bits_strb = lsu_io_axi_w_bits_strb; // @[quasar.scala 250:28]
  assign axi4_to_ahb_2_io_axi_b_ready = 1'h1; // @[quasar.scala 250:28]
  assign axi4_to_ahb_2_io_axi_ar_valid = lsu_io_axi_ar_valid; // @[quasar.scala 250:28]
  assign axi4_to_ahb_2_io_axi_ar_bits_addr = lsu_io_axi_ar_bits_addr; // @[quasar.scala 250:28]
  assign axi4_to_ahb_2_io_axi_ar_bits_size = lsu_io_axi_ar_bits_size; // @[quasar.scala 250:28]
  assign axi4_to_ahb_2_io_ahb_in_hready = io_lsu_ahb_in_hready; // @[quasar.scala 251:28]
  assign axi4_to_ahb_2_io_ahb_in_hresp = io_lsu_ahb_in_hresp; // @[quasar.scala 251:28]
  assign ahb_to_axi4_clock = clock;
  assign ahb_to_axi4_reset = reset;
  assign ahb_to_axi4_io_scan_mode = io_scan_mode; // @[quasar.scala 266:34]
  assign ahb_to_axi4_io_bus_clk_en = io_dma_bus_clk_en; // @[quasar.scala 267:35]
  assign ahb_to_axi4_io_axi_r_valid = dma_ctrl_io_dma_axi_r_valid; // @[quasar.scala 269:28]
  assign ahb_to_axi4_io_axi_r_bits_resp = dma_ctrl_io_dma_axi_r_bits_resp; // @[quasar.scala 269:28]
  assign ahb_to_axi4_io_ahb_sig_out_haddr = io_dma_ahb_sig_out_haddr; // @[quasar.scala 270:28]
  assign ahb_to_axi4_io_ahb_sig_out_hsize = io_dma_ahb_sig_out_hsize; // @[quasar.scala 270:28]
  assign ahb_to_axi4_io_ahb_sig_out_htrans = io_dma_ahb_sig_out_htrans; // @[quasar.scala 270:28]
  assign ahb_to_axi4_io_ahb_sig_out_hwrite = io_dma_ahb_sig_out_hwrite; // @[quasar.scala 270:28]
  assign ahb_to_axi4_io_ahb_hsel = io_dma_ahb_hsel; // @[quasar.scala 270:28]
  assign ahb_to_axi4_io_ahb_hreadyin = io_dma_ahb_hreadyin; // @[quasar.scala 270:28]
endmodule
module quasar_wrapper(
  input         clock,
  input         reset,
  input         io_dbg_rst_l,
  input  [30:0] io_rst_vec,
  input         io_nmi_int,
  input  [30:0] io_nmi_vec,
  input  [30:0] io_jtag_id,
  input  [63:0] io_lsu_brg_in_hrdata,
  input         io_lsu_brg_in_hready,
  input         io_lsu_brg_in_hresp,
  output [31:0] io_lsu_brg_out_haddr,
  output [2:0]  io_lsu_brg_out_hburst,
  output        io_lsu_brg_out_hmastlock,
  output [3:0]  io_lsu_brg_out_hprot,
  output [2:0]  io_lsu_brg_out_hsize,
  output [1:0]  io_lsu_brg_out_htrans,
  output        io_lsu_brg_out_hwrite,
  output [63:0] io_lsu_brg_out_hwdata,
  input  [63:0] io_ifu_brg_in_hrdata,
  input         io_ifu_brg_in_hready,
  input         io_ifu_brg_in_hresp,
  output [31:0] io_ifu_brg_out_haddr,
  output [2:0]  io_ifu_brg_out_hburst,
  output        io_ifu_brg_out_hmastlock,
  output [3:0]  io_ifu_brg_out_hprot,
  output [2:0]  io_ifu_brg_out_hsize,
  output [1:0]  io_ifu_brg_out_htrans,
  output        io_ifu_brg_out_hwrite,
  output [63:0] io_ifu_brg_out_hwdata,
  input  [63:0] io_sb_brg_in_hrdata,
  input         io_sb_brg_in_hready,
  input         io_sb_brg_in_hresp,
  output [31:0] io_sb_brg_out_haddr,
  output [2:0]  io_sb_brg_out_hburst,
  output        io_sb_brg_out_hmastlock,
  output [3:0]  io_sb_brg_out_hprot,
  output [2:0]  io_sb_brg_out_hsize,
  output [1:0]  io_sb_brg_out_htrans,
  output        io_sb_brg_out_hwrite,
  output [63:0] io_sb_brg_out_hwdata,
  output [63:0] io_dma_brg_sig_in_hrdata,
  output        io_dma_brg_sig_in_hready,
  output        io_dma_brg_sig_in_hresp,
  input  [31:0] io_dma_brg_sig_out_haddr,
  input  [2:0]  io_dma_brg_sig_out_hburst,
  input         io_dma_brg_sig_out_hmastlock,
  input  [3:0]  io_dma_brg_sig_out_hprot,
  input  [2:0]  io_dma_brg_sig_out_hsize,
  input  [1:0]  io_dma_brg_sig_out_htrans,
  input         io_dma_brg_sig_out_hwrite,
  input  [63:0] io_dma_brg_sig_out_hwdata,
  input         io_dma_brg_hsel,
  input         io_dma_brg_hreadyin,
  input         io_lsu_bus_clk_en,
  input         io_ifu_bus_clk_en,
  input         io_dbg_bus_clk_en,
  input         io_dma_bus_clk_en,
  input         io_timer_int,
  input         io_soft_int,
  input  [30:0] io_extintsrc_req,
  output        io_dec_tlu_perfcnt0,
  output        io_dec_tlu_perfcnt1,
  output        io_dec_tlu_perfcnt2,
  output        io_dec_tlu_perfcnt3,
  input         io_jtag_tck,
  input         io_jtag_tms,
  input         io_jtag_tdi,
  input         io_jtag_trst_n,
  output        io_jtag_tdo,
  input  [27:0] io_core_id,
  input         io_mpc_debug_halt_req,
  input         io_mpc_debug_run_req,
  input         io_mpc_reset_run_req,
  output        io_mpc_debug_halt_ack,
  output        io_mpc_debug_run_ack,
  output        io_debug_brkpt_status,
  input         io_i_cpu_halt_req,
  input         io_i_cpu_run_req,
  output        io_o_cpu_halt_ack,
  output        io_o_cpu_halt_status,
  output        io_o_debug_mode_status,
  output        io_o_cpu_run_ack,
  input         io_mbist_mode,
  output [1:0]  io_rv_trace_pkt_rv_i_valid_ip,
  output [31:0] io_rv_trace_pkt_rv_i_insn_ip,
  output [31:0] io_rv_trace_pkt_rv_i_address_ip,
  output [1:0]  io_rv_trace_pkt_rv_i_exception_ip,
  output [4:0]  io_rv_trace_pkt_rv_i_ecause_ip,
  output [1:0]  io_rv_trace_pkt_rv_i_interrupt_ip,
  output [31:0] io_rv_trace_pkt_rv_i_tval_ip,
  input         io_scan_mode
);
  wire  mem_clk; // @[quasar_wrapper.scala 63:19]
  wire  mem_rst_l; // @[quasar_wrapper.scala 63:19]
  wire  mem_dccm_clk_override; // @[quasar_wrapper.scala 63:19]
  wire  mem_icm_clk_override; // @[quasar_wrapper.scala 63:19]
  wire  mem_dec_tlu_core_ecc_disable; // @[quasar_wrapper.scala 63:19]
  wire  mem_dccm_wren; // @[quasar_wrapper.scala 63:19]
  wire  mem_dccm_rden; // @[quasar_wrapper.scala 63:19]
  wire [15:0] mem_dccm_wr_addr_lo; // @[quasar_wrapper.scala 63:19]
  wire [15:0] mem_dccm_wr_addr_hi; // @[quasar_wrapper.scala 63:19]
  wire [15:0] mem_dccm_rd_addr_lo; // @[quasar_wrapper.scala 63:19]
  wire [15:0] mem_dccm_rd_addr_hi; // @[quasar_wrapper.scala 63:19]
  wire [38:0] mem_dccm_wr_data_lo; // @[quasar_wrapper.scala 63:19]
  wire [38:0] mem_dccm_wr_data_hi; // @[quasar_wrapper.scala 63:19]
  wire [38:0] mem_dccm_rd_data_lo; // @[quasar_wrapper.scala 63:19]
  wire [38:0] mem_dccm_rd_data_hi; // @[quasar_wrapper.scala 63:19]
  wire [14:0] mem_iccm_rw_addr; // @[quasar_wrapper.scala 63:19]
  wire  mem_iccm_buf_correct_ecc; // @[quasar_wrapper.scala 63:19]
  wire  mem_iccm_correction_state; // @[quasar_wrapper.scala 63:19]
  wire  mem_iccm_wren; // @[quasar_wrapper.scala 63:19]
  wire  mem_iccm_rden; // @[quasar_wrapper.scala 63:19]
  wire [2:0] mem_iccm_wr_size; // @[quasar_wrapper.scala 63:19]
  wire [77:0] mem_iccm_wr_data; // @[quasar_wrapper.scala 63:19]
  wire [63:0] mem_iccm_rd_data; // @[quasar_wrapper.scala 63:19]
  wire [77:0] mem_iccm_rd_data_ecc; // @[quasar_wrapper.scala 63:19]
  wire [30:0] mem_ic_rw_addr; // @[quasar_wrapper.scala 63:19]
  wire [1:0] mem_ic_tag_valid; // @[quasar_wrapper.scala 63:19]
  wire [1:0] mem_ic_wr_en; // @[quasar_wrapper.scala 63:19]
  wire  mem_ic_rd_en; // @[quasar_wrapper.scala 63:19]
  wire [70:0] mem_ic_wr_data_0; // @[quasar_wrapper.scala 63:19]
  wire [70:0] mem_ic_wr_data_1; // @[quasar_wrapper.scala 63:19]
  wire [70:0] mem_ic_debug_wr_data; // @[quasar_wrapper.scala 63:19]
  wire [9:0] mem_ic_debug_addr; // @[quasar_wrapper.scala 63:19]
  wire [63:0] mem_ic_rd_data; // @[quasar_wrapper.scala 63:19]
  wire [70:0] mem_ic_debug_rd_data; // @[quasar_wrapper.scala 63:19]
  wire [25:0] mem_ic_tag_debug_rd_data; // @[quasar_wrapper.scala 63:19]
  wire [1:0] mem_ic_eccerr; // @[quasar_wrapper.scala 63:19]
  wire [1:0] mem_ic_parerr; // @[quasar_wrapper.scala 63:19]
  wire [1:0] mem_ic_rd_hit; // @[quasar_wrapper.scala 63:19]
  wire  mem_ic_tag_perr; // @[quasar_wrapper.scala 63:19]
  wire  mem_ic_debug_rd_en; // @[quasar_wrapper.scala 63:19]
  wire  mem_ic_debug_wr_en; // @[quasar_wrapper.scala 63:19]
  wire  mem_ic_debug_tag_array; // @[quasar_wrapper.scala 63:19]
  wire [1:0] mem_ic_debug_way; // @[quasar_wrapper.scala 63:19]
  wire [63:0] mem_ic_premux_data; // @[quasar_wrapper.scala 63:19]
  wire  mem_ic_sel_premux_data; // @[quasar_wrapper.scala 63:19]
  wire  mem_scan_mode; // @[quasar_wrapper.scala 63:19]
  wire  dmi_wrapper_trst_n; // @[quasar_wrapper.scala 64:27]
  wire  dmi_wrapper_tck; // @[quasar_wrapper.scala 64:27]
  wire  dmi_wrapper_tms; // @[quasar_wrapper.scala 64:27]
  wire  dmi_wrapper_tdi; // @[quasar_wrapper.scala 64:27]
  wire  dmi_wrapper_tdo; // @[quasar_wrapper.scala 64:27]
  wire  dmi_wrapper_tdoEnable; // @[quasar_wrapper.scala 64:27]
  wire  dmi_wrapper_core_rst_n; // @[quasar_wrapper.scala 64:27]
  wire  dmi_wrapper_core_clk; // @[quasar_wrapper.scala 64:27]
  wire [30:0] dmi_wrapper_jtag_id; // @[quasar_wrapper.scala 64:27]
  wire [31:0] dmi_wrapper_rd_data; // @[quasar_wrapper.scala 64:27]
  wire [31:0] dmi_wrapper_reg_wr_data; // @[quasar_wrapper.scala 64:27]
  wire [6:0] dmi_wrapper_reg_wr_addr; // @[quasar_wrapper.scala 64:27]
  wire  dmi_wrapper_reg_en; // @[quasar_wrapper.scala 64:27]
  wire  dmi_wrapper_reg_wr_en; // @[quasar_wrapper.scala 64:27]
  wire  dmi_wrapper_dmi_hard_reset; // @[quasar_wrapper.scala 64:27]
  wire  core_clock; // @[quasar_wrapper.scala 65:20]
  wire  core_reset; // @[quasar_wrapper.scala 65:20]
  wire  core_io_lsu_ahb_in_hready; // @[quasar_wrapper.scala 65:20]
  wire  core_io_lsu_ahb_in_hresp; // @[quasar_wrapper.scala 65:20]
  wire  core_io_ifu_ahb_in_hready; // @[quasar_wrapper.scala 65:20]
  wire  core_io_ifu_ahb_in_hresp; // @[quasar_wrapper.scala 65:20]
  wire  core_io_sb_ahb_in_hready; // @[quasar_wrapper.scala 65:20]
  wire  core_io_sb_ahb_in_hresp; // @[quasar_wrapper.scala 65:20]
  wire [31:0] core_io_dma_ahb_sig_out_haddr; // @[quasar_wrapper.scala 65:20]
  wire [2:0] core_io_dma_ahb_sig_out_hsize; // @[quasar_wrapper.scala 65:20]
  wire [1:0] core_io_dma_ahb_sig_out_htrans; // @[quasar_wrapper.scala 65:20]
  wire  core_io_dma_ahb_sig_out_hwrite; // @[quasar_wrapper.scala 65:20]
  wire  core_io_dma_ahb_hsel; // @[quasar_wrapper.scala 65:20]
  wire  core_io_dma_ahb_hreadyin; // @[quasar_wrapper.scala 65:20]
  wire  core_io_dbg_rst_l; // @[quasar_wrapper.scala 65:20]
  wire [30:0] core_io_rst_vec; // @[quasar_wrapper.scala 65:20]
  wire  core_io_nmi_int; // @[quasar_wrapper.scala 65:20]
  wire [30:0] core_io_nmi_vec; // @[quasar_wrapper.scala 65:20]
  wire  core_io_core_rst_l; // @[quasar_wrapper.scala 65:20]
  wire [1:0] core_io_rv_trace_pkt_rv_i_valid_ip; // @[quasar_wrapper.scala 65:20]
  wire [31:0] core_io_rv_trace_pkt_rv_i_insn_ip; // @[quasar_wrapper.scala 65:20]
  wire [31:0] core_io_rv_trace_pkt_rv_i_address_ip; // @[quasar_wrapper.scala 65:20]
  wire [1:0] core_io_rv_trace_pkt_rv_i_exception_ip; // @[quasar_wrapper.scala 65:20]
  wire [4:0] core_io_rv_trace_pkt_rv_i_ecause_ip; // @[quasar_wrapper.scala 65:20]
  wire [1:0] core_io_rv_trace_pkt_rv_i_interrupt_ip; // @[quasar_wrapper.scala 65:20]
  wire [31:0] core_io_rv_trace_pkt_rv_i_tval_ip; // @[quasar_wrapper.scala 65:20]
  wire  core_io_dccm_clk_override; // @[quasar_wrapper.scala 65:20]
  wire  core_io_icm_clk_override; // @[quasar_wrapper.scala 65:20]
  wire  core_io_dec_tlu_core_ecc_disable; // @[quasar_wrapper.scala 65:20]
  wire  core_io_i_cpu_halt_req; // @[quasar_wrapper.scala 65:20]
  wire  core_io_i_cpu_run_req; // @[quasar_wrapper.scala 65:20]
  wire  core_io_o_cpu_halt_ack; // @[quasar_wrapper.scala 65:20]
  wire  core_io_o_cpu_halt_status; // @[quasar_wrapper.scala 65:20]
  wire  core_io_o_cpu_run_ack; // @[quasar_wrapper.scala 65:20]
  wire  core_io_o_debug_mode_status; // @[quasar_wrapper.scala 65:20]
  wire [27:0] core_io_core_id; // @[quasar_wrapper.scala 65:20]
  wire  core_io_mpc_debug_halt_req; // @[quasar_wrapper.scala 65:20]
  wire  core_io_mpc_debug_run_req; // @[quasar_wrapper.scala 65:20]
  wire  core_io_mpc_reset_run_req; // @[quasar_wrapper.scala 65:20]
  wire  core_io_mpc_debug_halt_ack; // @[quasar_wrapper.scala 65:20]
  wire  core_io_mpc_debug_run_ack; // @[quasar_wrapper.scala 65:20]
  wire  core_io_debug_brkpt_status; // @[quasar_wrapper.scala 65:20]
  wire  core_io_dec_tlu_perfcnt0; // @[quasar_wrapper.scala 65:20]
  wire  core_io_dec_tlu_perfcnt1; // @[quasar_wrapper.scala 65:20]
  wire  core_io_dec_tlu_perfcnt2; // @[quasar_wrapper.scala 65:20]
  wire  core_io_dec_tlu_perfcnt3; // @[quasar_wrapper.scala 65:20]
  wire  core_io_dccm_wren; // @[quasar_wrapper.scala 65:20]
  wire  core_io_dccm_rden; // @[quasar_wrapper.scala 65:20]
  wire [15:0] core_io_dccm_wr_addr_lo; // @[quasar_wrapper.scala 65:20]
  wire [15:0] core_io_dccm_wr_addr_hi; // @[quasar_wrapper.scala 65:20]
  wire [15:0] core_io_dccm_rd_addr_lo; // @[quasar_wrapper.scala 65:20]
  wire [15:0] core_io_dccm_rd_addr_hi; // @[quasar_wrapper.scala 65:20]
  wire [38:0] core_io_dccm_wr_data_lo; // @[quasar_wrapper.scala 65:20]
  wire [38:0] core_io_dccm_wr_data_hi; // @[quasar_wrapper.scala 65:20]
  wire [38:0] core_io_dccm_rd_data_lo; // @[quasar_wrapper.scala 65:20]
  wire [38:0] core_io_dccm_rd_data_hi; // @[quasar_wrapper.scala 65:20]
  wire [30:0] core_io_ic_rw_addr; // @[quasar_wrapper.scala 65:20]
  wire [1:0] core_io_ic_tag_valid; // @[quasar_wrapper.scala 65:20]
  wire  core_io_ic_rd_en; // @[quasar_wrapper.scala 65:20]
  wire [70:0] core_io_ic_debug_wr_data; // @[quasar_wrapper.scala 65:20]
  wire [9:0] core_io_ic_debug_addr; // @[quasar_wrapper.scala 65:20]
  wire [63:0] core_io_ic_rd_data; // @[quasar_wrapper.scala 65:20]
  wire [70:0] core_io_ic_debug_rd_data; // @[quasar_wrapper.scala 65:20]
  wire [25:0] core_io_ic_tag_debug_rd_data; // @[quasar_wrapper.scala 65:20]
  wire [1:0] core_io_ic_eccerr; // @[quasar_wrapper.scala 65:20]
  wire [1:0] core_io_ic_rd_hit; // @[quasar_wrapper.scala 65:20]
  wire  core_io_ic_tag_perr; // @[quasar_wrapper.scala 65:20]
  wire  core_io_ic_debug_rd_en; // @[quasar_wrapper.scala 65:20]
  wire  core_io_ic_debug_wr_en; // @[quasar_wrapper.scala 65:20]
  wire  core_io_ic_debug_tag_array; // @[quasar_wrapper.scala 65:20]
  wire [1:0] core_io_ic_debug_way; // @[quasar_wrapper.scala 65:20]
  wire [63:0] core_io_ic_premux_data; // @[quasar_wrapper.scala 65:20]
  wire  core_io_ic_sel_premux_data; // @[quasar_wrapper.scala 65:20]
  wire [14:0] core_io_iccm_rw_addr; // @[quasar_wrapper.scala 65:20]
  wire  core_io_iccm_buf_correct_ecc; // @[quasar_wrapper.scala 65:20]
  wire  core_io_iccm_correction_state; // @[quasar_wrapper.scala 65:20]
  wire  core_io_iccm_wren; // @[quasar_wrapper.scala 65:20]
  wire  core_io_iccm_rden; // @[quasar_wrapper.scala 65:20]
  wire [2:0] core_io_iccm_wr_size; // @[quasar_wrapper.scala 65:20]
  wire [77:0] core_io_iccm_wr_data; // @[quasar_wrapper.scala 65:20]
  wire [63:0] core_io_iccm_rd_data; // @[quasar_wrapper.scala 65:20]
  wire [77:0] core_io_iccm_rd_data_ecc; // @[quasar_wrapper.scala 65:20]
  wire  core_io_lsu_bus_clk_en; // @[quasar_wrapper.scala 65:20]
  wire  core_io_ifu_bus_clk_en; // @[quasar_wrapper.scala 65:20]
  wire  core_io_dbg_bus_clk_en; // @[quasar_wrapper.scala 65:20]
  wire  core_io_dma_bus_clk_en; // @[quasar_wrapper.scala 65:20]
  wire  core_io_dmi_reg_en; // @[quasar_wrapper.scala 65:20]
  wire [6:0] core_io_dmi_reg_addr; // @[quasar_wrapper.scala 65:20]
  wire  core_io_dmi_reg_wr_en; // @[quasar_wrapper.scala 65:20]
  wire [31:0] core_io_dmi_reg_wdata; // @[quasar_wrapper.scala 65:20]
  wire [30:0] core_io_extintsrc_req; // @[quasar_wrapper.scala 65:20]
  wire  core_io_timer_int; // @[quasar_wrapper.scala 65:20]
  wire  core_io_soft_int; // @[quasar_wrapper.scala 65:20]
  wire  core_io_scan_mode; // @[quasar_wrapper.scala 65:20]
  mem #(.ICACHE_BEAT_BITS(3), .ICCM_BITS(16), .ICACHE_BANKS_WAY(2), .ICACHE_NUM_WAYS(2), .DCCM_BYTE_WIDTH(4), .ICCM_BANK_INDEX_LO(4), .ICACHE_BANK_BITS(1), .DCCM_BITS(16), .ICACHE_BEAT_ADDR_HI(5), .ICCM_INDEX_BITS(12), .ICCM_BANK_HI(3), .ICACHE_INDEX_HI(12), .DCCM_NUM_BANKS(4), .ICACHE_BANK_LO(3), .DCCM_ENABLE(1), .ICACHE_TAG_LO(13), .ICACHE_DATA_INDEX_LO(4), .ICCM_NUM_BANKS(4), .ICACHE_ECC(1), .ICACHE_ENABLE(1), .DCCM_BANK_BITS(2), .ICCM_ENABLE(1), .ICCM_BANK_BITS(2), .ICACHE_TAG_DEPTH(128), .ICACHE_WAYPACK(0), .DCCM_SIZE(64), .ICACHE_BANK_HI(3), .DCCM_FDATA_WIDTH(39), .ICACHE_TAG_INDEX_LO(6), .ICACHE_DATA_DEPTH(512)) mem ( // @[quasar_wrapper.scala 63:19]
    .clk(mem_clk),
    .rst_l(mem_rst_l),
    .dccm_clk_override(mem_dccm_clk_override),
    .icm_clk_override(mem_icm_clk_override),
    .dec_tlu_core_ecc_disable(mem_dec_tlu_core_ecc_disable),
    .dccm_wren(mem_dccm_wren),
    .dccm_rden(mem_dccm_rden),
    .dccm_wr_addr_lo(mem_dccm_wr_addr_lo),
    .dccm_wr_addr_hi(mem_dccm_wr_addr_hi),
    .dccm_rd_addr_lo(mem_dccm_rd_addr_lo),
    .dccm_rd_addr_hi(mem_dccm_rd_addr_hi),
    .dccm_wr_data_lo(mem_dccm_wr_data_lo),
    .dccm_wr_data_hi(mem_dccm_wr_data_hi),
    .dccm_rd_data_lo(mem_dccm_rd_data_lo),
    .dccm_rd_data_hi(mem_dccm_rd_data_hi),
    .iccm_rw_addr(mem_iccm_rw_addr),
    .iccm_buf_correct_ecc(mem_iccm_buf_correct_ecc),
    .iccm_correction_state(mem_iccm_correction_state),
    .iccm_wren(mem_iccm_wren),
    .iccm_rden(mem_iccm_rden),
    .iccm_wr_size(mem_iccm_wr_size),
    .iccm_wr_data(mem_iccm_wr_data),
    .iccm_rd_data(mem_iccm_rd_data),
    .iccm_rd_data_ecc(mem_iccm_rd_data_ecc),
    .ic_rw_addr(mem_ic_rw_addr),
    .ic_tag_valid(mem_ic_tag_valid),
    .ic_wr_en(mem_ic_wr_en),
    .ic_rd_en(mem_ic_rd_en),
    .ic_wr_data_0(mem_ic_wr_data_0),
    .ic_wr_data_1(mem_ic_wr_data_1),
    .ic_debug_wr_data(mem_ic_debug_wr_data),
    .ic_debug_addr(mem_ic_debug_addr),
    .ic_rd_data(mem_ic_rd_data),
    .ic_debug_rd_data(mem_ic_debug_rd_data),
    .ic_tag_debug_rd_data(mem_ic_tag_debug_rd_data),
    .ic_eccerr(mem_ic_eccerr),
    .ic_parerr(mem_ic_parerr),
    .ic_rd_hit(mem_ic_rd_hit),
    .ic_tag_perr(mem_ic_tag_perr),
    .ic_debug_rd_en(mem_ic_debug_rd_en),
    .ic_debug_wr_en(mem_ic_debug_wr_en),
    .ic_debug_tag_array(mem_ic_debug_tag_array),
    .ic_debug_way(mem_ic_debug_way),
    .ic_premux_data(mem_ic_premux_data),
    .ic_sel_premux_data(mem_ic_sel_premux_data),
    .scan_mode(mem_scan_mode)
  );
  dmi_wrapper dmi_wrapper ( // @[quasar_wrapper.scala 64:27]
    .trst_n(dmi_wrapper_trst_n),
    .tck(dmi_wrapper_tck),
    .tms(dmi_wrapper_tms),
    .tdi(dmi_wrapper_tdi),
    .tdo(dmi_wrapper_tdo),
    .tdoEnable(dmi_wrapper_tdoEnable),
    .core_rst_n(dmi_wrapper_core_rst_n),
    .core_clk(dmi_wrapper_core_clk),
    .jtag_id(dmi_wrapper_jtag_id),
    .rd_data(dmi_wrapper_rd_data),
    .reg_wr_data(dmi_wrapper_reg_wr_data),
    .reg_wr_addr(dmi_wrapper_reg_wr_addr),
    .reg_en(dmi_wrapper_reg_en),
    .reg_wr_en(dmi_wrapper_reg_wr_en),
    .dmi_hard_reset(dmi_wrapper_dmi_hard_reset)
  );
  quasar core ( // @[quasar_wrapper.scala 65:20]
    .clock(core_clock),
    .reset(core_reset),
    .io_lsu_ahb_in_hready(core_io_lsu_ahb_in_hready),
    .io_lsu_ahb_in_hresp(core_io_lsu_ahb_in_hresp),
    .io_ifu_ahb_in_hready(core_io_ifu_ahb_in_hready),
    .io_ifu_ahb_in_hresp(core_io_ifu_ahb_in_hresp),
    .io_sb_ahb_in_hready(core_io_sb_ahb_in_hready),
    .io_sb_ahb_in_hresp(core_io_sb_ahb_in_hresp),
    .io_dma_ahb_sig_out_haddr(core_io_dma_ahb_sig_out_haddr),
    .io_dma_ahb_sig_out_hsize(core_io_dma_ahb_sig_out_hsize),
    .io_dma_ahb_sig_out_htrans(core_io_dma_ahb_sig_out_htrans),
    .io_dma_ahb_sig_out_hwrite(core_io_dma_ahb_sig_out_hwrite),
    .io_dma_ahb_hsel(core_io_dma_ahb_hsel),
    .io_dma_ahb_hreadyin(core_io_dma_ahb_hreadyin),
    .io_dbg_rst_l(core_io_dbg_rst_l),
    .io_rst_vec(core_io_rst_vec),
    .io_nmi_int(core_io_nmi_int),
    .io_nmi_vec(core_io_nmi_vec),
    .io_core_rst_l(core_io_core_rst_l),
    .io_rv_trace_pkt_rv_i_valid_ip(core_io_rv_trace_pkt_rv_i_valid_ip),
    .io_rv_trace_pkt_rv_i_insn_ip(core_io_rv_trace_pkt_rv_i_insn_ip),
    .io_rv_trace_pkt_rv_i_address_ip(core_io_rv_trace_pkt_rv_i_address_ip),
    .io_rv_trace_pkt_rv_i_exception_ip(core_io_rv_trace_pkt_rv_i_exception_ip),
    .io_rv_trace_pkt_rv_i_ecause_ip(core_io_rv_trace_pkt_rv_i_ecause_ip),
    .io_rv_trace_pkt_rv_i_interrupt_ip(core_io_rv_trace_pkt_rv_i_interrupt_ip),
    .io_rv_trace_pkt_rv_i_tval_ip(core_io_rv_trace_pkt_rv_i_tval_ip),
    .io_dccm_clk_override(core_io_dccm_clk_override),
    .io_icm_clk_override(core_io_icm_clk_override),
    .io_dec_tlu_core_ecc_disable(core_io_dec_tlu_core_ecc_disable),
    .io_i_cpu_halt_req(core_io_i_cpu_halt_req),
    .io_i_cpu_run_req(core_io_i_cpu_run_req),
    .io_o_cpu_halt_ack(core_io_o_cpu_halt_ack),
    .io_o_cpu_halt_status(core_io_o_cpu_halt_status),
    .io_o_cpu_run_ack(core_io_o_cpu_run_ack),
    .io_o_debug_mode_status(core_io_o_debug_mode_status),
    .io_core_id(core_io_core_id),
    .io_mpc_debug_halt_req(core_io_mpc_debug_halt_req),
    .io_mpc_debug_run_req(core_io_mpc_debug_run_req),
    .io_mpc_reset_run_req(core_io_mpc_reset_run_req),
    .io_mpc_debug_halt_ack(core_io_mpc_debug_halt_ack),
    .io_mpc_debug_run_ack(core_io_mpc_debug_run_ack),
    .io_debug_brkpt_status(core_io_debug_brkpt_status),
    .io_dec_tlu_perfcnt0(core_io_dec_tlu_perfcnt0),
    .io_dec_tlu_perfcnt1(core_io_dec_tlu_perfcnt1),
    .io_dec_tlu_perfcnt2(core_io_dec_tlu_perfcnt2),
    .io_dec_tlu_perfcnt3(core_io_dec_tlu_perfcnt3),
    .io_dccm_wren(core_io_dccm_wren),
    .io_dccm_rden(core_io_dccm_rden),
    .io_dccm_wr_addr_lo(core_io_dccm_wr_addr_lo),
    .io_dccm_wr_addr_hi(core_io_dccm_wr_addr_hi),
    .io_dccm_rd_addr_lo(core_io_dccm_rd_addr_lo),
    .io_dccm_rd_addr_hi(core_io_dccm_rd_addr_hi),
    .io_dccm_wr_data_lo(core_io_dccm_wr_data_lo),
    .io_dccm_wr_data_hi(core_io_dccm_wr_data_hi),
    .io_dccm_rd_data_lo(core_io_dccm_rd_data_lo),
    .io_dccm_rd_data_hi(core_io_dccm_rd_data_hi),
    .io_ic_rw_addr(core_io_ic_rw_addr),
    .io_ic_tag_valid(core_io_ic_tag_valid),
    .io_ic_rd_en(core_io_ic_rd_en),
    .io_ic_debug_wr_data(core_io_ic_debug_wr_data),
    .io_ic_debug_addr(core_io_ic_debug_addr),
    .io_ic_rd_data(core_io_ic_rd_data),
    .io_ic_debug_rd_data(core_io_ic_debug_rd_data),
    .io_ic_tag_debug_rd_data(core_io_ic_tag_debug_rd_data),
    .io_ic_eccerr(core_io_ic_eccerr),
    .io_ic_rd_hit(core_io_ic_rd_hit),
    .io_ic_tag_perr(core_io_ic_tag_perr),
    .io_ic_debug_rd_en(core_io_ic_debug_rd_en),
    .io_ic_debug_wr_en(core_io_ic_debug_wr_en),
    .io_ic_debug_tag_array(core_io_ic_debug_tag_array),
    .io_ic_debug_way(core_io_ic_debug_way),
    .io_ic_premux_data(core_io_ic_premux_data),
    .io_ic_sel_premux_data(core_io_ic_sel_premux_data),
    .io_iccm_rw_addr(core_io_iccm_rw_addr),
    .io_iccm_buf_correct_ecc(core_io_iccm_buf_correct_ecc),
    .io_iccm_correction_state(core_io_iccm_correction_state),
    .io_iccm_wren(core_io_iccm_wren),
    .io_iccm_rden(core_io_iccm_rden),
    .io_iccm_wr_size(core_io_iccm_wr_size),
    .io_iccm_wr_data(core_io_iccm_wr_data),
    .io_iccm_rd_data(core_io_iccm_rd_data),
    .io_iccm_rd_data_ecc(core_io_iccm_rd_data_ecc),
    .io_lsu_bus_clk_en(core_io_lsu_bus_clk_en),
    .io_ifu_bus_clk_en(core_io_ifu_bus_clk_en),
    .io_dbg_bus_clk_en(core_io_dbg_bus_clk_en),
    .io_dma_bus_clk_en(core_io_dma_bus_clk_en),
    .io_dmi_reg_en(core_io_dmi_reg_en),
    .io_dmi_reg_addr(core_io_dmi_reg_addr),
    .io_dmi_reg_wr_en(core_io_dmi_reg_wr_en),
    .io_dmi_reg_wdata(core_io_dmi_reg_wdata),
    .io_extintsrc_req(core_io_extintsrc_req),
    .io_timer_int(core_io_timer_int),
    .io_soft_int(core_io_soft_int),
    .io_scan_mode(core_io_scan_mode)
  );
  assign io_lsu_brg_out_haddr = 32'h0; // @[quasar_wrapper.scala 111:21]
  assign io_lsu_brg_out_hburst = 3'h0; // @[quasar_wrapper.scala 111:21]
  assign io_lsu_brg_out_hmastlock = 1'h0; // @[quasar_wrapper.scala 111:21]
  assign io_lsu_brg_out_hprot = 4'h0; // @[quasar_wrapper.scala 111:21]
  assign io_lsu_brg_out_hsize = 3'h0; // @[quasar_wrapper.scala 111:21]
  assign io_lsu_brg_out_htrans = 2'h0; // @[quasar_wrapper.scala 111:21]
  assign io_lsu_brg_out_hwrite = 1'h0; // @[quasar_wrapper.scala 111:21]
  assign io_lsu_brg_out_hwdata = 64'h0; // @[quasar_wrapper.scala 111:21]
  assign io_ifu_brg_out_haddr = 32'h0; // @[quasar_wrapper.scala 110:21]
  assign io_ifu_brg_out_hburst = 3'h0; // @[quasar_wrapper.scala 110:21]
  assign io_ifu_brg_out_hmastlock = 1'h0; // @[quasar_wrapper.scala 110:21]
  assign io_ifu_brg_out_hprot = 4'h0; // @[quasar_wrapper.scala 110:21]
  assign io_ifu_brg_out_hsize = 3'h0; // @[quasar_wrapper.scala 110:21]
  assign io_ifu_brg_out_htrans = 2'h0; // @[quasar_wrapper.scala 110:21]
  assign io_ifu_brg_out_hwrite = 1'h0; // @[quasar_wrapper.scala 110:21]
  assign io_ifu_brg_out_hwdata = 64'h0; // @[quasar_wrapper.scala 110:21]
  assign io_sb_brg_out_haddr = 32'h0; // @[quasar_wrapper.scala 112:20]
  assign io_sb_brg_out_hburst = 3'h0; // @[quasar_wrapper.scala 112:20]
  assign io_sb_brg_out_hmastlock = 1'h0; // @[quasar_wrapper.scala 112:20]
  assign io_sb_brg_out_hprot = 4'h0; // @[quasar_wrapper.scala 112:20]
  assign io_sb_brg_out_hsize = 3'h0; // @[quasar_wrapper.scala 112:20]
  assign io_sb_brg_out_htrans = 2'h0; // @[quasar_wrapper.scala 112:20]
  assign io_sb_brg_out_hwrite = 1'h0; // @[quasar_wrapper.scala 112:20]
  assign io_sb_brg_out_hwdata = 64'h0; // @[quasar_wrapper.scala 112:20]
  assign io_dma_brg_sig_in_hrdata = 64'h0; // @[quasar_wrapper.scala 113:21]
  assign io_dma_brg_sig_in_hready = 1'h0; // @[quasar_wrapper.scala 113:21]
  assign io_dma_brg_sig_in_hresp = 1'h0; // @[quasar_wrapper.scala 113:21]
  assign io_dec_tlu_perfcnt0 = core_io_dec_tlu_perfcnt0; // @[quasar_wrapper.scala 159:23]
  assign io_dec_tlu_perfcnt1 = core_io_dec_tlu_perfcnt1; // @[quasar_wrapper.scala 160:23]
  assign io_dec_tlu_perfcnt2 = core_io_dec_tlu_perfcnt2; // @[quasar_wrapper.scala 161:23]
  assign io_dec_tlu_perfcnt3 = core_io_dec_tlu_perfcnt3; // @[quasar_wrapper.scala 162:23]
  assign io_jtag_tdo = dmi_wrapper_tdo; // @[quasar_wrapper.scala 82:15]
  assign io_mpc_debug_halt_ack = core_io_mpc_debug_halt_ack; // @[quasar_wrapper.scala 155:25]
  assign io_mpc_debug_run_ack = core_io_mpc_debug_run_ack; // @[quasar_wrapper.scala 156:24]
  assign io_debug_brkpt_status = core_io_debug_brkpt_status; // @[quasar_wrapper.scala 157:25]
  assign io_o_cpu_halt_ack = core_io_o_cpu_halt_ack; // @[quasar_wrapper.scala 150:21]
  assign io_o_cpu_halt_status = core_io_o_cpu_halt_status; // @[quasar_wrapper.scala 151:24]
  assign io_o_debug_mode_status = core_io_o_debug_mode_status; // @[quasar_wrapper.scala 153:26]
  assign io_o_cpu_run_ack = core_io_o_cpu_run_ack; // @[quasar_wrapper.scala 152:20]
  assign io_rv_trace_pkt_rv_i_valid_ip = core_io_rv_trace_pkt_rv_i_valid_ip; // @[quasar_wrapper.scala 147:19]
  assign io_rv_trace_pkt_rv_i_insn_ip = core_io_rv_trace_pkt_rv_i_insn_ip; // @[quasar_wrapper.scala 147:19]
  assign io_rv_trace_pkt_rv_i_address_ip = core_io_rv_trace_pkt_rv_i_address_ip; // @[quasar_wrapper.scala 147:19]
  assign io_rv_trace_pkt_rv_i_exception_ip = core_io_rv_trace_pkt_rv_i_exception_ip; // @[quasar_wrapper.scala 147:19]
  assign io_rv_trace_pkt_rv_i_ecause_ip = core_io_rv_trace_pkt_rv_i_ecause_ip; // @[quasar_wrapper.scala 147:19]
  assign io_rv_trace_pkt_rv_i_interrupt_ip = core_io_rv_trace_pkt_rv_i_interrupt_ip; // @[quasar_wrapper.scala 147:19]
  assign io_rv_trace_pkt_rv_i_tval_ip = core_io_rv_trace_pkt_rv_i_tval_ip; // @[quasar_wrapper.scala 147:19]
  assign mem_clk = clock; // @[quasar_wrapper.scala 90:14]
  assign mem_rst_l = reset; // @[quasar_wrapper.scala 89:16]
  assign mem_dccm_clk_override = core_io_dccm_clk_override; // @[quasar_wrapper.scala 85:28]
  assign mem_icm_clk_override = core_io_icm_clk_override; // @[quasar_wrapper.scala 86:27]
  assign mem_dec_tlu_core_ecc_disable = core_io_dec_tlu_core_ecc_disable; // @[quasar_wrapper.scala 87:35]
  assign mem_dccm_wren = core_io_dccm_wren; // @[quasar_wrapper.scala 88:15]
  assign mem_dccm_rden = core_io_dccm_rden; // @[quasar_wrapper.scala 88:15]
  assign mem_dccm_wr_addr_lo = core_io_dccm_wr_addr_lo; // @[quasar_wrapper.scala 88:15]
  assign mem_dccm_wr_addr_hi = core_io_dccm_wr_addr_hi; // @[quasar_wrapper.scala 88:15]
  assign mem_dccm_rd_addr_lo = core_io_dccm_rd_addr_lo; // @[quasar_wrapper.scala 88:15]
  assign mem_dccm_rd_addr_hi = core_io_dccm_rd_addr_hi; // @[quasar_wrapper.scala 88:15]
  assign mem_dccm_wr_data_lo = core_io_dccm_wr_data_lo; // @[quasar_wrapper.scala 88:15]
  assign mem_dccm_wr_data_hi = core_io_dccm_wr_data_hi; // @[quasar_wrapper.scala 88:15]
  assign mem_iccm_rw_addr = core_io_iccm_rw_addr; // @[quasar_wrapper.scala 95:16]
  assign mem_iccm_buf_correct_ecc = core_io_iccm_buf_correct_ecc; // @[quasar_wrapper.scala 95:16]
  assign mem_iccm_correction_state = core_io_iccm_correction_state; // @[quasar_wrapper.scala 95:16]
  assign mem_iccm_wren = core_io_iccm_wren; // @[quasar_wrapper.scala 95:16]
  assign mem_iccm_rden = core_io_iccm_rden; // @[quasar_wrapper.scala 95:16]
  assign mem_iccm_wr_size = core_io_iccm_wr_size; // @[quasar_wrapper.scala 95:16]
  assign mem_iccm_wr_data = core_io_iccm_wr_data; // @[quasar_wrapper.scala 95:16]
  assign mem_ic_rw_addr = core_io_ic_rw_addr; // @[quasar_wrapper.scala 94:14]
  assign mem_ic_tag_valid = core_io_ic_tag_valid; // @[quasar_wrapper.scala 94:14]
  assign mem_ic_wr_en = 2'h0; // @[quasar_wrapper.scala 94:14]
  assign mem_ic_rd_en = core_io_ic_rd_en; // @[quasar_wrapper.scala 94:14]
  assign mem_ic_wr_data_0 = 71'h0; // @[quasar_wrapper.scala 94:14]
  assign mem_ic_wr_data_1 = 71'h0; // @[quasar_wrapper.scala 94:14]
  assign mem_ic_debug_wr_data = core_io_ic_debug_wr_data; // @[quasar_wrapper.scala 94:14]
  assign mem_ic_debug_addr = core_io_ic_debug_addr; // @[quasar_wrapper.scala 94:14]
  assign mem_ic_debug_rd_en = core_io_ic_debug_rd_en; // @[quasar_wrapper.scala 94:14]
  assign mem_ic_debug_wr_en = core_io_ic_debug_wr_en; // @[quasar_wrapper.scala 94:14]
  assign mem_ic_debug_tag_array = core_io_ic_debug_tag_array; // @[quasar_wrapper.scala 94:14]
  assign mem_ic_debug_way = core_io_ic_debug_way; // @[quasar_wrapper.scala 94:14]
  assign mem_ic_premux_data = core_io_ic_premux_data; // @[quasar_wrapper.scala 94:14]
  assign mem_ic_sel_premux_data = core_io_ic_sel_premux_data; // @[quasar_wrapper.scala 94:14]
  assign mem_scan_mode = io_scan_mode; // @[quasar_wrapper.scala 91:20]
  assign dmi_wrapper_trst_n = io_jtag_trst_n; // @[quasar_wrapper.scala 67:25]
  assign dmi_wrapper_tck = io_jtag_tck; // @[quasar_wrapper.scala 68:22]
  assign dmi_wrapper_tms = io_jtag_tms; // @[quasar_wrapper.scala 69:22]
  assign dmi_wrapper_tdi = io_jtag_tdi; // @[quasar_wrapper.scala 70:22]
  assign dmi_wrapper_core_rst_n = io_dbg_rst_l; // @[quasar_wrapper.scala 76:29]
  assign dmi_wrapper_core_clk = clock; // @[quasar_wrapper.scala 71:27]
  assign dmi_wrapper_jtag_id = io_jtag_id; // @[quasar_wrapper.scala 72:26]
  assign dmi_wrapper_rd_data = 32'h0; // @[quasar_wrapper.scala 73:26]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_lsu_ahb_in_hready = io_lsu_brg_in_hready; // @[quasar_wrapper.scala 111:21]
  assign core_io_lsu_ahb_in_hresp = io_lsu_brg_in_hresp; // @[quasar_wrapper.scala 111:21]
  assign core_io_ifu_ahb_in_hready = io_ifu_brg_in_hready; // @[quasar_wrapper.scala 110:21]
  assign core_io_ifu_ahb_in_hresp = io_ifu_brg_in_hresp; // @[quasar_wrapper.scala 110:21]
  assign core_io_sb_ahb_in_hready = io_sb_brg_in_hready; // @[quasar_wrapper.scala 112:20]
  assign core_io_sb_ahb_in_hresp = io_sb_brg_in_hresp; // @[quasar_wrapper.scala 112:20]
  assign core_io_dma_ahb_sig_out_haddr = io_dma_brg_sig_out_haddr; // @[quasar_wrapper.scala 113:21]
  assign core_io_dma_ahb_sig_out_hsize = io_dma_brg_sig_out_hsize; // @[quasar_wrapper.scala 113:21]
  assign core_io_dma_ahb_sig_out_htrans = io_dma_brg_sig_out_htrans; // @[quasar_wrapper.scala 113:21]
  assign core_io_dma_ahb_sig_out_hwrite = io_dma_brg_sig_out_hwrite; // @[quasar_wrapper.scala 113:21]
  assign core_io_dma_ahb_hsel = io_dma_brg_hsel; // @[quasar_wrapper.scala 113:21]
  assign core_io_dma_ahb_hreadyin = io_dma_brg_hreadyin; // @[quasar_wrapper.scala 113:21]
  assign core_io_dbg_rst_l = io_dbg_rst_l; // @[quasar_wrapper.scala 93:21 quasar_wrapper.scala 121:21]
  assign core_io_rst_vec = io_rst_vec; // @[quasar_wrapper.scala 122:19]
  assign core_io_nmi_int = io_nmi_int; // @[quasar_wrapper.scala 123:19]
  assign core_io_nmi_vec = io_nmi_vec; // @[quasar_wrapper.scala 124:19]
  assign core_io_i_cpu_halt_req = io_i_cpu_halt_req; // @[quasar_wrapper.scala 127:26]
  assign core_io_i_cpu_run_req = io_i_cpu_run_req; // @[quasar_wrapper.scala 128:25]
  assign core_io_core_id = io_core_id; // @[quasar_wrapper.scala 129:19]
  assign core_io_mpc_debug_halt_req = io_mpc_debug_halt_req; // @[quasar_wrapper.scala 132:30]
  assign core_io_mpc_debug_run_req = io_mpc_debug_run_req; // @[quasar_wrapper.scala 133:29]
  assign core_io_mpc_reset_run_req = io_mpc_reset_run_req; // @[quasar_wrapper.scala 134:29]
  assign core_io_dccm_rd_data_lo = mem_dccm_rd_data_lo; // @[quasar_wrapper.scala 88:15]
  assign core_io_dccm_rd_data_hi = mem_dccm_rd_data_hi; // @[quasar_wrapper.scala 88:15]
  assign core_io_ic_rd_data = mem_ic_rd_data; // @[quasar_wrapper.scala 94:14]
  assign core_io_ic_debug_rd_data = mem_ic_debug_rd_data; // @[quasar_wrapper.scala 94:14]
  assign core_io_ic_tag_debug_rd_data = mem_ic_tag_debug_rd_data; // @[quasar_wrapper.scala 94:14]
  assign core_io_ic_eccerr = mem_ic_eccerr; // @[quasar_wrapper.scala 94:14]
  assign core_io_ic_rd_hit = mem_ic_rd_hit; // @[quasar_wrapper.scala 94:14]
  assign core_io_ic_tag_perr = mem_ic_tag_perr; // @[quasar_wrapper.scala 94:14]
  assign core_io_iccm_rd_data = mem_iccm_rd_data; // @[quasar_wrapper.scala 95:16]
  assign core_io_iccm_rd_data_ecc = mem_iccm_rd_data_ecc; // @[quasar_wrapper.scala 95:16]
  assign core_io_lsu_bus_clk_en = io_lsu_bus_clk_en; // @[quasar_wrapper.scala 136:26]
  assign core_io_ifu_bus_clk_en = io_ifu_bus_clk_en; // @[quasar_wrapper.scala 137:26]
  assign core_io_dbg_bus_clk_en = io_dbg_bus_clk_en; // @[quasar_wrapper.scala 138:26]
  assign core_io_dma_bus_clk_en = io_dma_bus_clk_en; // @[quasar_wrapper.scala 139:26]
  assign core_io_dmi_reg_en = dmi_wrapper_reg_en; // @[quasar_wrapper.scala 79:22]
  assign core_io_dmi_reg_addr = dmi_wrapper_reg_wr_addr; // @[quasar_wrapper.scala 78:24]
  assign core_io_dmi_reg_wr_en = dmi_wrapper_reg_wr_en; // @[quasar_wrapper.scala 80:25]
  assign core_io_dmi_reg_wdata = dmi_wrapper_reg_wr_data; // @[quasar_wrapper.scala 77:25]
  assign core_io_extintsrc_req = io_extintsrc_req; // @[quasar_wrapper.scala 143:25]
  assign core_io_timer_int = io_timer_int; // @[quasar_wrapper.scala 141:21]
  assign core_io_soft_int = io_soft_int; // @[quasar_wrapper.scala 142:20]
  assign core_io_scan_mode = io_scan_mode; // @[quasar_wrapper.scala 66:21]
endmodule
