module el2_ifu_mem_ctl(
  input         clock,
  input         reset,
  input         io_free_clk,
  input         io_active_clk,
  input         io_exu_flush_final,
  input         io_dec_tlu_flush_lower_wb,
  input         io_dec_tlu_flush_err_wb,
  input         io_dec_tlu_i0_commit_cmt,
  input         io_dec_tlu_force_halt,
  input  [30:0] io_ifc_fetch_addr_bf,
  input         io_ifc_fetch_uncacheable_bf,
  input         io_ifc_fetch_req_bf,
  input         io_ifc_fetch_req_bf_raw,
  input         io_ifc_iccm_access_bf,
  input         io_ifc_region_acc_fault_bf,
  input         io_ifc_dma_access_ok,
  input         io_dec_tlu_fence_i_wb,
  input         io_ifu_bp_hit_taken_f,
  input         io_ifu_bp_inst_mask_f,
  input         io_ifu_axi_arready,
  input         io_ifu_axi_rvalid,
  input  [2:0]  io_ifu_axi_rid,
  input  [63:0] io_ifu_axi_rdata,
  input  [1:0]  io_ifu_axi_rresp,
  input         io_ifu_bus_clk_en,
  input         io_dma_iccm_req,
  input  [31:0] io_dma_mem_addr,
  input  [2:0]  io_dma_mem_sz,
  input         io_dma_mem_write,
  input  [63:0] io_dma_mem_wdata,
  input  [2:0]  io_dma_mem_tag,
  input  [63:0] io_ic_rd_data,
  input  [70:0] io_ic_debug_rd_data,
  input  [25:0] io_ictag_debug_rd_data,
  input  [1:0]  io_ic_eccerr,
  input  [1:0]  io_ic_parerr,
  input  [1:0]  io_ic_rd_hit,
  input         io_ic_tag_perr,
  input  [63:0] io_iccm_rd_data,
  input  [77:0] io_iccm_rd_data_ecc,
  input  [1:0]  io_ifu_fetch_val,
  input  [70:0] io_dec_tlu_ic_diag_pkt_icache_wrdata,
  input  [16:0] io_dec_tlu_ic_diag_pkt_icache_dicawics,
  input         io_dec_tlu_ic_diag_pkt_icache_rd_valid,
  input         io_dec_tlu_ic_diag_pkt_icache_wr_valid,
  output        io_ifu_miss_state_idle,
  output        io_ifu_ic_mb_empty,
  output        io_ic_dma_active,
  output        io_ic_write_stall,
  output        io_ifu_pmu_ic_miss,
  output        io_ifu_pmu_ic_hit,
  output        io_ifu_pmu_bus_error,
  output        io_ifu_pmu_bus_busy,
  output        io_ifu_pmu_bus_trxn,
  output        io_ifu_axi_awvalid,
  output [2:0]  io_ifu_axi_awid,
  output [31:0] io_ifu_axi_awaddr,
  output [3:0]  io_ifu_axi_awregion,
  output [7:0]  io_ifu_axi_awlen,
  output [2:0]  io_ifu_axi_awsize,
  output [1:0]  io_ifu_axi_awburst,
  output        io_ifu_axi_awlock,
  output [3:0]  io_ifu_axi_awcache,
  output [2:0]  io_ifu_axi_awprot,
  output [3:0]  io_ifu_axi_awqos,
  output        io_ifu_axi_wvalid,
  output [63:0] io_ifu_axi_wdata,
  output [7:0]  io_ifu_axi_wstrb,
  output        io_ifu_axi_wlast,
  output        io_ifu_axi_bready,
  output        io_ifu_axi_arvalid,
  output [2:0]  io_ifu_axi_arid,
  output [31:0] io_ifu_axi_araddr,
  output [3:0]  io_ifu_axi_arregion,
  output [7:0]  io_ifu_axi_arlen,
  output [2:0]  io_ifu_axi_arsize,
  output [1:0]  io_ifu_axi_arburst,
  output        io_ifu_axi_arlock,
  output [3:0]  io_ifu_axi_arcache,
  output [2:0]  io_ifu_axi_arprot,
  output [3:0]  io_ifu_axi_arqos,
  output        io_ifu_axi_rready,
  output        io_iccm_dma_ecc_error,
  output        io_iccm_dma_rvalid,
  output [63:0] io_iccm_dma_rdata,
  output [2:0]  io_iccm_dma_rtag,
  output        io_iccm_ready,
  output [30:0] io_ic_rw_addr,
  output [1:0]  io_ic_wr_en,
  output        io_ic_rd_en,
  output [70:0] io_ic_wr_data_0,
  output [70:0] io_ic_wr_data_1,
  output [70:0] io_ic_debug_wr_data,
  output [70:0] io_ifu_ic_debug_rd_data,
  output [9:0]  io_ic_debug_addr,
  output        io_ic_debug_rd_en,
  output        io_ic_debug_wr_en,
  output        io_ic_debug_tag_array,
  output [1:0]  io_ic_debug_way,
  output [1:0]  io_ic_tag_valid,
  output [14:0] io_iccm_rw_addr,
  output        io_iccm_wren,
  output        io_iccm_rden,
  output [77:0] io_iccm_wr_data,
  output [2:0]  io_iccm_wr_size,
  output        io_ic_hit_f,
  output        io_ic_access_fault_f,
  output [1:0]  io_ic_access_fault_type_f,
  output        io_iccm_rd_ecc_single_err,
  output        io_iccm_rd_ecc_double_err,
  output        io_ic_error_start,
  output        io_ifu_async_error_start,
  output        io_iccm_dma_sb_error,
  output [1:0]  io_ic_fetch_val_f,
  output [31:0] io_ic_data_f,
  output [63:0] io_ic_premux_data,
  output        io_ic_sel_premux_data,
  input         io_dec_tlu_core_ecc_disable,
  output        io_ifu_ic_debug_rd_data_valid,
  output        io_iccm_buf_correct_ecc,
  output        io_iccm_correction_state,
  input         io_scan_mode,
  output [6:0]  io_test
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [63:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [95:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [63:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [63:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
`endif // RANDOMIZE_REG_INIT
  reg  flush_final_f; // @[el2_ifu_mem_ctl.scala 185:30]
  reg  ifc_fetch_req_f_raw; // @[el2_ifu_mem_ctl.scala 320:36]
  wire  _T_317 = ~io_exu_flush_final; // @[el2_ifu_mem_ctl.scala 321:44]
  wire  ifc_fetch_req_f = ifc_fetch_req_f_raw & _T_317; // @[el2_ifu_mem_ctl.scala 321:42]
  reg [2:0] miss_state; // @[Reg.scala 27:20]
  wire  miss_pending = miss_state != 3'h0; // @[el2_ifu_mem_ctl.scala 253:30]
  reg  scnd_miss_req_q; // @[el2_ifu_mem_ctl.scala 547:52]
  wire  scnd_miss_req = scnd_miss_req_q & _T_317; // @[el2_ifu_mem_ctl.scala 549:36]
  wire  debug_c1_clken = io_ic_debug_rd_en | io_ic_debug_wr_en; // @[el2_ifu_mem_ctl.scala 187:42]
  wire [3:0] ic_fetch_val_int_f = {2'h0,io_ic_fetch_val_f}; // @[Cat.scala 29:58]
  reg [30:0] ifu_fetch_addr_int_f; // @[el2_ifu_mem_ctl.scala 308:34]
  wire [4:0] _GEN_464 = {{1'd0}, ic_fetch_val_int_f}; // @[el2_ifu_mem_ctl.scala 665:53]
  wire [4:0] ic_fetch_val_shift_right = _GEN_464 << ifu_fetch_addr_int_f[0]; // @[el2_ifu_mem_ctl.scala 665:53]
  wire [1:0] _GEN_465 = {{1'd0}, _T_317}; // @[el2_ifu_mem_ctl.scala 668:91]
  wire [1:0] _T_3282 = ic_fetch_val_shift_right[3:2] & _GEN_465; // @[el2_ifu_mem_ctl.scala 668:91]
  reg  ifc_iccm_access_f; // @[el2_ifu_mem_ctl.scala 322:31]
  wire  fetch_req_iccm_f = ifc_fetch_req_f & ifc_iccm_access_f; // @[el2_ifu_mem_ctl.scala 275:46]
  wire [1:0] _GEN_466 = {{1'd0}, fetch_req_iccm_f}; // @[el2_ifu_mem_ctl.scala 668:113]
  wire [1:0] _T_3283 = _T_3282 & _GEN_466; // @[el2_ifu_mem_ctl.scala 668:113]
  reg  iccm_dma_rvalid_in; // @[el2_ifu_mem_ctl.scala 654:59]
  wire [1:0] _GEN_467 = {{1'd0}, iccm_dma_rvalid_in}; // @[el2_ifu_mem_ctl.scala 668:130]
  wire [1:0] _T_3284 = _T_3283 | _GEN_467; // @[el2_ifu_mem_ctl.scala 668:130]
  wire  _T_3285 = ~io_dec_tlu_core_ecc_disable; // @[el2_ifu_mem_ctl.scala 668:154]
  wire [1:0] _GEN_468 = {{1'd0}, _T_3285}; // @[el2_ifu_mem_ctl.scala 668:152]
  wire [1:0] _T_3286 = _T_3284 & _GEN_468; // @[el2_ifu_mem_ctl.scala 668:152]
  wire [1:0] _T_3275 = ic_fetch_val_shift_right[1:0] & _GEN_465; // @[el2_ifu_mem_ctl.scala 668:91]
  wire [1:0] _T_3276 = _T_3275 & _GEN_466; // @[el2_ifu_mem_ctl.scala 668:113]
  wire [1:0] _T_3277 = _T_3276 | _GEN_467; // @[el2_ifu_mem_ctl.scala 668:130]
  wire [1:0] _T_3279 = _T_3277 & _GEN_468; // @[el2_ifu_mem_ctl.scala 668:152]
  wire [3:0] iccm_ecc_word_enable = {_T_3286,_T_3279}; // @[Cat.scala 29:58]
  wire  _T_3386 = ^io_iccm_rd_data_ecc[31:0]; // @[el2_lib.scala 318:30]
  wire  _T_3387 = ^io_iccm_rd_data_ecc[38:32]; // @[el2_lib.scala 318:44]
  wire  _T_3388 = _T_3386 ^ _T_3387; // @[el2_lib.scala 318:35]
  wire [5:0] _T_3396 = {io_iccm_rd_data_ecc[31],io_iccm_rd_data_ecc[30],io_iccm_rd_data_ecc[29],io_iccm_rd_data_ecc[28],io_iccm_rd_data_ecc[27],io_iccm_rd_data_ecc[26]}; // @[el2_lib.scala 318:76]
  wire  _T_3397 = ^_T_3396; // @[el2_lib.scala 318:83]
  wire  _T_3398 = io_iccm_rd_data_ecc[37] ^ _T_3397; // @[el2_lib.scala 318:71]
  wire [6:0] _T_3405 = {io_iccm_rd_data_ecc[17],io_iccm_rd_data_ecc[16],io_iccm_rd_data_ecc[15],io_iccm_rd_data_ecc[14],io_iccm_rd_data_ecc[13],io_iccm_rd_data_ecc[12],io_iccm_rd_data_ecc[11]}; // @[el2_lib.scala 318:103]
  wire [14:0] _T_3413 = {io_iccm_rd_data_ecc[25],io_iccm_rd_data_ecc[24],io_iccm_rd_data_ecc[23],io_iccm_rd_data_ecc[22],io_iccm_rd_data_ecc[21],io_iccm_rd_data_ecc[20],io_iccm_rd_data_ecc[19],io_iccm_rd_data_ecc[18],_T_3405}; // @[el2_lib.scala 318:103]
  wire  _T_3414 = ^_T_3413; // @[el2_lib.scala 318:110]
  wire  _T_3415 = io_iccm_rd_data_ecc[36] ^ _T_3414; // @[el2_lib.scala 318:98]
  wire [6:0] _T_3422 = {io_iccm_rd_data_ecc[10],io_iccm_rd_data_ecc[9],io_iccm_rd_data_ecc[8],io_iccm_rd_data_ecc[7],io_iccm_rd_data_ecc[6],io_iccm_rd_data_ecc[5],io_iccm_rd_data_ecc[4]}; // @[el2_lib.scala 318:130]
  wire [14:0] _T_3430 = {io_iccm_rd_data_ecc[25],io_iccm_rd_data_ecc[24],io_iccm_rd_data_ecc[23],io_iccm_rd_data_ecc[22],io_iccm_rd_data_ecc[21],io_iccm_rd_data_ecc[20],io_iccm_rd_data_ecc[19],io_iccm_rd_data_ecc[18],_T_3422}; // @[el2_lib.scala 318:130]
  wire  _T_3431 = ^_T_3430; // @[el2_lib.scala 318:137]
  wire  _T_3432 = io_iccm_rd_data_ecc[35] ^ _T_3431; // @[el2_lib.scala 318:125]
  wire [8:0] _T_3441 = {io_iccm_rd_data_ecc[15],io_iccm_rd_data_ecc[14],io_iccm_rd_data_ecc[10],io_iccm_rd_data_ecc[9],io_iccm_rd_data_ecc[8],io_iccm_rd_data_ecc[7],io_iccm_rd_data_ecc[3],io_iccm_rd_data_ecc[2],io_iccm_rd_data_ecc[1]}; // @[el2_lib.scala 318:157]
  wire [17:0] _T_3450 = {io_iccm_rd_data_ecc[31],io_iccm_rd_data_ecc[30],io_iccm_rd_data_ecc[29],io_iccm_rd_data_ecc[25],io_iccm_rd_data_ecc[24],io_iccm_rd_data_ecc[23],io_iccm_rd_data_ecc[22],io_iccm_rd_data_ecc[17],io_iccm_rd_data_ecc[16],_T_3441}; // @[el2_lib.scala 318:157]
  wire  _T_3451 = ^_T_3450; // @[el2_lib.scala 318:164]
  wire  _T_3452 = io_iccm_rd_data_ecc[34] ^ _T_3451; // @[el2_lib.scala 318:152]
  wire [8:0] _T_3461 = {io_iccm_rd_data_ecc[13],io_iccm_rd_data_ecc[12],io_iccm_rd_data_ecc[10],io_iccm_rd_data_ecc[9],io_iccm_rd_data_ecc[6],io_iccm_rd_data_ecc[5],io_iccm_rd_data_ecc[3],io_iccm_rd_data_ecc[2],io_iccm_rd_data_ecc[0]}; // @[el2_lib.scala 318:184]
  wire [17:0] _T_3470 = {io_iccm_rd_data_ecc[31],io_iccm_rd_data_ecc[28],io_iccm_rd_data_ecc[27],io_iccm_rd_data_ecc[25],io_iccm_rd_data_ecc[24],io_iccm_rd_data_ecc[21],io_iccm_rd_data_ecc[20],io_iccm_rd_data_ecc[17],io_iccm_rd_data_ecc[16],_T_3461}; // @[el2_lib.scala 318:184]
  wire  _T_3471 = ^_T_3470; // @[el2_lib.scala 318:191]
  wire  _T_3472 = io_iccm_rd_data_ecc[33] ^ _T_3471; // @[el2_lib.scala 318:179]
  wire [8:0] _T_3481 = {io_iccm_rd_data_ecc[13],io_iccm_rd_data_ecc[11],io_iccm_rd_data_ecc[10],io_iccm_rd_data_ecc[8],io_iccm_rd_data_ecc[6],io_iccm_rd_data_ecc[4],io_iccm_rd_data_ecc[3],io_iccm_rd_data_ecc[1],io_iccm_rd_data_ecc[0]}; // @[el2_lib.scala 318:211]
  wire [17:0] _T_3490 = {io_iccm_rd_data_ecc[30],io_iccm_rd_data_ecc[28],io_iccm_rd_data_ecc[26],io_iccm_rd_data_ecc[25],io_iccm_rd_data_ecc[23],io_iccm_rd_data_ecc[21],io_iccm_rd_data_ecc[19],io_iccm_rd_data_ecc[17],io_iccm_rd_data_ecc[15],_T_3481}; // @[el2_lib.scala 318:211]
  wire  _T_3491 = ^_T_3490; // @[el2_lib.scala 318:218]
  wire  _T_3492 = io_iccm_rd_data_ecc[32] ^ _T_3491; // @[el2_lib.scala 318:206]
  wire [6:0] _T_3498 = {_T_3388,_T_3398,_T_3415,_T_3432,_T_3452,_T_3472,_T_3492}; // @[Cat.scala 29:58]
  wire  _T_3499 = _T_3498 != 7'h0; // @[el2_lib.scala 319:44]
  wire  _T_3500 = iccm_ecc_word_enable[0] & _T_3499; // @[el2_lib.scala 319:32]
  wire  _T_3502 = _T_3500 & _T_3498[6]; // @[el2_lib.scala 319:53]
  wire  _T_3771 = ^io_iccm_rd_data_ecc[70:39]; // @[el2_lib.scala 318:30]
  wire  _T_3772 = ^io_iccm_rd_data_ecc[77:71]; // @[el2_lib.scala 318:44]
  wire  _T_3773 = _T_3771 ^ _T_3772; // @[el2_lib.scala 318:35]
  wire [5:0] _T_3781 = {io_iccm_rd_data_ecc[70],io_iccm_rd_data_ecc[69],io_iccm_rd_data_ecc[68],io_iccm_rd_data_ecc[67],io_iccm_rd_data_ecc[66],io_iccm_rd_data_ecc[65]}; // @[el2_lib.scala 318:76]
  wire  _T_3782 = ^_T_3781; // @[el2_lib.scala 318:83]
  wire  _T_3783 = io_iccm_rd_data_ecc[76] ^ _T_3782; // @[el2_lib.scala 318:71]
  wire [6:0] _T_3790 = {io_iccm_rd_data_ecc[56],io_iccm_rd_data_ecc[55],io_iccm_rd_data_ecc[54],io_iccm_rd_data_ecc[53],io_iccm_rd_data_ecc[52],io_iccm_rd_data_ecc[51],io_iccm_rd_data_ecc[50]}; // @[el2_lib.scala 318:103]
  wire [14:0] _T_3798 = {io_iccm_rd_data_ecc[64],io_iccm_rd_data_ecc[63],io_iccm_rd_data_ecc[62],io_iccm_rd_data_ecc[61],io_iccm_rd_data_ecc[60],io_iccm_rd_data_ecc[59],io_iccm_rd_data_ecc[58],io_iccm_rd_data_ecc[57],_T_3790}; // @[el2_lib.scala 318:103]
  wire  _T_3799 = ^_T_3798; // @[el2_lib.scala 318:110]
  wire  _T_3800 = io_iccm_rd_data_ecc[75] ^ _T_3799; // @[el2_lib.scala 318:98]
  wire [6:0] _T_3807 = {io_iccm_rd_data_ecc[49],io_iccm_rd_data_ecc[48],io_iccm_rd_data_ecc[47],io_iccm_rd_data_ecc[46],io_iccm_rd_data_ecc[45],io_iccm_rd_data_ecc[44],io_iccm_rd_data_ecc[43]}; // @[el2_lib.scala 318:130]
  wire [14:0] _T_3815 = {io_iccm_rd_data_ecc[64],io_iccm_rd_data_ecc[63],io_iccm_rd_data_ecc[62],io_iccm_rd_data_ecc[61],io_iccm_rd_data_ecc[60],io_iccm_rd_data_ecc[59],io_iccm_rd_data_ecc[58],io_iccm_rd_data_ecc[57],_T_3807}; // @[el2_lib.scala 318:130]
  wire  _T_3816 = ^_T_3815; // @[el2_lib.scala 318:137]
  wire  _T_3817 = io_iccm_rd_data_ecc[74] ^ _T_3816; // @[el2_lib.scala 318:125]
  wire [8:0] _T_3826 = {io_iccm_rd_data_ecc[54],io_iccm_rd_data_ecc[53],io_iccm_rd_data_ecc[49],io_iccm_rd_data_ecc[48],io_iccm_rd_data_ecc[47],io_iccm_rd_data_ecc[46],io_iccm_rd_data_ecc[42],io_iccm_rd_data_ecc[41],io_iccm_rd_data_ecc[40]}; // @[el2_lib.scala 318:157]
  wire [17:0] _T_3835 = {io_iccm_rd_data_ecc[70],io_iccm_rd_data_ecc[69],io_iccm_rd_data_ecc[68],io_iccm_rd_data_ecc[64],io_iccm_rd_data_ecc[63],io_iccm_rd_data_ecc[62],io_iccm_rd_data_ecc[61],io_iccm_rd_data_ecc[56],io_iccm_rd_data_ecc[55],_T_3826}; // @[el2_lib.scala 318:157]
  wire  _T_3836 = ^_T_3835; // @[el2_lib.scala 318:164]
  wire  _T_3837 = io_iccm_rd_data_ecc[73] ^ _T_3836; // @[el2_lib.scala 318:152]
  wire [8:0] _T_3846 = {io_iccm_rd_data_ecc[52],io_iccm_rd_data_ecc[51],io_iccm_rd_data_ecc[49],io_iccm_rd_data_ecc[48],io_iccm_rd_data_ecc[45],io_iccm_rd_data_ecc[44],io_iccm_rd_data_ecc[42],io_iccm_rd_data_ecc[41],io_iccm_rd_data_ecc[39]}; // @[el2_lib.scala 318:184]
  wire [17:0] _T_3855 = {io_iccm_rd_data_ecc[70],io_iccm_rd_data_ecc[67],io_iccm_rd_data_ecc[66],io_iccm_rd_data_ecc[64],io_iccm_rd_data_ecc[63],io_iccm_rd_data_ecc[60],io_iccm_rd_data_ecc[59],io_iccm_rd_data_ecc[56],io_iccm_rd_data_ecc[55],_T_3846}; // @[el2_lib.scala 318:184]
  wire  _T_3856 = ^_T_3855; // @[el2_lib.scala 318:191]
  wire  _T_3857 = io_iccm_rd_data_ecc[72] ^ _T_3856; // @[el2_lib.scala 318:179]
  wire [8:0] _T_3866 = {io_iccm_rd_data_ecc[52],io_iccm_rd_data_ecc[50],io_iccm_rd_data_ecc[49],io_iccm_rd_data_ecc[47],io_iccm_rd_data_ecc[45],io_iccm_rd_data_ecc[43],io_iccm_rd_data_ecc[42],io_iccm_rd_data_ecc[40],io_iccm_rd_data_ecc[39]}; // @[el2_lib.scala 318:211]
  wire [17:0] _T_3875 = {io_iccm_rd_data_ecc[69],io_iccm_rd_data_ecc[67],io_iccm_rd_data_ecc[65],io_iccm_rd_data_ecc[64],io_iccm_rd_data_ecc[62],io_iccm_rd_data_ecc[60],io_iccm_rd_data_ecc[58],io_iccm_rd_data_ecc[56],io_iccm_rd_data_ecc[54],_T_3866}; // @[el2_lib.scala 318:211]
  wire  _T_3876 = ^_T_3875; // @[el2_lib.scala 318:218]
  wire  _T_3877 = io_iccm_rd_data_ecc[71] ^ _T_3876; // @[el2_lib.scala 318:206]
  wire [6:0] _T_3883 = {_T_3773,_T_3783,_T_3800,_T_3817,_T_3837,_T_3857,_T_3877}; // @[Cat.scala 29:58]
  wire  _T_3884 = _T_3883 != 7'h0; // @[el2_lib.scala 319:44]
  wire  _T_3885 = iccm_ecc_word_enable[1] & _T_3884; // @[el2_lib.scala 319:32]
  wire  _T_3887 = _T_3885 & _T_3883[6]; // @[el2_lib.scala 319:53]
  wire [1:0] iccm_single_ecc_error = {_T_3502,_T_3887}; // @[Cat.scala 29:58]
  wire  _T_3 = |iccm_single_ecc_error; // @[el2_ifu_mem_ctl.scala 190:52]
  reg  dma_iccm_req_f; // @[el2_ifu_mem_ctl.scala 631:51]
  wire  _T_6 = io_iccm_rd_ecc_single_err | io_ic_error_start; // @[el2_ifu_mem_ctl.scala 191:57]
  reg [2:0] perr_state; // @[Reg.scala 27:20]
  wire  _T_7 = perr_state == 3'h4; // @[el2_ifu_mem_ctl.scala 192:54]
  wire  iccm_correct_ecc = perr_state == 3'h3; // @[el2_ifu_mem_ctl.scala 476:34]
  wire  _T_8 = iccm_correct_ecc | _T_7; // @[el2_ifu_mem_ctl.scala 192:40]
  reg [1:0] err_stop_state; // @[Reg.scala 27:20]
  wire  _T_9 = err_stop_state == 2'h3; // @[el2_ifu_mem_ctl.scala 192:90]
  wire  _T_10 = _T_8 | _T_9; // @[el2_ifu_mem_ctl.scala 192:72]
  wire  _T_2490 = 2'h0 == err_stop_state; // @[Conditional.scala 37:30]
  wire  _T_2495 = 2'h1 == err_stop_state; // @[Conditional.scala 37:30]
  wire  _T_2515 = io_ifu_fetch_val == 2'h3; // @[el2_ifu_mem_ctl.scala 526:48]
  wire  two_byte_instr = io_ic_data_f[1:0] != 2'h3; // @[el2_ifu_mem_ctl.scala 390:42]
  wire  _T_2517 = io_ifu_fetch_val[0] & two_byte_instr; // @[el2_ifu_mem_ctl.scala 526:79]
  wire  _T_2518 = _T_2515 | _T_2517; // @[el2_ifu_mem_ctl.scala 526:56]
  wire  _T_2519 = io_exu_flush_final | io_dec_tlu_i0_commit_cmt; // @[el2_ifu_mem_ctl.scala 526:122]
  wire  _T_2520 = ~_T_2519; // @[el2_ifu_mem_ctl.scala 526:101]
  wire  _T_2521 = _T_2518 & _T_2520; // @[el2_ifu_mem_ctl.scala 526:99]
  wire  _T_2522 = 2'h2 == err_stop_state; // @[Conditional.scala 37:30]
  wire  _T_2536 = io_ifu_fetch_val[0] & _T_317; // @[el2_ifu_mem_ctl.scala 533:45]
  wire  _T_2537 = ~io_dec_tlu_i0_commit_cmt; // @[el2_ifu_mem_ctl.scala 533:69]
  wire  _T_2538 = _T_2536 & _T_2537; // @[el2_ifu_mem_ctl.scala 533:67]
  wire  _T_2539 = 2'h3 == err_stop_state; // @[Conditional.scala 37:30]
  wire  _GEN_55 = _T_2522 ? _T_2538 : _T_2539; // @[Conditional.scala 39:67]
  wire  _GEN_59 = _T_2495 ? _T_2521 : _GEN_55; // @[Conditional.scala 39:67]
  wire  err_stop_fetch = _T_2490 ? 1'h0 : _GEN_59; // @[Conditional.scala 40:58]
  wire  _T_11 = _T_10 | err_stop_fetch; // @[el2_ifu_mem_ctl.scala 192:112]
  wire  _T_13 = io_ifu_axi_rvalid & io_ifu_bus_clk_en; // @[el2_ifu_mem_ctl.scala 194:44]
  wire  _T_14 = _T_13 & io_ifu_axi_rready; // @[el2_ifu_mem_ctl.scala 194:65]
  wire  _T_227 = |io_ic_rd_hit; // @[el2_ifu_mem_ctl.scala 283:37]
  wire  _T_228 = ~_T_227; // @[el2_ifu_mem_ctl.scala 283:23]
  reg  reset_all_tags; // @[el2_ifu_mem_ctl.scala 700:53]
  wire  _T_229 = _T_228 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 283:41]
  wire  _T_207 = ~ifc_iccm_access_f; // @[el2_ifu_mem_ctl.scala 274:48]
  wire  _T_208 = ifc_fetch_req_f & _T_207; // @[el2_ifu_mem_ctl.scala 274:46]
  reg  ifc_region_acc_fault_final_f; // @[el2_ifu_mem_ctl.scala 324:42]
  wire  _T_209 = ~ifc_region_acc_fault_final_f; // @[el2_ifu_mem_ctl.scala 274:69]
  wire  fetch_req_icache_f = _T_208 & _T_209; // @[el2_ifu_mem_ctl.scala 274:67]
  wire  _T_230 = _T_229 & fetch_req_icache_f; // @[el2_ifu_mem_ctl.scala 283:59]
  wire  _T_231 = ~miss_pending; // @[el2_ifu_mem_ctl.scala 283:82]
  wire  _T_232 = _T_230 & _T_231; // @[el2_ifu_mem_ctl.scala 283:80]
  wire  _T_233 = _T_232 | scnd_miss_req; // @[el2_ifu_mem_ctl.scala 283:97]
  wire  ic_act_miss_f = _T_233 & _T_209; // @[el2_ifu_mem_ctl.scala 283:114]
  reg  ifu_bus_rvalid_unq_ff; // @[Reg.scala 27:20]
  reg  bus_ifu_bus_clk_en_ff; // @[el2_ifu_mem_ctl.scala 546:61]
  wire  ifu_bus_rvalid_ff = ifu_bus_rvalid_unq_ff & bus_ifu_bus_clk_en_ff; // @[el2_ifu_mem_ctl.scala 588:49]
  wire  bus_ifu_wr_en_ff = ifu_bus_rvalid_ff & miss_pending; // @[el2_ifu_mem_ctl.scala 615:41]
  reg  uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 310:33]
  reg [2:0] bus_data_beat_count; // @[el2_ifu_mem_ctl.scala 596:56]
  wire  _T_2641 = bus_data_beat_count == 3'h1; // @[el2_ifu_mem_ctl.scala 613:69]
  wire  _T_2642 = &bus_data_beat_count; // @[el2_ifu_mem_ctl.scala 613:101]
  wire  bus_last_data_beat = uncacheable_miss_ff ? _T_2641 : _T_2642; // @[el2_ifu_mem_ctl.scala 613:28]
  wire  _T_2588 = bus_ifu_wr_en_ff & bus_last_data_beat; // @[el2_ifu_mem_ctl.scala 592:68]
  wire  _T_2589 = ic_act_miss_f | _T_2588; // @[el2_ifu_mem_ctl.scala 592:48]
  wire  bus_reset_data_beat_cnt = _T_2589 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 592:91]
  wire  _T_2585 = ~bus_last_data_beat; // @[el2_ifu_mem_ctl.scala 591:50]
  wire  _T_2586 = bus_ifu_wr_en_ff & _T_2585; // @[el2_ifu_mem_ctl.scala 591:48]
  wire  _T_2587 = ~io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 591:72]
  wire  bus_inc_data_beat_cnt = _T_2586 & _T_2587; // @[el2_ifu_mem_ctl.scala 591:70]
  wire [2:0] _T_2593 = bus_data_beat_count + 3'h1; // @[el2_ifu_mem_ctl.scala 595:115]
  wire [2:0] _T_2595 = bus_inc_data_beat_cnt ? _T_2593 : 3'h0; // @[Mux.scala 27:72]
  wire  _T_2590 = ~bus_inc_data_beat_cnt; // @[el2_ifu_mem_ctl.scala 593:32]
  wire  _T_2591 = ~bus_reset_data_beat_cnt; // @[el2_ifu_mem_ctl.scala 593:57]
  wire  bus_hold_data_beat_cnt = _T_2590 & _T_2591; // @[el2_ifu_mem_ctl.scala 593:55]
  wire [2:0] _T_2596 = bus_hold_data_beat_cnt ? bus_data_beat_count : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] bus_new_data_beat_count = _T_2595 | _T_2596; // @[Mux.scala 27:72]
  wire  _T_15 = &bus_new_data_beat_count; // @[el2_ifu_mem_ctl.scala 194:112]
  wire  _T_16 = _T_14 & _T_15; // @[el2_ifu_mem_ctl.scala 194:85]
  wire  _T_17 = ~uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 195:5]
  wire  _T_18 = _T_16 & _T_17; // @[el2_ifu_mem_ctl.scala 194:118]
  wire  _T_19 = miss_state == 3'h5; // @[el2_ifu_mem_ctl.scala 195:41]
  wire  _T_24 = 3'h0 == miss_state; // @[Conditional.scala 37:30]
  wire  _T_26 = ic_act_miss_f & _T_317; // @[el2_ifu_mem_ctl.scala 201:43]
  wire [2:0] _T_28 = _T_26 ? 3'h1 : 3'h2; // @[el2_ifu_mem_ctl.scala 201:27]
  wire  _T_31 = 3'h1 == miss_state; // @[Conditional.scala 37:30]
  wire [4:0] byp_fetch_index = ifu_fetch_addr_int_f[4:0]; // @[el2_ifu_mem_ctl.scala 426:45]
  wire  _T_2120 = byp_fetch_index[4:2] == 3'h0; // @[el2_ifu_mem_ctl.scala 447:127]
  reg [7:0] ic_miss_buff_data_valid; // @[el2_ifu_mem_ctl.scala 403:60]
  wire  _T_2151 = _T_2120 & ic_miss_buff_data_valid[0]; // @[Mux.scala 27:72]
  wire  _T_2124 = byp_fetch_index[4:2] == 3'h1; // @[el2_ifu_mem_ctl.scala 447:127]
  wire  _T_2152 = _T_2124 & ic_miss_buff_data_valid[1]; // @[Mux.scala 27:72]
  wire  _T_2159 = _T_2151 | _T_2152; // @[Mux.scala 27:72]
  wire  _T_2128 = byp_fetch_index[4:2] == 3'h2; // @[el2_ifu_mem_ctl.scala 447:127]
  wire  _T_2153 = _T_2128 & ic_miss_buff_data_valid[2]; // @[Mux.scala 27:72]
  wire  _T_2160 = _T_2159 | _T_2153; // @[Mux.scala 27:72]
  wire  _T_2132 = byp_fetch_index[4:2] == 3'h3; // @[el2_ifu_mem_ctl.scala 447:127]
  wire  _T_2154 = _T_2132 & ic_miss_buff_data_valid[3]; // @[Mux.scala 27:72]
  wire  _T_2161 = _T_2160 | _T_2154; // @[Mux.scala 27:72]
  wire  _T_2136 = byp_fetch_index[4:2] == 3'h4; // @[el2_ifu_mem_ctl.scala 447:127]
  wire  _T_2155 = _T_2136 & ic_miss_buff_data_valid[4]; // @[Mux.scala 27:72]
  wire  _T_2162 = _T_2161 | _T_2155; // @[Mux.scala 27:72]
  wire  _T_2140 = byp_fetch_index[4:2] == 3'h5; // @[el2_ifu_mem_ctl.scala 447:127]
  wire  _T_2156 = _T_2140 & ic_miss_buff_data_valid[5]; // @[Mux.scala 27:72]
  wire  _T_2163 = _T_2162 | _T_2156; // @[Mux.scala 27:72]
  wire  _T_2144 = byp_fetch_index[4:2] == 3'h6; // @[el2_ifu_mem_ctl.scala 447:127]
  wire  _T_2157 = _T_2144 & ic_miss_buff_data_valid[6]; // @[Mux.scala 27:72]
  wire  _T_2164 = _T_2163 | _T_2157; // @[Mux.scala 27:72]
  wire  _T_2148 = byp_fetch_index[4:2] == 3'h7; // @[el2_ifu_mem_ctl.scala 447:127]
  wire  _T_2158 = _T_2148 & ic_miss_buff_data_valid[7]; // @[Mux.scala 27:72]
  wire  ic_miss_buff_data_valid_bypass_index = _T_2164 | _T_2158; // @[Mux.scala 27:72]
  wire  _T_2206 = ~byp_fetch_index[1]; // @[el2_ifu_mem_ctl.scala 449:69]
  wire  _T_2207 = ic_miss_buff_data_valid_bypass_index & _T_2206; // @[el2_ifu_mem_ctl.scala 449:67]
  wire  _T_2209 = ~byp_fetch_index[0]; // @[el2_ifu_mem_ctl.scala 449:91]
  wire  _T_2210 = _T_2207 & _T_2209; // @[el2_ifu_mem_ctl.scala 449:89]
  wire  _T_2215 = _T_2207 & byp_fetch_index[0]; // @[el2_ifu_mem_ctl.scala 450:65]
  wire  _T_2216 = _T_2210 | _T_2215; // @[el2_ifu_mem_ctl.scala 449:112]
  wire  _T_2218 = ic_miss_buff_data_valid_bypass_index & byp_fetch_index[1]; // @[el2_ifu_mem_ctl.scala 451:43]
  wire  _T_2221 = _T_2218 & _T_2209; // @[el2_ifu_mem_ctl.scala 451:65]
  wire  _T_2222 = _T_2216 | _T_2221; // @[el2_ifu_mem_ctl.scala 450:88]
  wire  _T_2226 = _T_2218 & byp_fetch_index[0]; // @[el2_ifu_mem_ctl.scala 452:65]
  wire [2:0] byp_fetch_index_inc = ifu_fetch_addr_int_f[4:2] + 3'h1; // @[el2_ifu_mem_ctl.scala 429:75]
  wire  _T_2166 = byp_fetch_index_inc == 3'h0; // @[el2_ifu_mem_ctl.scala 448:110]
  wire  _T_2190 = _T_2166 & ic_miss_buff_data_valid[0]; // @[Mux.scala 27:72]
  wire  _T_2169 = byp_fetch_index_inc == 3'h1; // @[el2_ifu_mem_ctl.scala 448:110]
  wire  _T_2191 = _T_2169 & ic_miss_buff_data_valid[1]; // @[Mux.scala 27:72]
  wire  _T_2198 = _T_2190 | _T_2191; // @[Mux.scala 27:72]
  wire  _T_2172 = byp_fetch_index_inc == 3'h2; // @[el2_ifu_mem_ctl.scala 448:110]
  wire  _T_2192 = _T_2172 & ic_miss_buff_data_valid[2]; // @[Mux.scala 27:72]
  wire  _T_2199 = _T_2198 | _T_2192; // @[Mux.scala 27:72]
  wire  _T_2175 = byp_fetch_index_inc == 3'h3; // @[el2_ifu_mem_ctl.scala 448:110]
  wire  _T_2193 = _T_2175 & ic_miss_buff_data_valid[3]; // @[Mux.scala 27:72]
  wire  _T_2200 = _T_2199 | _T_2193; // @[Mux.scala 27:72]
  wire  _T_2178 = byp_fetch_index_inc == 3'h4; // @[el2_ifu_mem_ctl.scala 448:110]
  wire  _T_2194 = _T_2178 & ic_miss_buff_data_valid[4]; // @[Mux.scala 27:72]
  wire  _T_2201 = _T_2200 | _T_2194; // @[Mux.scala 27:72]
  wire  _T_2181 = byp_fetch_index_inc == 3'h5; // @[el2_ifu_mem_ctl.scala 448:110]
  wire  _T_2195 = _T_2181 & ic_miss_buff_data_valid[5]; // @[Mux.scala 27:72]
  wire  _T_2202 = _T_2201 | _T_2195; // @[Mux.scala 27:72]
  wire  _T_2184 = byp_fetch_index_inc == 3'h6; // @[el2_ifu_mem_ctl.scala 448:110]
  wire  _T_2196 = _T_2184 & ic_miss_buff_data_valid[6]; // @[Mux.scala 27:72]
  wire  _T_2203 = _T_2202 | _T_2196; // @[Mux.scala 27:72]
  wire  _T_2187 = byp_fetch_index_inc == 3'h7; // @[el2_ifu_mem_ctl.scala 448:110]
  wire  _T_2197 = _T_2187 & ic_miss_buff_data_valid[7]; // @[Mux.scala 27:72]
  wire  ic_miss_buff_data_valid_inc_bypass_index = _T_2203 | _T_2197; // @[Mux.scala 27:72]
  wire  _T_2227 = _T_2226 & ic_miss_buff_data_valid_inc_bypass_index; // @[el2_ifu_mem_ctl.scala 452:87]
  wire  _T_2228 = _T_2222 | _T_2227; // @[el2_ifu_mem_ctl.scala 451:88]
  wire  _T_2232 = ic_miss_buff_data_valid_bypass_index & _T_2148; // @[el2_ifu_mem_ctl.scala 453:43]
  wire  miss_buff_hit_unq_f = _T_2228 | _T_2232; // @[el2_ifu_mem_ctl.scala 452:131]
  wire  _T_2248 = miss_state == 3'h4; // @[el2_ifu_mem_ctl.scala 458:55]
  wire  _T_2249 = miss_state == 3'h1; // @[el2_ifu_mem_ctl.scala 458:87]
  wire  _T_2250 = _T_2248 | _T_2249; // @[el2_ifu_mem_ctl.scala 458:74]
  wire  crit_byp_hit_f = miss_buff_hit_unq_f & _T_2250; // @[el2_ifu_mem_ctl.scala 458:41]
  wire  _T_2233 = miss_state == 3'h6; // @[el2_ifu_mem_ctl.scala 455:30]
  reg [30:0] imb_ff; // @[el2_ifu_mem_ctl.scala 311:20]
  wire  miss_wrap_f = imb_ff[5] != ifu_fetch_addr_int_f[5]; // @[el2_ifu_mem_ctl.scala 446:51]
  wire  _T_2234 = ~miss_wrap_f; // @[el2_ifu_mem_ctl.scala 455:68]
  wire  _T_2235 = miss_buff_hit_unq_f & _T_2234; // @[el2_ifu_mem_ctl.scala 455:66]
  wire  stream_hit_f = _T_2233 & _T_2235; // @[el2_ifu_mem_ctl.scala 455:43]
  wire  _T_215 = crit_byp_hit_f | stream_hit_f; // @[el2_ifu_mem_ctl.scala 278:35]
  wire  _T_216 = _T_215 & fetch_req_icache_f; // @[el2_ifu_mem_ctl.scala 278:52]
  wire  ic_byp_hit_f = _T_216 & miss_pending; // @[el2_ifu_mem_ctl.scala 278:73]
  reg  last_data_recieved_ff; // @[el2_ifu_mem_ctl.scala 598:58]
  wire  last_beat = bus_last_data_beat & bus_ifu_wr_en_ff; // @[el2_ifu_mem_ctl.scala 625:35]
  wire  _T_32 = bus_ifu_wr_en_ff & last_beat; // @[el2_ifu_mem_ctl.scala 205:113]
  wire  _T_33 = last_data_recieved_ff | _T_32; // @[el2_ifu_mem_ctl.scala 205:93]
  wire  _T_34 = ic_byp_hit_f & _T_33; // @[el2_ifu_mem_ctl.scala 205:67]
  wire  _T_35 = _T_34 & uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 205:127]
  wire  _T_36 = io_dec_tlu_force_halt | _T_35; // @[el2_ifu_mem_ctl.scala 205:51]
  wire  _T_38 = ~last_data_recieved_ff; // @[el2_ifu_mem_ctl.scala 206:30]
  wire  _T_39 = ic_byp_hit_f & _T_38; // @[el2_ifu_mem_ctl.scala 206:27]
  wire  _T_40 = _T_39 & uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 206:53]
  wire  _T_42 = ~ic_byp_hit_f; // @[el2_ifu_mem_ctl.scala 207:16]
  wire  _T_44 = _T_42 & _T_317; // @[el2_ifu_mem_ctl.scala 207:30]
  wire  _T_46 = _T_44 & _T_32; // @[el2_ifu_mem_ctl.scala 207:52]
  wire  _T_47 = _T_46 & uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 207:85]
  wire  _T_51 = _T_32 & _T_17; // @[el2_ifu_mem_ctl.scala 208:49]
  wire  _T_54 = ic_byp_hit_f & _T_317; // @[el2_ifu_mem_ctl.scala 209:33]
  wire  _T_56 = ~_T_32; // @[el2_ifu_mem_ctl.scala 209:57]
  wire  _T_57 = _T_54 & _T_56; // @[el2_ifu_mem_ctl.scala 209:55]
  wire  ifu_bp_hit_taken_q_f = io_ifu_bp_hit_taken_f & io_ic_hit_f; // @[el2_ifu_mem_ctl.scala 197:52]
  wire  _T_58 = ~ifu_bp_hit_taken_q_f; // @[el2_ifu_mem_ctl.scala 209:91]
  wire  _T_59 = _T_57 & _T_58; // @[el2_ifu_mem_ctl.scala 209:89]
  wire  _T_61 = _T_59 & _T_17; // @[el2_ifu_mem_ctl.scala 209:113]
  wire  _T_64 = bus_ifu_wr_en_ff & _T_317; // @[el2_ifu_mem_ctl.scala 210:39]
  wire  _T_67 = _T_64 & _T_56; // @[el2_ifu_mem_ctl.scala 210:61]
  wire  _T_69 = _T_67 & _T_58; // @[el2_ifu_mem_ctl.scala 210:95]
  wire  _T_71 = _T_69 & _T_17; // @[el2_ifu_mem_ctl.scala 210:119]
  wire  _T_79 = _T_46 & _T_17; // @[el2_ifu_mem_ctl.scala 211:100]
  wire  _T_81 = io_exu_flush_final | ifu_bp_hit_taken_q_f; // @[el2_ifu_mem_ctl.scala 212:44]
  wire  _T_84 = _T_81 & _T_56; // @[el2_ifu_mem_ctl.scala 212:68]
  wire [2:0] _T_86 = _T_84 ? 3'h2 : 3'h0; // @[el2_ifu_mem_ctl.scala 212:22]
  wire [2:0] _T_87 = _T_79 ? 3'h0 : _T_86; // @[el2_ifu_mem_ctl.scala 211:20]
  wire [2:0] _T_88 = _T_71 ? 3'h6 : _T_87; // @[el2_ifu_mem_ctl.scala 210:20]
  wire [2:0] _T_89 = _T_61 ? 3'h6 : _T_88; // @[el2_ifu_mem_ctl.scala 209:18]
  wire [2:0] _T_90 = _T_51 ? 3'h0 : _T_89; // @[el2_ifu_mem_ctl.scala 208:16]
  wire [2:0] _T_91 = _T_47 ? 3'h4 : _T_90; // @[el2_ifu_mem_ctl.scala 207:14]
  wire [2:0] _T_92 = _T_40 ? 3'h3 : _T_91; // @[el2_ifu_mem_ctl.scala 206:12]
  wire [2:0] _T_93 = _T_36 ? 3'h0 : _T_92; // @[el2_ifu_mem_ctl.scala 205:27]
  wire  _T_102 = 3'h4 == miss_state; // @[Conditional.scala 37:30]
  wire  _T_106 = 3'h6 == miss_state; // @[Conditional.scala 37:30]
  wire  _T_2245 = byp_fetch_index[4:1] == 4'hf; // @[el2_ifu_mem_ctl.scala 457:60]
  wire  _T_2246 = _T_2245 & ifc_fetch_req_f; // @[el2_ifu_mem_ctl.scala 457:94]
  wire  stream_eol_f = _T_2246 & stream_hit_f; // @[el2_ifu_mem_ctl.scala 457:112]
  wire  _T_108 = _T_81 | stream_eol_f; // @[el2_ifu_mem_ctl.scala 220:72]
  wire  _T_111 = _T_108 & _T_56; // @[el2_ifu_mem_ctl.scala 220:87]
  wire  _T_113 = _T_111 & _T_2587; // @[el2_ifu_mem_ctl.scala 220:122]
  wire [2:0] _T_115 = _T_113 ? 3'h2 : 3'h0; // @[el2_ifu_mem_ctl.scala 220:27]
  wire  _T_121 = 3'h3 == miss_state; // @[Conditional.scala 37:30]
  wire  _T_124 = io_exu_flush_final & _T_56; // @[el2_ifu_mem_ctl.scala 224:48]
  wire  _T_126 = _T_124 & _T_2587; // @[el2_ifu_mem_ctl.scala 224:82]
  wire [2:0] _T_128 = _T_126 ? 3'h2 : 3'h0; // @[el2_ifu_mem_ctl.scala 224:27]
  wire  _T_132 = 3'h2 == miss_state; // @[Conditional.scala 37:30]
  wire  _T_236 = io_ic_rd_hit == 2'h0; // @[el2_ifu_mem_ctl.scala 284:28]
  wire  _T_237 = _T_236 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 284:42]
  wire  _T_238 = _T_237 & fetch_req_icache_f; // @[el2_ifu_mem_ctl.scala 284:60]
  wire  _T_239 = miss_state == 3'h2; // @[el2_ifu_mem_ctl.scala 284:94]
  wire  _T_240 = _T_238 & _T_239; // @[el2_ifu_mem_ctl.scala 284:81]
  wire  _T_243 = imb_ff[30:5] != ifu_fetch_addr_int_f[30:5]; // @[el2_ifu_mem_ctl.scala 285:39]
  wire  _T_244 = _T_240 & _T_243; // @[el2_ifu_mem_ctl.scala 284:111]
  wire  _T_246 = _T_244 & _T_17; // @[el2_ifu_mem_ctl.scala 285:91]
  reg  sel_mb_addr_ff; // @[el2_ifu_mem_ctl.scala 338:51]
  wire  _T_247 = ~sel_mb_addr_ff; // @[el2_ifu_mem_ctl.scala 285:116]
  wire  _T_248 = _T_246 & _T_247; // @[el2_ifu_mem_ctl.scala 285:114]
  wire  ic_miss_under_miss_f = _T_248 & _T_209; // @[el2_ifu_mem_ctl.scala 285:132]
  wire  _T_135 = ic_miss_under_miss_f & _T_56; // @[el2_ifu_mem_ctl.scala 228:50]
  wire  _T_137 = _T_135 & _T_2587; // @[el2_ifu_mem_ctl.scala 228:84]
  wire  _T_256 = _T_230 & _T_239; // @[el2_ifu_mem_ctl.scala 286:85]
  wire  _T_259 = imb_ff[30:5] == ifu_fetch_addr_int_f[30:5]; // @[el2_ifu_mem_ctl.scala 287:39]
  wire  _T_260 = _T_259 | uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 287:91]
  wire  ic_ignore_2nd_miss_f = _T_256 & _T_260; // @[el2_ifu_mem_ctl.scala 286:117]
  wire  _T_141 = ic_ignore_2nd_miss_f & _T_56; // @[el2_ifu_mem_ctl.scala 229:35]
  wire  _T_143 = _T_141 & _T_2587; // @[el2_ifu_mem_ctl.scala 229:69]
  wire [2:0] _T_145 = _T_143 ? 3'h7 : 3'h0; // @[el2_ifu_mem_ctl.scala 229:12]
  wire [2:0] _T_146 = _T_137 ? 3'h5 : _T_145; // @[el2_ifu_mem_ctl.scala 228:27]
  wire  _T_151 = 3'h5 == miss_state; // @[Conditional.scala 37:30]
  wire [2:0] _T_154 = _T_32 ? 3'h0 : 3'h2; // @[el2_ifu_mem_ctl.scala 234:12]
  wire [2:0] _T_155 = io_exu_flush_final ? _T_154 : 3'h1; // @[el2_ifu_mem_ctl.scala 233:62]
  wire [2:0] _T_156 = io_dec_tlu_force_halt ? 3'h0 : _T_155; // @[el2_ifu_mem_ctl.scala 233:27]
  wire  _T_160 = 3'h7 == miss_state; // @[Conditional.scala 37:30]
  wire [2:0] _T_164 = io_exu_flush_final ? _T_154 : 3'h0; // @[el2_ifu_mem_ctl.scala 238:62]
  wire [2:0] _T_165 = io_dec_tlu_force_halt ? 3'h0 : _T_164; // @[el2_ifu_mem_ctl.scala 238:27]
  wire [2:0] _GEN_0 = _T_160 ? _T_165 : 3'h0; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_2 = _T_151 ? _T_156 : _GEN_0; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_4 = _T_132 ? _T_146 : _GEN_2; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_6 = _T_121 ? _T_128 : _GEN_4; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_8 = _T_106 ? _T_115 : _GEN_6; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_10 = _T_102 ? 3'h0 : _GEN_8; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_12 = _T_31 ? _T_93 : _GEN_10; // @[Conditional.scala 39:67]
  wire [2:0] miss_nxtstate = _T_24 ? _T_28 : _GEN_12; // @[Conditional.scala 40:58]
  wire  _T_20 = miss_nxtstate == 3'h5; // @[el2_ifu_mem_ctl.scala 195:73]
  wire  _T_21 = _T_19 | _T_20; // @[el2_ifu_mem_ctl.scala 195:57]
  wire  _T_22 = _T_18 & _T_21; // @[el2_ifu_mem_ctl.scala 195:26]
  wire  scnd_miss_req_in = _T_22 & _T_317; // @[el2_ifu_mem_ctl.scala 195:91]
  wire  _T_30 = ic_act_miss_f & _T_2587; // @[el2_ifu_mem_ctl.scala 202:38]
  wire  _T_94 = io_dec_tlu_force_halt | io_exu_flush_final; // @[el2_ifu_mem_ctl.scala 213:46]
  wire  _T_95 = _T_94 | ic_byp_hit_f; // @[el2_ifu_mem_ctl.scala 213:67]
  wire  _T_96 = _T_95 | ifu_bp_hit_taken_q_f; // @[el2_ifu_mem_ctl.scala 213:82]
  wire  _T_98 = _T_96 | _T_32; // @[el2_ifu_mem_ctl.scala 213:105]
  wire  _T_100 = bus_ifu_wr_en_ff & _T_17; // @[el2_ifu_mem_ctl.scala 213:158]
  wire  _T_101 = _T_98 | _T_100; // @[el2_ifu_mem_ctl.scala 213:138]
  wire  _T_103 = io_exu_flush_final | flush_final_f; // @[el2_ifu_mem_ctl.scala 217:43]
  wire  _T_104 = _T_103 | ic_byp_hit_f; // @[el2_ifu_mem_ctl.scala 217:59]
  wire  _T_105 = _T_104 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 217:74]
  wire  _T_119 = _T_108 | _T_32; // @[el2_ifu_mem_ctl.scala 221:84]
  wire  _T_120 = _T_119 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 221:118]
  wire  _T_130 = io_exu_flush_final | _T_32; // @[el2_ifu_mem_ctl.scala 225:43]
  wire  _T_131 = _T_130 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 225:76]
  wire  _T_148 = _T_32 | ic_miss_under_miss_f; // @[el2_ifu_mem_ctl.scala 230:55]
  wire  _T_149 = _T_148 | ic_ignore_2nd_miss_f; // @[el2_ifu_mem_ctl.scala 230:78]
  wire  _T_150 = _T_149 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 230:101]
  wire  _T_158 = _T_32 | io_exu_flush_final; // @[el2_ifu_mem_ctl.scala 235:55]
  wire  _T_159 = _T_158 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 235:76]
  wire  _GEN_1 = _T_160 & _T_159; // @[Conditional.scala 39:67]
  wire  _GEN_3 = _T_151 ? _T_159 : _GEN_1; // @[Conditional.scala 39:67]
  wire  _GEN_5 = _T_132 ? _T_150 : _GEN_3; // @[Conditional.scala 39:67]
  wire  _GEN_7 = _T_121 ? _T_131 : _GEN_5; // @[Conditional.scala 39:67]
  wire  _GEN_9 = _T_106 ? _T_120 : _GEN_7; // @[Conditional.scala 39:67]
  wire  _GEN_11 = _T_102 ? _T_105 : _GEN_9; // @[Conditional.scala 39:67]
  wire  _GEN_13 = _T_31 ? _T_101 : _GEN_11; // @[Conditional.scala 39:67]
  wire  miss_state_en = _T_24 ? _T_30 : _GEN_13; // @[Conditional.scala 40:58]
  wire  _T_174 = ~flush_final_f; // @[el2_ifu_mem_ctl.scala 254:95]
  wire  _T_175 = _T_2248 & _T_174; // @[el2_ifu_mem_ctl.scala 254:93]
  wire  crit_wd_byp_ok_ff = _T_2249 | _T_175; // @[el2_ifu_mem_ctl.scala 254:58]
  wire  _T_178 = miss_pending & _T_56; // @[el2_ifu_mem_ctl.scala 255:36]
  wire  _T_180 = _T_2248 & io_exu_flush_final; // @[el2_ifu_mem_ctl.scala 255:106]
  wire  _T_181 = ~_T_180; // @[el2_ifu_mem_ctl.scala 255:72]
  wire  _T_182 = _T_178 & _T_181; // @[el2_ifu_mem_ctl.scala 255:70]
  wire  _T_184 = _T_2248 & crit_byp_hit_f; // @[el2_ifu_mem_ctl.scala 256:57]
  wire  _T_185 = ~_T_184; // @[el2_ifu_mem_ctl.scala 256:23]
  wire  _T_186 = _T_182 & _T_185; // @[el2_ifu_mem_ctl.scala 255:128]
  wire  _T_187 = _T_186 | ic_act_miss_f; // @[el2_ifu_mem_ctl.scala 256:77]
  wire  _T_188 = miss_nxtstate == 3'h4; // @[el2_ifu_mem_ctl.scala 257:36]
  wire  _T_189 = miss_pending & _T_188; // @[el2_ifu_mem_ctl.scala 257:19]
  wire  sel_hold_imb = _T_187 | _T_189; // @[el2_ifu_mem_ctl.scala 256:93]
  wire  _T_191 = _T_19 | ic_miss_under_miss_f; // @[el2_ifu_mem_ctl.scala 259:57]
  wire  sel_hold_imb_scnd = _T_191 & _T_174; // @[el2_ifu_mem_ctl.scala 259:81]
  reg  way_status_mb_scnd_ff; // @[el2_ifu_mem_ctl.scala 267:35]
  reg [6:0] ifu_ic_rw_int_addr_ff; // @[el2_ifu_mem_ctl.scala 734:14]
  wire  _T_4950 = ifu_ic_rw_int_addr_ff == 7'h0; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_0; // @[Reg.scala 27:20]
  wire  _T_5078 = _T_4950 & way_status_out_0; // @[Mux.scala 27:72]
  wire  _T_4951 = ifu_ic_rw_int_addr_ff == 7'h1; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_1; // @[Reg.scala 27:20]
  wire  _T_5079 = _T_4951 & way_status_out_1; // @[Mux.scala 27:72]
  wire  _T_5206 = _T_5078 | _T_5079; // @[Mux.scala 27:72]
  wire  _T_4952 = ifu_ic_rw_int_addr_ff == 7'h2; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_2; // @[Reg.scala 27:20]
  wire  _T_5080 = _T_4952 & way_status_out_2; // @[Mux.scala 27:72]
  wire  _T_5207 = _T_5206 | _T_5080; // @[Mux.scala 27:72]
  wire  _T_4953 = ifu_ic_rw_int_addr_ff == 7'h3; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_3; // @[Reg.scala 27:20]
  wire  _T_5081 = _T_4953 & way_status_out_3; // @[Mux.scala 27:72]
  wire  _T_5208 = _T_5207 | _T_5081; // @[Mux.scala 27:72]
  wire  _T_4954 = ifu_ic_rw_int_addr_ff == 7'h4; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_4; // @[Reg.scala 27:20]
  wire  _T_5082 = _T_4954 & way_status_out_4; // @[Mux.scala 27:72]
  wire  _T_5209 = _T_5208 | _T_5082; // @[Mux.scala 27:72]
  wire  _T_4955 = ifu_ic_rw_int_addr_ff == 7'h5; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_5; // @[Reg.scala 27:20]
  wire  _T_5083 = _T_4955 & way_status_out_5; // @[Mux.scala 27:72]
  wire  _T_5210 = _T_5209 | _T_5083; // @[Mux.scala 27:72]
  wire  _T_4956 = ifu_ic_rw_int_addr_ff == 7'h6; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_6; // @[Reg.scala 27:20]
  wire  _T_5084 = _T_4956 & way_status_out_6; // @[Mux.scala 27:72]
  wire  _T_5211 = _T_5210 | _T_5084; // @[Mux.scala 27:72]
  wire  _T_4957 = ifu_ic_rw_int_addr_ff == 7'h7; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_7; // @[Reg.scala 27:20]
  wire  _T_5085 = _T_4957 & way_status_out_7; // @[Mux.scala 27:72]
  wire  _T_5212 = _T_5211 | _T_5085; // @[Mux.scala 27:72]
  wire  _T_4958 = ifu_ic_rw_int_addr_ff == 7'h8; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_8; // @[Reg.scala 27:20]
  wire  _T_5086 = _T_4958 & way_status_out_8; // @[Mux.scala 27:72]
  wire  _T_5213 = _T_5212 | _T_5086; // @[Mux.scala 27:72]
  wire  _T_4959 = ifu_ic_rw_int_addr_ff == 7'h9; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_9; // @[Reg.scala 27:20]
  wire  _T_5087 = _T_4959 & way_status_out_9; // @[Mux.scala 27:72]
  wire  _T_5214 = _T_5213 | _T_5087; // @[Mux.scala 27:72]
  wire  _T_4960 = ifu_ic_rw_int_addr_ff == 7'ha; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_10; // @[Reg.scala 27:20]
  wire  _T_5088 = _T_4960 & way_status_out_10; // @[Mux.scala 27:72]
  wire  _T_5215 = _T_5214 | _T_5088; // @[Mux.scala 27:72]
  wire  _T_4961 = ifu_ic_rw_int_addr_ff == 7'hb; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_11; // @[Reg.scala 27:20]
  wire  _T_5089 = _T_4961 & way_status_out_11; // @[Mux.scala 27:72]
  wire  _T_5216 = _T_5215 | _T_5089; // @[Mux.scala 27:72]
  wire  _T_4962 = ifu_ic_rw_int_addr_ff == 7'hc; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_12; // @[Reg.scala 27:20]
  wire  _T_5090 = _T_4962 & way_status_out_12; // @[Mux.scala 27:72]
  wire  _T_5217 = _T_5216 | _T_5090; // @[Mux.scala 27:72]
  wire  _T_4963 = ifu_ic_rw_int_addr_ff == 7'hd; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_13; // @[Reg.scala 27:20]
  wire  _T_5091 = _T_4963 & way_status_out_13; // @[Mux.scala 27:72]
  wire  _T_5218 = _T_5217 | _T_5091; // @[Mux.scala 27:72]
  wire  _T_4964 = ifu_ic_rw_int_addr_ff == 7'he; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_14; // @[Reg.scala 27:20]
  wire  _T_5092 = _T_4964 & way_status_out_14; // @[Mux.scala 27:72]
  wire  _T_5219 = _T_5218 | _T_5092; // @[Mux.scala 27:72]
  wire  _T_4965 = ifu_ic_rw_int_addr_ff == 7'hf; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_15; // @[Reg.scala 27:20]
  wire  _T_5093 = _T_4965 & way_status_out_15; // @[Mux.scala 27:72]
  wire  _T_5220 = _T_5219 | _T_5093; // @[Mux.scala 27:72]
  wire  _T_4966 = ifu_ic_rw_int_addr_ff == 7'h10; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_16; // @[Reg.scala 27:20]
  wire  _T_5094 = _T_4966 & way_status_out_16; // @[Mux.scala 27:72]
  wire  _T_5221 = _T_5220 | _T_5094; // @[Mux.scala 27:72]
  wire  _T_4967 = ifu_ic_rw_int_addr_ff == 7'h11; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_17; // @[Reg.scala 27:20]
  wire  _T_5095 = _T_4967 & way_status_out_17; // @[Mux.scala 27:72]
  wire  _T_5222 = _T_5221 | _T_5095; // @[Mux.scala 27:72]
  wire  _T_4968 = ifu_ic_rw_int_addr_ff == 7'h12; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_18; // @[Reg.scala 27:20]
  wire  _T_5096 = _T_4968 & way_status_out_18; // @[Mux.scala 27:72]
  wire  _T_5223 = _T_5222 | _T_5096; // @[Mux.scala 27:72]
  wire  _T_4969 = ifu_ic_rw_int_addr_ff == 7'h13; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_19; // @[Reg.scala 27:20]
  wire  _T_5097 = _T_4969 & way_status_out_19; // @[Mux.scala 27:72]
  wire  _T_5224 = _T_5223 | _T_5097; // @[Mux.scala 27:72]
  wire  _T_4970 = ifu_ic_rw_int_addr_ff == 7'h14; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_20; // @[Reg.scala 27:20]
  wire  _T_5098 = _T_4970 & way_status_out_20; // @[Mux.scala 27:72]
  wire  _T_5225 = _T_5224 | _T_5098; // @[Mux.scala 27:72]
  wire  _T_4971 = ifu_ic_rw_int_addr_ff == 7'h15; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_21; // @[Reg.scala 27:20]
  wire  _T_5099 = _T_4971 & way_status_out_21; // @[Mux.scala 27:72]
  wire  _T_5226 = _T_5225 | _T_5099; // @[Mux.scala 27:72]
  wire  _T_4972 = ifu_ic_rw_int_addr_ff == 7'h16; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_22; // @[Reg.scala 27:20]
  wire  _T_5100 = _T_4972 & way_status_out_22; // @[Mux.scala 27:72]
  wire  _T_5227 = _T_5226 | _T_5100; // @[Mux.scala 27:72]
  wire  _T_4973 = ifu_ic_rw_int_addr_ff == 7'h17; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_23; // @[Reg.scala 27:20]
  wire  _T_5101 = _T_4973 & way_status_out_23; // @[Mux.scala 27:72]
  wire  _T_5228 = _T_5227 | _T_5101; // @[Mux.scala 27:72]
  wire  _T_4974 = ifu_ic_rw_int_addr_ff == 7'h18; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_24; // @[Reg.scala 27:20]
  wire  _T_5102 = _T_4974 & way_status_out_24; // @[Mux.scala 27:72]
  wire  _T_5229 = _T_5228 | _T_5102; // @[Mux.scala 27:72]
  wire  _T_4975 = ifu_ic_rw_int_addr_ff == 7'h19; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_25; // @[Reg.scala 27:20]
  wire  _T_5103 = _T_4975 & way_status_out_25; // @[Mux.scala 27:72]
  wire  _T_5230 = _T_5229 | _T_5103; // @[Mux.scala 27:72]
  wire  _T_4976 = ifu_ic_rw_int_addr_ff == 7'h1a; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_26; // @[Reg.scala 27:20]
  wire  _T_5104 = _T_4976 & way_status_out_26; // @[Mux.scala 27:72]
  wire  _T_5231 = _T_5230 | _T_5104; // @[Mux.scala 27:72]
  wire  _T_4977 = ifu_ic_rw_int_addr_ff == 7'h1b; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_27; // @[Reg.scala 27:20]
  wire  _T_5105 = _T_4977 & way_status_out_27; // @[Mux.scala 27:72]
  wire  _T_5232 = _T_5231 | _T_5105; // @[Mux.scala 27:72]
  wire  _T_4978 = ifu_ic_rw_int_addr_ff == 7'h1c; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_28; // @[Reg.scala 27:20]
  wire  _T_5106 = _T_4978 & way_status_out_28; // @[Mux.scala 27:72]
  wire  _T_5233 = _T_5232 | _T_5106; // @[Mux.scala 27:72]
  wire  _T_4979 = ifu_ic_rw_int_addr_ff == 7'h1d; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_29; // @[Reg.scala 27:20]
  wire  _T_5107 = _T_4979 & way_status_out_29; // @[Mux.scala 27:72]
  wire  _T_5234 = _T_5233 | _T_5107; // @[Mux.scala 27:72]
  wire  _T_4980 = ifu_ic_rw_int_addr_ff == 7'h1e; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_30; // @[Reg.scala 27:20]
  wire  _T_5108 = _T_4980 & way_status_out_30; // @[Mux.scala 27:72]
  wire  _T_5235 = _T_5234 | _T_5108; // @[Mux.scala 27:72]
  wire  _T_4981 = ifu_ic_rw_int_addr_ff == 7'h1f; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_31; // @[Reg.scala 27:20]
  wire  _T_5109 = _T_4981 & way_status_out_31; // @[Mux.scala 27:72]
  wire  _T_5236 = _T_5235 | _T_5109; // @[Mux.scala 27:72]
  wire  _T_4982 = ifu_ic_rw_int_addr_ff == 7'h20; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_32; // @[Reg.scala 27:20]
  wire  _T_5110 = _T_4982 & way_status_out_32; // @[Mux.scala 27:72]
  wire  _T_5237 = _T_5236 | _T_5110; // @[Mux.scala 27:72]
  wire  _T_4983 = ifu_ic_rw_int_addr_ff == 7'h21; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_33; // @[Reg.scala 27:20]
  wire  _T_5111 = _T_4983 & way_status_out_33; // @[Mux.scala 27:72]
  wire  _T_5238 = _T_5237 | _T_5111; // @[Mux.scala 27:72]
  wire  _T_4984 = ifu_ic_rw_int_addr_ff == 7'h22; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_34; // @[Reg.scala 27:20]
  wire  _T_5112 = _T_4984 & way_status_out_34; // @[Mux.scala 27:72]
  wire  _T_5239 = _T_5238 | _T_5112; // @[Mux.scala 27:72]
  wire  _T_4985 = ifu_ic_rw_int_addr_ff == 7'h23; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_35; // @[Reg.scala 27:20]
  wire  _T_5113 = _T_4985 & way_status_out_35; // @[Mux.scala 27:72]
  wire  _T_5240 = _T_5239 | _T_5113; // @[Mux.scala 27:72]
  wire  _T_4986 = ifu_ic_rw_int_addr_ff == 7'h24; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_36; // @[Reg.scala 27:20]
  wire  _T_5114 = _T_4986 & way_status_out_36; // @[Mux.scala 27:72]
  wire  _T_5241 = _T_5240 | _T_5114; // @[Mux.scala 27:72]
  wire  _T_4987 = ifu_ic_rw_int_addr_ff == 7'h25; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_37; // @[Reg.scala 27:20]
  wire  _T_5115 = _T_4987 & way_status_out_37; // @[Mux.scala 27:72]
  wire  _T_5242 = _T_5241 | _T_5115; // @[Mux.scala 27:72]
  wire  _T_4988 = ifu_ic_rw_int_addr_ff == 7'h26; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_38; // @[Reg.scala 27:20]
  wire  _T_5116 = _T_4988 & way_status_out_38; // @[Mux.scala 27:72]
  wire  _T_5243 = _T_5242 | _T_5116; // @[Mux.scala 27:72]
  wire  _T_4989 = ifu_ic_rw_int_addr_ff == 7'h27; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_39; // @[Reg.scala 27:20]
  wire  _T_5117 = _T_4989 & way_status_out_39; // @[Mux.scala 27:72]
  wire  _T_5244 = _T_5243 | _T_5117; // @[Mux.scala 27:72]
  wire  _T_4990 = ifu_ic_rw_int_addr_ff == 7'h28; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_40; // @[Reg.scala 27:20]
  wire  _T_5118 = _T_4990 & way_status_out_40; // @[Mux.scala 27:72]
  wire  _T_5245 = _T_5244 | _T_5118; // @[Mux.scala 27:72]
  wire  _T_4991 = ifu_ic_rw_int_addr_ff == 7'h29; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_41; // @[Reg.scala 27:20]
  wire  _T_5119 = _T_4991 & way_status_out_41; // @[Mux.scala 27:72]
  wire  _T_5246 = _T_5245 | _T_5119; // @[Mux.scala 27:72]
  wire  _T_4992 = ifu_ic_rw_int_addr_ff == 7'h2a; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_42; // @[Reg.scala 27:20]
  wire  _T_5120 = _T_4992 & way_status_out_42; // @[Mux.scala 27:72]
  wire  _T_5247 = _T_5246 | _T_5120; // @[Mux.scala 27:72]
  wire  _T_4993 = ifu_ic_rw_int_addr_ff == 7'h2b; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_43; // @[Reg.scala 27:20]
  wire  _T_5121 = _T_4993 & way_status_out_43; // @[Mux.scala 27:72]
  wire  _T_5248 = _T_5247 | _T_5121; // @[Mux.scala 27:72]
  wire  _T_4994 = ifu_ic_rw_int_addr_ff == 7'h2c; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_44; // @[Reg.scala 27:20]
  wire  _T_5122 = _T_4994 & way_status_out_44; // @[Mux.scala 27:72]
  wire  _T_5249 = _T_5248 | _T_5122; // @[Mux.scala 27:72]
  wire  _T_4995 = ifu_ic_rw_int_addr_ff == 7'h2d; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_45; // @[Reg.scala 27:20]
  wire  _T_5123 = _T_4995 & way_status_out_45; // @[Mux.scala 27:72]
  wire  _T_5250 = _T_5249 | _T_5123; // @[Mux.scala 27:72]
  wire  _T_4996 = ifu_ic_rw_int_addr_ff == 7'h2e; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_46; // @[Reg.scala 27:20]
  wire  _T_5124 = _T_4996 & way_status_out_46; // @[Mux.scala 27:72]
  wire  _T_5251 = _T_5250 | _T_5124; // @[Mux.scala 27:72]
  wire  _T_4997 = ifu_ic_rw_int_addr_ff == 7'h2f; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_47; // @[Reg.scala 27:20]
  wire  _T_5125 = _T_4997 & way_status_out_47; // @[Mux.scala 27:72]
  wire  _T_5252 = _T_5251 | _T_5125; // @[Mux.scala 27:72]
  wire  _T_4998 = ifu_ic_rw_int_addr_ff == 7'h30; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_48; // @[Reg.scala 27:20]
  wire  _T_5126 = _T_4998 & way_status_out_48; // @[Mux.scala 27:72]
  wire  _T_5253 = _T_5252 | _T_5126; // @[Mux.scala 27:72]
  wire  _T_4999 = ifu_ic_rw_int_addr_ff == 7'h31; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_49; // @[Reg.scala 27:20]
  wire  _T_5127 = _T_4999 & way_status_out_49; // @[Mux.scala 27:72]
  wire  _T_5254 = _T_5253 | _T_5127; // @[Mux.scala 27:72]
  wire  _T_5000 = ifu_ic_rw_int_addr_ff == 7'h32; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_50; // @[Reg.scala 27:20]
  wire  _T_5128 = _T_5000 & way_status_out_50; // @[Mux.scala 27:72]
  wire  _T_5255 = _T_5254 | _T_5128; // @[Mux.scala 27:72]
  wire  _T_5001 = ifu_ic_rw_int_addr_ff == 7'h33; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_51; // @[Reg.scala 27:20]
  wire  _T_5129 = _T_5001 & way_status_out_51; // @[Mux.scala 27:72]
  wire  _T_5256 = _T_5255 | _T_5129; // @[Mux.scala 27:72]
  wire  _T_5002 = ifu_ic_rw_int_addr_ff == 7'h34; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_52; // @[Reg.scala 27:20]
  wire  _T_5130 = _T_5002 & way_status_out_52; // @[Mux.scala 27:72]
  wire  _T_5257 = _T_5256 | _T_5130; // @[Mux.scala 27:72]
  wire  _T_5003 = ifu_ic_rw_int_addr_ff == 7'h35; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_53; // @[Reg.scala 27:20]
  wire  _T_5131 = _T_5003 & way_status_out_53; // @[Mux.scala 27:72]
  wire  _T_5258 = _T_5257 | _T_5131; // @[Mux.scala 27:72]
  wire  _T_5004 = ifu_ic_rw_int_addr_ff == 7'h36; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_54; // @[Reg.scala 27:20]
  wire  _T_5132 = _T_5004 & way_status_out_54; // @[Mux.scala 27:72]
  wire  _T_5259 = _T_5258 | _T_5132; // @[Mux.scala 27:72]
  wire  _T_5005 = ifu_ic_rw_int_addr_ff == 7'h37; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_55; // @[Reg.scala 27:20]
  wire  _T_5133 = _T_5005 & way_status_out_55; // @[Mux.scala 27:72]
  wire  _T_5260 = _T_5259 | _T_5133; // @[Mux.scala 27:72]
  wire  _T_5006 = ifu_ic_rw_int_addr_ff == 7'h38; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_56; // @[Reg.scala 27:20]
  wire  _T_5134 = _T_5006 & way_status_out_56; // @[Mux.scala 27:72]
  wire  _T_5261 = _T_5260 | _T_5134; // @[Mux.scala 27:72]
  wire  _T_5007 = ifu_ic_rw_int_addr_ff == 7'h39; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_57; // @[Reg.scala 27:20]
  wire  _T_5135 = _T_5007 & way_status_out_57; // @[Mux.scala 27:72]
  wire  _T_5262 = _T_5261 | _T_5135; // @[Mux.scala 27:72]
  wire  _T_5008 = ifu_ic_rw_int_addr_ff == 7'h3a; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_58; // @[Reg.scala 27:20]
  wire  _T_5136 = _T_5008 & way_status_out_58; // @[Mux.scala 27:72]
  wire  _T_5263 = _T_5262 | _T_5136; // @[Mux.scala 27:72]
  wire  _T_5009 = ifu_ic_rw_int_addr_ff == 7'h3b; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_59; // @[Reg.scala 27:20]
  wire  _T_5137 = _T_5009 & way_status_out_59; // @[Mux.scala 27:72]
  wire  _T_5264 = _T_5263 | _T_5137; // @[Mux.scala 27:72]
  wire  _T_5010 = ifu_ic_rw_int_addr_ff == 7'h3c; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_60; // @[Reg.scala 27:20]
  wire  _T_5138 = _T_5010 & way_status_out_60; // @[Mux.scala 27:72]
  wire  _T_5265 = _T_5264 | _T_5138; // @[Mux.scala 27:72]
  wire  _T_5011 = ifu_ic_rw_int_addr_ff == 7'h3d; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_61; // @[Reg.scala 27:20]
  wire  _T_5139 = _T_5011 & way_status_out_61; // @[Mux.scala 27:72]
  wire  _T_5266 = _T_5265 | _T_5139; // @[Mux.scala 27:72]
  wire  _T_5012 = ifu_ic_rw_int_addr_ff == 7'h3e; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_62; // @[Reg.scala 27:20]
  wire  _T_5140 = _T_5012 & way_status_out_62; // @[Mux.scala 27:72]
  wire  _T_5267 = _T_5266 | _T_5140; // @[Mux.scala 27:72]
  wire  _T_5013 = ifu_ic_rw_int_addr_ff == 7'h3f; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_63; // @[Reg.scala 27:20]
  wire  _T_5141 = _T_5013 & way_status_out_63; // @[Mux.scala 27:72]
  wire  _T_5268 = _T_5267 | _T_5141; // @[Mux.scala 27:72]
  wire  _T_5014 = ifu_ic_rw_int_addr_ff == 7'h40; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_64; // @[Reg.scala 27:20]
  wire  _T_5142 = _T_5014 & way_status_out_64; // @[Mux.scala 27:72]
  wire  _T_5269 = _T_5268 | _T_5142; // @[Mux.scala 27:72]
  wire  _T_5015 = ifu_ic_rw_int_addr_ff == 7'h41; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_65; // @[Reg.scala 27:20]
  wire  _T_5143 = _T_5015 & way_status_out_65; // @[Mux.scala 27:72]
  wire  _T_5270 = _T_5269 | _T_5143; // @[Mux.scala 27:72]
  wire  _T_5016 = ifu_ic_rw_int_addr_ff == 7'h42; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_66; // @[Reg.scala 27:20]
  wire  _T_5144 = _T_5016 & way_status_out_66; // @[Mux.scala 27:72]
  wire  _T_5271 = _T_5270 | _T_5144; // @[Mux.scala 27:72]
  wire  _T_5017 = ifu_ic_rw_int_addr_ff == 7'h43; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_67; // @[Reg.scala 27:20]
  wire  _T_5145 = _T_5017 & way_status_out_67; // @[Mux.scala 27:72]
  wire  _T_5272 = _T_5271 | _T_5145; // @[Mux.scala 27:72]
  wire  _T_5018 = ifu_ic_rw_int_addr_ff == 7'h44; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_68; // @[Reg.scala 27:20]
  wire  _T_5146 = _T_5018 & way_status_out_68; // @[Mux.scala 27:72]
  wire  _T_5273 = _T_5272 | _T_5146; // @[Mux.scala 27:72]
  wire  _T_5019 = ifu_ic_rw_int_addr_ff == 7'h45; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_69; // @[Reg.scala 27:20]
  wire  _T_5147 = _T_5019 & way_status_out_69; // @[Mux.scala 27:72]
  wire  _T_5274 = _T_5273 | _T_5147; // @[Mux.scala 27:72]
  wire  _T_5020 = ifu_ic_rw_int_addr_ff == 7'h46; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_70; // @[Reg.scala 27:20]
  wire  _T_5148 = _T_5020 & way_status_out_70; // @[Mux.scala 27:72]
  wire  _T_5275 = _T_5274 | _T_5148; // @[Mux.scala 27:72]
  wire  _T_5021 = ifu_ic_rw_int_addr_ff == 7'h47; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_71; // @[Reg.scala 27:20]
  wire  _T_5149 = _T_5021 & way_status_out_71; // @[Mux.scala 27:72]
  wire  _T_5276 = _T_5275 | _T_5149; // @[Mux.scala 27:72]
  wire  _T_5022 = ifu_ic_rw_int_addr_ff == 7'h48; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_72; // @[Reg.scala 27:20]
  wire  _T_5150 = _T_5022 & way_status_out_72; // @[Mux.scala 27:72]
  wire  _T_5277 = _T_5276 | _T_5150; // @[Mux.scala 27:72]
  wire  _T_5023 = ifu_ic_rw_int_addr_ff == 7'h49; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_73; // @[Reg.scala 27:20]
  wire  _T_5151 = _T_5023 & way_status_out_73; // @[Mux.scala 27:72]
  wire  _T_5278 = _T_5277 | _T_5151; // @[Mux.scala 27:72]
  wire  _T_5024 = ifu_ic_rw_int_addr_ff == 7'h4a; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_74; // @[Reg.scala 27:20]
  wire  _T_5152 = _T_5024 & way_status_out_74; // @[Mux.scala 27:72]
  wire  _T_5279 = _T_5278 | _T_5152; // @[Mux.scala 27:72]
  wire  _T_5025 = ifu_ic_rw_int_addr_ff == 7'h4b; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_75; // @[Reg.scala 27:20]
  wire  _T_5153 = _T_5025 & way_status_out_75; // @[Mux.scala 27:72]
  wire  _T_5280 = _T_5279 | _T_5153; // @[Mux.scala 27:72]
  wire  _T_5026 = ifu_ic_rw_int_addr_ff == 7'h4c; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_76; // @[Reg.scala 27:20]
  wire  _T_5154 = _T_5026 & way_status_out_76; // @[Mux.scala 27:72]
  wire  _T_5281 = _T_5280 | _T_5154; // @[Mux.scala 27:72]
  wire  _T_5027 = ifu_ic_rw_int_addr_ff == 7'h4d; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_77; // @[Reg.scala 27:20]
  wire  _T_5155 = _T_5027 & way_status_out_77; // @[Mux.scala 27:72]
  wire  _T_5282 = _T_5281 | _T_5155; // @[Mux.scala 27:72]
  wire  _T_5028 = ifu_ic_rw_int_addr_ff == 7'h4e; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_78; // @[Reg.scala 27:20]
  wire  _T_5156 = _T_5028 & way_status_out_78; // @[Mux.scala 27:72]
  wire  _T_5283 = _T_5282 | _T_5156; // @[Mux.scala 27:72]
  wire  _T_5029 = ifu_ic_rw_int_addr_ff == 7'h4f; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_79; // @[Reg.scala 27:20]
  wire  _T_5157 = _T_5029 & way_status_out_79; // @[Mux.scala 27:72]
  wire  _T_5284 = _T_5283 | _T_5157; // @[Mux.scala 27:72]
  wire  _T_5030 = ifu_ic_rw_int_addr_ff == 7'h50; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_80; // @[Reg.scala 27:20]
  wire  _T_5158 = _T_5030 & way_status_out_80; // @[Mux.scala 27:72]
  wire  _T_5285 = _T_5284 | _T_5158; // @[Mux.scala 27:72]
  wire  _T_5031 = ifu_ic_rw_int_addr_ff == 7'h51; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_81; // @[Reg.scala 27:20]
  wire  _T_5159 = _T_5031 & way_status_out_81; // @[Mux.scala 27:72]
  wire  _T_5286 = _T_5285 | _T_5159; // @[Mux.scala 27:72]
  wire  _T_5032 = ifu_ic_rw_int_addr_ff == 7'h52; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_82; // @[Reg.scala 27:20]
  wire  _T_5160 = _T_5032 & way_status_out_82; // @[Mux.scala 27:72]
  wire  _T_5287 = _T_5286 | _T_5160; // @[Mux.scala 27:72]
  wire  _T_5033 = ifu_ic_rw_int_addr_ff == 7'h53; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_83; // @[Reg.scala 27:20]
  wire  _T_5161 = _T_5033 & way_status_out_83; // @[Mux.scala 27:72]
  wire  _T_5288 = _T_5287 | _T_5161; // @[Mux.scala 27:72]
  wire  _T_5034 = ifu_ic_rw_int_addr_ff == 7'h54; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_84; // @[Reg.scala 27:20]
  wire  _T_5162 = _T_5034 & way_status_out_84; // @[Mux.scala 27:72]
  wire  _T_5289 = _T_5288 | _T_5162; // @[Mux.scala 27:72]
  wire  _T_5035 = ifu_ic_rw_int_addr_ff == 7'h55; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_85; // @[Reg.scala 27:20]
  wire  _T_5163 = _T_5035 & way_status_out_85; // @[Mux.scala 27:72]
  wire  _T_5290 = _T_5289 | _T_5163; // @[Mux.scala 27:72]
  wire  _T_5036 = ifu_ic_rw_int_addr_ff == 7'h56; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_86; // @[Reg.scala 27:20]
  wire  _T_5164 = _T_5036 & way_status_out_86; // @[Mux.scala 27:72]
  wire  _T_5291 = _T_5290 | _T_5164; // @[Mux.scala 27:72]
  wire  _T_5037 = ifu_ic_rw_int_addr_ff == 7'h57; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_87; // @[Reg.scala 27:20]
  wire  _T_5165 = _T_5037 & way_status_out_87; // @[Mux.scala 27:72]
  wire  _T_5292 = _T_5291 | _T_5165; // @[Mux.scala 27:72]
  wire  _T_5038 = ifu_ic_rw_int_addr_ff == 7'h58; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_88; // @[Reg.scala 27:20]
  wire  _T_5166 = _T_5038 & way_status_out_88; // @[Mux.scala 27:72]
  wire  _T_5293 = _T_5292 | _T_5166; // @[Mux.scala 27:72]
  wire  _T_5039 = ifu_ic_rw_int_addr_ff == 7'h59; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_89; // @[Reg.scala 27:20]
  wire  _T_5167 = _T_5039 & way_status_out_89; // @[Mux.scala 27:72]
  wire  _T_5294 = _T_5293 | _T_5167; // @[Mux.scala 27:72]
  wire  _T_5040 = ifu_ic_rw_int_addr_ff == 7'h5a; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_90; // @[Reg.scala 27:20]
  wire  _T_5168 = _T_5040 & way_status_out_90; // @[Mux.scala 27:72]
  wire  _T_5295 = _T_5294 | _T_5168; // @[Mux.scala 27:72]
  wire  _T_5041 = ifu_ic_rw_int_addr_ff == 7'h5b; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_91; // @[Reg.scala 27:20]
  wire  _T_5169 = _T_5041 & way_status_out_91; // @[Mux.scala 27:72]
  wire  _T_5296 = _T_5295 | _T_5169; // @[Mux.scala 27:72]
  wire  _T_5042 = ifu_ic_rw_int_addr_ff == 7'h5c; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_92; // @[Reg.scala 27:20]
  wire  _T_5170 = _T_5042 & way_status_out_92; // @[Mux.scala 27:72]
  wire  _T_5297 = _T_5296 | _T_5170; // @[Mux.scala 27:72]
  wire  _T_5043 = ifu_ic_rw_int_addr_ff == 7'h5d; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_93; // @[Reg.scala 27:20]
  wire  _T_5171 = _T_5043 & way_status_out_93; // @[Mux.scala 27:72]
  wire  _T_5298 = _T_5297 | _T_5171; // @[Mux.scala 27:72]
  wire  _T_5044 = ifu_ic_rw_int_addr_ff == 7'h5e; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_94; // @[Reg.scala 27:20]
  wire  _T_5172 = _T_5044 & way_status_out_94; // @[Mux.scala 27:72]
  wire  _T_5299 = _T_5298 | _T_5172; // @[Mux.scala 27:72]
  wire  _T_5045 = ifu_ic_rw_int_addr_ff == 7'h5f; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_95; // @[Reg.scala 27:20]
  wire  _T_5173 = _T_5045 & way_status_out_95; // @[Mux.scala 27:72]
  wire  _T_5300 = _T_5299 | _T_5173; // @[Mux.scala 27:72]
  wire  _T_5046 = ifu_ic_rw_int_addr_ff == 7'h60; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_96; // @[Reg.scala 27:20]
  wire  _T_5174 = _T_5046 & way_status_out_96; // @[Mux.scala 27:72]
  wire  _T_5301 = _T_5300 | _T_5174; // @[Mux.scala 27:72]
  wire  _T_5047 = ifu_ic_rw_int_addr_ff == 7'h61; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_97; // @[Reg.scala 27:20]
  wire  _T_5175 = _T_5047 & way_status_out_97; // @[Mux.scala 27:72]
  wire  _T_5302 = _T_5301 | _T_5175; // @[Mux.scala 27:72]
  wire  _T_5048 = ifu_ic_rw_int_addr_ff == 7'h62; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_98; // @[Reg.scala 27:20]
  wire  _T_5176 = _T_5048 & way_status_out_98; // @[Mux.scala 27:72]
  wire  _T_5303 = _T_5302 | _T_5176; // @[Mux.scala 27:72]
  wire  _T_5049 = ifu_ic_rw_int_addr_ff == 7'h63; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_99; // @[Reg.scala 27:20]
  wire  _T_5177 = _T_5049 & way_status_out_99; // @[Mux.scala 27:72]
  wire  _T_5304 = _T_5303 | _T_5177; // @[Mux.scala 27:72]
  wire  _T_5050 = ifu_ic_rw_int_addr_ff == 7'h64; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_100; // @[Reg.scala 27:20]
  wire  _T_5178 = _T_5050 & way_status_out_100; // @[Mux.scala 27:72]
  wire  _T_5305 = _T_5304 | _T_5178; // @[Mux.scala 27:72]
  wire  _T_5051 = ifu_ic_rw_int_addr_ff == 7'h65; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_101; // @[Reg.scala 27:20]
  wire  _T_5179 = _T_5051 & way_status_out_101; // @[Mux.scala 27:72]
  wire  _T_5306 = _T_5305 | _T_5179; // @[Mux.scala 27:72]
  wire  _T_5052 = ifu_ic_rw_int_addr_ff == 7'h66; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_102; // @[Reg.scala 27:20]
  wire  _T_5180 = _T_5052 & way_status_out_102; // @[Mux.scala 27:72]
  wire  _T_5307 = _T_5306 | _T_5180; // @[Mux.scala 27:72]
  wire  _T_5053 = ifu_ic_rw_int_addr_ff == 7'h67; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_103; // @[Reg.scala 27:20]
  wire  _T_5181 = _T_5053 & way_status_out_103; // @[Mux.scala 27:72]
  wire  _T_5308 = _T_5307 | _T_5181; // @[Mux.scala 27:72]
  wire  _T_5054 = ifu_ic_rw_int_addr_ff == 7'h68; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_104; // @[Reg.scala 27:20]
  wire  _T_5182 = _T_5054 & way_status_out_104; // @[Mux.scala 27:72]
  wire  _T_5309 = _T_5308 | _T_5182; // @[Mux.scala 27:72]
  wire  _T_5055 = ifu_ic_rw_int_addr_ff == 7'h69; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_105; // @[Reg.scala 27:20]
  wire  _T_5183 = _T_5055 & way_status_out_105; // @[Mux.scala 27:72]
  wire  _T_5310 = _T_5309 | _T_5183; // @[Mux.scala 27:72]
  wire  _T_5056 = ifu_ic_rw_int_addr_ff == 7'h6a; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_106; // @[Reg.scala 27:20]
  wire  _T_5184 = _T_5056 & way_status_out_106; // @[Mux.scala 27:72]
  wire  _T_5311 = _T_5310 | _T_5184; // @[Mux.scala 27:72]
  wire  _T_5057 = ifu_ic_rw_int_addr_ff == 7'h6b; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_107; // @[Reg.scala 27:20]
  wire  _T_5185 = _T_5057 & way_status_out_107; // @[Mux.scala 27:72]
  wire  _T_5312 = _T_5311 | _T_5185; // @[Mux.scala 27:72]
  wire  _T_5058 = ifu_ic_rw_int_addr_ff == 7'h6c; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_108; // @[Reg.scala 27:20]
  wire  _T_5186 = _T_5058 & way_status_out_108; // @[Mux.scala 27:72]
  wire  _T_5313 = _T_5312 | _T_5186; // @[Mux.scala 27:72]
  wire  _T_5059 = ifu_ic_rw_int_addr_ff == 7'h6d; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_109; // @[Reg.scala 27:20]
  wire  _T_5187 = _T_5059 & way_status_out_109; // @[Mux.scala 27:72]
  wire  _T_5314 = _T_5313 | _T_5187; // @[Mux.scala 27:72]
  wire  _T_5060 = ifu_ic_rw_int_addr_ff == 7'h6e; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_110; // @[Reg.scala 27:20]
  wire  _T_5188 = _T_5060 & way_status_out_110; // @[Mux.scala 27:72]
  wire  _T_5315 = _T_5314 | _T_5188; // @[Mux.scala 27:72]
  wire  _T_5061 = ifu_ic_rw_int_addr_ff == 7'h6f; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_111; // @[Reg.scala 27:20]
  wire  _T_5189 = _T_5061 & way_status_out_111; // @[Mux.scala 27:72]
  wire  _T_5316 = _T_5315 | _T_5189; // @[Mux.scala 27:72]
  wire  _T_5062 = ifu_ic_rw_int_addr_ff == 7'h70; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_112; // @[Reg.scala 27:20]
  wire  _T_5190 = _T_5062 & way_status_out_112; // @[Mux.scala 27:72]
  wire  _T_5317 = _T_5316 | _T_5190; // @[Mux.scala 27:72]
  wire  _T_5063 = ifu_ic_rw_int_addr_ff == 7'h71; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_113; // @[Reg.scala 27:20]
  wire  _T_5191 = _T_5063 & way_status_out_113; // @[Mux.scala 27:72]
  wire  _T_5318 = _T_5317 | _T_5191; // @[Mux.scala 27:72]
  wire  _T_5064 = ifu_ic_rw_int_addr_ff == 7'h72; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_114; // @[Reg.scala 27:20]
  wire  _T_5192 = _T_5064 & way_status_out_114; // @[Mux.scala 27:72]
  wire  _T_5319 = _T_5318 | _T_5192; // @[Mux.scala 27:72]
  wire  _T_5065 = ifu_ic_rw_int_addr_ff == 7'h73; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_115; // @[Reg.scala 27:20]
  wire  _T_5193 = _T_5065 & way_status_out_115; // @[Mux.scala 27:72]
  wire  _T_5320 = _T_5319 | _T_5193; // @[Mux.scala 27:72]
  wire  _T_5066 = ifu_ic_rw_int_addr_ff == 7'h74; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_116; // @[Reg.scala 27:20]
  wire  _T_5194 = _T_5066 & way_status_out_116; // @[Mux.scala 27:72]
  wire  _T_5321 = _T_5320 | _T_5194; // @[Mux.scala 27:72]
  wire  _T_5067 = ifu_ic_rw_int_addr_ff == 7'h75; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_117; // @[Reg.scala 27:20]
  wire  _T_5195 = _T_5067 & way_status_out_117; // @[Mux.scala 27:72]
  wire  _T_5322 = _T_5321 | _T_5195; // @[Mux.scala 27:72]
  wire  _T_5068 = ifu_ic_rw_int_addr_ff == 7'h76; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_118; // @[Reg.scala 27:20]
  wire  _T_5196 = _T_5068 & way_status_out_118; // @[Mux.scala 27:72]
  wire  _T_5323 = _T_5322 | _T_5196; // @[Mux.scala 27:72]
  wire  _T_5069 = ifu_ic_rw_int_addr_ff == 7'h77; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_119; // @[Reg.scala 27:20]
  wire  _T_5197 = _T_5069 & way_status_out_119; // @[Mux.scala 27:72]
  wire  _T_5324 = _T_5323 | _T_5197; // @[Mux.scala 27:72]
  wire  _T_5070 = ifu_ic_rw_int_addr_ff == 7'h78; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_120; // @[Reg.scala 27:20]
  wire  _T_5198 = _T_5070 & way_status_out_120; // @[Mux.scala 27:72]
  wire  _T_5325 = _T_5324 | _T_5198; // @[Mux.scala 27:72]
  wire  _T_5071 = ifu_ic_rw_int_addr_ff == 7'h79; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_121; // @[Reg.scala 27:20]
  wire  _T_5199 = _T_5071 & way_status_out_121; // @[Mux.scala 27:72]
  wire  _T_5326 = _T_5325 | _T_5199; // @[Mux.scala 27:72]
  wire  _T_5072 = ifu_ic_rw_int_addr_ff == 7'h7a; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_122; // @[Reg.scala 27:20]
  wire  _T_5200 = _T_5072 & way_status_out_122; // @[Mux.scala 27:72]
  wire  _T_5327 = _T_5326 | _T_5200; // @[Mux.scala 27:72]
  wire  _T_5073 = ifu_ic_rw_int_addr_ff == 7'h7b; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_123; // @[Reg.scala 27:20]
  wire  _T_5201 = _T_5073 & way_status_out_123; // @[Mux.scala 27:72]
  wire  _T_5328 = _T_5327 | _T_5201; // @[Mux.scala 27:72]
  wire  _T_5074 = ifu_ic_rw_int_addr_ff == 7'h7c; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_124; // @[Reg.scala 27:20]
  wire  _T_5202 = _T_5074 & way_status_out_124; // @[Mux.scala 27:72]
  wire  _T_5329 = _T_5328 | _T_5202; // @[Mux.scala 27:72]
  wire  _T_5075 = ifu_ic_rw_int_addr_ff == 7'h7d; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_125; // @[Reg.scala 27:20]
  wire  _T_5203 = _T_5075 & way_status_out_125; // @[Mux.scala 27:72]
  wire  _T_5330 = _T_5329 | _T_5203; // @[Mux.scala 27:72]
  wire  _T_5076 = ifu_ic_rw_int_addr_ff == 7'h7e; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_126; // @[Reg.scala 27:20]
  wire  _T_5204 = _T_5076 & way_status_out_126; // @[Mux.scala 27:72]
  wire  _T_5331 = _T_5330 | _T_5204; // @[Mux.scala 27:72]
  wire  _T_5077 = ifu_ic_rw_int_addr_ff == 7'h7f; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_127; // @[Reg.scala 27:20]
  wire  _T_5205 = _T_5077 & way_status_out_127; // @[Mux.scala 27:72]
  wire  way_status = _T_5331 | _T_5205; // @[Mux.scala 27:72]
  wire  _T_195 = ~reset_all_tags; // @[el2_ifu_mem_ctl.scala 262:96]
  wire [1:0] _T_197 = _T_195 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [1:0] _T_198 = _T_197 & io_ic_tag_valid; // @[el2_ifu_mem_ctl.scala 262:113]
  reg [1:0] tagv_mb_scnd_ff; // @[el2_ifu_mem_ctl.scala 268:29]
  reg  uncacheable_miss_scnd_ff; // @[el2_ifu_mem_ctl.scala 264:38]
  reg [30:0] imb_scnd_ff; // @[el2_ifu_mem_ctl.scala 266:25]
  wire [2:0] _T_206 = bus_ifu_wr_en_ff ? 3'h7 : 3'h0; // @[Bitwise.scala 72:12]
  reg [2:0] ifu_bus_rid_ff; // @[Reg.scala 27:20]
  wire [2:0] ic_wr_addr_bits_hi_3 = ifu_bus_rid_ff & _T_206; // @[el2_ifu_mem_ctl.scala 271:45]
  wire  _T_212 = _T_231 | _T_239; // @[el2_ifu_mem_ctl.scala 276:59]
  wire  _T_214 = _T_212 | _T_2233; // @[el2_ifu_mem_ctl.scala 276:91]
  wire  ic_iccm_hit_f = fetch_req_iccm_f & _T_214; // @[el2_ifu_mem_ctl.scala 276:41]
  wire  _T_219 = _T_227 & fetch_req_icache_f; // @[el2_ifu_mem_ctl.scala 282:39]
  wire  _T_221 = _T_219 & _T_195; // @[el2_ifu_mem_ctl.scala 282:60]
  wire  _T_225 = _T_221 & _T_212; // @[el2_ifu_mem_ctl.scala 282:78]
  wire  ic_act_hit_f = _T_225 & _T_247; // @[el2_ifu_mem_ctl.scala 282:126]
  wire  _T_262 = ic_act_hit_f | ic_byp_hit_f; // @[el2_ifu_mem_ctl.scala 289:31]
  wire  _T_263 = _T_262 | ic_iccm_hit_f; // @[el2_ifu_mem_ctl.scala 289:46]
  wire  _T_264 = ifc_region_acc_fault_final_f & ifc_fetch_req_f; // @[el2_ifu_mem_ctl.scala 289:94]
  wire  _T_268 = sel_hold_imb ? uncacheable_miss_ff : io_ifc_fetch_uncacheable_bf; // @[el2_ifu_mem_ctl.scala 290:84]
  wire  uncacheable_miss_in = scnd_miss_req ? uncacheable_miss_scnd_ff : _T_268; // @[el2_ifu_mem_ctl.scala 290:32]
  wire  _T_274 = imb_ff[11:5] == imb_scnd_ff[11:5]; // @[el2_ifu_mem_ctl.scala 293:79]
  wire  _T_275 = _T_274 & scnd_miss_req; // @[el2_ifu_mem_ctl.scala 293:135]
  reg [1:0] ifu_bus_rresp_ff; // @[Reg.scala 27:20]
  wire  _T_2662 = |ifu_bus_rresp_ff; // @[el2_ifu_mem_ctl.scala 621:48]
  wire  _T_2663 = _T_2662 & ifu_bus_rvalid_ff; // @[el2_ifu_mem_ctl.scala 621:52]
  wire  bus_ifu_wr_data_error_ff = _T_2663 & miss_pending; // @[el2_ifu_mem_ctl.scala 621:73]
  reg  ifu_wr_data_comb_err_ff; // @[el2_ifu_mem_ctl.scala 366:61]
  wire  ifu_wr_cumulative_err_data = bus_ifu_wr_data_error_ff | ifu_wr_data_comb_err_ff; // @[el2_ifu_mem_ctl.scala 365:55]
  wire  _T_276 = ~ifu_wr_cumulative_err_data; // @[el2_ifu_mem_ctl.scala 293:153]
  wire  scnd_miss_index_match = _T_275 & _T_276; // @[el2_ifu_mem_ctl.scala 293:151]
  wire  _T_277 = ~scnd_miss_index_match; // @[el2_ifu_mem_ctl.scala 296:47]
  wire  _T_278 = scnd_miss_req & _T_277; // @[el2_ifu_mem_ctl.scala 296:45]
  wire  _T_280 = scnd_miss_req & scnd_miss_index_match; // @[el2_ifu_mem_ctl.scala 297:26]
  reg  way_status_mb_ff; // @[el2_ifu_mem_ctl.scala 316:30]
  wire  _T_10539 = ~way_status_mb_ff; // @[el2_ifu_mem_ctl.scala 786:33]
  reg [1:0] tagv_mb_ff; // @[el2_ifu_mem_ctl.scala 317:24]
  wire  _T_10541 = _T_10539 & tagv_mb_ff[0]; // @[el2_ifu_mem_ctl.scala 786:51]
  wire  _T_10543 = _T_10541 & tagv_mb_ff[1]; // @[el2_ifu_mem_ctl.scala 786:67]
  wire  _T_10545 = ~tagv_mb_ff[0]; // @[el2_ifu_mem_ctl.scala 786:86]
  wire  replace_way_mb_any_0 = _T_10543 | _T_10545; // @[el2_ifu_mem_ctl.scala 786:84]
  wire [1:0] _T_287 = scnd_miss_index_match ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire  _T_10548 = way_status_mb_ff & tagv_mb_ff[0]; // @[el2_ifu_mem_ctl.scala 787:50]
  wire  _T_10550 = _T_10548 & tagv_mb_ff[1]; // @[el2_ifu_mem_ctl.scala 787:66]
  wire  _T_10552 = ~tagv_mb_ff[1]; // @[el2_ifu_mem_ctl.scala 787:85]
  wire  _T_10554 = _T_10552 & tagv_mb_ff[0]; // @[el2_ifu_mem_ctl.scala 787:100]
  wire  replace_way_mb_any_1 = _T_10550 | _T_10554; // @[el2_ifu_mem_ctl.scala 787:83]
  wire [1:0] _T_288 = {replace_way_mb_any_1,replace_way_mb_any_0}; // @[Cat.scala 29:58]
  wire [1:0] _T_289 = _T_287 & _T_288; // @[el2_ifu_mem_ctl.scala 301:110]
  wire [1:0] _T_290 = tagv_mb_scnd_ff | _T_289; // @[el2_ifu_mem_ctl.scala 301:62]
  wire [1:0] _T_295 = io_ic_tag_valid & _T_197; // @[el2_ifu_mem_ctl.scala 302:56]
  wire  _T_297 = ~scnd_miss_req_q; // @[el2_ifu_mem_ctl.scala 305:36]
  wire  _T_298 = miss_pending & _T_297; // @[el2_ifu_mem_ctl.scala 305:34]
  reg  reset_ic_ff; // @[el2_ifu_mem_ctl.scala 306:25]
  wire  _T_299 = reset_all_tags | reset_ic_ff; // @[el2_ifu_mem_ctl.scala 305:72]
  wire  reset_ic_in = _T_298 & _T_299; // @[el2_ifu_mem_ctl.scala 305:53]
  reg  fetch_uncacheable_ff; // @[el2_ifu_mem_ctl.scala 307:37]
  reg [25:0] miss_addr; // @[el2_ifu_mem_ctl.scala 315:23]
  wire  _T_313 = _T_2248 & flush_final_f; // @[el2_ifu_mem_ctl.scala 319:87]
  wire  _T_314 = ~_T_313; // @[el2_ifu_mem_ctl.scala 319:55]
  wire  _T_315 = io_ifc_fetch_req_bf & _T_314; // @[el2_ifu_mem_ctl.scala 319:53]
  wire  _T_2240 = ~_T_2235; // @[el2_ifu_mem_ctl.scala 456:46]
  wire  _T_2241 = _T_2233 & _T_2240; // @[el2_ifu_mem_ctl.scala 456:44]
  wire  stream_miss_f = _T_2241 & ifc_fetch_req_f; // @[el2_ifu_mem_ctl.scala 456:84]
  wire  _T_316 = ~stream_miss_f; // @[el2_ifu_mem_ctl.scala 319:106]
  wire  ifc_fetch_req_qual_bf = _T_315 & _T_316; // @[el2_ifu_mem_ctl.scala 319:104]
  reg  ifc_region_acc_fault_f; // @[el2_ifu_mem_ctl.scala 325:39]
  reg [2:0] bus_rd_addr_count; // @[Reg.scala 27:20]
  wire [28:0] ifu_ic_req_addr_f = {miss_addr,bus_rd_addr_count}; // @[Cat.scala 29:58]
  wire  _T_323 = _T_239 | _T_2233; // @[el2_ifu_mem_ctl.scala 327:55]
  wire  _T_326 = _T_323 & _T_56; // @[el2_ifu_mem_ctl.scala 327:82]
  wire  _T_2254 = ~ifu_bus_rid_ff[0]; // @[el2_ifu_mem_ctl.scala 461:55]
  wire [2:0] other_tag = {ifu_bus_rid_ff[2:1],_T_2254}; // @[Cat.scala 29:58]
  wire  _T_2255 = other_tag == 3'h0; // @[el2_ifu_mem_ctl.scala 462:81]
  wire  _T_2279 = _T_2255 & ic_miss_buff_data_valid[0]; // @[Mux.scala 27:72]
  wire  _T_2258 = other_tag == 3'h1; // @[el2_ifu_mem_ctl.scala 462:81]
  wire  _T_2280 = _T_2258 & ic_miss_buff_data_valid[1]; // @[Mux.scala 27:72]
  wire  _T_2287 = _T_2279 | _T_2280; // @[Mux.scala 27:72]
  wire  _T_2261 = other_tag == 3'h2; // @[el2_ifu_mem_ctl.scala 462:81]
  wire  _T_2281 = _T_2261 & ic_miss_buff_data_valid[2]; // @[Mux.scala 27:72]
  wire  _T_2288 = _T_2287 | _T_2281; // @[Mux.scala 27:72]
  wire  _T_2264 = other_tag == 3'h3; // @[el2_ifu_mem_ctl.scala 462:81]
  wire  _T_2282 = _T_2264 & ic_miss_buff_data_valid[3]; // @[Mux.scala 27:72]
  wire  _T_2289 = _T_2288 | _T_2282; // @[Mux.scala 27:72]
  wire  _T_2267 = other_tag == 3'h4; // @[el2_ifu_mem_ctl.scala 462:81]
  wire  _T_2283 = _T_2267 & ic_miss_buff_data_valid[4]; // @[Mux.scala 27:72]
  wire  _T_2290 = _T_2289 | _T_2283; // @[Mux.scala 27:72]
  wire  _T_2270 = other_tag == 3'h5; // @[el2_ifu_mem_ctl.scala 462:81]
  wire  _T_2284 = _T_2270 & ic_miss_buff_data_valid[5]; // @[Mux.scala 27:72]
  wire  _T_2291 = _T_2290 | _T_2284; // @[Mux.scala 27:72]
  wire  _T_2273 = other_tag == 3'h6; // @[el2_ifu_mem_ctl.scala 462:81]
  wire  _T_2285 = _T_2273 & ic_miss_buff_data_valid[6]; // @[Mux.scala 27:72]
  wire  _T_2292 = _T_2291 | _T_2285; // @[Mux.scala 27:72]
  wire  _T_2276 = other_tag == 3'h7; // @[el2_ifu_mem_ctl.scala 462:81]
  wire  _T_2286 = _T_2276 & ic_miss_buff_data_valid[7]; // @[Mux.scala 27:72]
  wire  second_half_available = _T_2292 | _T_2286; // @[Mux.scala 27:72]
  wire  write_ic_16_bytes = second_half_available & bus_ifu_wr_en_ff; // @[el2_ifu_mem_ctl.scala 463:46]
  wire  _T_330 = miss_pending & write_ic_16_bytes; // @[el2_ifu_mem_ctl.scala 331:35]
  wire  _T_332 = _T_330 & _T_17; // @[el2_ifu_mem_ctl.scala 331:55]
  reg  ic_act_miss_f_delayed; // @[el2_ifu_mem_ctl.scala 618:61]
  wire  _T_2656 = ic_act_miss_f_delayed & _T_2249; // @[el2_ifu_mem_ctl.scala 619:53]
  wire  reset_tag_valid_for_miss = _T_2656 & _T_17; // @[el2_ifu_mem_ctl.scala 619:84]
  wire  sel_mb_addr = _T_332 | reset_tag_valid_for_miss; // @[el2_ifu_mem_ctl.scala 331:79]
  wire [30:0] _T_336 = {imb_ff[30:5],ic_wr_addr_bits_hi_3,imb_ff[1:0]}; // @[Cat.scala 29:58]
  wire  _T_337 = ~sel_mb_addr; // @[el2_ifu_mem_ctl.scala 333:37]
  wire [30:0] _T_338 = sel_mb_addr ? _T_336 : 31'h0; // @[Mux.scala 27:72]
  wire [30:0] _T_339 = _T_337 ? io_ifc_fetch_addr_bf : 31'h0; // @[Mux.scala 27:72]
  wire [30:0] ifu_ic_rw_int_addr = _T_338 | _T_339; // @[Mux.scala 27:72]
  wire  _T_344 = _T_332 & last_beat; // @[el2_ifu_mem_ctl.scala 335:84]
  wire  _T_2650 = ~_T_2662; // @[el2_ifu_mem_ctl.scala 616:84]
  wire  _T_2651 = _T_100 & _T_2650; // @[el2_ifu_mem_ctl.scala 616:82]
  wire  bus_ifu_wr_en_ff_q = _T_2651 & write_ic_16_bytes; // @[el2_ifu_mem_ctl.scala 616:108]
  wire  sel_mb_status_addr = _T_344 & bus_ifu_wr_en_ff_q; // @[el2_ifu_mem_ctl.scala 335:96]
  wire [30:0] ifu_status_wr_addr = sel_mb_status_addr ? _T_336 : ifu_fetch_addr_int_f; // @[el2_ifu_mem_ctl.scala 336:31]
  reg [63:0] ifu_bus_rdata_ff; // @[Reg.scala 27:20]
  wire [6:0] _T_567 = {ifu_bus_rdata_ff[63],ifu_bus_rdata_ff[62],ifu_bus_rdata_ff[61],ifu_bus_rdata_ff[60],ifu_bus_rdata_ff[59],ifu_bus_rdata_ff[58],ifu_bus_rdata_ff[57]}; // @[el2_lib.scala 401:13]
  wire  _T_568 = ^_T_567; // @[el2_lib.scala 401:20]
  wire [6:0] _T_574 = {ifu_bus_rdata_ff[32],ifu_bus_rdata_ff[31],ifu_bus_rdata_ff[30],ifu_bus_rdata_ff[29],ifu_bus_rdata_ff[28],ifu_bus_rdata_ff[27],ifu_bus_rdata_ff[26]}; // @[el2_lib.scala 401:30]
  wire [7:0] _T_581 = {ifu_bus_rdata_ff[40],ifu_bus_rdata_ff[39],ifu_bus_rdata_ff[38],ifu_bus_rdata_ff[37],ifu_bus_rdata_ff[36],ifu_bus_rdata_ff[35],ifu_bus_rdata_ff[34],ifu_bus_rdata_ff[33]}; // @[el2_lib.scala 401:30]
  wire [14:0] _T_582 = {ifu_bus_rdata_ff[40],ifu_bus_rdata_ff[39],ifu_bus_rdata_ff[38],ifu_bus_rdata_ff[37],ifu_bus_rdata_ff[36],ifu_bus_rdata_ff[35],ifu_bus_rdata_ff[34],ifu_bus_rdata_ff[33],_T_574}; // @[el2_lib.scala 401:30]
  wire [7:0] _T_589 = {ifu_bus_rdata_ff[48],ifu_bus_rdata_ff[47],ifu_bus_rdata_ff[46],ifu_bus_rdata_ff[45],ifu_bus_rdata_ff[44],ifu_bus_rdata_ff[43],ifu_bus_rdata_ff[42],ifu_bus_rdata_ff[41]}; // @[el2_lib.scala 401:30]
  wire [30:0] _T_598 = {ifu_bus_rdata_ff[56],ifu_bus_rdata_ff[55],ifu_bus_rdata_ff[54],ifu_bus_rdata_ff[53],ifu_bus_rdata_ff[52],ifu_bus_rdata_ff[51],ifu_bus_rdata_ff[50],ifu_bus_rdata_ff[49],_T_589,_T_582}; // @[el2_lib.scala 401:30]
  wire  _T_599 = ^_T_598; // @[el2_lib.scala 401:37]
  wire [6:0] _T_605 = {ifu_bus_rdata_ff[17],ifu_bus_rdata_ff[16],ifu_bus_rdata_ff[15],ifu_bus_rdata_ff[14],ifu_bus_rdata_ff[13],ifu_bus_rdata_ff[12],ifu_bus_rdata_ff[11]}; // @[el2_lib.scala 401:47]
  wire [14:0] _T_613 = {ifu_bus_rdata_ff[25],ifu_bus_rdata_ff[24],ifu_bus_rdata_ff[23],ifu_bus_rdata_ff[22],ifu_bus_rdata_ff[21],ifu_bus_rdata_ff[20],ifu_bus_rdata_ff[19],ifu_bus_rdata_ff[18],_T_605}; // @[el2_lib.scala 401:47]
  wire [30:0] _T_629 = {ifu_bus_rdata_ff[56],ifu_bus_rdata_ff[55],ifu_bus_rdata_ff[54],ifu_bus_rdata_ff[53],ifu_bus_rdata_ff[52],ifu_bus_rdata_ff[51],ifu_bus_rdata_ff[50],ifu_bus_rdata_ff[49],_T_589,_T_613}; // @[el2_lib.scala 401:47]
  wire  _T_630 = ^_T_629; // @[el2_lib.scala 401:54]
  wire [6:0] _T_636 = {ifu_bus_rdata_ff[10],ifu_bus_rdata_ff[9],ifu_bus_rdata_ff[8],ifu_bus_rdata_ff[7],ifu_bus_rdata_ff[6],ifu_bus_rdata_ff[5],ifu_bus_rdata_ff[4]}; // @[el2_lib.scala 401:64]
  wire [14:0] _T_644 = {ifu_bus_rdata_ff[25],ifu_bus_rdata_ff[24],ifu_bus_rdata_ff[23],ifu_bus_rdata_ff[22],ifu_bus_rdata_ff[21],ifu_bus_rdata_ff[20],ifu_bus_rdata_ff[19],ifu_bus_rdata_ff[18],_T_636}; // @[el2_lib.scala 401:64]
  wire [30:0] _T_660 = {ifu_bus_rdata_ff[56],ifu_bus_rdata_ff[55],ifu_bus_rdata_ff[54],ifu_bus_rdata_ff[53],ifu_bus_rdata_ff[52],ifu_bus_rdata_ff[51],ifu_bus_rdata_ff[50],ifu_bus_rdata_ff[49],_T_581,_T_644}; // @[el2_lib.scala 401:64]
  wire  _T_661 = ^_T_660; // @[el2_lib.scala 401:71]
  wire [7:0] _T_668 = {ifu_bus_rdata_ff[14],ifu_bus_rdata_ff[10],ifu_bus_rdata_ff[9],ifu_bus_rdata_ff[8],ifu_bus_rdata_ff[7],ifu_bus_rdata_ff[3],ifu_bus_rdata_ff[2],ifu_bus_rdata_ff[1]}; // @[el2_lib.scala 401:81]
  wire [16:0] _T_677 = {ifu_bus_rdata_ff[30],ifu_bus_rdata_ff[29],ifu_bus_rdata_ff[25],ifu_bus_rdata_ff[24],ifu_bus_rdata_ff[23],ifu_bus_rdata_ff[22],ifu_bus_rdata_ff[17],ifu_bus_rdata_ff[16],ifu_bus_rdata_ff[15],_T_668}; // @[el2_lib.scala 401:81]
  wire [8:0] _T_685 = {ifu_bus_rdata_ff[47],ifu_bus_rdata_ff[46],ifu_bus_rdata_ff[45],ifu_bus_rdata_ff[40],ifu_bus_rdata_ff[39],ifu_bus_rdata_ff[38],ifu_bus_rdata_ff[37],ifu_bus_rdata_ff[32],ifu_bus_rdata_ff[31]}; // @[el2_lib.scala 401:81]
  wire [17:0] _T_694 = {ifu_bus_rdata_ff[63],ifu_bus_rdata_ff[62],ifu_bus_rdata_ff[61],ifu_bus_rdata_ff[60],ifu_bus_rdata_ff[56],ifu_bus_rdata_ff[55],ifu_bus_rdata_ff[54],ifu_bus_rdata_ff[53],ifu_bus_rdata_ff[48],_T_685}; // @[el2_lib.scala 401:81]
  wire [34:0] _T_695 = {_T_694,_T_677}; // @[el2_lib.scala 401:81]
  wire  _T_696 = ^_T_695; // @[el2_lib.scala 401:88]
  wire [7:0] _T_703 = {ifu_bus_rdata_ff[12],ifu_bus_rdata_ff[10],ifu_bus_rdata_ff[9],ifu_bus_rdata_ff[6],ifu_bus_rdata_ff[5],ifu_bus_rdata_ff[3],ifu_bus_rdata_ff[2],ifu_bus_rdata_ff[0]}; // @[el2_lib.scala 401:98]
  wire [16:0] _T_712 = {ifu_bus_rdata_ff[28],ifu_bus_rdata_ff[27],ifu_bus_rdata_ff[25],ifu_bus_rdata_ff[24],ifu_bus_rdata_ff[21],ifu_bus_rdata_ff[20],ifu_bus_rdata_ff[17],ifu_bus_rdata_ff[16],ifu_bus_rdata_ff[13],_T_703}; // @[el2_lib.scala 401:98]
  wire [8:0] _T_720 = {ifu_bus_rdata_ff[47],ifu_bus_rdata_ff[44],ifu_bus_rdata_ff[43],ifu_bus_rdata_ff[40],ifu_bus_rdata_ff[39],ifu_bus_rdata_ff[36],ifu_bus_rdata_ff[35],ifu_bus_rdata_ff[32],ifu_bus_rdata_ff[31]}; // @[el2_lib.scala 401:98]
  wire [17:0] _T_729 = {ifu_bus_rdata_ff[63],ifu_bus_rdata_ff[62],ifu_bus_rdata_ff[59],ifu_bus_rdata_ff[58],ifu_bus_rdata_ff[56],ifu_bus_rdata_ff[55],ifu_bus_rdata_ff[52],ifu_bus_rdata_ff[51],ifu_bus_rdata_ff[48],_T_720}; // @[el2_lib.scala 401:98]
  wire [34:0] _T_730 = {_T_729,_T_712}; // @[el2_lib.scala 401:98]
  wire  _T_731 = ^_T_730; // @[el2_lib.scala 401:105]
  wire [7:0] _T_738 = {ifu_bus_rdata_ff[11],ifu_bus_rdata_ff[10],ifu_bus_rdata_ff[8],ifu_bus_rdata_ff[6],ifu_bus_rdata_ff[4],ifu_bus_rdata_ff[3],ifu_bus_rdata_ff[1],ifu_bus_rdata_ff[0]}; // @[el2_lib.scala 401:115]
  wire [16:0] _T_747 = {ifu_bus_rdata_ff[28],ifu_bus_rdata_ff[26],ifu_bus_rdata_ff[25],ifu_bus_rdata_ff[23],ifu_bus_rdata_ff[21],ifu_bus_rdata_ff[19],ifu_bus_rdata_ff[17],ifu_bus_rdata_ff[15],ifu_bus_rdata_ff[13],_T_738}; // @[el2_lib.scala 401:115]
  wire [8:0] _T_755 = {ifu_bus_rdata_ff[46],ifu_bus_rdata_ff[44],ifu_bus_rdata_ff[42],ifu_bus_rdata_ff[40],ifu_bus_rdata_ff[38],ifu_bus_rdata_ff[36],ifu_bus_rdata_ff[34],ifu_bus_rdata_ff[32],ifu_bus_rdata_ff[30]}; // @[el2_lib.scala 401:115]
  wire [17:0] _T_764 = {ifu_bus_rdata_ff[63],ifu_bus_rdata_ff[61],ifu_bus_rdata_ff[59],ifu_bus_rdata_ff[57],ifu_bus_rdata_ff[56],ifu_bus_rdata_ff[54],ifu_bus_rdata_ff[52],ifu_bus_rdata_ff[50],ifu_bus_rdata_ff[48],_T_755}; // @[el2_lib.scala 401:115]
  wire [34:0] _T_765 = {_T_764,_T_747}; // @[el2_lib.scala 401:115]
  wire  _T_766 = ^_T_765; // @[el2_lib.scala 401:122]
  wire [3:0] _T_2295 = {ifu_bus_rid_ff[2:1],_T_2254,1'h1}; // @[Cat.scala 29:58]
  wire  _T_2296 = _T_2295 == 4'h0; // @[el2_ifu_mem_ctl.scala 464:89]
  reg [31:0] ic_miss_buff_data_0; // @[Reg.scala 27:20]
  wire [31:0] _T_2343 = _T_2296 ? ic_miss_buff_data_0 : 32'h0; // @[Mux.scala 27:72]
  wire  _T_2299 = _T_2295 == 4'h1; // @[el2_ifu_mem_ctl.scala 464:89]
  reg [31:0] ic_miss_buff_data_1; // @[Reg.scala 27:20]
  wire [31:0] _T_2344 = _T_2299 ? ic_miss_buff_data_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2359 = _T_2343 | _T_2344; // @[Mux.scala 27:72]
  wire  _T_2302 = _T_2295 == 4'h2; // @[el2_ifu_mem_ctl.scala 464:89]
  reg [31:0] ic_miss_buff_data_2; // @[Reg.scala 27:20]
  wire [31:0] _T_2345 = _T_2302 ? ic_miss_buff_data_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2360 = _T_2359 | _T_2345; // @[Mux.scala 27:72]
  wire  _T_2305 = _T_2295 == 4'h3; // @[el2_ifu_mem_ctl.scala 464:89]
  reg [31:0] ic_miss_buff_data_3; // @[Reg.scala 27:20]
  wire [31:0] _T_2346 = _T_2305 ? ic_miss_buff_data_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2361 = _T_2360 | _T_2346; // @[Mux.scala 27:72]
  wire  _T_2308 = _T_2295 == 4'h4; // @[el2_ifu_mem_ctl.scala 464:89]
  reg [31:0] ic_miss_buff_data_4; // @[Reg.scala 27:20]
  wire [31:0] _T_2347 = _T_2308 ? ic_miss_buff_data_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2362 = _T_2361 | _T_2347; // @[Mux.scala 27:72]
  wire  _T_2311 = _T_2295 == 4'h5; // @[el2_ifu_mem_ctl.scala 464:89]
  reg [31:0] ic_miss_buff_data_5; // @[Reg.scala 27:20]
  wire [31:0] _T_2348 = _T_2311 ? ic_miss_buff_data_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2363 = _T_2362 | _T_2348; // @[Mux.scala 27:72]
  wire  _T_2314 = _T_2295 == 4'h6; // @[el2_ifu_mem_ctl.scala 464:89]
  reg [31:0] ic_miss_buff_data_6; // @[Reg.scala 27:20]
  wire [31:0] _T_2349 = _T_2314 ? ic_miss_buff_data_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2364 = _T_2363 | _T_2349; // @[Mux.scala 27:72]
  wire  _T_2317 = _T_2295 == 4'h7; // @[el2_ifu_mem_ctl.scala 464:89]
  reg [31:0] ic_miss_buff_data_7; // @[Reg.scala 27:20]
  wire [31:0] _T_2350 = _T_2317 ? ic_miss_buff_data_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2365 = _T_2364 | _T_2350; // @[Mux.scala 27:72]
  wire  _T_2320 = _T_2295 == 4'h8; // @[el2_ifu_mem_ctl.scala 464:89]
  reg [31:0] ic_miss_buff_data_8; // @[Reg.scala 27:20]
  wire [31:0] _T_2351 = _T_2320 ? ic_miss_buff_data_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2366 = _T_2365 | _T_2351; // @[Mux.scala 27:72]
  wire  _T_2323 = _T_2295 == 4'h9; // @[el2_ifu_mem_ctl.scala 464:89]
  reg [31:0] ic_miss_buff_data_9; // @[Reg.scala 27:20]
  wire [31:0] _T_2352 = _T_2323 ? ic_miss_buff_data_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2367 = _T_2366 | _T_2352; // @[Mux.scala 27:72]
  wire  _T_2326 = _T_2295 == 4'ha; // @[el2_ifu_mem_ctl.scala 464:89]
  reg [31:0] ic_miss_buff_data_10; // @[Reg.scala 27:20]
  wire [31:0] _T_2353 = _T_2326 ? ic_miss_buff_data_10 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2368 = _T_2367 | _T_2353; // @[Mux.scala 27:72]
  wire  _T_2329 = _T_2295 == 4'hb; // @[el2_ifu_mem_ctl.scala 464:89]
  reg [31:0] ic_miss_buff_data_11; // @[Reg.scala 27:20]
  wire [31:0] _T_2354 = _T_2329 ? ic_miss_buff_data_11 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2369 = _T_2368 | _T_2354; // @[Mux.scala 27:72]
  wire  _T_2332 = _T_2295 == 4'hc; // @[el2_ifu_mem_ctl.scala 464:89]
  reg [31:0] ic_miss_buff_data_12; // @[Reg.scala 27:20]
  wire [31:0] _T_2355 = _T_2332 ? ic_miss_buff_data_12 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2370 = _T_2369 | _T_2355; // @[Mux.scala 27:72]
  wire  _T_2335 = _T_2295 == 4'hd; // @[el2_ifu_mem_ctl.scala 464:89]
  reg [31:0] ic_miss_buff_data_13; // @[Reg.scala 27:20]
  wire [31:0] _T_2356 = _T_2335 ? ic_miss_buff_data_13 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2371 = _T_2370 | _T_2356; // @[Mux.scala 27:72]
  wire  _T_2338 = _T_2295 == 4'he; // @[el2_ifu_mem_ctl.scala 464:89]
  reg [31:0] ic_miss_buff_data_14; // @[Reg.scala 27:20]
  wire [31:0] _T_2357 = _T_2338 ? ic_miss_buff_data_14 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2372 = _T_2371 | _T_2357; // @[Mux.scala 27:72]
  wire  _T_2341 = _T_2295 == 4'hf; // @[el2_ifu_mem_ctl.scala 464:89]
  reg [31:0] ic_miss_buff_data_15; // @[Reg.scala 27:20]
  wire [31:0] _T_2358 = _T_2341 ? ic_miss_buff_data_15 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2373 = _T_2372 | _T_2358; // @[Mux.scala 27:72]
  wire [3:0] _T_2375 = {ifu_bus_rid_ff[2:1],_T_2254,1'h0}; // @[Cat.scala 29:58]
  wire  _T_2376 = _T_2375 == 4'h0; // @[el2_ifu_mem_ctl.scala 465:66]
  wire [31:0] _T_2423 = _T_2376 ? ic_miss_buff_data_0 : 32'h0; // @[Mux.scala 27:72]
  wire  _T_2379 = _T_2375 == 4'h1; // @[el2_ifu_mem_ctl.scala 465:66]
  wire [31:0] _T_2424 = _T_2379 ? ic_miss_buff_data_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2439 = _T_2423 | _T_2424; // @[Mux.scala 27:72]
  wire  _T_2382 = _T_2375 == 4'h2; // @[el2_ifu_mem_ctl.scala 465:66]
  wire [31:0] _T_2425 = _T_2382 ? ic_miss_buff_data_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2440 = _T_2439 | _T_2425; // @[Mux.scala 27:72]
  wire  _T_2385 = _T_2375 == 4'h3; // @[el2_ifu_mem_ctl.scala 465:66]
  wire [31:0] _T_2426 = _T_2385 ? ic_miss_buff_data_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2441 = _T_2440 | _T_2426; // @[Mux.scala 27:72]
  wire  _T_2388 = _T_2375 == 4'h4; // @[el2_ifu_mem_ctl.scala 465:66]
  wire [31:0] _T_2427 = _T_2388 ? ic_miss_buff_data_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2442 = _T_2441 | _T_2427; // @[Mux.scala 27:72]
  wire  _T_2391 = _T_2375 == 4'h5; // @[el2_ifu_mem_ctl.scala 465:66]
  wire [31:0] _T_2428 = _T_2391 ? ic_miss_buff_data_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2443 = _T_2442 | _T_2428; // @[Mux.scala 27:72]
  wire  _T_2394 = _T_2375 == 4'h6; // @[el2_ifu_mem_ctl.scala 465:66]
  wire [31:0] _T_2429 = _T_2394 ? ic_miss_buff_data_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2444 = _T_2443 | _T_2429; // @[Mux.scala 27:72]
  wire  _T_2397 = _T_2375 == 4'h7; // @[el2_ifu_mem_ctl.scala 465:66]
  wire [31:0] _T_2430 = _T_2397 ? ic_miss_buff_data_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2445 = _T_2444 | _T_2430; // @[Mux.scala 27:72]
  wire  _T_2400 = _T_2375 == 4'h8; // @[el2_ifu_mem_ctl.scala 465:66]
  wire [31:0] _T_2431 = _T_2400 ? ic_miss_buff_data_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2446 = _T_2445 | _T_2431; // @[Mux.scala 27:72]
  wire  _T_2403 = _T_2375 == 4'h9; // @[el2_ifu_mem_ctl.scala 465:66]
  wire [31:0] _T_2432 = _T_2403 ? ic_miss_buff_data_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2447 = _T_2446 | _T_2432; // @[Mux.scala 27:72]
  wire  _T_2406 = _T_2375 == 4'ha; // @[el2_ifu_mem_ctl.scala 465:66]
  wire [31:0] _T_2433 = _T_2406 ? ic_miss_buff_data_10 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2448 = _T_2447 | _T_2433; // @[Mux.scala 27:72]
  wire  _T_2409 = _T_2375 == 4'hb; // @[el2_ifu_mem_ctl.scala 465:66]
  wire [31:0] _T_2434 = _T_2409 ? ic_miss_buff_data_11 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2449 = _T_2448 | _T_2434; // @[Mux.scala 27:72]
  wire  _T_2412 = _T_2375 == 4'hc; // @[el2_ifu_mem_ctl.scala 465:66]
  wire [31:0] _T_2435 = _T_2412 ? ic_miss_buff_data_12 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2450 = _T_2449 | _T_2435; // @[Mux.scala 27:72]
  wire  _T_2415 = _T_2375 == 4'hd; // @[el2_ifu_mem_ctl.scala 465:66]
  wire [31:0] _T_2436 = _T_2415 ? ic_miss_buff_data_13 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2451 = _T_2450 | _T_2436; // @[Mux.scala 27:72]
  wire  _T_2418 = _T_2375 == 4'he; // @[el2_ifu_mem_ctl.scala 465:66]
  wire [31:0] _T_2437 = _T_2418 ? ic_miss_buff_data_14 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2452 = _T_2451 | _T_2437; // @[Mux.scala 27:72]
  wire  _T_2421 = _T_2375 == 4'hf; // @[el2_ifu_mem_ctl.scala 465:66]
  wire [31:0] _T_2438 = _T_2421 ? ic_miss_buff_data_15 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2453 = _T_2452 | _T_2438; // @[Mux.scala 27:72]
  wire [63:0] ic_miss_buff_half = {_T_2373,_T_2453}; // @[Cat.scala 29:58]
  wire [6:0] _T_989 = {ic_miss_buff_half[63],ic_miss_buff_half[62],ic_miss_buff_half[61],ic_miss_buff_half[60],ic_miss_buff_half[59],ic_miss_buff_half[58],ic_miss_buff_half[57]}; // @[el2_lib.scala 401:13]
  wire  _T_990 = ^_T_989; // @[el2_lib.scala 401:20]
  wire [6:0] _T_996 = {ic_miss_buff_half[32],ic_miss_buff_half[31],ic_miss_buff_half[30],ic_miss_buff_half[29],ic_miss_buff_half[28],ic_miss_buff_half[27],ic_miss_buff_half[26]}; // @[el2_lib.scala 401:30]
  wire [7:0] _T_1003 = {ic_miss_buff_half[40],ic_miss_buff_half[39],ic_miss_buff_half[38],ic_miss_buff_half[37],ic_miss_buff_half[36],ic_miss_buff_half[35],ic_miss_buff_half[34],ic_miss_buff_half[33]}; // @[el2_lib.scala 401:30]
  wire [14:0] _T_1004 = {ic_miss_buff_half[40],ic_miss_buff_half[39],ic_miss_buff_half[38],ic_miss_buff_half[37],ic_miss_buff_half[36],ic_miss_buff_half[35],ic_miss_buff_half[34],ic_miss_buff_half[33],_T_996}; // @[el2_lib.scala 401:30]
  wire [7:0] _T_1011 = {ic_miss_buff_half[48],ic_miss_buff_half[47],ic_miss_buff_half[46],ic_miss_buff_half[45],ic_miss_buff_half[44],ic_miss_buff_half[43],ic_miss_buff_half[42],ic_miss_buff_half[41]}; // @[el2_lib.scala 401:30]
  wire [30:0] _T_1020 = {ic_miss_buff_half[56],ic_miss_buff_half[55],ic_miss_buff_half[54],ic_miss_buff_half[53],ic_miss_buff_half[52],ic_miss_buff_half[51],ic_miss_buff_half[50],ic_miss_buff_half[49],_T_1011,_T_1004}; // @[el2_lib.scala 401:30]
  wire  _T_1021 = ^_T_1020; // @[el2_lib.scala 401:37]
  wire [6:0] _T_1027 = {ic_miss_buff_half[17],ic_miss_buff_half[16],ic_miss_buff_half[15],ic_miss_buff_half[14],ic_miss_buff_half[13],ic_miss_buff_half[12],ic_miss_buff_half[11]}; // @[el2_lib.scala 401:47]
  wire [14:0] _T_1035 = {ic_miss_buff_half[25],ic_miss_buff_half[24],ic_miss_buff_half[23],ic_miss_buff_half[22],ic_miss_buff_half[21],ic_miss_buff_half[20],ic_miss_buff_half[19],ic_miss_buff_half[18],_T_1027}; // @[el2_lib.scala 401:47]
  wire [30:0] _T_1051 = {ic_miss_buff_half[56],ic_miss_buff_half[55],ic_miss_buff_half[54],ic_miss_buff_half[53],ic_miss_buff_half[52],ic_miss_buff_half[51],ic_miss_buff_half[50],ic_miss_buff_half[49],_T_1011,_T_1035}; // @[el2_lib.scala 401:47]
  wire  _T_1052 = ^_T_1051; // @[el2_lib.scala 401:54]
  wire [6:0] _T_1058 = {ic_miss_buff_half[10],ic_miss_buff_half[9],ic_miss_buff_half[8],ic_miss_buff_half[7],ic_miss_buff_half[6],ic_miss_buff_half[5],ic_miss_buff_half[4]}; // @[el2_lib.scala 401:64]
  wire [14:0] _T_1066 = {ic_miss_buff_half[25],ic_miss_buff_half[24],ic_miss_buff_half[23],ic_miss_buff_half[22],ic_miss_buff_half[21],ic_miss_buff_half[20],ic_miss_buff_half[19],ic_miss_buff_half[18],_T_1058}; // @[el2_lib.scala 401:64]
  wire [30:0] _T_1082 = {ic_miss_buff_half[56],ic_miss_buff_half[55],ic_miss_buff_half[54],ic_miss_buff_half[53],ic_miss_buff_half[52],ic_miss_buff_half[51],ic_miss_buff_half[50],ic_miss_buff_half[49],_T_1003,_T_1066}; // @[el2_lib.scala 401:64]
  wire  _T_1083 = ^_T_1082; // @[el2_lib.scala 401:71]
  wire [7:0] _T_1090 = {ic_miss_buff_half[14],ic_miss_buff_half[10],ic_miss_buff_half[9],ic_miss_buff_half[8],ic_miss_buff_half[7],ic_miss_buff_half[3],ic_miss_buff_half[2],ic_miss_buff_half[1]}; // @[el2_lib.scala 401:81]
  wire [16:0] _T_1099 = {ic_miss_buff_half[30],ic_miss_buff_half[29],ic_miss_buff_half[25],ic_miss_buff_half[24],ic_miss_buff_half[23],ic_miss_buff_half[22],ic_miss_buff_half[17],ic_miss_buff_half[16],ic_miss_buff_half[15],_T_1090}; // @[el2_lib.scala 401:81]
  wire [8:0] _T_1107 = {ic_miss_buff_half[47],ic_miss_buff_half[46],ic_miss_buff_half[45],ic_miss_buff_half[40],ic_miss_buff_half[39],ic_miss_buff_half[38],ic_miss_buff_half[37],ic_miss_buff_half[32],ic_miss_buff_half[31]}; // @[el2_lib.scala 401:81]
  wire [17:0] _T_1116 = {ic_miss_buff_half[63],ic_miss_buff_half[62],ic_miss_buff_half[61],ic_miss_buff_half[60],ic_miss_buff_half[56],ic_miss_buff_half[55],ic_miss_buff_half[54],ic_miss_buff_half[53],ic_miss_buff_half[48],_T_1107}; // @[el2_lib.scala 401:81]
  wire [34:0] _T_1117 = {_T_1116,_T_1099}; // @[el2_lib.scala 401:81]
  wire  _T_1118 = ^_T_1117; // @[el2_lib.scala 401:88]
  wire [7:0] _T_1125 = {ic_miss_buff_half[12],ic_miss_buff_half[10],ic_miss_buff_half[9],ic_miss_buff_half[6],ic_miss_buff_half[5],ic_miss_buff_half[3],ic_miss_buff_half[2],ic_miss_buff_half[0]}; // @[el2_lib.scala 401:98]
  wire [16:0] _T_1134 = {ic_miss_buff_half[28],ic_miss_buff_half[27],ic_miss_buff_half[25],ic_miss_buff_half[24],ic_miss_buff_half[21],ic_miss_buff_half[20],ic_miss_buff_half[17],ic_miss_buff_half[16],ic_miss_buff_half[13],_T_1125}; // @[el2_lib.scala 401:98]
  wire [8:0] _T_1142 = {ic_miss_buff_half[47],ic_miss_buff_half[44],ic_miss_buff_half[43],ic_miss_buff_half[40],ic_miss_buff_half[39],ic_miss_buff_half[36],ic_miss_buff_half[35],ic_miss_buff_half[32],ic_miss_buff_half[31]}; // @[el2_lib.scala 401:98]
  wire [17:0] _T_1151 = {ic_miss_buff_half[63],ic_miss_buff_half[62],ic_miss_buff_half[59],ic_miss_buff_half[58],ic_miss_buff_half[56],ic_miss_buff_half[55],ic_miss_buff_half[52],ic_miss_buff_half[51],ic_miss_buff_half[48],_T_1142}; // @[el2_lib.scala 401:98]
  wire [34:0] _T_1152 = {_T_1151,_T_1134}; // @[el2_lib.scala 401:98]
  wire  _T_1153 = ^_T_1152; // @[el2_lib.scala 401:105]
  wire [7:0] _T_1160 = {ic_miss_buff_half[11],ic_miss_buff_half[10],ic_miss_buff_half[8],ic_miss_buff_half[6],ic_miss_buff_half[4],ic_miss_buff_half[3],ic_miss_buff_half[1],ic_miss_buff_half[0]}; // @[el2_lib.scala 401:115]
  wire [16:0] _T_1169 = {ic_miss_buff_half[28],ic_miss_buff_half[26],ic_miss_buff_half[25],ic_miss_buff_half[23],ic_miss_buff_half[21],ic_miss_buff_half[19],ic_miss_buff_half[17],ic_miss_buff_half[15],ic_miss_buff_half[13],_T_1160}; // @[el2_lib.scala 401:115]
  wire [8:0] _T_1177 = {ic_miss_buff_half[46],ic_miss_buff_half[44],ic_miss_buff_half[42],ic_miss_buff_half[40],ic_miss_buff_half[38],ic_miss_buff_half[36],ic_miss_buff_half[34],ic_miss_buff_half[32],ic_miss_buff_half[30]}; // @[el2_lib.scala 401:115]
  wire [17:0] _T_1186 = {ic_miss_buff_half[63],ic_miss_buff_half[61],ic_miss_buff_half[59],ic_miss_buff_half[57],ic_miss_buff_half[56],ic_miss_buff_half[54],ic_miss_buff_half[52],ic_miss_buff_half[50],ic_miss_buff_half[48],_T_1177}; // @[el2_lib.scala 401:115]
  wire [34:0] _T_1187 = {_T_1186,_T_1169}; // @[el2_lib.scala 401:115]
  wire  _T_1188 = ^_T_1187; // @[el2_lib.scala 401:122]
  wire [70:0] _T_1233 = {_T_568,_T_599,_T_630,_T_661,_T_696,_T_731,_T_766,ifu_bus_rdata_ff}; // @[Cat.scala 29:58]
  wire [70:0] _T_1232 = {_T_990,_T_1021,_T_1052,_T_1083,_T_1118,_T_1153,_T_1188,_T_2373,_T_2453}; // @[Cat.scala 29:58]
  wire [141:0] _T_1234 = {_T_568,_T_599,_T_630,_T_661,_T_696,_T_731,_T_766,ifu_bus_rdata_ff,_T_1232}; // @[Cat.scala 29:58]
  wire [141:0] _T_1237 = {_T_990,_T_1021,_T_1052,_T_1083,_T_1118,_T_1153,_T_1188,_T_2373,_T_2453,_T_1233}; // @[Cat.scala 29:58]
  wire [141:0] ic_wr_16bytes_data = ifu_bus_rid_ff[0] ? _T_1234 : _T_1237; // @[el2_ifu_mem_ctl.scala 357:28]
  wire  _T_1196 = |io_ic_eccerr; // @[el2_ifu_mem_ctl.scala 347:56]
  wire  _T_1197 = _T_1196 & ic_act_hit_f; // @[el2_ifu_mem_ctl.scala 347:83]
  wire [4:0] bypass_index = imb_ff[4:0]; // @[el2_ifu_mem_ctl.scala 411:28]
  wire  _T_1413 = bypass_index[4:2] == 3'h0; // @[el2_ifu_mem_ctl.scala 413:114]
  wire  bus_ifu_wr_en = _T_13 & miss_pending; // @[el2_ifu_mem_ctl.scala 614:35]
  wire  _T_1282 = io_ifu_axi_rid == 3'h0; // @[el2_ifu_mem_ctl.scala 396:91]
  wire  write_fill_data_0 = bus_ifu_wr_en & _T_1282; // @[el2_ifu_mem_ctl.scala 396:73]
  wire  _T_1339 = ~ic_act_miss_f; // @[el2_ifu_mem_ctl.scala 402:118]
  wire  _T_1340 = ic_miss_buff_data_valid[0] & _T_1339; // @[el2_ifu_mem_ctl.scala 402:116]
  wire  ic_miss_buff_data_valid_in_0 = write_fill_data_0 | _T_1340; // @[el2_ifu_mem_ctl.scala 402:88]
  wire  _T_1436 = _T_1413 & ic_miss_buff_data_valid_in_0; // @[Mux.scala 27:72]
  wire  _T_1416 = bypass_index[4:2] == 3'h1; // @[el2_ifu_mem_ctl.scala 413:114]
  wire  _T_1283 = io_ifu_axi_rid == 3'h1; // @[el2_ifu_mem_ctl.scala 396:91]
  wire  write_fill_data_1 = bus_ifu_wr_en & _T_1283; // @[el2_ifu_mem_ctl.scala 396:73]
  wire  _T_1343 = ic_miss_buff_data_valid[1] & _T_1339; // @[el2_ifu_mem_ctl.scala 402:116]
  wire  ic_miss_buff_data_valid_in_1 = write_fill_data_1 | _T_1343; // @[el2_ifu_mem_ctl.scala 402:88]
  wire  _T_1437 = _T_1416 & ic_miss_buff_data_valid_in_1; // @[Mux.scala 27:72]
  wire  _T_1444 = _T_1436 | _T_1437; // @[Mux.scala 27:72]
  wire  _T_1419 = bypass_index[4:2] == 3'h2; // @[el2_ifu_mem_ctl.scala 413:114]
  wire  _T_1284 = io_ifu_axi_rid == 3'h2; // @[el2_ifu_mem_ctl.scala 396:91]
  wire  write_fill_data_2 = bus_ifu_wr_en & _T_1284; // @[el2_ifu_mem_ctl.scala 396:73]
  wire  _T_1346 = ic_miss_buff_data_valid[2] & _T_1339; // @[el2_ifu_mem_ctl.scala 402:116]
  wire  ic_miss_buff_data_valid_in_2 = write_fill_data_2 | _T_1346; // @[el2_ifu_mem_ctl.scala 402:88]
  wire  _T_1438 = _T_1419 & ic_miss_buff_data_valid_in_2; // @[Mux.scala 27:72]
  wire  _T_1445 = _T_1444 | _T_1438; // @[Mux.scala 27:72]
  wire  _T_1422 = bypass_index[4:2] == 3'h3; // @[el2_ifu_mem_ctl.scala 413:114]
  wire  _T_1285 = io_ifu_axi_rid == 3'h3; // @[el2_ifu_mem_ctl.scala 396:91]
  wire  write_fill_data_3 = bus_ifu_wr_en & _T_1285; // @[el2_ifu_mem_ctl.scala 396:73]
  wire  _T_1349 = ic_miss_buff_data_valid[3] & _T_1339; // @[el2_ifu_mem_ctl.scala 402:116]
  wire  ic_miss_buff_data_valid_in_3 = write_fill_data_3 | _T_1349; // @[el2_ifu_mem_ctl.scala 402:88]
  wire  _T_1439 = _T_1422 & ic_miss_buff_data_valid_in_3; // @[Mux.scala 27:72]
  wire  _T_1446 = _T_1445 | _T_1439; // @[Mux.scala 27:72]
  wire  _T_1425 = bypass_index[4:2] == 3'h4; // @[el2_ifu_mem_ctl.scala 413:114]
  wire  _T_1286 = io_ifu_axi_rid == 3'h4; // @[el2_ifu_mem_ctl.scala 396:91]
  wire  write_fill_data_4 = bus_ifu_wr_en & _T_1286; // @[el2_ifu_mem_ctl.scala 396:73]
  wire  _T_1352 = ic_miss_buff_data_valid[4] & _T_1339; // @[el2_ifu_mem_ctl.scala 402:116]
  wire  ic_miss_buff_data_valid_in_4 = write_fill_data_4 | _T_1352; // @[el2_ifu_mem_ctl.scala 402:88]
  wire  _T_1440 = _T_1425 & ic_miss_buff_data_valid_in_4; // @[Mux.scala 27:72]
  wire  _T_1447 = _T_1446 | _T_1440; // @[Mux.scala 27:72]
  wire  _T_1428 = bypass_index[4:2] == 3'h5; // @[el2_ifu_mem_ctl.scala 413:114]
  wire  _T_1287 = io_ifu_axi_rid == 3'h5; // @[el2_ifu_mem_ctl.scala 396:91]
  wire  write_fill_data_5 = bus_ifu_wr_en & _T_1287; // @[el2_ifu_mem_ctl.scala 396:73]
  wire  _T_1355 = ic_miss_buff_data_valid[5] & _T_1339; // @[el2_ifu_mem_ctl.scala 402:116]
  wire  ic_miss_buff_data_valid_in_5 = write_fill_data_5 | _T_1355; // @[el2_ifu_mem_ctl.scala 402:88]
  wire  _T_1441 = _T_1428 & ic_miss_buff_data_valid_in_5; // @[Mux.scala 27:72]
  wire  _T_1448 = _T_1447 | _T_1441; // @[Mux.scala 27:72]
  wire  _T_1431 = bypass_index[4:2] == 3'h6; // @[el2_ifu_mem_ctl.scala 413:114]
  wire  _T_1288 = io_ifu_axi_rid == 3'h6; // @[el2_ifu_mem_ctl.scala 396:91]
  wire  write_fill_data_6 = bus_ifu_wr_en & _T_1288; // @[el2_ifu_mem_ctl.scala 396:73]
  wire  _T_1358 = ic_miss_buff_data_valid[6] & _T_1339; // @[el2_ifu_mem_ctl.scala 402:116]
  wire  ic_miss_buff_data_valid_in_6 = write_fill_data_6 | _T_1358; // @[el2_ifu_mem_ctl.scala 402:88]
  wire  _T_1442 = _T_1431 & ic_miss_buff_data_valid_in_6; // @[Mux.scala 27:72]
  wire  _T_1449 = _T_1448 | _T_1442; // @[Mux.scala 27:72]
  wire  _T_1434 = bypass_index[4:2] == 3'h7; // @[el2_ifu_mem_ctl.scala 413:114]
  wire  _T_1289 = io_ifu_axi_rid == 3'h7; // @[el2_ifu_mem_ctl.scala 396:91]
  wire  write_fill_data_7 = bus_ifu_wr_en & _T_1289; // @[el2_ifu_mem_ctl.scala 396:73]
  wire  _T_1361 = ic_miss_buff_data_valid[7] & _T_1339; // @[el2_ifu_mem_ctl.scala 402:116]
  wire  ic_miss_buff_data_valid_in_7 = write_fill_data_7 | _T_1361; // @[el2_ifu_mem_ctl.scala 402:88]
  wire  _T_1443 = _T_1434 & ic_miss_buff_data_valid_in_7; // @[Mux.scala 27:72]
  wire  bypass_valid_value_check = _T_1449 | _T_1443; // @[Mux.scala 27:72]
  wire  _T_1452 = ~bypass_index[1]; // @[el2_ifu_mem_ctl.scala 414:58]
  wire  _T_1453 = bypass_valid_value_check & _T_1452; // @[el2_ifu_mem_ctl.scala 414:56]
  wire  _T_1455 = ~bypass_index[0]; // @[el2_ifu_mem_ctl.scala 414:77]
  wire  _T_1456 = _T_1453 & _T_1455; // @[el2_ifu_mem_ctl.scala 414:75]
  wire  _T_1461 = _T_1453 & bypass_index[0]; // @[el2_ifu_mem_ctl.scala 415:75]
  wire  _T_1462 = _T_1456 | _T_1461; // @[el2_ifu_mem_ctl.scala 414:95]
  wire  _T_1464 = bypass_valid_value_check & bypass_index[1]; // @[el2_ifu_mem_ctl.scala 416:56]
  wire  _T_1467 = _T_1464 & _T_1455; // @[el2_ifu_mem_ctl.scala 416:74]
  wire  _T_1468 = _T_1462 | _T_1467; // @[el2_ifu_mem_ctl.scala 415:94]
  wire  _T_1472 = _T_1464 & bypass_index[0]; // @[el2_ifu_mem_ctl.scala 417:51]
  wire [2:0] bypass_index_5_3_inc = bypass_index[4:2] + 3'h1; // @[el2_ifu_mem_ctl.scala 412:70]
  wire  _T_1473 = bypass_index_5_3_inc == 3'h0; // @[el2_ifu_mem_ctl.scala 417:132]
  wire  _T_1489 = _T_1473 & ic_miss_buff_data_valid_in_0; // @[Mux.scala 27:72]
  wire  _T_1475 = bypass_index_5_3_inc == 3'h1; // @[el2_ifu_mem_ctl.scala 417:132]
  wire  _T_1490 = _T_1475 & ic_miss_buff_data_valid_in_1; // @[Mux.scala 27:72]
  wire  _T_1497 = _T_1489 | _T_1490; // @[Mux.scala 27:72]
  wire  _T_1477 = bypass_index_5_3_inc == 3'h2; // @[el2_ifu_mem_ctl.scala 417:132]
  wire  _T_1491 = _T_1477 & ic_miss_buff_data_valid_in_2; // @[Mux.scala 27:72]
  wire  _T_1498 = _T_1497 | _T_1491; // @[Mux.scala 27:72]
  wire  _T_1479 = bypass_index_5_3_inc == 3'h3; // @[el2_ifu_mem_ctl.scala 417:132]
  wire  _T_1492 = _T_1479 & ic_miss_buff_data_valid_in_3; // @[Mux.scala 27:72]
  wire  _T_1499 = _T_1498 | _T_1492; // @[Mux.scala 27:72]
  wire  _T_1481 = bypass_index_5_3_inc == 3'h4; // @[el2_ifu_mem_ctl.scala 417:132]
  wire  _T_1493 = _T_1481 & ic_miss_buff_data_valid_in_4; // @[Mux.scala 27:72]
  wire  _T_1500 = _T_1499 | _T_1493; // @[Mux.scala 27:72]
  wire  _T_1483 = bypass_index_5_3_inc == 3'h5; // @[el2_ifu_mem_ctl.scala 417:132]
  wire  _T_1494 = _T_1483 & ic_miss_buff_data_valid_in_5; // @[Mux.scala 27:72]
  wire  _T_1501 = _T_1500 | _T_1494; // @[Mux.scala 27:72]
  wire  _T_1485 = bypass_index_5_3_inc == 3'h6; // @[el2_ifu_mem_ctl.scala 417:132]
  wire  _T_1495 = _T_1485 & ic_miss_buff_data_valid_in_6; // @[Mux.scala 27:72]
  wire  _T_1502 = _T_1501 | _T_1495; // @[Mux.scala 27:72]
  wire  _T_1487 = bypass_index_5_3_inc == 3'h7; // @[el2_ifu_mem_ctl.scala 417:132]
  wire  _T_1496 = _T_1487 & ic_miss_buff_data_valid_in_7; // @[Mux.scala 27:72]
  wire  _T_1503 = _T_1502 | _T_1496; // @[Mux.scala 27:72]
  wire  _T_1505 = _T_1472 & _T_1503; // @[el2_ifu_mem_ctl.scala 417:69]
  wire  _T_1506 = _T_1468 | _T_1505; // @[el2_ifu_mem_ctl.scala 416:94]
  wire [4:0] _GEN_473 = {{2'd0}, bypass_index[4:2]}; // @[el2_ifu_mem_ctl.scala 418:95]
  wire  _T_1509 = _GEN_473 == 5'h1f; // @[el2_ifu_mem_ctl.scala 418:95]
  wire  _T_1510 = bypass_valid_value_check & _T_1509; // @[el2_ifu_mem_ctl.scala 418:56]
  wire  bypass_data_ready_in = _T_1506 | _T_1510; // @[el2_ifu_mem_ctl.scala 417:181]
  wire  _T_1511 = bypass_data_ready_in & crit_wd_byp_ok_ff; // @[el2_ifu_mem_ctl.scala 422:53]
  wire  _T_1512 = _T_1511 & uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 422:73]
  wire  _T_1514 = _T_1512 & _T_317; // @[el2_ifu_mem_ctl.scala 422:96]
  wire  _T_1516 = _T_1514 & _T_58; // @[el2_ifu_mem_ctl.scala 422:118]
  wire  _T_1518 = crit_wd_byp_ok_ff & _T_17; // @[el2_ifu_mem_ctl.scala 423:73]
  wire  _T_1520 = _T_1518 & _T_317; // @[el2_ifu_mem_ctl.scala 423:96]
  wire  _T_1522 = _T_1520 & _T_58; // @[el2_ifu_mem_ctl.scala 423:118]
  wire  _T_1523 = _T_1516 | _T_1522; // @[el2_ifu_mem_ctl.scala 422:143]
  reg  ic_crit_wd_rdy_new_ff; // @[el2_ifu_mem_ctl.scala 425:58]
  wire  _T_1524 = ic_crit_wd_rdy_new_ff & crit_wd_byp_ok_ff; // @[el2_ifu_mem_ctl.scala 424:54]
  wire  _T_1525 = ~fetch_req_icache_f; // @[el2_ifu_mem_ctl.scala 424:76]
  wire  _T_1526 = _T_1524 & _T_1525; // @[el2_ifu_mem_ctl.scala 424:74]
  wire  _T_1528 = _T_1526 & _T_317; // @[el2_ifu_mem_ctl.scala 424:96]
  wire  ic_crit_wd_rdy_new_in = _T_1523 | _T_1528; // @[el2_ifu_mem_ctl.scala 423:143]
  wire  ic_crit_wd_rdy = ic_crit_wd_rdy_new_in | ic_crit_wd_rdy_new_ff; // @[el2_ifu_mem_ctl.scala 624:43]
  wire  _T_1249 = ic_crit_wd_rdy | _T_2233; // @[el2_ifu_mem_ctl.scala 370:38]
  wire  _T_1251 = _T_1249 | _T_2249; // @[el2_ifu_mem_ctl.scala 370:64]
  wire  _T_1252 = ~_T_1251; // @[el2_ifu_mem_ctl.scala 370:21]
  wire  _T_1253 = ~fetch_req_iccm_f; // @[el2_ifu_mem_ctl.scala 370:98]
  wire  sel_ic_data = _T_1252 & _T_1253; // @[el2_ifu_mem_ctl.scala 370:96]
  wire  _T_2456 = io_ic_tag_perr & sel_ic_data; // @[el2_ifu_mem_ctl.scala 469:44]
  wire  _T_1622 = ifu_fetch_addr_int_f[1] & ifu_fetch_addr_int_f[0]; // @[el2_ifu_mem_ctl.scala 436:31]
  reg [7:0] ic_miss_buff_data_error; // @[el2_ifu_mem_ctl.scala 408:60]
  wire  _T_1566 = _T_1413 & ic_miss_buff_data_error[0]; // @[Mux.scala 27:72]
  wire  _T_1567 = _T_1416 & ic_miss_buff_data_error[1]; // @[Mux.scala 27:72]
  wire  _T_1574 = _T_1566 | _T_1567; // @[Mux.scala 27:72]
  wire  _T_1568 = _T_1419 & ic_miss_buff_data_error[2]; // @[Mux.scala 27:72]
  wire  _T_1575 = _T_1574 | _T_1568; // @[Mux.scala 27:72]
  wire  _T_1569 = _T_1422 & ic_miss_buff_data_error[3]; // @[Mux.scala 27:72]
  wire  _T_1576 = _T_1575 | _T_1569; // @[Mux.scala 27:72]
  wire  _T_1570 = _T_1425 & ic_miss_buff_data_error[4]; // @[Mux.scala 27:72]
  wire  _T_1577 = _T_1576 | _T_1570; // @[Mux.scala 27:72]
  wire  _T_1571 = _T_1428 & ic_miss_buff_data_error[5]; // @[Mux.scala 27:72]
  wire  _T_1578 = _T_1577 | _T_1571; // @[Mux.scala 27:72]
  wire  _T_1572 = _T_1431 & ic_miss_buff_data_error[6]; // @[Mux.scala 27:72]
  wire  _T_1579 = _T_1578 | _T_1572; // @[Mux.scala 27:72]
  wire  _T_1573 = _T_1434 & ic_miss_buff_data_error[7]; // @[Mux.scala 27:72]
  wire  ic_miss_buff_data_error_bypass = _T_1579 | _T_1573; // @[Mux.scala 27:72]
  wire  _T_1605 = _T_2166 & ic_miss_buff_data_error[0]; // @[Mux.scala 27:72]
  wire  _T_1606 = _T_2169 & ic_miss_buff_data_error[1]; // @[Mux.scala 27:72]
  wire  _T_1613 = _T_1605 | _T_1606; // @[Mux.scala 27:72]
  wire  _T_1607 = _T_2172 & ic_miss_buff_data_error[2]; // @[Mux.scala 27:72]
  wire  _T_1614 = _T_1613 | _T_1607; // @[Mux.scala 27:72]
  wire  _T_1608 = _T_2175 & ic_miss_buff_data_error[3]; // @[Mux.scala 27:72]
  wire  _T_1615 = _T_1614 | _T_1608; // @[Mux.scala 27:72]
  wire  _T_1609 = _T_2178 & ic_miss_buff_data_error[4]; // @[Mux.scala 27:72]
  wire  _T_1616 = _T_1615 | _T_1609; // @[Mux.scala 27:72]
  wire  _T_1610 = _T_2181 & ic_miss_buff_data_error[5]; // @[Mux.scala 27:72]
  wire  _T_1617 = _T_1616 | _T_1610; // @[Mux.scala 27:72]
  wire  _T_1611 = _T_2184 & ic_miss_buff_data_error[6]; // @[Mux.scala 27:72]
  wire  _T_1618 = _T_1617 | _T_1611; // @[Mux.scala 27:72]
  wire  _T_1612 = _T_2187 & ic_miss_buff_data_error[7]; // @[Mux.scala 27:72]
  wire  ic_miss_buff_data_error_bypass_inc = _T_1618 | _T_1612; // @[Mux.scala 27:72]
  wire  _T_1623 = ic_miss_buff_data_error_bypass | ic_miss_buff_data_error_bypass_inc; // @[el2_ifu_mem_ctl.scala 438:70]
  wire  ifu_byp_data_err_new = _T_1622 ? ic_miss_buff_data_error_bypass : _T_1623; // @[el2_ifu_mem_ctl.scala 436:56]
  wire  ifc_bus_acc_fault_f = ic_byp_hit_f & ifu_byp_data_err_new; // @[el2_ifu_mem_ctl.scala 381:42]
  wire  _T_2457 = ifc_region_acc_fault_final_f | ifc_bus_acc_fault_f; // @[el2_ifu_mem_ctl.scala 469:91]
  wire  _T_2458 = ~_T_2457; // @[el2_ifu_mem_ctl.scala 469:60]
  wire  ic_rd_parity_final_err = _T_2456 & _T_2458; // @[el2_ifu_mem_ctl.scala 469:58]
  reg  ic_debug_ict_array_sel_ff; // @[Reg.scala 27:20]
  reg  ic_tag_valid_out_1_0; // @[Reg.scala 27:20]
  wire  _T_10157 = _T_4950 & ic_tag_valid_out_1_0; // @[el2_ifu_mem_ctl.scala 761:10]
  reg  ic_tag_valid_out_1_1; // @[Reg.scala 27:20]
  wire  _T_10159 = _T_4951 & ic_tag_valid_out_1_1; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10412 = _T_10157 | _T_10159; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_2; // @[Reg.scala 27:20]
  wire  _T_10161 = _T_4952 & ic_tag_valid_out_1_2; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10413 = _T_10412 | _T_10161; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_3; // @[Reg.scala 27:20]
  wire  _T_10163 = _T_4953 & ic_tag_valid_out_1_3; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10414 = _T_10413 | _T_10163; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_4; // @[Reg.scala 27:20]
  wire  _T_10165 = _T_4954 & ic_tag_valid_out_1_4; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10415 = _T_10414 | _T_10165; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_5; // @[Reg.scala 27:20]
  wire  _T_10167 = _T_4955 & ic_tag_valid_out_1_5; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10416 = _T_10415 | _T_10167; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_6; // @[Reg.scala 27:20]
  wire  _T_10169 = _T_4956 & ic_tag_valid_out_1_6; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10417 = _T_10416 | _T_10169; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_7; // @[Reg.scala 27:20]
  wire  _T_10171 = _T_4957 & ic_tag_valid_out_1_7; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10418 = _T_10417 | _T_10171; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_8; // @[Reg.scala 27:20]
  wire  _T_10173 = _T_4958 & ic_tag_valid_out_1_8; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10419 = _T_10418 | _T_10173; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_9; // @[Reg.scala 27:20]
  wire  _T_10175 = _T_4959 & ic_tag_valid_out_1_9; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10420 = _T_10419 | _T_10175; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_10; // @[Reg.scala 27:20]
  wire  _T_10177 = _T_4960 & ic_tag_valid_out_1_10; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10421 = _T_10420 | _T_10177; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_11; // @[Reg.scala 27:20]
  wire  _T_10179 = _T_4961 & ic_tag_valid_out_1_11; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10422 = _T_10421 | _T_10179; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_12; // @[Reg.scala 27:20]
  wire  _T_10181 = _T_4962 & ic_tag_valid_out_1_12; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10423 = _T_10422 | _T_10181; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_13; // @[Reg.scala 27:20]
  wire  _T_10183 = _T_4963 & ic_tag_valid_out_1_13; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10424 = _T_10423 | _T_10183; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_14; // @[Reg.scala 27:20]
  wire  _T_10185 = _T_4964 & ic_tag_valid_out_1_14; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10425 = _T_10424 | _T_10185; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_15; // @[Reg.scala 27:20]
  wire  _T_10187 = _T_4965 & ic_tag_valid_out_1_15; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10426 = _T_10425 | _T_10187; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_16; // @[Reg.scala 27:20]
  wire  _T_10189 = _T_4966 & ic_tag_valid_out_1_16; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10427 = _T_10426 | _T_10189; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_17; // @[Reg.scala 27:20]
  wire  _T_10191 = _T_4967 & ic_tag_valid_out_1_17; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10428 = _T_10427 | _T_10191; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_18; // @[Reg.scala 27:20]
  wire  _T_10193 = _T_4968 & ic_tag_valid_out_1_18; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10429 = _T_10428 | _T_10193; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_19; // @[Reg.scala 27:20]
  wire  _T_10195 = _T_4969 & ic_tag_valid_out_1_19; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10430 = _T_10429 | _T_10195; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_20; // @[Reg.scala 27:20]
  wire  _T_10197 = _T_4970 & ic_tag_valid_out_1_20; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10431 = _T_10430 | _T_10197; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_21; // @[Reg.scala 27:20]
  wire  _T_10199 = _T_4971 & ic_tag_valid_out_1_21; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10432 = _T_10431 | _T_10199; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_22; // @[Reg.scala 27:20]
  wire  _T_10201 = _T_4972 & ic_tag_valid_out_1_22; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10433 = _T_10432 | _T_10201; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_23; // @[Reg.scala 27:20]
  wire  _T_10203 = _T_4973 & ic_tag_valid_out_1_23; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10434 = _T_10433 | _T_10203; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_24; // @[Reg.scala 27:20]
  wire  _T_10205 = _T_4974 & ic_tag_valid_out_1_24; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10435 = _T_10434 | _T_10205; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_25; // @[Reg.scala 27:20]
  wire  _T_10207 = _T_4975 & ic_tag_valid_out_1_25; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10436 = _T_10435 | _T_10207; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_26; // @[Reg.scala 27:20]
  wire  _T_10209 = _T_4976 & ic_tag_valid_out_1_26; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10437 = _T_10436 | _T_10209; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_27; // @[Reg.scala 27:20]
  wire  _T_10211 = _T_4977 & ic_tag_valid_out_1_27; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10438 = _T_10437 | _T_10211; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_28; // @[Reg.scala 27:20]
  wire  _T_10213 = _T_4978 & ic_tag_valid_out_1_28; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10439 = _T_10438 | _T_10213; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_29; // @[Reg.scala 27:20]
  wire  _T_10215 = _T_4979 & ic_tag_valid_out_1_29; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10440 = _T_10439 | _T_10215; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_30; // @[Reg.scala 27:20]
  wire  _T_10217 = _T_4980 & ic_tag_valid_out_1_30; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10441 = _T_10440 | _T_10217; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_31; // @[Reg.scala 27:20]
  wire  _T_10219 = _T_4981 & ic_tag_valid_out_1_31; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10442 = _T_10441 | _T_10219; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_32; // @[Reg.scala 27:20]
  wire  _T_10221 = _T_4982 & ic_tag_valid_out_1_32; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10443 = _T_10442 | _T_10221; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_33; // @[Reg.scala 27:20]
  wire  _T_10223 = _T_4983 & ic_tag_valid_out_1_33; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10444 = _T_10443 | _T_10223; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_34; // @[Reg.scala 27:20]
  wire  _T_10225 = _T_4984 & ic_tag_valid_out_1_34; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10445 = _T_10444 | _T_10225; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_35; // @[Reg.scala 27:20]
  wire  _T_10227 = _T_4985 & ic_tag_valid_out_1_35; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10446 = _T_10445 | _T_10227; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_36; // @[Reg.scala 27:20]
  wire  _T_10229 = _T_4986 & ic_tag_valid_out_1_36; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10447 = _T_10446 | _T_10229; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_37; // @[Reg.scala 27:20]
  wire  _T_10231 = _T_4987 & ic_tag_valid_out_1_37; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10448 = _T_10447 | _T_10231; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_38; // @[Reg.scala 27:20]
  wire  _T_10233 = _T_4988 & ic_tag_valid_out_1_38; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10449 = _T_10448 | _T_10233; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_39; // @[Reg.scala 27:20]
  wire  _T_10235 = _T_4989 & ic_tag_valid_out_1_39; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10450 = _T_10449 | _T_10235; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_40; // @[Reg.scala 27:20]
  wire  _T_10237 = _T_4990 & ic_tag_valid_out_1_40; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10451 = _T_10450 | _T_10237; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_41; // @[Reg.scala 27:20]
  wire  _T_10239 = _T_4991 & ic_tag_valid_out_1_41; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10452 = _T_10451 | _T_10239; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_42; // @[Reg.scala 27:20]
  wire  _T_10241 = _T_4992 & ic_tag_valid_out_1_42; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10453 = _T_10452 | _T_10241; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_43; // @[Reg.scala 27:20]
  wire  _T_10243 = _T_4993 & ic_tag_valid_out_1_43; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10454 = _T_10453 | _T_10243; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_44; // @[Reg.scala 27:20]
  wire  _T_10245 = _T_4994 & ic_tag_valid_out_1_44; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10455 = _T_10454 | _T_10245; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_45; // @[Reg.scala 27:20]
  wire  _T_10247 = _T_4995 & ic_tag_valid_out_1_45; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10456 = _T_10455 | _T_10247; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_46; // @[Reg.scala 27:20]
  wire  _T_10249 = _T_4996 & ic_tag_valid_out_1_46; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10457 = _T_10456 | _T_10249; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_47; // @[Reg.scala 27:20]
  wire  _T_10251 = _T_4997 & ic_tag_valid_out_1_47; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10458 = _T_10457 | _T_10251; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_48; // @[Reg.scala 27:20]
  wire  _T_10253 = _T_4998 & ic_tag_valid_out_1_48; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10459 = _T_10458 | _T_10253; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_49; // @[Reg.scala 27:20]
  wire  _T_10255 = _T_4999 & ic_tag_valid_out_1_49; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10460 = _T_10459 | _T_10255; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_50; // @[Reg.scala 27:20]
  wire  _T_10257 = _T_5000 & ic_tag_valid_out_1_50; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10461 = _T_10460 | _T_10257; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_51; // @[Reg.scala 27:20]
  wire  _T_10259 = _T_5001 & ic_tag_valid_out_1_51; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10462 = _T_10461 | _T_10259; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_52; // @[Reg.scala 27:20]
  wire  _T_10261 = _T_5002 & ic_tag_valid_out_1_52; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10463 = _T_10462 | _T_10261; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_53; // @[Reg.scala 27:20]
  wire  _T_10263 = _T_5003 & ic_tag_valid_out_1_53; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10464 = _T_10463 | _T_10263; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_54; // @[Reg.scala 27:20]
  wire  _T_10265 = _T_5004 & ic_tag_valid_out_1_54; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10465 = _T_10464 | _T_10265; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_55; // @[Reg.scala 27:20]
  wire  _T_10267 = _T_5005 & ic_tag_valid_out_1_55; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10466 = _T_10465 | _T_10267; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_56; // @[Reg.scala 27:20]
  wire  _T_10269 = _T_5006 & ic_tag_valid_out_1_56; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10467 = _T_10466 | _T_10269; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_57; // @[Reg.scala 27:20]
  wire  _T_10271 = _T_5007 & ic_tag_valid_out_1_57; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10468 = _T_10467 | _T_10271; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_58; // @[Reg.scala 27:20]
  wire  _T_10273 = _T_5008 & ic_tag_valid_out_1_58; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10469 = _T_10468 | _T_10273; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_59; // @[Reg.scala 27:20]
  wire  _T_10275 = _T_5009 & ic_tag_valid_out_1_59; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10470 = _T_10469 | _T_10275; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_60; // @[Reg.scala 27:20]
  wire  _T_10277 = _T_5010 & ic_tag_valid_out_1_60; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10471 = _T_10470 | _T_10277; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_61; // @[Reg.scala 27:20]
  wire  _T_10279 = _T_5011 & ic_tag_valid_out_1_61; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10472 = _T_10471 | _T_10279; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_62; // @[Reg.scala 27:20]
  wire  _T_10281 = _T_5012 & ic_tag_valid_out_1_62; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10473 = _T_10472 | _T_10281; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_63; // @[Reg.scala 27:20]
  wire  _T_10283 = _T_5013 & ic_tag_valid_out_1_63; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10474 = _T_10473 | _T_10283; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_64; // @[Reg.scala 27:20]
  wire  _T_10285 = _T_5014 & ic_tag_valid_out_1_64; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10475 = _T_10474 | _T_10285; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_65; // @[Reg.scala 27:20]
  wire  _T_10287 = _T_5015 & ic_tag_valid_out_1_65; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10476 = _T_10475 | _T_10287; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_66; // @[Reg.scala 27:20]
  wire  _T_10289 = _T_5016 & ic_tag_valid_out_1_66; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10477 = _T_10476 | _T_10289; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_67; // @[Reg.scala 27:20]
  wire  _T_10291 = _T_5017 & ic_tag_valid_out_1_67; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10478 = _T_10477 | _T_10291; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_68; // @[Reg.scala 27:20]
  wire  _T_10293 = _T_5018 & ic_tag_valid_out_1_68; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10479 = _T_10478 | _T_10293; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_69; // @[Reg.scala 27:20]
  wire  _T_10295 = _T_5019 & ic_tag_valid_out_1_69; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10480 = _T_10479 | _T_10295; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_70; // @[Reg.scala 27:20]
  wire  _T_10297 = _T_5020 & ic_tag_valid_out_1_70; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10481 = _T_10480 | _T_10297; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_71; // @[Reg.scala 27:20]
  wire  _T_10299 = _T_5021 & ic_tag_valid_out_1_71; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10482 = _T_10481 | _T_10299; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_72; // @[Reg.scala 27:20]
  wire  _T_10301 = _T_5022 & ic_tag_valid_out_1_72; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10483 = _T_10482 | _T_10301; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_73; // @[Reg.scala 27:20]
  wire  _T_10303 = _T_5023 & ic_tag_valid_out_1_73; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10484 = _T_10483 | _T_10303; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_74; // @[Reg.scala 27:20]
  wire  _T_10305 = _T_5024 & ic_tag_valid_out_1_74; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10485 = _T_10484 | _T_10305; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_75; // @[Reg.scala 27:20]
  wire  _T_10307 = _T_5025 & ic_tag_valid_out_1_75; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10486 = _T_10485 | _T_10307; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_76; // @[Reg.scala 27:20]
  wire  _T_10309 = _T_5026 & ic_tag_valid_out_1_76; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10487 = _T_10486 | _T_10309; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_77; // @[Reg.scala 27:20]
  wire  _T_10311 = _T_5027 & ic_tag_valid_out_1_77; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10488 = _T_10487 | _T_10311; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_78; // @[Reg.scala 27:20]
  wire  _T_10313 = _T_5028 & ic_tag_valid_out_1_78; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10489 = _T_10488 | _T_10313; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_79; // @[Reg.scala 27:20]
  wire  _T_10315 = _T_5029 & ic_tag_valid_out_1_79; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10490 = _T_10489 | _T_10315; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_80; // @[Reg.scala 27:20]
  wire  _T_10317 = _T_5030 & ic_tag_valid_out_1_80; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10491 = _T_10490 | _T_10317; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_81; // @[Reg.scala 27:20]
  wire  _T_10319 = _T_5031 & ic_tag_valid_out_1_81; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10492 = _T_10491 | _T_10319; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_82; // @[Reg.scala 27:20]
  wire  _T_10321 = _T_5032 & ic_tag_valid_out_1_82; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10493 = _T_10492 | _T_10321; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_83; // @[Reg.scala 27:20]
  wire  _T_10323 = _T_5033 & ic_tag_valid_out_1_83; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10494 = _T_10493 | _T_10323; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_84; // @[Reg.scala 27:20]
  wire  _T_10325 = _T_5034 & ic_tag_valid_out_1_84; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10495 = _T_10494 | _T_10325; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_85; // @[Reg.scala 27:20]
  wire  _T_10327 = _T_5035 & ic_tag_valid_out_1_85; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10496 = _T_10495 | _T_10327; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_86; // @[Reg.scala 27:20]
  wire  _T_10329 = _T_5036 & ic_tag_valid_out_1_86; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10497 = _T_10496 | _T_10329; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_87; // @[Reg.scala 27:20]
  wire  _T_10331 = _T_5037 & ic_tag_valid_out_1_87; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10498 = _T_10497 | _T_10331; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_88; // @[Reg.scala 27:20]
  wire  _T_10333 = _T_5038 & ic_tag_valid_out_1_88; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10499 = _T_10498 | _T_10333; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_89; // @[Reg.scala 27:20]
  wire  _T_10335 = _T_5039 & ic_tag_valid_out_1_89; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10500 = _T_10499 | _T_10335; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_90; // @[Reg.scala 27:20]
  wire  _T_10337 = _T_5040 & ic_tag_valid_out_1_90; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10501 = _T_10500 | _T_10337; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_91; // @[Reg.scala 27:20]
  wire  _T_10339 = _T_5041 & ic_tag_valid_out_1_91; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10502 = _T_10501 | _T_10339; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_92; // @[Reg.scala 27:20]
  wire  _T_10341 = _T_5042 & ic_tag_valid_out_1_92; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10503 = _T_10502 | _T_10341; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_93; // @[Reg.scala 27:20]
  wire  _T_10343 = _T_5043 & ic_tag_valid_out_1_93; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10504 = _T_10503 | _T_10343; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_94; // @[Reg.scala 27:20]
  wire  _T_10345 = _T_5044 & ic_tag_valid_out_1_94; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10505 = _T_10504 | _T_10345; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_95; // @[Reg.scala 27:20]
  wire  _T_10347 = _T_5045 & ic_tag_valid_out_1_95; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10506 = _T_10505 | _T_10347; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_96; // @[Reg.scala 27:20]
  wire  _T_10349 = _T_5046 & ic_tag_valid_out_1_96; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10507 = _T_10506 | _T_10349; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_97; // @[Reg.scala 27:20]
  wire  _T_10351 = _T_5047 & ic_tag_valid_out_1_97; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10508 = _T_10507 | _T_10351; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_98; // @[Reg.scala 27:20]
  wire  _T_10353 = _T_5048 & ic_tag_valid_out_1_98; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10509 = _T_10508 | _T_10353; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_99; // @[Reg.scala 27:20]
  wire  _T_10355 = _T_5049 & ic_tag_valid_out_1_99; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10510 = _T_10509 | _T_10355; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_100; // @[Reg.scala 27:20]
  wire  _T_10357 = _T_5050 & ic_tag_valid_out_1_100; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10511 = _T_10510 | _T_10357; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_101; // @[Reg.scala 27:20]
  wire  _T_10359 = _T_5051 & ic_tag_valid_out_1_101; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10512 = _T_10511 | _T_10359; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_102; // @[Reg.scala 27:20]
  wire  _T_10361 = _T_5052 & ic_tag_valid_out_1_102; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10513 = _T_10512 | _T_10361; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_103; // @[Reg.scala 27:20]
  wire  _T_10363 = _T_5053 & ic_tag_valid_out_1_103; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10514 = _T_10513 | _T_10363; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_104; // @[Reg.scala 27:20]
  wire  _T_10365 = _T_5054 & ic_tag_valid_out_1_104; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10515 = _T_10514 | _T_10365; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_105; // @[Reg.scala 27:20]
  wire  _T_10367 = _T_5055 & ic_tag_valid_out_1_105; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10516 = _T_10515 | _T_10367; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_106; // @[Reg.scala 27:20]
  wire  _T_10369 = _T_5056 & ic_tag_valid_out_1_106; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10517 = _T_10516 | _T_10369; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_107; // @[Reg.scala 27:20]
  wire  _T_10371 = _T_5057 & ic_tag_valid_out_1_107; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10518 = _T_10517 | _T_10371; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_108; // @[Reg.scala 27:20]
  wire  _T_10373 = _T_5058 & ic_tag_valid_out_1_108; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10519 = _T_10518 | _T_10373; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_109; // @[Reg.scala 27:20]
  wire  _T_10375 = _T_5059 & ic_tag_valid_out_1_109; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10520 = _T_10519 | _T_10375; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_110; // @[Reg.scala 27:20]
  wire  _T_10377 = _T_5060 & ic_tag_valid_out_1_110; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10521 = _T_10520 | _T_10377; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_111; // @[Reg.scala 27:20]
  wire  _T_10379 = _T_5061 & ic_tag_valid_out_1_111; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10522 = _T_10521 | _T_10379; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_112; // @[Reg.scala 27:20]
  wire  _T_10381 = _T_5062 & ic_tag_valid_out_1_112; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10523 = _T_10522 | _T_10381; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_113; // @[Reg.scala 27:20]
  wire  _T_10383 = _T_5063 & ic_tag_valid_out_1_113; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10524 = _T_10523 | _T_10383; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_114; // @[Reg.scala 27:20]
  wire  _T_10385 = _T_5064 & ic_tag_valid_out_1_114; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10525 = _T_10524 | _T_10385; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_115; // @[Reg.scala 27:20]
  wire  _T_10387 = _T_5065 & ic_tag_valid_out_1_115; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10526 = _T_10525 | _T_10387; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_116; // @[Reg.scala 27:20]
  wire  _T_10389 = _T_5066 & ic_tag_valid_out_1_116; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10527 = _T_10526 | _T_10389; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_117; // @[Reg.scala 27:20]
  wire  _T_10391 = _T_5067 & ic_tag_valid_out_1_117; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10528 = _T_10527 | _T_10391; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_118; // @[Reg.scala 27:20]
  wire  _T_10393 = _T_5068 & ic_tag_valid_out_1_118; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10529 = _T_10528 | _T_10393; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_119; // @[Reg.scala 27:20]
  wire  _T_10395 = _T_5069 & ic_tag_valid_out_1_119; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10530 = _T_10529 | _T_10395; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_120; // @[Reg.scala 27:20]
  wire  _T_10397 = _T_5070 & ic_tag_valid_out_1_120; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10531 = _T_10530 | _T_10397; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_121; // @[Reg.scala 27:20]
  wire  _T_10399 = _T_5071 & ic_tag_valid_out_1_121; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10532 = _T_10531 | _T_10399; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_122; // @[Reg.scala 27:20]
  wire  _T_10401 = _T_5072 & ic_tag_valid_out_1_122; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10533 = _T_10532 | _T_10401; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_123; // @[Reg.scala 27:20]
  wire  _T_10403 = _T_5073 & ic_tag_valid_out_1_123; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10534 = _T_10533 | _T_10403; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_124; // @[Reg.scala 27:20]
  wire  _T_10405 = _T_5074 & ic_tag_valid_out_1_124; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10535 = _T_10534 | _T_10405; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_125; // @[Reg.scala 27:20]
  wire  _T_10407 = _T_5075 & ic_tag_valid_out_1_125; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10536 = _T_10535 | _T_10407; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_126; // @[Reg.scala 27:20]
  wire  _T_10409 = _T_5076 & ic_tag_valid_out_1_126; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10537 = _T_10536 | _T_10409; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_127; // @[Reg.scala 27:20]
  wire  _T_10411 = _T_5077 & ic_tag_valid_out_1_127; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10538 = _T_10537 | _T_10411; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_0; // @[Reg.scala 27:20]
  wire  _T_9774 = _T_4950 & ic_tag_valid_out_0_0; // @[el2_ifu_mem_ctl.scala 761:10]
  reg  ic_tag_valid_out_0_1; // @[Reg.scala 27:20]
  wire  _T_9776 = _T_4951 & ic_tag_valid_out_0_1; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10029 = _T_9774 | _T_9776; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_2; // @[Reg.scala 27:20]
  wire  _T_9778 = _T_4952 & ic_tag_valid_out_0_2; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10030 = _T_10029 | _T_9778; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_3; // @[Reg.scala 27:20]
  wire  _T_9780 = _T_4953 & ic_tag_valid_out_0_3; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10031 = _T_10030 | _T_9780; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_4; // @[Reg.scala 27:20]
  wire  _T_9782 = _T_4954 & ic_tag_valid_out_0_4; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10032 = _T_10031 | _T_9782; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_5; // @[Reg.scala 27:20]
  wire  _T_9784 = _T_4955 & ic_tag_valid_out_0_5; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10033 = _T_10032 | _T_9784; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_6; // @[Reg.scala 27:20]
  wire  _T_9786 = _T_4956 & ic_tag_valid_out_0_6; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10034 = _T_10033 | _T_9786; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_7; // @[Reg.scala 27:20]
  wire  _T_9788 = _T_4957 & ic_tag_valid_out_0_7; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10035 = _T_10034 | _T_9788; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_8; // @[Reg.scala 27:20]
  wire  _T_9790 = _T_4958 & ic_tag_valid_out_0_8; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10036 = _T_10035 | _T_9790; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_9; // @[Reg.scala 27:20]
  wire  _T_9792 = _T_4959 & ic_tag_valid_out_0_9; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10037 = _T_10036 | _T_9792; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_10; // @[Reg.scala 27:20]
  wire  _T_9794 = _T_4960 & ic_tag_valid_out_0_10; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10038 = _T_10037 | _T_9794; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_11; // @[Reg.scala 27:20]
  wire  _T_9796 = _T_4961 & ic_tag_valid_out_0_11; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10039 = _T_10038 | _T_9796; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_12; // @[Reg.scala 27:20]
  wire  _T_9798 = _T_4962 & ic_tag_valid_out_0_12; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10040 = _T_10039 | _T_9798; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_13; // @[Reg.scala 27:20]
  wire  _T_9800 = _T_4963 & ic_tag_valid_out_0_13; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10041 = _T_10040 | _T_9800; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_14; // @[Reg.scala 27:20]
  wire  _T_9802 = _T_4964 & ic_tag_valid_out_0_14; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10042 = _T_10041 | _T_9802; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_15; // @[Reg.scala 27:20]
  wire  _T_9804 = _T_4965 & ic_tag_valid_out_0_15; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10043 = _T_10042 | _T_9804; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_16; // @[Reg.scala 27:20]
  wire  _T_9806 = _T_4966 & ic_tag_valid_out_0_16; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10044 = _T_10043 | _T_9806; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_17; // @[Reg.scala 27:20]
  wire  _T_9808 = _T_4967 & ic_tag_valid_out_0_17; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10045 = _T_10044 | _T_9808; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_18; // @[Reg.scala 27:20]
  wire  _T_9810 = _T_4968 & ic_tag_valid_out_0_18; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10046 = _T_10045 | _T_9810; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_19; // @[Reg.scala 27:20]
  wire  _T_9812 = _T_4969 & ic_tag_valid_out_0_19; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10047 = _T_10046 | _T_9812; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_20; // @[Reg.scala 27:20]
  wire  _T_9814 = _T_4970 & ic_tag_valid_out_0_20; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10048 = _T_10047 | _T_9814; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_21; // @[Reg.scala 27:20]
  wire  _T_9816 = _T_4971 & ic_tag_valid_out_0_21; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10049 = _T_10048 | _T_9816; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_22; // @[Reg.scala 27:20]
  wire  _T_9818 = _T_4972 & ic_tag_valid_out_0_22; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10050 = _T_10049 | _T_9818; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_23; // @[Reg.scala 27:20]
  wire  _T_9820 = _T_4973 & ic_tag_valid_out_0_23; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10051 = _T_10050 | _T_9820; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_24; // @[Reg.scala 27:20]
  wire  _T_9822 = _T_4974 & ic_tag_valid_out_0_24; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10052 = _T_10051 | _T_9822; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_25; // @[Reg.scala 27:20]
  wire  _T_9824 = _T_4975 & ic_tag_valid_out_0_25; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10053 = _T_10052 | _T_9824; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_26; // @[Reg.scala 27:20]
  wire  _T_9826 = _T_4976 & ic_tag_valid_out_0_26; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10054 = _T_10053 | _T_9826; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_27; // @[Reg.scala 27:20]
  wire  _T_9828 = _T_4977 & ic_tag_valid_out_0_27; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10055 = _T_10054 | _T_9828; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_28; // @[Reg.scala 27:20]
  wire  _T_9830 = _T_4978 & ic_tag_valid_out_0_28; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10056 = _T_10055 | _T_9830; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_29; // @[Reg.scala 27:20]
  wire  _T_9832 = _T_4979 & ic_tag_valid_out_0_29; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10057 = _T_10056 | _T_9832; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_30; // @[Reg.scala 27:20]
  wire  _T_9834 = _T_4980 & ic_tag_valid_out_0_30; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10058 = _T_10057 | _T_9834; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_31; // @[Reg.scala 27:20]
  wire  _T_9836 = _T_4981 & ic_tag_valid_out_0_31; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10059 = _T_10058 | _T_9836; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_32; // @[Reg.scala 27:20]
  wire  _T_9838 = _T_4982 & ic_tag_valid_out_0_32; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10060 = _T_10059 | _T_9838; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_33; // @[Reg.scala 27:20]
  wire  _T_9840 = _T_4983 & ic_tag_valid_out_0_33; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10061 = _T_10060 | _T_9840; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_34; // @[Reg.scala 27:20]
  wire  _T_9842 = _T_4984 & ic_tag_valid_out_0_34; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10062 = _T_10061 | _T_9842; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_35; // @[Reg.scala 27:20]
  wire  _T_9844 = _T_4985 & ic_tag_valid_out_0_35; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10063 = _T_10062 | _T_9844; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_36; // @[Reg.scala 27:20]
  wire  _T_9846 = _T_4986 & ic_tag_valid_out_0_36; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10064 = _T_10063 | _T_9846; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_37; // @[Reg.scala 27:20]
  wire  _T_9848 = _T_4987 & ic_tag_valid_out_0_37; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10065 = _T_10064 | _T_9848; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_38; // @[Reg.scala 27:20]
  wire  _T_9850 = _T_4988 & ic_tag_valid_out_0_38; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10066 = _T_10065 | _T_9850; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_39; // @[Reg.scala 27:20]
  wire  _T_9852 = _T_4989 & ic_tag_valid_out_0_39; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10067 = _T_10066 | _T_9852; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_40; // @[Reg.scala 27:20]
  wire  _T_9854 = _T_4990 & ic_tag_valid_out_0_40; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10068 = _T_10067 | _T_9854; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_41; // @[Reg.scala 27:20]
  wire  _T_9856 = _T_4991 & ic_tag_valid_out_0_41; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10069 = _T_10068 | _T_9856; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_42; // @[Reg.scala 27:20]
  wire  _T_9858 = _T_4992 & ic_tag_valid_out_0_42; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10070 = _T_10069 | _T_9858; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_43; // @[Reg.scala 27:20]
  wire  _T_9860 = _T_4993 & ic_tag_valid_out_0_43; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10071 = _T_10070 | _T_9860; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_44; // @[Reg.scala 27:20]
  wire  _T_9862 = _T_4994 & ic_tag_valid_out_0_44; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10072 = _T_10071 | _T_9862; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_45; // @[Reg.scala 27:20]
  wire  _T_9864 = _T_4995 & ic_tag_valid_out_0_45; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10073 = _T_10072 | _T_9864; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_46; // @[Reg.scala 27:20]
  wire  _T_9866 = _T_4996 & ic_tag_valid_out_0_46; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10074 = _T_10073 | _T_9866; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_47; // @[Reg.scala 27:20]
  wire  _T_9868 = _T_4997 & ic_tag_valid_out_0_47; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10075 = _T_10074 | _T_9868; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_48; // @[Reg.scala 27:20]
  wire  _T_9870 = _T_4998 & ic_tag_valid_out_0_48; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10076 = _T_10075 | _T_9870; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_49; // @[Reg.scala 27:20]
  wire  _T_9872 = _T_4999 & ic_tag_valid_out_0_49; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10077 = _T_10076 | _T_9872; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_50; // @[Reg.scala 27:20]
  wire  _T_9874 = _T_5000 & ic_tag_valid_out_0_50; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10078 = _T_10077 | _T_9874; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_51; // @[Reg.scala 27:20]
  wire  _T_9876 = _T_5001 & ic_tag_valid_out_0_51; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10079 = _T_10078 | _T_9876; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_52; // @[Reg.scala 27:20]
  wire  _T_9878 = _T_5002 & ic_tag_valid_out_0_52; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10080 = _T_10079 | _T_9878; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_53; // @[Reg.scala 27:20]
  wire  _T_9880 = _T_5003 & ic_tag_valid_out_0_53; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10081 = _T_10080 | _T_9880; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_54; // @[Reg.scala 27:20]
  wire  _T_9882 = _T_5004 & ic_tag_valid_out_0_54; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10082 = _T_10081 | _T_9882; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_55; // @[Reg.scala 27:20]
  wire  _T_9884 = _T_5005 & ic_tag_valid_out_0_55; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10083 = _T_10082 | _T_9884; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_56; // @[Reg.scala 27:20]
  wire  _T_9886 = _T_5006 & ic_tag_valid_out_0_56; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10084 = _T_10083 | _T_9886; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_57; // @[Reg.scala 27:20]
  wire  _T_9888 = _T_5007 & ic_tag_valid_out_0_57; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10085 = _T_10084 | _T_9888; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_58; // @[Reg.scala 27:20]
  wire  _T_9890 = _T_5008 & ic_tag_valid_out_0_58; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10086 = _T_10085 | _T_9890; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_59; // @[Reg.scala 27:20]
  wire  _T_9892 = _T_5009 & ic_tag_valid_out_0_59; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10087 = _T_10086 | _T_9892; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_60; // @[Reg.scala 27:20]
  wire  _T_9894 = _T_5010 & ic_tag_valid_out_0_60; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10088 = _T_10087 | _T_9894; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_61; // @[Reg.scala 27:20]
  wire  _T_9896 = _T_5011 & ic_tag_valid_out_0_61; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10089 = _T_10088 | _T_9896; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_62; // @[Reg.scala 27:20]
  wire  _T_9898 = _T_5012 & ic_tag_valid_out_0_62; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10090 = _T_10089 | _T_9898; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_63; // @[Reg.scala 27:20]
  wire  _T_9900 = _T_5013 & ic_tag_valid_out_0_63; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10091 = _T_10090 | _T_9900; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_64; // @[Reg.scala 27:20]
  wire  _T_9902 = _T_5014 & ic_tag_valid_out_0_64; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10092 = _T_10091 | _T_9902; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_65; // @[Reg.scala 27:20]
  wire  _T_9904 = _T_5015 & ic_tag_valid_out_0_65; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10093 = _T_10092 | _T_9904; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_66; // @[Reg.scala 27:20]
  wire  _T_9906 = _T_5016 & ic_tag_valid_out_0_66; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10094 = _T_10093 | _T_9906; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_67; // @[Reg.scala 27:20]
  wire  _T_9908 = _T_5017 & ic_tag_valid_out_0_67; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10095 = _T_10094 | _T_9908; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_68; // @[Reg.scala 27:20]
  wire  _T_9910 = _T_5018 & ic_tag_valid_out_0_68; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10096 = _T_10095 | _T_9910; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_69; // @[Reg.scala 27:20]
  wire  _T_9912 = _T_5019 & ic_tag_valid_out_0_69; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10097 = _T_10096 | _T_9912; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_70; // @[Reg.scala 27:20]
  wire  _T_9914 = _T_5020 & ic_tag_valid_out_0_70; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10098 = _T_10097 | _T_9914; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_71; // @[Reg.scala 27:20]
  wire  _T_9916 = _T_5021 & ic_tag_valid_out_0_71; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10099 = _T_10098 | _T_9916; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_72; // @[Reg.scala 27:20]
  wire  _T_9918 = _T_5022 & ic_tag_valid_out_0_72; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10100 = _T_10099 | _T_9918; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_73; // @[Reg.scala 27:20]
  wire  _T_9920 = _T_5023 & ic_tag_valid_out_0_73; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10101 = _T_10100 | _T_9920; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_74; // @[Reg.scala 27:20]
  wire  _T_9922 = _T_5024 & ic_tag_valid_out_0_74; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10102 = _T_10101 | _T_9922; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_75; // @[Reg.scala 27:20]
  wire  _T_9924 = _T_5025 & ic_tag_valid_out_0_75; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10103 = _T_10102 | _T_9924; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_76; // @[Reg.scala 27:20]
  wire  _T_9926 = _T_5026 & ic_tag_valid_out_0_76; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10104 = _T_10103 | _T_9926; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_77; // @[Reg.scala 27:20]
  wire  _T_9928 = _T_5027 & ic_tag_valid_out_0_77; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10105 = _T_10104 | _T_9928; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_78; // @[Reg.scala 27:20]
  wire  _T_9930 = _T_5028 & ic_tag_valid_out_0_78; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10106 = _T_10105 | _T_9930; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_79; // @[Reg.scala 27:20]
  wire  _T_9932 = _T_5029 & ic_tag_valid_out_0_79; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10107 = _T_10106 | _T_9932; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_80; // @[Reg.scala 27:20]
  wire  _T_9934 = _T_5030 & ic_tag_valid_out_0_80; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10108 = _T_10107 | _T_9934; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_81; // @[Reg.scala 27:20]
  wire  _T_9936 = _T_5031 & ic_tag_valid_out_0_81; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10109 = _T_10108 | _T_9936; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_82; // @[Reg.scala 27:20]
  wire  _T_9938 = _T_5032 & ic_tag_valid_out_0_82; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10110 = _T_10109 | _T_9938; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_83; // @[Reg.scala 27:20]
  wire  _T_9940 = _T_5033 & ic_tag_valid_out_0_83; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10111 = _T_10110 | _T_9940; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_84; // @[Reg.scala 27:20]
  wire  _T_9942 = _T_5034 & ic_tag_valid_out_0_84; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10112 = _T_10111 | _T_9942; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_85; // @[Reg.scala 27:20]
  wire  _T_9944 = _T_5035 & ic_tag_valid_out_0_85; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10113 = _T_10112 | _T_9944; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_86; // @[Reg.scala 27:20]
  wire  _T_9946 = _T_5036 & ic_tag_valid_out_0_86; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10114 = _T_10113 | _T_9946; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_87; // @[Reg.scala 27:20]
  wire  _T_9948 = _T_5037 & ic_tag_valid_out_0_87; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10115 = _T_10114 | _T_9948; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_88; // @[Reg.scala 27:20]
  wire  _T_9950 = _T_5038 & ic_tag_valid_out_0_88; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10116 = _T_10115 | _T_9950; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_89; // @[Reg.scala 27:20]
  wire  _T_9952 = _T_5039 & ic_tag_valid_out_0_89; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10117 = _T_10116 | _T_9952; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_90; // @[Reg.scala 27:20]
  wire  _T_9954 = _T_5040 & ic_tag_valid_out_0_90; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10118 = _T_10117 | _T_9954; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_91; // @[Reg.scala 27:20]
  wire  _T_9956 = _T_5041 & ic_tag_valid_out_0_91; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10119 = _T_10118 | _T_9956; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_92; // @[Reg.scala 27:20]
  wire  _T_9958 = _T_5042 & ic_tag_valid_out_0_92; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10120 = _T_10119 | _T_9958; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_93; // @[Reg.scala 27:20]
  wire  _T_9960 = _T_5043 & ic_tag_valid_out_0_93; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10121 = _T_10120 | _T_9960; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_94; // @[Reg.scala 27:20]
  wire  _T_9962 = _T_5044 & ic_tag_valid_out_0_94; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10122 = _T_10121 | _T_9962; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_95; // @[Reg.scala 27:20]
  wire  _T_9964 = _T_5045 & ic_tag_valid_out_0_95; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10123 = _T_10122 | _T_9964; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_96; // @[Reg.scala 27:20]
  wire  _T_9966 = _T_5046 & ic_tag_valid_out_0_96; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10124 = _T_10123 | _T_9966; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_97; // @[Reg.scala 27:20]
  wire  _T_9968 = _T_5047 & ic_tag_valid_out_0_97; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10125 = _T_10124 | _T_9968; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_98; // @[Reg.scala 27:20]
  wire  _T_9970 = _T_5048 & ic_tag_valid_out_0_98; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10126 = _T_10125 | _T_9970; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_99; // @[Reg.scala 27:20]
  wire  _T_9972 = _T_5049 & ic_tag_valid_out_0_99; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10127 = _T_10126 | _T_9972; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_100; // @[Reg.scala 27:20]
  wire  _T_9974 = _T_5050 & ic_tag_valid_out_0_100; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10128 = _T_10127 | _T_9974; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_101; // @[Reg.scala 27:20]
  wire  _T_9976 = _T_5051 & ic_tag_valid_out_0_101; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10129 = _T_10128 | _T_9976; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_102; // @[Reg.scala 27:20]
  wire  _T_9978 = _T_5052 & ic_tag_valid_out_0_102; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10130 = _T_10129 | _T_9978; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_103; // @[Reg.scala 27:20]
  wire  _T_9980 = _T_5053 & ic_tag_valid_out_0_103; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10131 = _T_10130 | _T_9980; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_104; // @[Reg.scala 27:20]
  wire  _T_9982 = _T_5054 & ic_tag_valid_out_0_104; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10132 = _T_10131 | _T_9982; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_105; // @[Reg.scala 27:20]
  wire  _T_9984 = _T_5055 & ic_tag_valid_out_0_105; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10133 = _T_10132 | _T_9984; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_106; // @[Reg.scala 27:20]
  wire  _T_9986 = _T_5056 & ic_tag_valid_out_0_106; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10134 = _T_10133 | _T_9986; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_107; // @[Reg.scala 27:20]
  wire  _T_9988 = _T_5057 & ic_tag_valid_out_0_107; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10135 = _T_10134 | _T_9988; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_108; // @[Reg.scala 27:20]
  wire  _T_9990 = _T_5058 & ic_tag_valid_out_0_108; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10136 = _T_10135 | _T_9990; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_109; // @[Reg.scala 27:20]
  wire  _T_9992 = _T_5059 & ic_tag_valid_out_0_109; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10137 = _T_10136 | _T_9992; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_110; // @[Reg.scala 27:20]
  wire  _T_9994 = _T_5060 & ic_tag_valid_out_0_110; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10138 = _T_10137 | _T_9994; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_111; // @[Reg.scala 27:20]
  wire  _T_9996 = _T_5061 & ic_tag_valid_out_0_111; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10139 = _T_10138 | _T_9996; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_112; // @[Reg.scala 27:20]
  wire  _T_9998 = _T_5062 & ic_tag_valid_out_0_112; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10140 = _T_10139 | _T_9998; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_113; // @[Reg.scala 27:20]
  wire  _T_10000 = _T_5063 & ic_tag_valid_out_0_113; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10141 = _T_10140 | _T_10000; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_114; // @[Reg.scala 27:20]
  wire  _T_10002 = _T_5064 & ic_tag_valid_out_0_114; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10142 = _T_10141 | _T_10002; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_115; // @[Reg.scala 27:20]
  wire  _T_10004 = _T_5065 & ic_tag_valid_out_0_115; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10143 = _T_10142 | _T_10004; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_116; // @[Reg.scala 27:20]
  wire  _T_10006 = _T_5066 & ic_tag_valid_out_0_116; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10144 = _T_10143 | _T_10006; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_117; // @[Reg.scala 27:20]
  wire  _T_10008 = _T_5067 & ic_tag_valid_out_0_117; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10145 = _T_10144 | _T_10008; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_118; // @[Reg.scala 27:20]
  wire  _T_10010 = _T_5068 & ic_tag_valid_out_0_118; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10146 = _T_10145 | _T_10010; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_119; // @[Reg.scala 27:20]
  wire  _T_10012 = _T_5069 & ic_tag_valid_out_0_119; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10147 = _T_10146 | _T_10012; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_120; // @[Reg.scala 27:20]
  wire  _T_10014 = _T_5070 & ic_tag_valid_out_0_120; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10148 = _T_10147 | _T_10014; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_121; // @[Reg.scala 27:20]
  wire  _T_10016 = _T_5071 & ic_tag_valid_out_0_121; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10149 = _T_10148 | _T_10016; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_122; // @[Reg.scala 27:20]
  wire  _T_10018 = _T_5072 & ic_tag_valid_out_0_122; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10150 = _T_10149 | _T_10018; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_123; // @[Reg.scala 27:20]
  wire  _T_10020 = _T_5073 & ic_tag_valid_out_0_123; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10151 = _T_10150 | _T_10020; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_124; // @[Reg.scala 27:20]
  wire  _T_10022 = _T_5074 & ic_tag_valid_out_0_124; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10152 = _T_10151 | _T_10022; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_125; // @[Reg.scala 27:20]
  wire  _T_10024 = _T_5075 & ic_tag_valid_out_0_125; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10153 = _T_10152 | _T_10024; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_126; // @[Reg.scala 27:20]
  wire  _T_10026 = _T_5076 & ic_tag_valid_out_0_126; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10154 = _T_10153 | _T_10026; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_127; // @[Reg.scala 27:20]
  wire  _T_10028 = _T_5077 & ic_tag_valid_out_0_127; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10155 = _T_10154 | _T_10028; // @[el2_ifu_mem_ctl.scala 761:91]
  wire [1:0] ic_tag_valid_unq = {_T_10538,_T_10155}; // @[Cat.scala 29:58]
  reg [1:0] ic_debug_way_ff; // @[Reg.scala 27:20]
  reg  ic_debug_rd_en_ff; // @[el2_ifu_mem_ctl.scala 835:54]
  wire [1:0] _T_10578 = ic_debug_rd_en_ff ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [1:0] _T_10579 = ic_debug_way_ff & _T_10578; // @[el2_ifu_mem_ctl.scala 816:67]
  wire [1:0] _T_10580 = ic_tag_valid_unq & _T_10579; // @[el2_ifu_mem_ctl.scala 816:48]
  wire  ic_debug_tag_val_rd_out = |_T_10580; // @[el2_ifu_mem_ctl.scala 816:115]
  wire [65:0] _T_1208 = {2'h0,io_ictag_debug_rd_data[25:21],32'h0,io_ictag_debug_rd_data[20:0],1'h0,way_status,3'h0,ic_debug_tag_val_rd_out}; // @[Cat.scala 29:58]
  reg [70:0] _T_1209; // @[Reg.scala 27:20]
  wire  ifu_wr_cumulative_err = ifu_wr_cumulative_err_data & _T_2591; // @[el2_ifu_mem_ctl.scala 364:80]
  wire  _T_1247 = ~ifu_byp_data_err_new; // @[el2_ifu_mem_ctl.scala 369:98]
  wire  sel_byp_data = _T_1251 & _T_1247; // @[el2_ifu_mem_ctl.scala 369:96]
  wire [63:0] _T_1258 = fetch_req_iccm_f ? 64'hffffffffffffffff : 64'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_1259 = _T_1258 & io_iccm_rd_data; // @[el2_ifu_mem_ctl.scala 376:69]
  wire [63:0] _T_1261 = sel_byp_data ? 64'hffffffffffffffff : 64'h0; // @[Bitwise.scala 72:12]
  wire  _T_2113 = ~ifu_fetch_addr_int_f[0]; // @[el2_ifu_mem_ctl.scala 444:31]
  wire  _T_1626 = ~ifu_fetch_addr_int_f[1]; // @[el2_ifu_mem_ctl.scala 440:38]
  wire [3:0] byp_fetch_index_inc_0 = {byp_fetch_index_inc,1'h0}; // @[Cat.scala 29:58]
  wire  _T_1627 = byp_fetch_index_inc_0 == 4'h0; // @[el2_ifu_mem_ctl.scala 441:73]
  wire [15:0] _T_1675 = _T_1627 ? ic_miss_buff_data_0[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire  _T_1630 = byp_fetch_index_inc_0 == 4'h1; // @[el2_ifu_mem_ctl.scala 441:73]
  wire [15:0] _T_1676 = _T_1630 ? ic_miss_buff_data_1[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1691 = _T_1675 | _T_1676; // @[Mux.scala 27:72]
  wire  _T_1633 = byp_fetch_index_inc_0 == 4'h2; // @[el2_ifu_mem_ctl.scala 441:73]
  wire [15:0] _T_1677 = _T_1633 ? ic_miss_buff_data_2[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1692 = _T_1691 | _T_1677; // @[Mux.scala 27:72]
  wire  _T_1636 = byp_fetch_index_inc_0 == 4'h3; // @[el2_ifu_mem_ctl.scala 441:73]
  wire [15:0] _T_1678 = _T_1636 ? ic_miss_buff_data_3[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1693 = _T_1692 | _T_1678; // @[Mux.scala 27:72]
  wire  _T_1639 = byp_fetch_index_inc_0 == 4'h4; // @[el2_ifu_mem_ctl.scala 441:73]
  wire [15:0] _T_1679 = _T_1639 ? ic_miss_buff_data_4[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1694 = _T_1693 | _T_1679; // @[Mux.scala 27:72]
  wire  _T_1642 = byp_fetch_index_inc_0 == 4'h5; // @[el2_ifu_mem_ctl.scala 441:73]
  wire [15:0] _T_1680 = _T_1642 ? ic_miss_buff_data_5[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1695 = _T_1694 | _T_1680; // @[Mux.scala 27:72]
  wire  _T_1645 = byp_fetch_index_inc_0 == 4'h6; // @[el2_ifu_mem_ctl.scala 441:73]
  wire [15:0] _T_1681 = _T_1645 ? ic_miss_buff_data_6[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1696 = _T_1695 | _T_1681; // @[Mux.scala 27:72]
  wire  _T_1648 = byp_fetch_index_inc_0 == 4'h7; // @[el2_ifu_mem_ctl.scala 441:73]
  wire [15:0] _T_1682 = _T_1648 ? ic_miss_buff_data_7[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1697 = _T_1696 | _T_1682; // @[Mux.scala 27:72]
  wire  _T_1651 = byp_fetch_index_inc_0 == 4'h8; // @[el2_ifu_mem_ctl.scala 441:73]
  wire [15:0] _T_1683 = _T_1651 ? ic_miss_buff_data_8[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1698 = _T_1697 | _T_1683; // @[Mux.scala 27:72]
  wire  _T_1654 = byp_fetch_index_inc_0 == 4'h9; // @[el2_ifu_mem_ctl.scala 441:73]
  wire [15:0] _T_1684 = _T_1654 ? ic_miss_buff_data_9[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1699 = _T_1698 | _T_1684; // @[Mux.scala 27:72]
  wire  _T_1657 = byp_fetch_index_inc_0 == 4'ha; // @[el2_ifu_mem_ctl.scala 441:73]
  wire [15:0] _T_1685 = _T_1657 ? ic_miss_buff_data_10[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1700 = _T_1699 | _T_1685; // @[Mux.scala 27:72]
  wire  _T_1660 = byp_fetch_index_inc_0 == 4'hb; // @[el2_ifu_mem_ctl.scala 441:73]
  wire [15:0] _T_1686 = _T_1660 ? ic_miss_buff_data_11[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1701 = _T_1700 | _T_1686; // @[Mux.scala 27:72]
  wire  _T_1663 = byp_fetch_index_inc_0 == 4'hc; // @[el2_ifu_mem_ctl.scala 441:73]
  wire [15:0] _T_1687 = _T_1663 ? ic_miss_buff_data_12[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1702 = _T_1701 | _T_1687; // @[Mux.scala 27:72]
  wire  _T_1666 = byp_fetch_index_inc_0 == 4'hd; // @[el2_ifu_mem_ctl.scala 441:73]
  wire [15:0] _T_1688 = _T_1666 ? ic_miss_buff_data_13[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1703 = _T_1702 | _T_1688; // @[Mux.scala 27:72]
  wire  _T_1669 = byp_fetch_index_inc_0 == 4'he; // @[el2_ifu_mem_ctl.scala 441:73]
  wire [15:0] _T_1689 = _T_1669 ? ic_miss_buff_data_14[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1704 = _T_1703 | _T_1689; // @[Mux.scala 27:72]
  wire  _T_1672 = byp_fetch_index_inc_0 == 4'hf; // @[el2_ifu_mem_ctl.scala 441:73]
  wire [15:0] _T_1690 = _T_1672 ? ic_miss_buff_data_15[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1705 = _T_1704 | _T_1690; // @[Mux.scala 27:72]
  wire [3:0] byp_fetch_index_1 = {ifu_fetch_addr_int_f[4:2],1'h1}; // @[Cat.scala 29:58]
  wire  _T_1707 = byp_fetch_index_1 == 4'h0; // @[el2_ifu_mem_ctl.scala 441:179]
  wire [31:0] _T_1755 = _T_1707 ? ic_miss_buff_data_0 : 32'h0; // @[Mux.scala 27:72]
  wire  _T_1710 = byp_fetch_index_1 == 4'h1; // @[el2_ifu_mem_ctl.scala 441:179]
  wire [31:0] _T_1756 = _T_1710 ? ic_miss_buff_data_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1771 = _T_1755 | _T_1756; // @[Mux.scala 27:72]
  wire  _T_1713 = byp_fetch_index_1 == 4'h2; // @[el2_ifu_mem_ctl.scala 441:179]
  wire [31:0] _T_1757 = _T_1713 ? ic_miss_buff_data_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1772 = _T_1771 | _T_1757; // @[Mux.scala 27:72]
  wire  _T_1716 = byp_fetch_index_1 == 4'h3; // @[el2_ifu_mem_ctl.scala 441:179]
  wire [31:0] _T_1758 = _T_1716 ? ic_miss_buff_data_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1773 = _T_1772 | _T_1758; // @[Mux.scala 27:72]
  wire  _T_1719 = byp_fetch_index_1 == 4'h4; // @[el2_ifu_mem_ctl.scala 441:179]
  wire [31:0] _T_1759 = _T_1719 ? ic_miss_buff_data_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1774 = _T_1773 | _T_1759; // @[Mux.scala 27:72]
  wire  _T_1722 = byp_fetch_index_1 == 4'h5; // @[el2_ifu_mem_ctl.scala 441:179]
  wire [31:0] _T_1760 = _T_1722 ? ic_miss_buff_data_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1775 = _T_1774 | _T_1760; // @[Mux.scala 27:72]
  wire  _T_1725 = byp_fetch_index_1 == 4'h6; // @[el2_ifu_mem_ctl.scala 441:179]
  wire [31:0] _T_1761 = _T_1725 ? ic_miss_buff_data_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1776 = _T_1775 | _T_1761; // @[Mux.scala 27:72]
  wire  _T_1728 = byp_fetch_index_1 == 4'h7; // @[el2_ifu_mem_ctl.scala 441:179]
  wire [31:0] _T_1762 = _T_1728 ? ic_miss_buff_data_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1777 = _T_1776 | _T_1762; // @[Mux.scala 27:72]
  wire  _T_1731 = byp_fetch_index_1 == 4'h8; // @[el2_ifu_mem_ctl.scala 441:179]
  wire [31:0] _T_1763 = _T_1731 ? ic_miss_buff_data_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1778 = _T_1777 | _T_1763; // @[Mux.scala 27:72]
  wire  _T_1734 = byp_fetch_index_1 == 4'h9; // @[el2_ifu_mem_ctl.scala 441:179]
  wire [31:0] _T_1764 = _T_1734 ? ic_miss_buff_data_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1779 = _T_1778 | _T_1764; // @[Mux.scala 27:72]
  wire  _T_1737 = byp_fetch_index_1 == 4'ha; // @[el2_ifu_mem_ctl.scala 441:179]
  wire [31:0] _T_1765 = _T_1737 ? ic_miss_buff_data_10 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1780 = _T_1779 | _T_1765; // @[Mux.scala 27:72]
  wire  _T_1740 = byp_fetch_index_1 == 4'hb; // @[el2_ifu_mem_ctl.scala 441:179]
  wire [31:0] _T_1766 = _T_1740 ? ic_miss_buff_data_11 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1781 = _T_1780 | _T_1766; // @[Mux.scala 27:72]
  wire  _T_1743 = byp_fetch_index_1 == 4'hc; // @[el2_ifu_mem_ctl.scala 441:179]
  wire [31:0] _T_1767 = _T_1743 ? ic_miss_buff_data_12 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1782 = _T_1781 | _T_1767; // @[Mux.scala 27:72]
  wire  _T_1746 = byp_fetch_index_1 == 4'hd; // @[el2_ifu_mem_ctl.scala 441:179]
  wire [31:0] _T_1768 = _T_1746 ? ic_miss_buff_data_13 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1783 = _T_1782 | _T_1768; // @[Mux.scala 27:72]
  wire  _T_1749 = byp_fetch_index_1 == 4'he; // @[el2_ifu_mem_ctl.scala 441:179]
  wire [31:0] _T_1769 = _T_1749 ? ic_miss_buff_data_14 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1784 = _T_1783 | _T_1769; // @[Mux.scala 27:72]
  wire  _T_1752 = byp_fetch_index_1 == 4'hf; // @[el2_ifu_mem_ctl.scala 441:179]
  wire [31:0] _T_1770 = _T_1752 ? ic_miss_buff_data_15 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1785 = _T_1784 | _T_1770; // @[Mux.scala 27:72]
  wire [3:0] byp_fetch_index_0 = {ifu_fetch_addr_int_f[4:2],1'h0}; // @[Cat.scala 29:58]
  wire  _T_1787 = byp_fetch_index_0 == 4'h0; // @[el2_ifu_mem_ctl.scala 441:285]
  wire [31:0] _T_1835 = _T_1787 ? ic_miss_buff_data_0 : 32'h0; // @[Mux.scala 27:72]
  wire  _T_1790 = byp_fetch_index_0 == 4'h1; // @[el2_ifu_mem_ctl.scala 441:285]
  wire [31:0] _T_1836 = _T_1790 ? ic_miss_buff_data_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1851 = _T_1835 | _T_1836; // @[Mux.scala 27:72]
  wire  _T_1793 = byp_fetch_index_0 == 4'h2; // @[el2_ifu_mem_ctl.scala 441:285]
  wire [31:0] _T_1837 = _T_1793 ? ic_miss_buff_data_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1852 = _T_1851 | _T_1837; // @[Mux.scala 27:72]
  wire  _T_1796 = byp_fetch_index_0 == 4'h3; // @[el2_ifu_mem_ctl.scala 441:285]
  wire [31:0] _T_1838 = _T_1796 ? ic_miss_buff_data_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1853 = _T_1852 | _T_1838; // @[Mux.scala 27:72]
  wire  _T_1799 = byp_fetch_index_0 == 4'h4; // @[el2_ifu_mem_ctl.scala 441:285]
  wire [31:0] _T_1839 = _T_1799 ? ic_miss_buff_data_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1854 = _T_1853 | _T_1839; // @[Mux.scala 27:72]
  wire  _T_1802 = byp_fetch_index_0 == 4'h5; // @[el2_ifu_mem_ctl.scala 441:285]
  wire [31:0] _T_1840 = _T_1802 ? ic_miss_buff_data_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1855 = _T_1854 | _T_1840; // @[Mux.scala 27:72]
  wire  _T_1805 = byp_fetch_index_0 == 4'h6; // @[el2_ifu_mem_ctl.scala 441:285]
  wire [31:0] _T_1841 = _T_1805 ? ic_miss_buff_data_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1856 = _T_1855 | _T_1841; // @[Mux.scala 27:72]
  wire  _T_1808 = byp_fetch_index_0 == 4'h7; // @[el2_ifu_mem_ctl.scala 441:285]
  wire [31:0] _T_1842 = _T_1808 ? ic_miss_buff_data_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1857 = _T_1856 | _T_1842; // @[Mux.scala 27:72]
  wire  _T_1811 = byp_fetch_index_0 == 4'h8; // @[el2_ifu_mem_ctl.scala 441:285]
  wire [31:0] _T_1843 = _T_1811 ? ic_miss_buff_data_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1858 = _T_1857 | _T_1843; // @[Mux.scala 27:72]
  wire  _T_1814 = byp_fetch_index_0 == 4'h9; // @[el2_ifu_mem_ctl.scala 441:285]
  wire [31:0] _T_1844 = _T_1814 ? ic_miss_buff_data_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1859 = _T_1858 | _T_1844; // @[Mux.scala 27:72]
  wire  _T_1817 = byp_fetch_index_0 == 4'ha; // @[el2_ifu_mem_ctl.scala 441:285]
  wire [31:0] _T_1845 = _T_1817 ? ic_miss_buff_data_10 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1860 = _T_1859 | _T_1845; // @[Mux.scala 27:72]
  wire  _T_1820 = byp_fetch_index_0 == 4'hb; // @[el2_ifu_mem_ctl.scala 441:285]
  wire [31:0] _T_1846 = _T_1820 ? ic_miss_buff_data_11 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1861 = _T_1860 | _T_1846; // @[Mux.scala 27:72]
  wire  _T_1823 = byp_fetch_index_0 == 4'hc; // @[el2_ifu_mem_ctl.scala 441:285]
  wire [31:0] _T_1847 = _T_1823 ? ic_miss_buff_data_12 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1862 = _T_1861 | _T_1847; // @[Mux.scala 27:72]
  wire  _T_1826 = byp_fetch_index_0 == 4'hd; // @[el2_ifu_mem_ctl.scala 441:285]
  wire [31:0] _T_1848 = _T_1826 ? ic_miss_buff_data_13 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1863 = _T_1862 | _T_1848; // @[Mux.scala 27:72]
  wire  _T_1829 = byp_fetch_index_0 == 4'he; // @[el2_ifu_mem_ctl.scala 441:285]
  wire [31:0] _T_1849 = _T_1829 ? ic_miss_buff_data_14 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1864 = _T_1863 | _T_1849; // @[Mux.scala 27:72]
  wire  _T_1832 = byp_fetch_index_0 == 4'hf; // @[el2_ifu_mem_ctl.scala 441:285]
  wire [31:0] _T_1850 = _T_1832 ? ic_miss_buff_data_15 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1865 = _T_1864 | _T_1850; // @[Mux.scala 27:72]
  wire [79:0] _T_1868 = {_T_1705,_T_1785,_T_1865}; // @[Cat.scala 29:58]
  wire [3:0] byp_fetch_index_inc_1 = {byp_fetch_index_inc,1'h1}; // @[Cat.scala 29:58]
  wire  _T_1869 = byp_fetch_index_inc_1 == 4'h0; // @[el2_ifu_mem_ctl.scala 442:73]
  wire [15:0] _T_1917 = _T_1869 ? ic_miss_buff_data_0[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire  _T_1872 = byp_fetch_index_inc_1 == 4'h1; // @[el2_ifu_mem_ctl.scala 442:73]
  wire [15:0] _T_1918 = _T_1872 ? ic_miss_buff_data_1[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1933 = _T_1917 | _T_1918; // @[Mux.scala 27:72]
  wire  _T_1875 = byp_fetch_index_inc_1 == 4'h2; // @[el2_ifu_mem_ctl.scala 442:73]
  wire [15:0] _T_1919 = _T_1875 ? ic_miss_buff_data_2[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1934 = _T_1933 | _T_1919; // @[Mux.scala 27:72]
  wire  _T_1878 = byp_fetch_index_inc_1 == 4'h3; // @[el2_ifu_mem_ctl.scala 442:73]
  wire [15:0] _T_1920 = _T_1878 ? ic_miss_buff_data_3[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1935 = _T_1934 | _T_1920; // @[Mux.scala 27:72]
  wire  _T_1881 = byp_fetch_index_inc_1 == 4'h4; // @[el2_ifu_mem_ctl.scala 442:73]
  wire [15:0] _T_1921 = _T_1881 ? ic_miss_buff_data_4[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1936 = _T_1935 | _T_1921; // @[Mux.scala 27:72]
  wire  _T_1884 = byp_fetch_index_inc_1 == 4'h5; // @[el2_ifu_mem_ctl.scala 442:73]
  wire [15:0] _T_1922 = _T_1884 ? ic_miss_buff_data_5[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1937 = _T_1936 | _T_1922; // @[Mux.scala 27:72]
  wire  _T_1887 = byp_fetch_index_inc_1 == 4'h6; // @[el2_ifu_mem_ctl.scala 442:73]
  wire [15:0] _T_1923 = _T_1887 ? ic_miss_buff_data_6[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1938 = _T_1937 | _T_1923; // @[Mux.scala 27:72]
  wire  _T_1890 = byp_fetch_index_inc_1 == 4'h7; // @[el2_ifu_mem_ctl.scala 442:73]
  wire [15:0] _T_1924 = _T_1890 ? ic_miss_buff_data_7[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1939 = _T_1938 | _T_1924; // @[Mux.scala 27:72]
  wire  _T_1893 = byp_fetch_index_inc_1 == 4'h8; // @[el2_ifu_mem_ctl.scala 442:73]
  wire [15:0] _T_1925 = _T_1893 ? ic_miss_buff_data_8[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1940 = _T_1939 | _T_1925; // @[Mux.scala 27:72]
  wire  _T_1896 = byp_fetch_index_inc_1 == 4'h9; // @[el2_ifu_mem_ctl.scala 442:73]
  wire [15:0] _T_1926 = _T_1896 ? ic_miss_buff_data_9[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1941 = _T_1940 | _T_1926; // @[Mux.scala 27:72]
  wire  _T_1899 = byp_fetch_index_inc_1 == 4'ha; // @[el2_ifu_mem_ctl.scala 442:73]
  wire [15:0] _T_1927 = _T_1899 ? ic_miss_buff_data_10[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1942 = _T_1941 | _T_1927; // @[Mux.scala 27:72]
  wire  _T_1902 = byp_fetch_index_inc_1 == 4'hb; // @[el2_ifu_mem_ctl.scala 442:73]
  wire [15:0] _T_1928 = _T_1902 ? ic_miss_buff_data_11[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1943 = _T_1942 | _T_1928; // @[Mux.scala 27:72]
  wire  _T_1905 = byp_fetch_index_inc_1 == 4'hc; // @[el2_ifu_mem_ctl.scala 442:73]
  wire [15:0] _T_1929 = _T_1905 ? ic_miss_buff_data_12[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1944 = _T_1943 | _T_1929; // @[Mux.scala 27:72]
  wire  _T_1908 = byp_fetch_index_inc_1 == 4'hd; // @[el2_ifu_mem_ctl.scala 442:73]
  wire [15:0] _T_1930 = _T_1908 ? ic_miss_buff_data_13[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1945 = _T_1944 | _T_1930; // @[Mux.scala 27:72]
  wire  _T_1911 = byp_fetch_index_inc_1 == 4'he; // @[el2_ifu_mem_ctl.scala 442:73]
  wire [15:0] _T_1931 = _T_1911 ? ic_miss_buff_data_14[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1946 = _T_1945 | _T_1931; // @[Mux.scala 27:72]
  wire  _T_1914 = byp_fetch_index_inc_1 == 4'hf; // @[el2_ifu_mem_ctl.scala 442:73]
  wire [15:0] _T_1932 = _T_1914 ? ic_miss_buff_data_15[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1947 = _T_1946 | _T_1932; // @[Mux.scala 27:72]
  wire [31:0] _T_1997 = _T_1627 ? ic_miss_buff_data_0 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1998 = _T_1630 ? ic_miss_buff_data_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2013 = _T_1997 | _T_1998; // @[Mux.scala 27:72]
  wire [31:0] _T_1999 = _T_1633 ? ic_miss_buff_data_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2014 = _T_2013 | _T_1999; // @[Mux.scala 27:72]
  wire [31:0] _T_2000 = _T_1636 ? ic_miss_buff_data_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2015 = _T_2014 | _T_2000; // @[Mux.scala 27:72]
  wire [31:0] _T_2001 = _T_1639 ? ic_miss_buff_data_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2016 = _T_2015 | _T_2001; // @[Mux.scala 27:72]
  wire [31:0] _T_2002 = _T_1642 ? ic_miss_buff_data_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2017 = _T_2016 | _T_2002; // @[Mux.scala 27:72]
  wire [31:0] _T_2003 = _T_1645 ? ic_miss_buff_data_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2018 = _T_2017 | _T_2003; // @[Mux.scala 27:72]
  wire [31:0] _T_2004 = _T_1648 ? ic_miss_buff_data_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2019 = _T_2018 | _T_2004; // @[Mux.scala 27:72]
  wire [31:0] _T_2005 = _T_1651 ? ic_miss_buff_data_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2020 = _T_2019 | _T_2005; // @[Mux.scala 27:72]
  wire [31:0] _T_2006 = _T_1654 ? ic_miss_buff_data_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2021 = _T_2020 | _T_2006; // @[Mux.scala 27:72]
  wire [31:0] _T_2007 = _T_1657 ? ic_miss_buff_data_10 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2022 = _T_2021 | _T_2007; // @[Mux.scala 27:72]
  wire [31:0] _T_2008 = _T_1660 ? ic_miss_buff_data_11 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2023 = _T_2022 | _T_2008; // @[Mux.scala 27:72]
  wire [31:0] _T_2009 = _T_1663 ? ic_miss_buff_data_12 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2024 = _T_2023 | _T_2009; // @[Mux.scala 27:72]
  wire [31:0] _T_2010 = _T_1666 ? ic_miss_buff_data_13 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2025 = _T_2024 | _T_2010; // @[Mux.scala 27:72]
  wire [31:0] _T_2011 = _T_1669 ? ic_miss_buff_data_14 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2026 = _T_2025 | _T_2011; // @[Mux.scala 27:72]
  wire [31:0] _T_2012 = _T_1672 ? ic_miss_buff_data_15 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2027 = _T_2026 | _T_2012; // @[Mux.scala 27:72]
  wire [79:0] _T_2110 = {_T_1947,_T_2027,_T_1785}; // @[Cat.scala 29:58]
  wire [79:0] ic_byp_data_only_pre_new = _T_1626 ? _T_1868 : _T_2110; // @[el2_ifu_mem_ctl.scala 440:37]
  wire [79:0] _T_2115 = {16'h0,ic_byp_data_only_pre_new[79:16]}; // @[Cat.scala 29:58]
  wire [79:0] ic_byp_data_only_new = _T_2113 ? ic_byp_data_only_pre_new : _T_2115; // @[el2_ifu_mem_ctl.scala 444:30]
  wire [79:0] _GEN_474 = {{16'd0}, _T_1261}; // @[el2_ifu_mem_ctl.scala 376:114]
  wire [79:0] _T_1262 = _GEN_474 & ic_byp_data_only_new; // @[el2_ifu_mem_ctl.scala 376:114]
  wire [79:0] _GEN_475 = {{16'd0}, _T_1259}; // @[el2_ifu_mem_ctl.scala 376:88]
  wire [79:0] ic_premux_data_temp = _GEN_475 | _T_1262; // @[el2_ifu_mem_ctl.scala 376:88]
  wire  fetch_req_f_qual = io_ic_hit_f & _T_317; // @[el2_ifu_mem_ctl.scala 383:38]
  wire [1:0] _T_1271 = ifc_region_acc_fault_f ? 2'h2 : 2'h0; // @[el2_ifu_mem_ctl.scala 387:8]
  wire  _T_1273 = fetch_req_f_qual & io_ifu_bp_inst_mask_f; // @[el2_ifu_mem_ctl.scala 389:45]
  wire  _T_1275 = byp_fetch_index == 5'h1f; // @[el2_ifu_mem_ctl.scala 389:80]
  wire  _T_1276 = ~_T_1275; // @[el2_ifu_mem_ctl.scala 389:71]
  wire  _T_1277 = _T_1273 & _T_1276; // @[el2_ifu_mem_ctl.scala 389:69]
  wire  _T_1278 = err_stop_state != 2'h2; // @[el2_ifu_mem_ctl.scala 389:131]
  wire  _T_1279 = _T_1277 & _T_1278; // @[el2_ifu_mem_ctl.scala 389:114]
  wire [7:0] _T_1368 = {ic_miss_buff_data_valid_in_7,ic_miss_buff_data_valid_in_6,ic_miss_buff_data_valid_in_5,ic_miss_buff_data_valid_in_4,ic_miss_buff_data_valid_in_3,ic_miss_buff_data_valid_in_2,ic_miss_buff_data_valid_in_1,ic_miss_buff_data_valid_in_0}; // @[Cat.scala 29:58]
  wire  _T_1373 = ic_miss_buff_data_error[0] & _T_1339; // @[el2_ifu_mem_ctl.scala 407:32]
  wire  _T_2659 = |io_ifu_axi_rresp; // @[el2_ifu_mem_ctl.scala 620:47]
  wire  _T_2660 = _T_2659 & _T_13; // @[el2_ifu_mem_ctl.scala 620:50]
  wire  bus_ifu_wr_data_error = _T_2660 & miss_pending; // @[el2_ifu_mem_ctl.scala 620:68]
  wire  ic_miss_buff_data_error_in_0 = write_fill_data_0 ? bus_ifu_wr_data_error : _T_1373; // @[el2_ifu_mem_ctl.scala 406:72]
  wire  _T_1377 = ic_miss_buff_data_error[1] & _T_1339; // @[el2_ifu_mem_ctl.scala 407:32]
  wire  ic_miss_buff_data_error_in_1 = write_fill_data_1 ? bus_ifu_wr_data_error : _T_1377; // @[el2_ifu_mem_ctl.scala 406:72]
  wire  _T_1381 = ic_miss_buff_data_error[2] & _T_1339; // @[el2_ifu_mem_ctl.scala 407:32]
  wire  ic_miss_buff_data_error_in_2 = write_fill_data_2 ? bus_ifu_wr_data_error : _T_1381; // @[el2_ifu_mem_ctl.scala 406:72]
  wire  _T_1385 = ic_miss_buff_data_error[3] & _T_1339; // @[el2_ifu_mem_ctl.scala 407:32]
  wire  ic_miss_buff_data_error_in_3 = write_fill_data_3 ? bus_ifu_wr_data_error : _T_1385; // @[el2_ifu_mem_ctl.scala 406:72]
  wire  _T_1389 = ic_miss_buff_data_error[4] & _T_1339; // @[el2_ifu_mem_ctl.scala 407:32]
  wire  ic_miss_buff_data_error_in_4 = write_fill_data_4 ? bus_ifu_wr_data_error : _T_1389; // @[el2_ifu_mem_ctl.scala 406:72]
  wire  _T_1393 = ic_miss_buff_data_error[5] & _T_1339; // @[el2_ifu_mem_ctl.scala 407:32]
  wire  ic_miss_buff_data_error_in_5 = write_fill_data_5 ? bus_ifu_wr_data_error : _T_1393; // @[el2_ifu_mem_ctl.scala 406:72]
  wire  _T_1397 = ic_miss_buff_data_error[6] & _T_1339; // @[el2_ifu_mem_ctl.scala 407:32]
  wire  ic_miss_buff_data_error_in_6 = write_fill_data_6 ? bus_ifu_wr_data_error : _T_1397; // @[el2_ifu_mem_ctl.scala 406:72]
  wire  _T_1401 = ic_miss_buff_data_error[7] & _T_1339; // @[el2_ifu_mem_ctl.scala 407:32]
  wire  ic_miss_buff_data_error_in_7 = write_fill_data_7 ? bus_ifu_wr_data_error : _T_1401; // @[el2_ifu_mem_ctl.scala 406:72]
  wire [7:0] _T_1408 = {ic_miss_buff_data_error_in_7,ic_miss_buff_data_error_in_6,ic_miss_buff_data_error_in_5,ic_miss_buff_data_error_in_4,ic_miss_buff_data_error_in_3,ic_miss_buff_data_error_in_2,ic_miss_buff_data_error_in_1,ic_miss_buff_data_error_in_0}; // @[Cat.scala 29:58]
  reg [6:0] perr_ic_index_ff; // @[Reg.scala 27:20]
  wire  _T_2465 = 3'h0 == perr_state; // @[Conditional.scala 37:30]
  wire  _T_2473 = _T_6 & _T_317; // @[el2_ifu_mem_ctl.scala 489:65]
  wire  _T_2474 = _T_2473 | io_iccm_dma_sb_error; // @[el2_ifu_mem_ctl.scala 489:88]
  wire  _T_2476 = _T_2474 & _T_2587; // @[el2_ifu_mem_ctl.scala 489:112]
  wire  _T_2477 = 3'h1 == perr_state; // @[Conditional.scala 37:30]
  wire  _T_2478 = io_dec_tlu_flush_lower_wb | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 494:50]
  wire  _T_2480 = 3'h2 == perr_state; // @[Conditional.scala 37:30]
  wire  _T_2486 = 3'h4 == perr_state; // @[Conditional.scala 37:30]
  wire  _T_2488 = 3'h3 == perr_state; // @[Conditional.scala 37:30]
  wire  _GEN_39 = _T_2486 | _T_2488; // @[Conditional.scala 39:67]
  wire  _GEN_41 = _T_2480 ? _T_2478 : _GEN_39; // @[Conditional.scala 39:67]
  wire  _GEN_43 = _T_2477 ? _T_2478 : _GEN_41; // @[Conditional.scala 39:67]
  wire  perr_state_en = _T_2465 ? _T_2476 : _GEN_43; // @[Conditional.scala 40:58]
  wire  perr_sb_write_status = _T_2465 & perr_state_en; // @[Conditional.scala 40:58]
  wire  _T_2479 = io_dec_tlu_flush_lower_wb & io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 495:56]
  wire  _GEN_44 = _T_2477 & _T_2479; // @[Conditional.scala 39:67]
  wire  perr_sel_invalidate = _T_2465 ? 1'h0 : _GEN_44; // @[Conditional.scala 40:58]
  wire [1:0] perr_err_inv_way = perr_sel_invalidate ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  reg  dma_sb_err_state_ff; // @[el2_ifu_mem_ctl.scala 480:58]
  wire  _T_2462 = ~dma_sb_err_state_ff; // @[el2_ifu_mem_ctl.scala 479:49]
  wire  _T_2467 = io_ic_error_start & _T_317; // @[el2_ifu_mem_ctl.scala 488:87]
  wire  _T_2481 = io_dec_tlu_flush_err_wb & io_dec_tlu_flush_lower_wb; // @[el2_ifu_mem_ctl.scala 498:54]
  wire  _T_2482 = _T_2481 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 498:84]
  wire  _T_2491 = perr_state == 3'h2; // @[el2_ifu_mem_ctl.scala 519:66]
  wire  _T_2492 = io_dec_tlu_flush_err_wb & _T_2491; // @[el2_ifu_mem_ctl.scala 519:52]
  wire  _T_2494 = _T_2492 & _T_2587; // @[el2_ifu_mem_ctl.scala 519:81]
  wire  _T_2496 = io_dec_tlu_flush_lower_wb | io_dec_tlu_i0_commit_cmt; // @[el2_ifu_mem_ctl.scala 522:59]
  wire  _T_2497 = _T_2496 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 522:86]
  wire  _T_2511 = _T_2496 | io_ifu_fetch_val[0]; // @[el2_ifu_mem_ctl.scala 525:81]
  wire  _T_2512 = _T_2511 | ifu_bp_hit_taken_q_f; // @[el2_ifu_mem_ctl.scala 525:103]
  wire  _T_2513 = _T_2512 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 525:126]
  wire  _T_2533 = _T_2511 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 532:103]
  wire  _T_2540 = ~io_dec_tlu_flush_err_wb; // @[el2_ifu_mem_ctl.scala 537:62]
  wire  _T_2541 = io_dec_tlu_flush_lower_wb & _T_2540; // @[el2_ifu_mem_ctl.scala 537:60]
  wire  _T_2542 = _T_2541 | io_dec_tlu_i0_commit_cmt; // @[el2_ifu_mem_ctl.scala 537:88]
  wire  _T_2543 = _T_2542 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 537:115]
  wire  _GEN_51 = _T_2539 & _T_2497; // @[Conditional.scala 39:67]
  wire  _GEN_54 = _T_2522 ? _T_2533 : _GEN_51; // @[Conditional.scala 39:67]
  wire  _GEN_56 = _T_2522 | _T_2539; // @[Conditional.scala 39:67]
  wire  _GEN_58 = _T_2495 ? _T_2513 : _GEN_54; // @[Conditional.scala 39:67]
  wire  _GEN_60 = _T_2495 | _GEN_56; // @[Conditional.scala 39:67]
  wire  err_stop_state_en = _T_2490 ? _T_2494 : _GEN_58; // @[Conditional.scala 40:58]
  reg  ifu_bus_cmd_valid; // @[Reg.scala 27:20]
  wire  _T_2555 = ic_act_miss_f | ifu_bus_cmd_valid; // @[el2_ifu_mem_ctl.scala 554:64]
  wire  _T_2557 = _T_2555 & _T_2587; // @[el2_ifu_mem_ctl.scala 554:85]
  reg [2:0] bus_cmd_beat_count; // @[Reg.scala 27:20]
  wire  _T_2559 = bus_cmd_beat_count == 3'h7; // @[el2_ifu_mem_ctl.scala 554:133]
  wire  _T_2560 = _T_2559 & ifu_bus_cmd_valid; // @[el2_ifu_mem_ctl.scala 554:164]
  wire  _T_2561 = _T_2560 & io_ifu_axi_arready; // @[el2_ifu_mem_ctl.scala 554:184]
  wire  _T_2562 = _T_2561 & miss_pending; // @[el2_ifu_mem_ctl.scala 554:204]
  wire  _T_2563 = ~_T_2562; // @[el2_ifu_mem_ctl.scala 554:112]
  wire  ifc_bus_ic_req_ff_in = _T_2557 & _T_2563; // @[el2_ifu_mem_ctl.scala 554:110]
  wire  _T_2564 = io_ifu_bus_clk_en | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 555:80]
  wire  ifu_bus_arready = io_ifu_axi_arready & io_ifu_bus_clk_en; // @[el2_ifu_mem_ctl.scala 586:45]
  wire  _T_2581 = io_ifu_axi_arvalid & ifu_bus_arready; // @[el2_ifu_mem_ctl.scala 589:35]
  wire  _T_2582 = _T_2581 & miss_pending; // @[el2_ifu_mem_ctl.scala 589:53]
  wire  bus_cmd_sent = _T_2582 & _T_2587; // @[el2_ifu_mem_ctl.scala 589:68]
  wire [2:0] _T_2572 = ifu_bus_cmd_valid ? 3'h7 : 3'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_2574 = {miss_addr,bus_rd_addr_count,3'h0}; // @[Cat.scala 29:58]
  wire [31:0] _T_2576 = ifu_bus_cmd_valid ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  reg  ifu_bus_arready_unq_ff; // @[Reg.scala 27:20]
  reg  ifu_bus_arvalid_ff; // @[Reg.scala 27:20]
  wire  ifu_bus_arready_ff = ifu_bus_arready_unq_ff & bus_ifu_bus_clk_en_ff; // @[el2_ifu_mem_ctl.scala 587:51]
  wire  _T_2602 = ~scnd_miss_req; // @[el2_ifu_mem_ctl.scala 597:73]
  wire  _T_2603 = _T_2588 & _T_2602; // @[el2_ifu_mem_ctl.scala 597:71]
  wire  _T_2605 = last_data_recieved_ff & _T_1339; // @[el2_ifu_mem_ctl.scala 597:114]
  wire  last_data_recieved_in = _T_2603 | _T_2605; // @[el2_ifu_mem_ctl.scala 597:89]
  wire [2:0] _T_2611 = bus_rd_addr_count + 3'h1; // @[el2_ifu_mem_ctl.scala 602:45]
  wire  _T_2614 = io_ifu_bus_clk_en | ic_act_miss_f; // @[el2_ifu_mem_ctl.scala 603:81]
  wire  _T_2615 = _T_2614 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 603:97]
  wire  _T_2617 = ifu_bus_cmd_valid & io_ifu_axi_arready; // @[el2_ifu_mem_ctl.scala 605:48]
  wire  _T_2618 = _T_2617 & miss_pending; // @[el2_ifu_mem_ctl.scala 605:68]
  wire  bus_inc_cmd_beat_cnt = _T_2618 & _T_2587; // @[el2_ifu_mem_ctl.scala 605:83]
  wire  bus_reset_cmd_beat_cnt_secondlast = ic_act_miss_f & uncacheable_miss_in; // @[el2_ifu_mem_ctl.scala 607:57]
  wire  _T_2622 = ~bus_inc_cmd_beat_cnt; // @[el2_ifu_mem_ctl.scala 608:31]
  wire  _T_2623 = ic_act_miss_f | scnd_miss_req; // @[el2_ifu_mem_ctl.scala 608:71]
  wire  _T_2624 = _T_2623 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 608:87]
  wire  _T_2625 = ~_T_2624; // @[el2_ifu_mem_ctl.scala 608:55]
  wire  bus_hold_cmd_beat_cnt = _T_2622 & _T_2625; // @[el2_ifu_mem_ctl.scala 608:53]
  wire  _T_2626 = bus_inc_cmd_beat_cnt | ic_act_miss_f; // @[el2_ifu_mem_ctl.scala 609:46]
  wire  bus_cmd_beat_en = _T_2626 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 609:62]
  wire [2:0] _T_2629 = bus_cmd_beat_count + 3'h1; // @[el2_ifu_mem_ctl.scala 611:46]
  wire [2:0] _T_2631 = bus_reset_cmd_beat_cnt_secondlast ? 3'h6 : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_2632 = bus_inc_cmd_beat_cnt ? _T_2629 : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_2633 = bus_hold_cmd_beat_cnt ? bus_cmd_beat_count : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_2635 = _T_2631 | _T_2632; // @[Mux.scala 27:72]
  wire [2:0] bus_new_cmd_beat_count = _T_2635 | _T_2633; // @[Mux.scala 27:72]
  wire  _T_2639 = _T_2615 & bus_cmd_beat_en; // @[el2_ifu_mem_ctl.scala 612:125]
  reg  ifc_dma_access_ok_prev; // @[el2_ifu_mem_ctl.scala 623:62]
  wire  _T_2667 = ~iccm_correct_ecc; // @[el2_ifu_mem_ctl.scala 628:50]
  wire  _T_2668 = io_ifc_dma_access_ok & _T_2667; // @[el2_ifu_mem_ctl.scala 628:47]
  wire  _T_2669 = ~io_iccm_dma_sb_error; // @[el2_ifu_mem_ctl.scala 628:70]
  wire  ifc_dma_access_ok_d = _T_2668 & _T_2669; // @[el2_ifu_mem_ctl.scala 628:68]
  wire  _T_2673 = _T_2668 & ifc_dma_access_ok_prev; // @[el2_ifu_mem_ctl.scala 629:72]
  wire  _T_2674 = perr_state == 3'h0; // @[el2_ifu_mem_ctl.scala 629:111]
  wire  _T_2675 = _T_2673 & _T_2674; // @[el2_ifu_mem_ctl.scala 629:97]
  wire  ifc_dma_access_q_ok = _T_2675 & _T_2669; // @[el2_ifu_mem_ctl.scala 629:127]
  wire  _T_2678 = ifc_dma_access_q_ok & io_dma_iccm_req; // @[el2_ifu_mem_ctl.scala 632:40]
  wire  _T_2679 = _T_2678 & io_dma_mem_write; // @[el2_ifu_mem_ctl.scala 632:58]
  wire  _T_2682 = ~io_dma_mem_write; // @[el2_ifu_mem_ctl.scala 633:60]
  wire  _T_2683 = _T_2678 & _T_2682; // @[el2_ifu_mem_ctl.scala 633:58]
  wire  _T_2684 = io_ifc_iccm_access_bf & io_ifc_fetch_req_bf; // @[el2_ifu_mem_ctl.scala 633:104]
  wire [2:0] _T_2689 = io_dma_iccm_req ? 3'h7 : 3'h0; // @[Bitwise.scala 72:12]
  wire  _T_2710 = io_dma_mem_wdata[0] ^ io_dma_mem_wdata[1]; // @[el2_lib.scala 244:74]
  wire  _T_2711 = _T_2710 ^ io_dma_mem_wdata[3]; // @[el2_lib.scala 244:74]
  wire  _T_2712 = _T_2711 ^ io_dma_mem_wdata[4]; // @[el2_lib.scala 244:74]
  wire  _T_2713 = _T_2712 ^ io_dma_mem_wdata[6]; // @[el2_lib.scala 244:74]
  wire  _T_2714 = _T_2713 ^ io_dma_mem_wdata[8]; // @[el2_lib.scala 244:74]
  wire  _T_2715 = _T_2714 ^ io_dma_mem_wdata[10]; // @[el2_lib.scala 244:74]
  wire  _T_2716 = _T_2715 ^ io_dma_mem_wdata[11]; // @[el2_lib.scala 244:74]
  wire  _T_2717 = _T_2716 ^ io_dma_mem_wdata[13]; // @[el2_lib.scala 244:74]
  wire  _T_2718 = _T_2717 ^ io_dma_mem_wdata[15]; // @[el2_lib.scala 244:74]
  wire  _T_2719 = _T_2718 ^ io_dma_mem_wdata[17]; // @[el2_lib.scala 244:74]
  wire  _T_2720 = _T_2719 ^ io_dma_mem_wdata[19]; // @[el2_lib.scala 244:74]
  wire  _T_2721 = _T_2720 ^ io_dma_mem_wdata[21]; // @[el2_lib.scala 244:74]
  wire  _T_2722 = _T_2721 ^ io_dma_mem_wdata[23]; // @[el2_lib.scala 244:74]
  wire  _T_2723 = _T_2722 ^ io_dma_mem_wdata[25]; // @[el2_lib.scala 244:74]
  wire  _T_2724 = _T_2723 ^ io_dma_mem_wdata[26]; // @[el2_lib.scala 244:74]
  wire  _T_2725 = _T_2724 ^ io_dma_mem_wdata[28]; // @[el2_lib.scala 244:74]
  wire  _T_2726 = _T_2725 ^ io_dma_mem_wdata[30]; // @[el2_lib.scala 244:74]
  wire  _T_2745 = io_dma_mem_wdata[0] ^ io_dma_mem_wdata[2]; // @[el2_lib.scala 244:74]
  wire  _T_2746 = _T_2745 ^ io_dma_mem_wdata[3]; // @[el2_lib.scala 244:74]
  wire  _T_2747 = _T_2746 ^ io_dma_mem_wdata[5]; // @[el2_lib.scala 244:74]
  wire  _T_2748 = _T_2747 ^ io_dma_mem_wdata[6]; // @[el2_lib.scala 244:74]
  wire  _T_2749 = _T_2748 ^ io_dma_mem_wdata[9]; // @[el2_lib.scala 244:74]
  wire  _T_2750 = _T_2749 ^ io_dma_mem_wdata[10]; // @[el2_lib.scala 244:74]
  wire  _T_2751 = _T_2750 ^ io_dma_mem_wdata[12]; // @[el2_lib.scala 244:74]
  wire  _T_2752 = _T_2751 ^ io_dma_mem_wdata[13]; // @[el2_lib.scala 244:74]
  wire  _T_2753 = _T_2752 ^ io_dma_mem_wdata[16]; // @[el2_lib.scala 244:74]
  wire  _T_2754 = _T_2753 ^ io_dma_mem_wdata[17]; // @[el2_lib.scala 244:74]
  wire  _T_2755 = _T_2754 ^ io_dma_mem_wdata[20]; // @[el2_lib.scala 244:74]
  wire  _T_2756 = _T_2755 ^ io_dma_mem_wdata[21]; // @[el2_lib.scala 244:74]
  wire  _T_2757 = _T_2756 ^ io_dma_mem_wdata[24]; // @[el2_lib.scala 244:74]
  wire  _T_2758 = _T_2757 ^ io_dma_mem_wdata[25]; // @[el2_lib.scala 244:74]
  wire  _T_2759 = _T_2758 ^ io_dma_mem_wdata[27]; // @[el2_lib.scala 244:74]
  wire  _T_2760 = _T_2759 ^ io_dma_mem_wdata[28]; // @[el2_lib.scala 244:74]
  wire  _T_2761 = _T_2760 ^ io_dma_mem_wdata[31]; // @[el2_lib.scala 244:74]
  wire  _T_2780 = io_dma_mem_wdata[1] ^ io_dma_mem_wdata[2]; // @[el2_lib.scala 244:74]
  wire  _T_2781 = _T_2780 ^ io_dma_mem_wdata[3]; // @[el2_lib.scala 244:74]
  wire  _T_2782 = _T_2781 ^ io_dma_mem_wdata[7]; // @[el2_lib.scala 244:74]
  wire  _T_2783 = _T_2782 ^ io_dma_mem_wdata[8]; // @[el2_lib.scala 244:74]
  wire  _T_2784 = _T_2783 ^ io_dma_mem_wdata[9]; // @[el2_lib.scala 244:74]
  wire  _T_2785 = _T_2784 ^ io_dma_mem_wdata[10]; // @[el2_lib.scala 244:74]
  wire  _T_2786 = _T_2785 ^ io_dma_mem_wdata[14]; // @[el2_lib.scala 244:74]
  wire  _T_2787 = _T_2786 ^ io_dma_mem_wdata[15]; // @[el2_lib.scala 244:74]
  wire  _T_2788 = _T_2787 ^ io_dma_mem_wdata[16]; // @[el2_lib.scala 244:74]
  wire  _T_2789 = _T_2788 ^ io_dma_mem_wdata[17]; // @[el2_lib.scala 244:74]
  wire  _T_2790 = _T_2789 ^ io_dma_mem_wdata[22]; // @[el2_lib.scala 244:74]
  wire  _T_2791 = _T_2790 ^ io_dma_mem_wdata[23]; // @[el2_lib.scala 244:74]
  wire  _T_2792 = _T_2791 ^ io_dma_mem_wdata[24]; // @[el2_lib.scala 244:74]
  wire  _T_2793 = _T_2792 ^ io_dma_mem_wdata[25]; // @[el2_lib.scala 244:74]
  wire  _T_2794 = _T_2793 ^ io_dma_mem_wdata[29]; // @[el2_lib.scala 244:74]
  wire  _T_2795 = _T_2794 ^ io_dma_mem_wdata[30]; // @[el2_lib.scala 244:74]
  wire  _T_2796 = _T_2795 ^ io_dma_mem_wdata[31]; // @[el2_lib.scala 244:74]
  wire  _T_2812 = io_dma_mem_wdata[4] ^ io_dma_mem_wdata[5]; // @[el2_lib.scala 244:74]
  wire  _T_2813 = _T_2812 ^ io_dma_mem_wdata[6]; // @[el2_lib.scala 244:74]
  wire  _T_2814 = _T_2813 ^ io_dma_mem_wdata[7]; // @[el2_lib.scala 244:74]
  wire  _T_2815 = _T_2814 ^ io_dma_mem_wdata[8]; // @[el2_lib.scala 244:74]
  wire  _T_2816 = _T_2815 ^ io_dma_mem_wdata[9]; // @[el2_lib.scala 244:74]
  wire  _T_2817 = _T_2816 ^ io_dma_mem_wdata[10]; // @[el2_lib.scala 244:74]
  wire  _T_2818 = _T_2817 ^ io_dma_mem_wdata[18]; // @[el2_lib.scala 244:74]
  wire  _T_2819 = _T_2818 ^ io_dma_mem_wdata[19]; // @[el2_lib.scala 244:74]
  wire  _T_2820 = _T_2819 ^ io_dma_mem_wdata[20]; // @[el2_lib.scala 244:74]
  wire  _T_2821 = _T_2820 ^ io_dma_mem_wdata[21]; // @[el2_lib.scala 244:74]
  wire  _T_2822 = _T_2821 ^ io_dma_mem_wdata[22]; // @[el2_lib.scala 244:74]
  wire  _T_2823 = _T_2822 ^ io_dma_mem_wdata[23]; // @[el2_lib.scala 244:74]
  wire  _T_2824 = _T_2823 ^ io_dma_mem_wdata[24]; // @[el2_lib.scala 244:74]
  wire  _T_2825 = _T_2824 ^ io_dma_mem_wdata[25]; // @[el2_lib.scala 244:74]
  wire  _T_2841 = io_dma_mem_wdata[11] ^ io_dma_mem_wdata[12]; // @[el2_lib.scala 244:74]
  wire  _T_2842 = _T_2841 ^ io_dma_mem_wdata[13]; // @[el2_lib.scala 244:74]
  wire  _T_2843 = _T_2842 ^ io_dma_mem_wdata[14]; // @[el2_lib.scala 244:74]
  wire  _T_2844 = _T_2843 ^ io_dma_mem_wdata[15]; // @[el2_lib.scala 244:74]
  wire  _T_2845 = _T_2844 ^ io_dma_mem_wdata[16]; // @[el2_lib.scala 244:74]
  wire  _T_2846 = _T_2845 ^ io_dma_mem_wdata[17]; // @[el2_lib.scala 244:74]
  wire  _T_2847 = _T_2846 ^ io_dma_mem_wdata[18]; // @[el2_lib.scala 244:74]
  wire  _T_2848 = _T_2847 ^ io_dma_mem_wdata[19]; // @[el2_lib.scala 244:74]
  wire  _T_2849 = _T_2848 ^ io_dma_mem_wdata[20]; // @[el2_lib.scala 244:74]
  wire  _T_2850 = _T_2849 ^ io_dma_mem_wdata[21]; // @[el2_lib.scala 244:74]
  wire  _T_2851 = _T_2850 ^ io_dma_mem_wdata[22]; // @[el2_lib.scala 244:74]
  wire  _T_2852 = _T_2851 ^ io_dma_mem_wdata[23]; // @[el2_lib.scala 244:74]
  wire  _T_2853 = _T_2852 ^ io_dma_mem_wdata[24]; // @[el2_lib.scala 244:74]
  wire  _T_2854 = _T_2853 ^ io_dma_mem_wdata[25]; // @[el2_lib.scala 244:74]
  wire  _T_2861 = io_dma_mem_wdata[26] ^ io_dma_mem_wdata[27]; // @[el2_lib.scala 244:74]
  wire  _T_2862 = _T_2861 ^ io_dma_mem_wdata[28]; // @[el2_lib.scala 244:74]
  wire  _T_2863 = _T_2862 ^ io_dma_mem_wdata[29]; // @[el2_lib.scala 244:74]
  wire  _T_2864 = _T_2863 ^ io_dma_mem_wdata[30]; // @[el2_lib.scala 244:74]
  wire  _T_2865 = _T_2864 ^ io_dma_mem_wdata[31]; // @[el2_lib.scala 244:74]
  wire [5:0] _T_2870 = {_T_2865,_T_2854,_T_2825,_T_2796,_T_2761,_T_2726}; // @[Cat.scala 29:58]
  wire  _T_2871 = ^io_dma_mem_wdata[31:0]; // @[el2_lib.scala 252:13]
  wire  _T_2872 = ^_T_2870; // @[el2_lib.scala 252:23]
  wire  _T_2873 = _T_2871 ^ _T_2872; // @[el2_lib.scala 252:18]
  wire [6:0] _T_2874 = {_T_2873,_T_2865,_T_2854,_T_2825,_T_2796,_T_2761,_T_2726}; // @[Cat.scala 29:58]
  wire  _T_2894 = io_dma_mem_wdata[32] ^ io_dma_mem_wdata[33]; // @[el2_lib.scala 244:74]
  wire  _T_2895 = _T_2894 ^ io_dma_mem_wdata[35]; // @[el2_lib.scala 244:74]
  wire  _T_2896 = _T_2895 ^ io_dma_mem_wdata[36]; // @[el2_lib.scala 244:74]
  wire  _T_2897 = _T_2896 ^ io_dma_mem_wdata[38]; // @[el2_lib.scala 244:74]
  wire  _T_2898 = _T_2897 ^ io_dma_mem_wdata[40]; // @[el2_lib.scala 244:74]
  wire  _T_2899 = _T_2898 ^ io_dma_mem_wdata[42]; // @[el2_lib.scala 244:74]
  wire  _T_2900 = _T_2899 ^ io_dma_mem_wdata[43]; // @[el2_lib.scala 244:74]
  wire  _T_2901 = _T_2900 ^ io_dma_mem_wdata[45]; // @[el2_lib.scala 244:74]
  wire  _T_2902 = _T_2901 ^ io_dma_mem_wdata[47]; // @[el2_lib.scala 244:74]
  wire  _T_2903 = _T_2902 ^ io_dma_mem_wdata[49]; // @[el2_lib.scala 244:74]
  wire  _T_2904 = _T_2903 ^ io_dma_mem_wdata[51]; // @[el2_lib.scala 244:74]
  wire  _T_2905 = _T_2904 ^ io_dma_mem_wdata[53]; // @[el2_lib.scala 244:74]
  wire  _T_2906 = _T_2905 ^ io_dma_mem_wdata[55]; // @[el2_lib.scala 244:74]
  wire  _T_2907 = _T_2906 ^ io_dma_mem_wdata[57]; // @[el2_lib.scala 244:74]
  wire  _T_2908 = _T_2907 ^ io_dma_mem_wdata[58]; // @[el2_lib.scala 244:74]
  wire  _T_2909 = _T_2908 ^ io_dma_mem_wdata[60]; // @[el2_lib.scala 244:74]
  wire  _T_2910 = _T_2909 ^ io_dma_mem_wdata[62]; // @[el2_lib.scala 244:74]
  wire  _T_2929 = io_dma_mem_wdata[32] ^ io_dma_mem_wdata[34]; // @[el2_lib.scala 244:74]
  wire  _T_2930 = _T_2929 ^ io_dma_mem_wdata[35]; // @[el2_lib.scala 244:74]
  wire  _T_2931 = _T_2930 ^ io_dma_mem_wdata[37]; // @[el2_lib.scala 244:74]
  wire  _T_2932 = _T_2931 ^ io_dma_mem_wdata[38]; // @[el2_lib.scala 244:74]
  wire  _T_2933 = _T_2932 ^ io_dma_mem_wdata[41]; // @[el2_lib.scala 244:74]
  wire  _T_2934 = _T_2933 ^ io_dma_mem_wdata[42]; // @[el2_lib.scala 244:74]
  wire  _T_2935 = _T_2934 ^ io_dma_mem_wdata[44]; // @[el2_lib.scala 244:74]
  wire  _T_2936 = _T_2935 ^ io_dma_mem_wdata[45]; // @[el2_lib.scala 244:74]
  wire  _T_2937 = _T_2936 ^ io_dma_mem_wdata[48]; // @[el2_lib.scala 244:74]
  wire  _T_2938 = _T_2937 ^ io_dma_mem_wdata[49]; // @[el2_lib.scala 244:74]
  wire  _T_2939 = _T_2938 ^ io_dma_mem_wdata[52]; // @[el2_lib.scala 244:74]
  wire  _T_2940 = _T_2939 ^ io_dma_mem_wdata[53]; // @[el2_lib.scala 244:74]
  wire  _T_2941 = _T_2940 ^ io_dma_mem_wdata[56]; // @[el2_lib.scala 244:74]
  wire  _T_2942 = _T_2941 ^ io_dma_mem_wdata[57]; // @[el2_lib.scala 244:74]
  wire  _T_2943 = _T_2942 ^ io_dma_mem_wdata[59]; // @[el2_lib.scala 244:74]
  wire  _T_2944 = _T_2943 ^ io_dma_mem_wdata[60]; // @[el2_lib.scala 244:74]
  wire  _T_2945 = _T_2944 ^ io_dma_mem_wdata[63]; // @[el2_lib.scala 244:74]
  wire  _T_2964 = io_dma_mem_wdata[33] ^ io_dma_mem_wdata[34]; // @[el2_lib.scala 244:74]
  wire  _T_2965 = _T_2964 ^ io_dma_mem_wdata[35]; // @[el2_lib.scala 244:74]
  wire  _T_2966 = _T_2965 ^ io_dma_mem_wdata[39]; // @[el2_lib.scala 244:74]
  wire  _T_2967 = _T_2966 ^ io_dma_mem_wdata[40]; // @[el2_lib.scala 244:74]
  wire  _T_2968 = _T_2967 ^ io_dma_mem_wdata[41]; // @[el2_lib.scala 244:74]
  wire  _T_2969 = _T_2968 ^ io_dma_mem_wdata[42]; // @[el2_lib.scala 244:74]
  wire  _T_2970 = _T_2969 ^ io_dma_mem_wdata[46]; // @[el2_lib.scala 244:74]
  wire  _T_2971 = _T_2970 ^ io_dma_mem_wdata[47]; // @[el2_lib.scala 244:74]
  wire  _T_2972 = _T_2971 ^ io_dma_mem_wdata[48]; // @[el2_lib.scala 244:74]
  wire  _T_2973 = _T_2972 ^ io_dma_mem_wdata[49]; // @[el2_lib.scala 244:74]
  wire  _T_2974 = _T_2973 ^ io_dma_mem_wdata[54]; // @[el2_lib.scala 244:74]
  wire  _T_2975 = _T_2974 ^ io_dma_mem_wdata[55]; // @[el2_lib.scala 244:74]
  wire  _T_2976 = _T_2975 ^ io_dma_mem_wdata[56]; // @[el2_lib.scala 244:74]
  wire  _T_2977 = _T_2976 ^ io_dma_mem_wdata[57]; // @[el2_lib.scala 244:74]
  wire  _T_2978 = _T_2977 ^ io_dma_mem_wdata[61]; // @[el2_lib.scala 244:74]
  wire  _T_2979 = _T_2978 ^ io_dma_mem_wdata[62]; // @[el2_lib.scala 244:74]
  wire  _T_2980 = _T_2979 ^ io_dma_mem_wdata[63]; // @[el2_lib.scala 244:74]
  wire  _T_2996 = io_dma_mem_wdata[36] ^ io_dma_mem_wdata[37]; // @[el2_lib.scala 244:74]
  wire  _T_2997 = _T_2996 ^ io_dma_mem_wdata[38]; // @[el2_lib.scala 244:74]
  wire  _T_2998 = _T_2997 ^ io_dma_mem_wdata[39]; // @[el2_lib.scala 244:74]
  wire  _T_2999 = _T_2998 ^ io_dma_mem_wdata[40]; // @[el2_lib.scala 244:74]
  wire  _T_3000 = _T_2999 ^ io_dma_mem_wdata[41]; // @[el2_lib.scala 244:74]
  wire  _T_3001 = _T_3000 ^ io_dma_mem_wdata[42]; // @[el2_lib.scala 244:74]
  wire  _T_3002 = _T_3001 ^ io_dma_mem_wdata[50]; // @[el2_lib.scala 244:74]
  wire  _T_3003 = _T_3002 ^ io_dma_mem_wdata[51]; // @[el2_lib.scala 244:74]
  wire  _T_3004 = _T_3003 ^ io_dma_mem_wdata[52]; // @[el2_lib.scala 244:74]
  wire  _T_3005 = _T_3004 ^ io_dma_mem_wdata[53]; // @[el2_lib.scala 244:74]
  wire  _T_3006 = _T_3005 ^ io_dma_mem_wdata[54]; // @[el2_lib.scala 244:74]
  wire  _T_3007 = _T_3006 ^ io_dma_mem_wdata[55]; // @[el2_lib.scala 244:74]
  wire  _T_3008 = _T_3007 ^ io_dma_mem_wdata[56]; // @[el2_lib.scala 244:74]
  wire  _T_3009 = _T_3008 ^ io_dma_mem_wdata[57]; // @[el2_lib.scala 244:74]
  wire  _T_3025 = io_dma_mem_wdata[43] ^ io_dma_mem_wdata[44]; // @[el2_lib.scala 244:74]
  wire  _T_3026 = _T_3025 ^ io_dma_mem_wdata[45]; // @[el2_lib.scala 244:74]
  wire  _T_3027 = _T_3026 ^ io_dma_mem_wdata[46]; // @[el2_lib.scala 244:74]
  wire  _T_3028 = _T_3027 ^ io_dma_mem_wdata[47]; // @[el2_lib.scala 244:74]
  wire  _T_3029 = _T_3028 ^ io_dma_mem_wdata[48]; // @[el2_lib.scala 244:74]
  wire  _T_3030 = _T_3029 ^ io_dma_mem_wdata[49]; // @[el2_lib.scala 244:74]
  wire  _T_3031 = _T_3030 ^ io_dma_mem_wdata[50]; // @[el2_lib.scala 244:74]
  wire  _T_3032 = _T_3031 ^ io_dma_mem_wdata[51]; // @[el2_lib.scala 244:74]
  wire  _T_3033 = _T_3032 ^ io_dma_mem_wdata[52]; // @[el2_lib.scala 244:74]
  wire  _T_3034 = _T_3033 ^ io_dma_mem_wdata[53]; // @[el2_lib.scala 244:74]
  wire  _T_3035 = _T_3034 ^ io_dma_mem_wdata[54]; // @[el2_lib.scala 244:74]
  wire  _T_3036 = _T_3035 ^ io_dma_mem_wdata[55]; // @[el2_lib.scala 244:74]
  wire  _T_3037 = _T_3036 ^ io_dma_mem_wdata[56]; // @[el2_lib.scala 244:74]
  wire  _T_3038 = _T_3037 ^ io_dma_mem_wdata[57]; // @[el2_lib.scala 244:74]
  wire  _T_3045 = io_dma_mem_wdata[58] ^ io_dma_mem_wdata[59]; // @[el2_lib.scala 244:74]
  wire  _T_3046 = _T_3045 ^ io_dma_mem_wdata[60]; // @[el2_lib.scala 244:74]
  wire  _T_3047 = _T_3046 ^ io_dma_mem_wdata[61]; // @[el2_lib.scala 244:74]
  wire  _T_3048 = _T_3047 ^ io_dma_mem_wdata[62]; // @[el2_lib.scala 244:74]
  wire  _T_3049 = _T_3048 ^ io_dma_mem_wdata[63]; // @[el2_lib.scala 244:74]
  wire [5:0] _T_3054 = {_T_3049,_T_3038,_T_3009,_T_2980,_T_2945,_T_2910}; // @[Cat.scala 29:58]
  wire  _T_3055 = ^io_dma_mem_wdata[63:32]; // @[el2_lib.scala 252:13]
  wire  _T_3056 = ^_T_3054; // @[el2_lib.scala 252:23]
  wire  _T_3057 = _T_3055 ^ _T_3056; // @[el2_lib.scala 252:18]
  wire [13:0] dma_mem_ecc = {_T_3057,_T_3049,_T_3038,_T_3009,_T_2980,_T_2945,_T_2910,_T_2874}; // @[Cat.scala 29:58]
  wire  _T_3244 = ~_T_2678; // @[el2_ifu_mem_ctl.scala 639:45]
  wire  _T_3245 = iccm_correct_ecc & _T_3244; // @[el2_ifu_mem_ctl.scala 639:43]
  reg [38:0] iccm_ecc_corr_data_ff; // @[Reg.scala 27:20]
  wire [77:0] _T_3246 = {iccm_ecc_corr_data_ff,iccm_ecc_corr_data_ff}; // @[Cat.scala 29:58]
  wire [77:0] _T_3253 = {dma_mem_ecc[13:7],io_dma_mem_wdata[63:32],dma_mem_ecc[6:0],io_dma_mem_wdata[31:0]}; // @[Cat.scala 29:58]
  reg [1:0] dma_mem_addr_ff; // @[el2_ifu_mem_ctl.scala 653:53]
  wire  _T_3586 = _T_3498[5:0] == 6'h27; // @[el2_lib.scala 324:41]
  wire  _T_3584 = _T_3498[5:0] == 6'h26; // @[el2_lib.scala 324:41]
  wire  _T_3582 = _T_3498[5:0] == 6'h25; // @[el2_lib.scala 324:41]
  wire  _T_3580 = _T_3498[5:0] == 6'h24; // @[el2_lib.scala 324:41]
  wire  _T_3578 = _T_3498[5:0] == 6'h23; // @[el2_lib.scala 324:41]
  wire  _T_3576 = _T_3498[5:0] == 6'h22; // @[el2_lib.scala 324:41]
  wire  _T_3574 = _T_3498[5:0] == 6'h21; // @[el2_lib.scala 324:41]
  wire  _T_3572 = _T_3498[5:0] == 6'h20; // @[el2_lib.scala 324:41]
  wire  _T_3570 = _T_3498[5:0] == 6'h1f; // @[el2_lib.scala 324:41]
  wire  _T_3568 = _T_3498[5:0] == 6'h1e; // @[el2_lib.scala 324:41]
  wire [9:0] _T_3644 = {_T_3586,_T_3584,_T_3582,_T_3580,_T_3578,_T_3576,_T_3574,_T_3572,_T_3570,_T_3568}; // @[el2_lib.scala 327:69]
  wire  _T_3566 = _T_3498[5:0] == 6'h1d; // @[el2_lib.scala 324:41]
  wire  _T_3564 = _T_3498[5:0] == 6'h1c; // @[el2_lib.scala 324:41]
  wire  _T_3562 = _T_3498[5:0] == 6'h1b; // @[el2_lib.scala 324:41]
  wire  _T_3560 = _T_3498[5:0] == 6'h1a; // @[el2_lib.scala 324:41]
  wire  _T_3558 = _T_3498[5:0] == 6'h19; // @[el2_lib.scala 324:41]
  wire  _T_3556 = _T_3498[5:0] == 6'h18; // @[el2_lib.scala 324:41]
  wire  _T_3554 = _T_3498[5:0] == 6'h17; // @[el2_lib.scala 324:41]
  wire  _T_3552 = _T_3498[5:0] == 6'h16; // @[el2_lib.scala 324:41]
  wire  _T_3550 = _T_3498[5:0] == 6'h15; // @[el2_lib.scala 324:41]
  wire  _T_3548 = _T_3498[5:0] == 6'h14; // @[el2_lib.scala 324:41]
  wire [9:0] _T_3635 = {_T_3566,_T_3564,_T_3562,_T_3560,_T_3558,_T_3556,_T_3554,_T_3552,_T_3550,_T_3548}; // @[el2_lib.scala 327:69]
  wire  _T_3546 = _T_3498[5:0] == 6'h13; // @[el2_lib.scala 324:41]
  wire  _T_3544 = _T_3498[5:0] == 6'h12; // @[el2_lib.scala 324:41]
  wire  _T_3542 = _T_3498[5:0] == 6'h11; // @[el2_lib.scala 324:41]
  wire  _T_3540 = _T_3498[5:0] == 6'h10; // @[el2_lib.scala 324:41]
  wire  _T_3538 = _T_3498[5:0] == 6'hf; // @[el2_lib.scala 324:41]
  wire  _T_3536 = _T_3498[5:0] == 6'he; // @[el2_lib.scala 324:41]
  wire  _T_3534 = _T_3498[5:0] == 6'hd; // @[el2_lib.scala 324:41]
  wire  _T_3532 = _T_3498[5:0] == 6'hc; // @[el2_lib.scala 324:41]
  wire  _T_3530 = _T_3498[5:0] == 6'hb; // @[el2_lib.scala 324:41]
  wire  _T_3528 = _T_3498[5:0] == 6'ha; // @[el2_lib.scala 324:41]
  wire [9:0] _T_3625 = {_T_3546,_T_3544,_T_3542,_T_3540,_T_3538,_T_3536,_T_3534,_T_3532,_T_3530,_T_3528}; // @[el2_lib.scala 327:69]
  wire  _T_3526 = _T_3498[5:0] == 6'h9; // @[el2_lib.scala 324:41]
  wire  _T_3524 = _T_3498[5:0] == 6'h8; // @[el2_lib.scala 324:41]
  wire  _T_3522 = _T_3498[5:0] == 6'h7; // @[el2_lib.scala 324:41]
  wire  _T_3520 = _T_3498[5:0] == 6'h6; // @[el2_lib.scala 324:41]
  wire  _T_3518 = _T_3498[5:0] == 6'h5; // @[el2_lib.scala 324:41]
  wire  _T_3516 = _T_3498[5:0] == 6'h4; // @[el2_lib.scala 324:41]
  wire  _T_3514 = _T_3498[5:0] == 6'h3; // @[el2_lib.scala 324:41]
  wire  _T_3512 = _T_3498[5:0] == 6'h2; // @[el2_lib.scala 324:41]
  wire  _T_3510 = _T_3498[5:0] == 6'h1; // @[el2_lib.scala 324:41]
  wire [18:0] _T_3626 = {_T_3625,_T_3526,_T_3524,_T_3522,_T_3520,_T_3518,_T_3516,_T_3514,_T_3512,_T_3510}; // @[el2_lib.scala 327:69]
  wire [38:0] _T_3646 = {_T_3644,_T_3635,_T_3626}; // @[el2_lib.scala 327:69]
  wire [7:0] _T_3601 = {io_iccm_rd_data_ecc[35],io_iccm_rd_data_ecc[3:1],io_iccm_rd_data_ecc[34],io_iccm_rd_data_ecc[0],io_iccm_rd_data_ecc[33:32]}; // @[Cat.scala 29:58]
  wire [38:0] _T_3607 = {io_iccm_rd_data_ecc[38],io_iccm_rd_data_ecc[31:26],io_iccm_rd_data_ecc[37],io_iccm_rd_data_ecc[25:11],io_iccm_rd_data_ecc[36],io_iccm_rd_data_ecc[10:4],_T_3601}; // @[Cat.scala 29:58]
  wire [38:0] _T_3647 = _T_3646 ^ _T_3607; // @[el2_lib.scala 327:76]
  wire [38:0] _T_3648 = _T_3502 ? _T_3647 : _T_3607; // @[el2_lib.scala 327:31]
  wire [31:0] iccm_corrected_data_0 = {_T_3648[37:32],_T_3648[30:16],_T_3648[14:8],_T_3648[6:4],_T_3648[2]}; // @[Cat.scala 29:58]
  wire  _T_3971 = _T_3883[5:0] == 6'h27; // @[el2_lib.scala 324:41]
  wire  _T_3969 = _T_3883[5:0] == 6'h26; // @[el2_lib.scala 324:41]
  wire  _T_3967 = _T_3883[5:0] == 6'h25; // @[el2_lib.scala 324:41]
  wire  _T_3965 = _T_3883[5:0] == 6'h24; // @[el2_lib.scala 324:41]
  wire  _T_3963 = _T_3883[5:0] == 6'h23; // @[el2_lib.scala 324:41]
  wire  _T_3961 = _T_3883[5:0] == 6'h22; // @[el2_lib.scala 324:41]
  wire  _T_3959 = _T_3883[5:0] == 6'h21; // @[el2_lib.scala 324:41]
  wire  _T_3957 = _T_3883[5:0] == 6'h20; // @[el2_lib.scala 324:41]
  wire  _T_3955 = _T_3883[5:0] == 6'h1f; // @[el2_lib.scala 324:41]
  wire  _T_3953 = _T_3883[5:0] == 6'h1e; // @[el2_lib.scala 324:41]
  wire [9:0] _T_4029 = {_T_3971,_T_3969,_T_3967,_T_3965,_T_3963,_T_3961,_T_3959,_T_3957,_T_3955,_T_3953}; // @[el2_lib.scala 327:69]
  wire  _T_3951 = _T_3883[5:0] == 6'h1d; // @[el2_lib.scala 324:41]
  wire  _T_3949 = _T_3883[5:0] == 6'h1c; // @[el2_lib.scala 324:41]
  wire  _T_3947 = _T_3883[5:0] == 6'h1b; // @[el2_lib.scala 324:41]
  wire  _T_3945 = _T_3883[5:0] == 6'h1a; // @[el2_lib.scala 324:41]
  wire  _T_3943 = _T_3883[5:0] == 6'h19; // @[el2_lib.scala 324:41]
  wire  _T_3941 = _T_3883[5:0] == 6'h18; // @[el2_lib.scala 324:41]
  wire  _T_3939 = _T_3883[5:0] == 6'h17; // @[el2_lib.scala 324:41]
  wire  _T_3937 = _T_3883[5:0] == 6'h16; // @[el2_lib.scala 324:41]
  wire  _T_3935 = _T_3883[5:0] == 6'h15; // @[el2_lib.scala 324:41]
  wire  _T_3933 = _T_3883[5:0] == 6'h14; // @[el2_lib.scala 324:41]
  wire [9:0] _T_4020 = {_T_3951,_T_3949,_T_3947,_T_3945,_T_3943,_T_3941,_T_3939,_T_3937,_T_3935,_T_3933}; // @[el2_lib.scala 327:69]
  wire  _T_3931 = _T_3883[5:0] == 6'h13; // @[el2_lib.scala 324:41]
  wire  _T_3929 = _T_3883[5:0] == 6'h12; // @[el2_lib.scala 324:41]
  wire  _T_3927 = _T_3883[5:0] == 6'h11; // @[el2_lib.scala 324:41]
  wire  _T_3925 = _T_3883[5:0] == 6'h10; // @[el2_lib.scala 324:41]
  wire  _T_3923 = _T_3883[5:0] == 6'hf; // @[el2_lib.scala 324:41]
  wire  _T_3921 = _T_3883[5:0] == 6'he; // @[el2_lib.scala 324:41]
  wire  _T_3919 = _T_3883[5:0] == 6'hd; // @[el2_lib.scala 324:41]
  wire  _T_3917 = _T_3883[5:0] == 6'hc; // @[el2_lib.scala 324:41]
  wire  _T_3915 = _T_3883[5:0] == 6'hb; // @[el2_lib.scala 324:41]
  wire  _T_3913 = _T_3883[5:0] == 6'ha; // @[el2_lib.scala 324:41]
  wire [9:0] _T_4010 = {_T_3931,_T_3929,_T_3927,_T_3925,_T_3923,_T_3921,_T_3919,_T_3917,_T_3915,_T_3913}; // @[el2_lib.scala 327:69]
  wire  _T_3911 = _T_3883[5:0] == 6'h9; // @[el2_lib.scala 324:41]
  wire  _T_3909 = _T_3883[5:0] == 6'h8; // @[el2_lib.scala 324:41]
  wire  _T_3907 = _T_3883[5:0] == 6'h7; // @[el2_lib.scala 324:41]
  wire  _T_3905 = _T_3883[5:0] == 6'h6; // @[el2_lib.scala 324:41]
  wire  _T_3903 = _T_3883[5:0] == 6'h5; // @[el2_lib.scala 324:41]
  wire  _T_3901 = _T_3883[5:0] == 6'h4; // @[el2_lib.scala 324:41]
  wire  _T_3899 = _T_3883[5:0] == 6'h3; // @[el2_lib.scala 324:41]
  wire  _T_3897 = _T_3883[5:0] == 6'h2; // @[el2_lib.scala 324:41]
  wire  _T_3895 = _T_3883[5:0] == 6'h1; // @[el2_lib.scala 324:41]
  wire [18:0] _T_4011 = {_T_4010,_T_3911,_T_3909,_T_3907,_T_3905,_T_3903,_T_3901,_T_3899,_T_3897,_T_3895}; // @[el2_lib.scala 327:69]
  wire [38:0] _T_4031 = {_T_4029,_T_4020,_T_4011}; // @[el2_lib.scala 327:69]
  wire [7:0] _T_3986 = {io_iccm_rd_data_ecc[74],io_iccm_rd_data_ecc[42:40],io_iccm_rd_data_ecc[73],io_iccm_rd_data_ecc[39],io_iccm_rd_data_ecc[72:71]}; // @[Cat.scala 29:58]
  wire [38:0] _T_3992 = {io_iccm_rd_data_ecc[77],io_iccm_rd_data_ecc[70:65],io_iccm_rd_data_ecc[76],io_iccm_rd_data_ecc[64:50],io_iccm_rd_data_ecc[75],io_iccm_rd_data_ecc[49:43],_T_3986}; // @[Cat.scala 29:58]
  wire [38:0] _T_4032 = _T_4031 ^ _T_3992; // @[el2_lib.scala 327:76]
  wire [38:0] _T_4033 = _T_3887 ? _T_4032 : _T_3992; // @[el2_lib.scala 327:31]
  wire [31:0] iccm_corrected_data_1 = {_T_4033[37:32],_T_4033[30:16],_T_4033[14:8],_T_4033[6:4],_T_4033[2]}; // @[Cat.scala 29:58]
  wire [31:0] iccm_dma_rdata_1_muxed = dma_mem_addr_ff[0] ? iccm_corrected_data_0 : iccm_corrected_data_1; // @[el2_ifu_mem_ctl.scala 645:35]
  wire  _T_3506 = ~_T_3498[6]; // @[el2_lib.scala 320:55]
  wire  _T_3507 = _T_3500 & _T_3506; // @[el2_lib.scala 320:53]
  wire  _T_3891 = ~_T_3883[6]; // @[el2_lib.scala 320:55]
  wire  _T_3892 = _T_3885 & _T_3891; // @[el2_lib.scala 320:53]
  wire [1:0] iccm_double_ecc_error = {_T_3507,_T_3892}; // @[Cat.scala 29:58]
  wire  iccm_dma_ecc_error_in = |iccm_double_ecc_error; // @[el2_ifu_mem_ctl.scala 647:53]
  wire [63:0] _T_3257 = {io_dma_mem_addr,io_dma_mem_addr}; // @[Cat.scala 29:58]
  wire [63:0] _T_3258 = {iccm_dma_rdata_1_muxed,_T_3648[37:32],_T_3648[30:16],_T_3648[14:8],_T_3648[6:4],_T_3648[2]}; // @[Cat.scala 29:58]
  reg [2:0] dma_mem_tag_ff; // @[el2_ifu_mem_ctl.scala 649:54]
  reg [2:0] iccm_dma_rtag_temp; // @[el2_ifu_mem_ctl.scala 650:74]
  reg  iccm_dma_rvalid_temp; // @[el2_ifu_mem_ctl.scala 655:76]
  reg [63:0] iccm_dma_rdata_temp; // @[el2_ifu_mem_ctl.scala 659:75]
  wire  _T_3263 = _T_2678 & _T_2667; // @[el2_ifu_mem_ctl.scala 662:65]
  wire  _T_3267 = _T_3244 & iccm_correct_ecc; // @[el2_ifu_mem_ctl.scala 663:50]
  reg [13:0] iccm_ecc_corr_index_ff; // @[Reg.scala 27:20]
  wire [14:0] _T_3268 = {iccm_ecc_corr_index_ff,1'h0}; // @[Cat.scala 29:58]
  wire [14:0] _T_3270 = _T_3267 ? _T_3268 : io_ifc_fetch_addr_bf[14:0]; // @[el2_ifu_mem_ctl.scala 663:8]
  wire  _T_3660 = _T_3498 == 7'h40; // @[el2_lib.scala 330:62]
  wire  _T_3661 = _T_3648[38] ^ _T_3660; // @[el2_lib.scala 330:44]
  wire [6:0] iccm_corrected_ecc_0 = {_T_3661,_T_3648[31],_T_3648[15],_T_3648[7],_T_3648[3],_T_3648[1:0]}; // @[Cat.scala 29:58]
  wire  _T_4045 = _T_3883 == 7'h40; // @[el2_lib.scala 330:62]
  wire  _T_4046 = _T_4033[38] ^ _T_4045; // @[el2_lib.scala 330:44]
  wire [6:0] iccm_corrected_ecc_1 = {_T_4046,_T_4033[31],_T_4033[15],_T_4033[7],_T_4033[3],_T_4033[1:0]}; // @[Cat.scala 29:58]
  wire  _T_4062 = _T_3 & ifc_iccm_access_f; // @[el2_ifu_mem_ctl.scala 675:58]
  wire [31:0] iccm_corrected_data_f_mux = iccm_single_ecc_error[0] ? iccm_corrected_data_0 : iccm_corrected_data_1; // @[el2_ifu_mem_ctl.scala 677:38]
  wire [6:0] iccm_corrected_ecc_f_mux = iccm_single_ecc_error[0] ? iccm_corrected_ecc_0 : iccm_corrected_ecc_1; // @[el2_ifu_mem_ctl.scala 678:37]
  reg  iccm_rd_ecc_single_err_ff; // @[el2_ifu_mem_ctl.scala 686:62]
  wire  _T_4070 = ~iccm_rd_ecc_single_err_ff; // @[el2_ifu_mem_ctl.scala 680:76]
  wire  _T_4071 = io_iccm_rd_ecc_single_err & _T_4070; // @[el2_ifu_mem_ctl.scala 680:74]
  wire  _T_4073 = _T_4071 & _T_317; // @[el2_ifu_mem_ctl.scala 680:104]
  wire  iccm_ecc_write_status = _T_4073 | io_iccm_dma_sb_error; // @[el2_ifu_mem_ctl.scala 680:127]
  wire  _T_4074 = io_iccm_rd_ecc_single_err | iccm_rd_ecc_single_err_ff; // @[el2_ifu_mem_ctl.scala 681:67]
  wire  iccm_rd_ecc_single_err_hold_in = _T_4074 & _T_317; // @[el2_ifu_mem_ctl.scala 681:96]
  reg [13:0] iccm_rw_addr_f; // @[el2_ifu_mem_ctl.scala 685:51]
  wire [13:0] _T_4079 = iccm_rw_addr_f + 14'h1; // @[el2_ifu_mem_ctl.scala 684:102]
  wire [38:0] _T_4083 = {iccm_corrected_ecc_f_mux,iccm_corrected_data_f_mux}; // @[Cat.scala 29:58]
  wire  _T_4088 = ~io_ifc_fetch_uncacheable_bf; // @[el2_ifu_mem_ctl.scala 689:41]
  wire  _T_4089 = io_ifc_fetch_req_bf & _T_4088; // @[el2_ifu_mem_ctl.scala 689:39]
  wire  _T_4090 = ~io_ifc_iccm_access_bf; // @[el2_ifu_mem_ctl.scala 689:72]
  wire  _T_4091 = _T_4089 & _T_4090; // @[el2_ifu_mem_ctl.scala 689:70]
  wire  _T_4093 = ~miss_state_en; // @[el2_ifu_mem_ctl.scala 690:34]
  wire  _T_4094 = _T_2233 & _T_4093; // @[el2_ifu_mem_ctl.scala 690:32]
  wire  _T_4097 = _T_2249 & _T_4093; // @[el2_ifu_mem_ctl.scala 691:37]
  wire  _T_4098 = _T_4094 | _T_4097; // @[el2_ifu_mem_ctl.scala 690:88]
  wire  _T_4099 = miss_state == 3'h7; // @[el2_ifu_mem_ctl.scala 692:19]
  wire  _T_4101 = _T_4099 & _T_4093; // @[el2_ifu_mem_ctl.scala 692:41]
  wire  _T_4102 = _T_4098 | _T_4101; // @[el2_ifu_mem_ctl.scala 691:88]
  wire  _T_4103 = miss_state == 3'h3; // @[el2_ifu_mem_ctl.scala 693:19]
  wire  _T_4105 = _T_4103 & _T_4093; // @[el2_ifu_mem_ctl.scala 693:35]
  wire  _T_4106 = _T_4102 | _T_4105; // @[el2_ifu_mem_ctl.scala 692:88]
  wire  _T_4109 = _T_2248 & _T_4093; // @[el2_ifu_mem_ctl.scala 694:38]
  wire  _T_4110 = _T_4106 | _T_4109; // @[el2_ifu_mem_ctl.scala 693:88]
  wire  _T_4112 = _T_2249 & miss_state_en; // @[el2_ifu_mem_ctl.scala 695:37]
  wire  _T_4113 = miss_nxtstate == 3'h3; // @[el2_ifu_mem_ctl.scala 695:71]
  wire  _T_4114 = _T_4112 & _T_4113; // @[el2_ifu_mem_ctl.scala 695:54]
  wire  _T_4115 = _T_4110 | _T_4114; // @[el2_ifu_mem_ctl.scala 694:57]
  wire  _T_4116 = ~_T_4115; // @[el2_ifu_mem_ctl.scala 690:5]
  wire  _T_4117 = _T_4091 & _T_4116; // @[el2_ifu_mem_ctl.scala 689:96]
  wire  _T_4118 = io_ifc_fetch_req_bf & io_exu_flush_final; // @[el2_ifu_mem_ctl.scala 696:28]
  wire  _T_4120 = _T_4118 & _T_4088; // @[el2_ifu_mem_ctl.scala 696:50]
  wire  _T_4122 = _T_4120 & _T_4090; // @[el2_ifu_mem_ctl.scala 696:81]
  wire [1:0] _T_4125 = write_ic_16_bytes ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire  _T_10563 = bus_ifu_wr_en_ff_q & replace_way_mb_any_1; // @[el2_ifu_mem_ctl.scala 793:74]
  wire  bus_wren_1 = _T_10563 & miss_pending; // @[el2_ifu_mem_ctl.scala 793:98]
  wire  _T_10562 = bus_ifu_wr_en_ff_q & replace_way_mb_any_0; // @[el2_ifu_mem_ctl.scala 793:74]
  wire  bus_wren_0 = _T_10562 & miss_pending; // @[el2_ifu_mem_ctl.scala 793:98]
  wire [1:0] bus_ic_wr_en = {bus_wren_1,bus_wren_0}; // @[Cat.scala 29:58]
  wire  _T_4131 = ~_T_108; // @[el2_ifu_mem_ctl.scala 699:106]
  wire  _T_4132 = _T_2233 & _T_4131; // @[el2_ifu_mem_ctl.scala 699:104]
  wire  _T_4133 = _T_2249 | _T_4132; // @[el2_ifu_mem_ctl.scala 699:77]
  wire  _T_4137 = ~_T_51; // @[el2_ifu_mem_ctl.scala 699:172]
  wire  _T_4138 = _T_4133 & _T_4137; // @[el2_ifu_mem_ctl.scala 699:170]
  wire  _T_4139 = ~_T_4138; // @[el2_ifu_mem_ctl.scala 699:44]
  wire  _T_4143 = reset_ic_in | reset_ic_ff; // @[el2_ifu_mem_ctl.scala 702:64]
  wire  _T_4144 = ~_T_4143; // @[el2_ifu_mem_ctl.scala 702:50]
  wire  _T_4145 = _T_276 & _T_4144; // @[el2_ifu_mem_ctl.scala 702:48]
  wire  _T_4146 = ~reset_tag_valid_for_miss; // @[el2_ifu_mem_ctl.scala 702:81]
  wire  ic_valid = _T_4145 & _T_4146; // @[el2_ifu_mem_ctl.scala 702:79]
  wire  _T_4148 = debug_c1_clken & io_ic_debug_tag_array; // @[el2_ifu_mem_ctl.scala 703:82]
  reg [6:0] ifu_status_wr_addr_ff; // @[el2_ifu_mem_ctl.scala 706:14]
  wire  _T_4151 = io_ic_debug_wr_en & io_ic_debug_tag_array; // @[el2_ifu_mem_ctl.scala 709:74]
  wire  _T_10560 = bus_ifu_wr_en_ff_q & last_beat; // @[el2_ifu_mem_ctl.scala 792:45]
  wire  way_status_wr_en = _T_10560 | ic_act_hit_f; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  way_status_wr_en_w_debug = way_status_wr_en | _T_4151; // @[el2_ifu_mem_ctl.scala 709:53]
  reg  way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 711:14]
  wire  way_status_hit_new = io_ic_rd_hit[0]; // @[el2_ifu_mem_ctl.scala 788:41]
  reg  way_status_new_ff; // @[el2_ifu_mem_ctl.scala 719:14]
  wire  way_status_clken_0 = ifu_status_wr_addr_ff[6:3] == 4'h0; // @[el2_ifu_mem_ctl.scala 721:132]
  wire  way_status_clken_1 = ifu_status_wr_addr_ff[6:3] == 4'h1; // @[el2_ifu_mem_ctl.scala 721:132]
  wire  way_status_clken_2 = ifu_status_wr_addr_ff[6:3] == 4'h2; // @[el2_ifu_mem_ctl.scala 721:132]
  wire  way_status_clken_3 = ifu_status_wr_addr_ff[6:3] == 4'h3; // @[el2_ifu_mem_ctl.scala 721:132]
  wire  way_status_clken_4 = ifu_status_wr_addr_ff[6:3] == 4'h4; // @[el2_ifu_mem_ctl.scala 721:132]
  wire  way_status_clken_5 = ifu_status_wr_addr_ff[6:3] == 4'h5; // @[el2_ifu_mem_ctl.scala 721:132]
  wire  way_status_clken_6 = ifu_status_wr_addr_ff[6:3] == 4'h6; // @[el2_ifu_mem_ctl.scala 721:132]
  wire  way_status_clken_7 = ifu_status_wr_addr_ff[6:3] == 4'h7; // @[el2_ifu_mem_ctl.scala 721:132]
  wire  way_status_clken_8 = ifu_status_wr_addr_ff[6:3] == 4'h8; // @[el2_ifu_mem_ctl.scala 721:132]
  wire  way_status_clken_9 = ifu_status_wr_addr_ff[6:3] == 4'h9; // @[el2_ifu_mem_ctl.scala 721:132]
  wire  way_status_clken_10 = ifu_status_wr_addr_ff[6:3] == 4'ha; // @[el2_ifu_mem_ctl.scala 721:132]
  wire  way_status_clken_11 = ifu_status_wr_addr_ff[6:3] == 4'hb; // @[el2_ifu_mem_ctl.scala 721:132]
  wire  way_status_clken_12 = ifu_status_wr_addr_ff[6:3] == 4'hc; // @[el2_ifu_mem_ctl.scala 721:132]
  wire  way_status_clken_13 = ifu_status_wr_addr_ff[6:3] == 4'hd; // @[el2_ifu_mem_ctl.scala 721:132]
  wire  way_status_clken_14 = ifu_status_wr_addr_ff[6:3] == 4'he; // @[el2_ifu_mem_ctl.scala 721:132]
  wire  way_status_clken_15 = ifu_status_wr_addr_ff[6:3] == 4'hf; // @[el2_ifu_mem_ctl.scala 721:132]
  wire  _T_4171 = ifu_status_wr_addr_ff[2:0] == 3'h0; // @[el2_ifu_mem_ctl.scala 725:100]
  wire  _T_4172 = _T_4171 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 725:108]
  wire  _T_4173 = _T_4172 & way_status_clken_0; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4176 = ifu_status_wr_addr_ff[2:0] == 3'h1; // @[el2_ifu_mem_ctl.scala 725:100]
  wire  _T_4177 = _T_4176 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 725:108]
  wire  _T_4178 = _T_4177 & way_status_clken_0; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4181 = ifu_status_wr_addr_ff[2:0] == 3'h2; // @[el2_ifu_mem_ctl.scala 725:100]
  wire  _T_4182 = _T_4181 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 725:108]
  wire  _T_4183 = _T_4182 & way_status_clken_0; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4186 = ifu_status_wr_addr_ff[2:0] == 3'h3; // @[el2_ifu_mem_ctl.scala 725:100]
  wire  _T_4187 = _T_4186 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 725:108]
  wire  _T_4188 = _T_4187 & way_status_clken_0; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4191 = ifu_status_wr_addr_ff[2:0] == 3'h4; // @[el2_ifu_mem_ctl.scala 725:100]
  wire  _T_4192 = _T_4191 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 725:108]
  wire  _T_4193 = _T_4192 & way_status_clken_0; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4196 = ifu_status_wr_addr_ff[2:0] == 3'h5; // @[el2_ifu_mem_ctl.scala 725:100]
  wire  _T_4197 = _T_4196 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 725:108]
  wire  _T_4198 = _T_4197 & way_status_clken_0; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4201 = ifu_status_wr_addr_ff[2:0] == 3'h6; // @[el2_ifu_mem_ctl.scala 725:100]
  wire  _T_4202 = _T_4201 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 725:108]
  wire  _T_4203 = _T_4202 & way_status_clken_0; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4206 = ifu_status_wr_addr_ff[2:0] == 3'h7; // @[el2_ifu_mem_ctl.scala 725:100]
  wire  _T_4207 = _T_4206 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 725:108]
  wire  _T_4208 = _T_4207 & way_status_clken_0; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4213 = _T_4172 & way_status_clken_1; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4218 = _T_4177 & way_status_clken_1; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4223 = _T_4182 & way_status_clken_1; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4228 = _T_4187 & way_status_clken_1; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4233 = _T_4192 & way_status_clken_1; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4238 = _T_4197 & way_status_clken_1; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4243 = _T_4202 & way_status_clken_1; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4248 = _T_4207 & way_status_clken_1; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4253 = _T_4172 & way_status_clken_2; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4258 = _T_4177 & way_status_clken_2; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4263 = _T_4182 & way_status_clken_2; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4268 = _T_4187 & way_status_clken_2; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4273 = _T_4192 & way_status_clken_2; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4278 = _T_4197 & way_status_clken_2; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4283 = _T_4202 & way_status_clken_2; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4288 = _T_4207 & way_status_clken_2; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4293 = _T_4172 & way_status_clken_3; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4298 = _T_4177 & way_status_clken_3; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4303 = _T_4182 & way_status_clken_3; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4308 = _T_4187 & way_status_clken_3; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4313 = _T_4192 & way_status_clken_3; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4318 = _T_4197 & way_status_clken_3; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4323 = _T_4202 & way_status_clken_3; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4328 = _T_4207 & way_status_clken_3; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4333 = _T_4172 & way_status_clken_4; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4338 = _T_4177 & way_status_clken_4; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4343 = _T_4182 & way_status_clken_4; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4348 = _T_4187 & way_status_clken_4; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4353 = _T_4192 & way_status_clken_4; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4358 = _T_4197 & way_status_clken_4; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4363 = _T_4202 & way_status_clken_4; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4368 = _T_4207 & way_status_clken_4; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4373 = _T_4172 & way_status_clken_5; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4378 = _T_4177 & way_status_clken_5; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4383 = _T_4182 & way_status_clken_5; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4388 = _T_4187 & way_status_clken_5; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4393 = _T_4192 & way_status_clken_5; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4398 = _T_4197 & way_status_clken_5; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4403 = _T_4202 & way_status_clken_5; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4408 = _T_4207 & way_status_clken_5; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4413 = _T_4172 & way_status_clken_6; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4418 = _T_4177 & way_status_clken_6; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4423 = _T_4182 & way_status_clken_6; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4428 = _T_4187 & way_status_clken_6; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4433 = _T_4192 & way_status_clken_6; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4438 = _T_4197 & way_status_clken_6; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4443 = _T_4202 & way_status_clken_6; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4448 = _T_4207 & way_status_clken_6; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4453 = _T_4172 & way_status_clken_7; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4458 = _T_4177 & way_status_clken_7; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4463 = _T_4182 & way_status_clken_7; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4468 = _T_4187 & way_status_clken_7; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4473 = _T_4192 & way_status_clken_7; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4478 = _T_4197 & way_status_clken_7; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4483 = _T_4202 & way_status_clken_7; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4488 = _T_4207 & way_status_clken_7; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4493 = _T_4172 & way_status_clken_8; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4498 = _T_4177 & way_status_clken_8; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4503 = _T_4182 & way_status_clken_8; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4508 = _T_4187 & way_status_clken_8; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4513 = _T_4192 & way_status_clken_8; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4518 = _T_4197 & way_status_clken_8; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4523 = _T_4202 & way_status_clken_8; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4528 = _T_4207 & way_status_clken_8; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4533 = _T_4172 & way_status_clken_9; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4538 = _T_4177 & way_status_clken_9; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4543 = _T_4182 & way_status_clken_9; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4548 = _T_4187 & way_status_clken_9; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4553 = _T_4192 & way_status_clken_9; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4558 = _T_4197 & way_status_clken_9; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4563 = _T_4202 & way_status_clken_9; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4568 = _T_4207 & way_status_clken_9; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4573 = _T_4172 & way_status_clken_10; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4578 = _T_4177 & way_status_clken_10; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4583 = _T_4182 & way_status_clken_10; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4588 = _T_4187 & way_status_clken_10; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4593 = _T_4192 & way_status_clken_10; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4598 = _T_4197 & way_status_clken_10; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4603 = _T_4202 & way_status_clken_10; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4608 = _T_4207 & way_status_clken_10; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4613 = _T_4172 & way_status_clken_11; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4618 = _T_4177 & way_status_clken_11; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4623 = _T_4182 & way_status_clken_11; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4628 = _T_4187 & way_status_clken_11; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4633 = _T_4192 & way_status_clken_11; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4638 = _T_4197 & way_status_clken_11; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4643 = _T_4202 & way_status_clken_11; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4648 = _T_4207 & way_status_clken_11; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4653 = _T_4172 & way_status_clken_12; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4658 = _T_4177 & way_status_clken_12; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4663 = _T_4182 & way_status_clken_12; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4668 = _T_4187 & way_status_clken_12; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4673 = _T_4192 & way_status_clken_12; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4678 = _T_4197 & way_status_clken_12; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4683 = _T_4202 & way_status_clken_12; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4688 = _T_4207 & way_status_clken_12; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4693 = _T_4172 & way_status_clken_13; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4698 = _T_4177 & way_status_clken_13; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4703 = _T_4182 & way_status_clken_13; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4708 = _T_4187 & way_status_clken_13; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4713 = _T_4192 & way_status_clken_13; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4718 = _T_4197 & way_status_clken_13; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4723 = _T_4202 & way_status_clken_13; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4728 = _T_4207 & way_status_clken_13; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4733 = _T_4172 & way_status_clken_14; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4738 = _T_4177 & way_status_clken_14; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4743 = _T_4182 & way_status_clken_14; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4748 = _T_4187 & way_status_clken_14; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4753 = _T_4192 & way_status_clken_14; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4758 = _T_4197 & way_status_clken_14; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4763 = _T_4202 & way_status_clken_14; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4768 = _T_4207 & way_status_clken_14; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4773 = _T_4172 & way_status_clken_15; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4778 = _T_4177 & way_status_clken_15; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4783 = _T_4182 & way_status_clken_15; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4788 = _T_4187 & way_status_clken_15; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4793 = _T_4192 & way_status_clken_15; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4798 = _T_4197 & way_status_clken_15; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4803 = _T_4202 & way_status_clken_15; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4808 = _T_4207 & way_status_clken_15; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_10566 = _T_100 & replace_way_mb_any_1; // @[el2_ifu_mem_ctl.scala 795:84]
  wire  _T_10567 = _T_10566 & miss_pending; // @[el2_ifu_mem_ctl.scala 795:108]
  wire  bus_wren_last_1 = _T_10567 & bus_last_data_beat; // @[el2_ifu_mem_ctl.scala 795:123]
  wire  wren_reset_miss_1 = replace_way_mb_any_1 & reset_tag_valid_for_miss; // @[el2_ifu_mem_ctl.scala 796:84]
  wire  _T_10569 = bus_wren_last_1 | wren_reset_miss_1; // @[el2_ifu_mem_ctl.scala 797:73]
  wire  _T_10564 = _T_100 & replace_way_mb_any_0; // @[el2_ifu_mem_ctl.scala 795:84]
  wire  _T_10565 = _T_10564 & miss_pending; // @[el2_ifu_mem_ctl.scala 795:108]
  wire  bus_wren_last_0 = _T_10565 & bus_last_data_beat; // @[el2_ifu_mem_ctl.scala 795:123]
  wire  wren_reset_miss_0 = replace_way_mb_any_0 & reset_tag_valid_for_miss; // @[el2_ifu_mem_ctl.scala 796:84]
  wire  _T_10568 = bus_wren_last_0 | wren_reset_miss_0; // @[el2_ifu_mem_ctl.scala 797:73]
  wire [1:0] ifu_tag_wren = {_T_10569,_T_10568}; // @[Cat.scala 29:58]
  wire [1:0] _T_10604 = _T_4151 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [1:0] ic_debug_tag_wr_en = _T_10604 & io_ic_debug_way; // @[el2_ifu_mem_ctl.scala 831:90]
  wire [1:0] ifu_tag_wren_w_debug = ifu_tag_wren | ic_debug_tag_wr_en; // @[el2_ifu_mem_ctl.scala 738:45]
  reg [1:0] ifu_tag_wren_ff; // @[el2_ifu_mem_ctl.scala 740:14]
  reg  ic_valid_ff; // @[el2_ifu_mem_ctl.scala 744:14]
  wire  _T_5342 = ifu_ic_rw_int_addr_ff[6:5] == 2'h0; // @[el2_ifu_mem_ctl.scala 748:78]
  wire  _T_5344 = _T_5342 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 748:87]
  wire  _T_5346 = perr_ic_index_ff[6:5] == 2'h0; // @[el2_ifu_mem_ctl.scala 749:70]
  wire  _T_5348 = _T_5346 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:79]
  wire  _T_5349 = _T_5344 | _T_5348; // @[el2_ifu_mem_ctl.scala 748:109]
  wire  _T_5350 = _T_5349 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:102]
  wire  _T_5354 = _T_5342 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 748:87]
  wire  _T_5358 = _T_5346 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:79]
  wire  _T_5359 = _T_5354 | _T_5358; // @[el2_ifu_mem_ctl.scala 748:109]
  wire  _T_5360 = _T_5359 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:102]
  wire [1:0] tag_valid_clken_0 = {_T_5360,_T_5350}; // @[Cat.scala 29:58]
  wire  _T_5362 = ifu_ic_rw_int_addr_ff[6:5] == 2'h1; // @[el2_ifu_mem_ctl.scala 748:78]
  wire  _T_5364 = _T_5362 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 748:87]
  wire  _T_5366 = perr_ic_index_ff[6:5] == 2'h1; // @[el2_ifu_mem_ctl.scala 749:70]
  wire  _T_5368 = _T_5366 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:79]
  wire  _T_5369 = _T_5364 | _T_5368; // @[el2_ifu_mem_ctl.scala 748:109]
  wire  _T_5370 = _T_5369 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:102]
  wire  _T_5374 = _T_5362 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 748:87]
  wire  _T_5378 = _T_5366 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:79]
  wire  _T_5379 = _T_5374 | _T_5378; // @[el2_ifu_mem_ctl.scala 748:109]
  wire  _T_5380 = _T_5379 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:102]
  wire [1:0] tag_valid_clken_1 = {_T_5380,_T_5370}; // @[Cat.scala 29:58]
  wire  _T_5382 = ifu_ic_rw_int_addr_ff[6:5] == 2'h2; // @[el2_ifu_mem_ctl.scala 748:78]
  wire  _T_5384 = _T_5382 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 748:87]
  wire  _T_5386 = perr_ic_index_ff[6:5] == 2'h2; // @[el2_ifu_mem_ctl.scala 749:70]
  wire  _T_5388 = _T_5386 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:79]
  wire  _T_5389 = _T_5384 | _T_5388; // @[el2_ifu_mem_ctl.scala 748:109]
  wire  _T_5390 = _T_5389 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:102]
  wire  _T_5394 = _T_5382 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 748:87]
  wire  _T_5398 = _T_5386 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:79]
  wire  _T_5399 = _T_5394 | _T_5398; // @[el2_ifu_mem_ctl.scala 748:109]
  wire  _T_5400 = _T_5399 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:102]
  wire [1:0] tag_valid_clken_2 = {_T_5400,_T_5390}; // @[Cat.scala 29:58]
  wire  _T_5402 = ifu_ic_rw_int_addr_ff[6:5] == 2'h3; // @[el2_ifu_mem_ctl.scala 748:78]
  wire  _T_5404 = _T_5402 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 748:87]
  wire  _T_5406 = perr_ic_index_ff[6:5] == 2'h3; // @[el2_ifu_mem_ctl.scala 749:70]
  wire  _T_5408 = _T_5406 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:79]
  wire  _T_5409 = _T_5404 | _T_5408; // @[el2_ifu_mem_ctl.scala 748:109]
  wire  _T_5410 = _T_5409 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:102]
  wire  _T_5414 = _T_5402 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 748:87]
  wire  _T_5418 = _T_5406 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:79]
  wire  _T_5419 = _T_5414 | _T_5418; // @[el2_ifu_mem_ctl.scala 748:109]
  wire  _T_5420 = _T_5419 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:102]
  wire [1:0] tag_valid_clken_3 = {_T_5420,_T_5410}; // @[Cat.scala 29:58]
  wire  _T_5423 = ic_valid_ff & _T_195; // @[el2_ifu_mem_ctl.scala 757:66]
  wire  _T_5424 = ~perr_sel_invalidate; // @[el2_ifu_mem_ctl.scala 757:93]
  wire  _T_5425 = _T_5423 & _T_5424; // @[el2_ifu_mem_ctl.scala 757:91]
  wire  _T_5428 = _T_4950 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_5429 = perr_ic_index_ff == 7'h0; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_5431 = _T_5429 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_5432 = _T_5428 | _T_5431; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_5433 = _T_5432 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_5435 = _T_5433 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_5445 = _T_4951 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_5446 = perr_ic_index_ff == 7'h1; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_5448 = _T_5446 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_5449 = _T_5445 | _T_5448; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_5450 = _T_5449 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_5452 = _T_5450 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_5462 = _T_4952 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_5463 = perr_ic_index_ff == 7'h2; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_5465 = _T_5463 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_5466 = _T_5462 | _T_5465; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_5467 = _T_5466 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_5469 = _T_5467 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_5479 = _T_4953 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_5480 = perr_ic_index_ff == 7'h3; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_5482 = _T_5480 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_5483 = _T_5479 | _T_5482; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_5484 = _T_5483 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_5486 = _T_5484 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_5496 = _T_4954 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_5497 = perr_ic_index_ff == 7'h4; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_5499 = _T_5497 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_5500 = _T_5496 | _T_5499; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_5501 = _T_5500 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_5503 = _T_5501 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_5513 = _T_4955 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_5514 = perr_ic_index_ff == 7'h5; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_5516 = _T_5514 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_5517 = _T_5513 | _T_5516; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_5518 = _T_5517 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_5520 = _T_5518 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_5530 = _T_4956 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_5531 = perr_ic_index_ff == 7'h6; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_5533 = _T_5531 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_5534 = _T_5530 | _T_5533; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_5535 = _T_5534 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_5537 = _T_5535 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_5547 = _T_4957 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_5548 = perr_ic_index_ff == 7'h7; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_5550 = _T_5548 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_5551 = _T_5547 | _T_5550; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_5552 = _T_5551 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_5554 = _T_5552 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_5564 = _T_4958 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_5565 = perr_ic_index_ff == 7'h8; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_5567 = _T_5565 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_5568 = _T_5564 | _T_5567; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_5569 = _T_5568 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_5571 = _T_5569 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_5581 = _T_4959 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_5582 = perr_ic_index_ff == 7'h9; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_5584 = _T_5582 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_5585 = _T_5581 | _T_5584; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_5586 = _T_5585 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_5588 = _T_5586 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_5598 = _T_4960 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_5599 = perr_ic_index_ff == 7'ha; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_5601 = _T_5599 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_5602 = _T_5598 | _T_5601; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_5603 = _T_5602 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_5605 = _T_5603 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_5615 = _T_4961 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_5616 = perr_ic_index_ff == 7'hb; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_5618 = _T_5616 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_5619 = _T_5615 | _T_5618; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_5620 = _T_5619 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_5622 = _T_5620 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_5632 = _T_4962 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_5633 = perr_ic_index_ff == 7'hc; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_5635 = _T_5633 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_5636 = _T_5632 | _T_5635; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_5637 = _T_5636 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_5639 = _T_5637 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_5649 = _T_4963 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_5650 = perr_ic_index_ff == 7'hd; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_5652 = _T_5650 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_5653 = _T_5649 | _T_5652; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_5654 = _T_5653 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_5656 = _T_5654 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_5666 = _T_4964 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_5667 = perr_ic_index_ff == 7'he; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_5669 = _T_5667 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_5670 = _T_5666 | _T_5669; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_5671 = _T_5670 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_5673 = _T_5671 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_5683 = _T_4965 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_5684 = perr_ic_index_ff == 7'hf; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_5686 = _T_5684 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_5687 = _T_5683 | _T_5686; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_5688 = _T_5687 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_5690 = _T_5688 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_5700 = _T_4966 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_5701 = perr_ic_index_ff == 7'h10; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_5703 = _T_5701 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_5704 = _T_5700 | _T_5703; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_5705 = _T_5704 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_5707 = _T_5705 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_5717 = _T_4967 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_5718 = perr_ic_index_ff == 7'h11; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_5720 = _T_5718 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_5721 = _T_5717 | _T_5720; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_5722 = _T_5721 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_5724 = _T_5722 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_5734 = _T_4968 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_5735 = perr_ic_index_ff == 7'h12; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_5737 = _T_5735 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_5738 = _T_5734 | _T_5737; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_5739 = _T_5738 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_5741 = _T_5739 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_5751 = _T_4969 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_5752 = perr_ic_index_ff == 7'h13; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_5754 = _T_5752 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_5755 = _T_5751 | _T_5754; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_5756 = _T_5755 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_5758 = _T_5756 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_5768 = _T_4970 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_5769 = perr_ic_index_ff == 7'h14; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_5771 = _T_5769 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_5772 = _T_5768 | _T_5771; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_5773 = _T_5772 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_5775 = _T_5773 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_5785 = _T_4971 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_5786 = perr_ic_index_ff == 7'h15; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_5788 = _T_5786 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_5789 = _T_5785 | _T_5788; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_5790 = _T_5789 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_5792 = _T_5790 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_5802 = _T_4972 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_5803 = perr_ic_index_ff == 7'h16; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_5805 = _T_5803 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_5806 = _T_5802 | _T_5805; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_5807 = _T_5806 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_5809 = _T_5807 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_5819 = _T_4973 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_5820 = perr_ic_index_ff == 7'h17; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_5822 = _T_5820 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_5823 = _T_5819 | _T_5822; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_5824 = _T_5823 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_5826 = _T_5824 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_5836 = _T_4974 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_5837 = perr_ic_index_ff == 7'h18; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_5839 = _T_5837 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_5840 = _T_5836 | _T_5839; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_5841 = _T_5840 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_5843 = _T_5841 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_5853 = _T_4975 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_5854 = perr_ic_index_ff == 7'h19; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_5856 = _T_5854 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_5857 = _T_5853 | _T_5856; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_5858 = _T_5857 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_5860 = _T_5858 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_5870 = _T_4976 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_5871 = perr_ic_index_ff == 7'h1a; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_5873 = _T_5871 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_5874 = _T_5870 | _T_5873; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_5875 = _T_5874 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_5877 = _T_5875 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_5887 = _T_4977 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_5888 = perr_ic_index_ff == 7'h1b; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_5890 = _T_5888 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_5891 = _T_5887 | _T_5890; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_5892 = _T_5891 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_5894 = _T_5892 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_5904 = _T_4978 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_5905 = perr_ic_index_ff == 7'h1c; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_5907 = _T_5905 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_5908 = _T_5904 | _T_5907; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_5909 = _T_5908 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_5911 = _T_5909 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_5921 = _T_4979 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_5922 = perr_ic_index_ff == 7'h1d; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_5924 = _T_5922 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_5925 = _T_5921 | _T_5924; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_5926 = _T_5925 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_5928 = _T_5926 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_5938 = _T_4980 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_5939 = perr_ic_index_ff == 7'h1e; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_5941 = _T_5939 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_5942 = _T_5938 | _T_5941; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_5943 = _T_5942 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_5945 = _T_5943 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_5955 = _T_4981 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_5956 = perr_ic_index_ff == 7'h1f; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_5958 = _T_5956 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_5959 = _T_5955 | _T_5958; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_5960 = _T_5959 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_5962 = _T_5960 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_5972 = _T_4950 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_5975 = _T_5429 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_5976 = _T_5972 | _T_5975; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_5977 = _T_5976 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_5979 = _T_5977 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_5989 = _T_4951 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_5992 = _T_5446 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_5993 = _T_5989 | _T_5992; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_5994 = _T_5993 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_5996 = _T_5994 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6006 = _T_4952 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6009 = _T_5463 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6010 = _T_6006 | _T_6009; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6011 = _T_6010 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6013 = _T_6011 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6023 = _T_4953 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6026 = _T_5480 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6027 = _T_6023 | _T_6026; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6028 = _T_6027 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6030 = _T_6028 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6040 = _T_4954 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6043 = _T_5497 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6044 = _T_6040 | _T_6043; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6045 = _T_6044 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6047 = _T_6045 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6057 = _T_4955 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6060 = _T_5514 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6061 = _T_6057 | _T_6060; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6062 = _T_6061 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6064 = _T_6062 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6074 = _T_4956 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6077 = _T_5531 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6078 = _T_6074 | _T_6077; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6079 = _T_6078 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6081 = _T_6079 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6091 = _T_4957 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6094 = _T_5548 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6095 = _T_6091 | _T_6094; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6096 = _T_6095 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6098 = _T_6096 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6108 = _T_4958 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6111 = _T_5565 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6112 = _T_6108 | _T_6111; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6113 = _T_6112 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6115 = _T_6113 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6125 = _T_4959 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6128 = _T_5582 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6129 = _T_6125 | _T_6128; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6130 = _T_6129 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6132 = _T_6130 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6142 = _T_4960 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6145 = _T_5599 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6146 = _T_6142 | _T_6145; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6147 = _T_6146 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6149 = _T_6147 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6159 = _T_4961 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6162 = _T_5616 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6163 = _T_6159 | _T_6162; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6164 = _T_6163 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6166 = _T_6164 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6176 = _T_4962 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6179 = _T_5633 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6180 = _T_6176 | _T_6179; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6181 = _T_6180 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6183 = _T_6181 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6193 = _T_4963 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6196 = _T_5650 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6197 = _T_6193 | _T_6196; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6198 = _T_6197 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6200 = _T_6198 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6210 = _T_4964 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6213 = _T_5667 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6214 = _T_6210 | _T_6213; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6215 = _T_6214 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6217 = _T_6215 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6227 = _T_4965 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6230 = _T_5684 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6231 = _T_6227 | _T_6230; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6232 = _T_6231 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6234 = _T_6232 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6244 = _T_4966 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6247 = _T_5701 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6248 = _T_6244 | _T_6247; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6249 = _T_6248 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6251 = _T_6249 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6261 = _T_4967 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6264 = _T_5718 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6265 = _T_6261 | _T_6264; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6266 = _T_6265 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6268 = _T_6266 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6278 = _T_4968 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6281 = _T_5735 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6282 = _T_6278 | _T_6281; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6283 = _T_6282 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6285 = _T_6283 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6295 = _T_4969 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6298 = _T_5752 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6299 = _T_6295 | _T_6298; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6300 = _T_6299 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6302 = _T_6300 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6312 = _T_4970 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6315 = _T_5769 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6316 = _T_6312 | _T_6315; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6317 = _T_6316 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6319 = _T_6317 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6329 = _T_4971 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6332 = _T_5786 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6333 = _T_6329 | _T_6332; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6334 = _T_6333 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6336 = _T_6334 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6346 = _T_4972 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6349 = _T_5803 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6350 = _T_6346 | _T_6349; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6351 = _T_6350 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6353 = _T_6351 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6363 = _T_4973 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6366 = _T_5820 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6367 = _T_6363 | _T_6366; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6368 = _T_6367 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6370 = _T_6368 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6380 = _T_4974 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6383 = _T_5837 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6384 = _T_6380 | _T_6383; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6385 = _T_6384 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6387 = _T_6385 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6397 = _T_4975 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6400 = _T_5854 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6401 = _T_6397 | _T_6400; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6402 = _T_6401 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6404 = _T_6402 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6414 = _T_4976 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6417 = _T_5871 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6418 = _T_6414 | _T_6417; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6419 = _T_6418 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6421 = _T_6419 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6431 = _T_4977 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6434 = _T_5888 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6435 = _T_6431 | _T_6434; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6436 = _T_6435 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6438 = _T_6436 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6448 = _T_4978 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6451 = _T_5905 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6452 = _T_6448 | _T_6451; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6453 = _T_6452 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6455 = _T_6453 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6465 = _T_4979 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6468 = _T_5922 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6469 = _T_6465 | _T_6468; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6470 = _T_6469 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6472 = _T_6470 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6482 = _T_4980 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6485 = _T_5939 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6486 = _T_6482 | _T_6485; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6487 = _T_6486 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6489 = _T_6487 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6499 = _T_4981 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6502 = _T_5956 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6503 = _T_6499 | _T_6502; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6504 = _T_6503 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6506 = _T_6504 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6516 = _T_4982 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6517 = perr_ic_index_ff == 7'h20; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_6519 = _T_6517 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6520 = _T_6516 | _T_6519; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6521 = _T_6520 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6523 = _T_6521 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6533 = _T_4983 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6534 = perr_ic_index_ff == 7'h21; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_6536 = _T_6534 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6537 = _T_6533 | _T_6536; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6538 = _T_6537 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6540 = _T_6538 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6550 = _T_4984 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6551 = perr_ic_index_ff == 7'h22; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_6553 = _T_6551 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6554 = _T_6550 | _T_6553; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6555 = _T_6554 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6557 = _T_6555 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6567 = _T_4985 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6568 = perr_ic_index_ff == 7'h23; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_6570 = _T_6568 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6571 = _T_6567 | _T_6570; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6572 = _T_6571 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6574 = _T_6572 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6584 = _T_4986 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6585 = perr_ic_index_ff == 7'h24; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_6587 = _T_6585 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6588 = _T_6584 | _T_6587; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6589 = _T_6588 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6591 = _T_6589 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6601 = _T_4987 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6602 = perr_ic_index_ff == 7'h25; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_6604 = _T_6602 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6605 = _T_6601 | _T_6604; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6606 = _T_6605 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6608 = _T_6606 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6618 = _T_4988 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6619 = perr_ic_index_ff == 7'h26; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_6621 = _T_6619 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6622 = _T_6618 | _T_6621; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6623 = _T_6622 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6625 = _T_6623 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6635 = _T_4989 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6636 = perr_ic_index_ff == 7'h27; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_6638 = _T_6636 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6639 = _T_6635 | _T_6638; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6640 = _T_6639 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6642 = _T_6640 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6652 = _T_4990 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6653 = perr_ic_index_ff == 7'h28; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_6655 = _T_6653 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6656 = _T_6652 | _T_6655; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6657 = _T_6656 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6659 = _T_6657 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6669 = _T_4991 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6670 = perr_ic_index_ff == 7'h29; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_6672 = _T_6670 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6673 = _T_6669 | _T_6672; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6674 = _T_6673 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6676 = _T_6674 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6686 = _T_4992 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6687 = perr_ic_index_ff == 7'h2a; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_6689 = _T_6687 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6690 = _T_6686 | _T_6689; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6691 = _T_6690 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6693 = _T_6691 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6703 = _T_4993 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6704 = perr_ic_index_ff == 7'h2b; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_6706 = _T_6704 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6707 = _T_6703 | _T_6706; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6708 = _T_6707 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6710 = _T_6708 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6720 = _T_4994 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6721 = perr_ic_index_ff == 7'h2c; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_6723 = _T_6721 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6724 = _T_6720 | _T_6723; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6725 = _T_6724 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6727 = _T_6725 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6737 = _T_4995 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6738 = perr_ic_index_ff == 7'h2d; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_6740 = _T_6738 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6741 = _T_6737 | _T_6740; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6742 = _T_6741 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6744 = _T_6742 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6754 = _T_4996 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6755 = perr_ic_index_ff == 7'h2e; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_6757 = _T_6755 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6758 = _T_6754 | _T_6757; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6759 = _T_6758 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6761 = _T_6759 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6771 = _T_4997 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6772 = perr_ic_index_ff == 7'h2f; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_6774 = _T_6772 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6775 = _T_6771 | _T_6774; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6776 = _T_6775 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6778 = _T_6776 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6788 = _T_4998 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6789 = perr_ic_index_ff == 7'h30; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_6791 = _T_6789 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6792 = _T_6788 | _T_6791; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6793 = _T_6792 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6795 = _T_6793 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6805 = _T_4999 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6806 = perr_ic_index_ff == 7'h31; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_6808 = _T_6806 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6809 = _T_6805 | _T_6808; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6810 = _T_6809 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6812 = _T_6810 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6822 = _T_5000 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6823 = perr_ic_index_ff == 7'h32; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_6825 = _T_6823 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6826 = _T_6822 | _T_6825; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6827 = _T_6826 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6829 = _T_6827 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6839 = _T_5001 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6840 = perr_ic_index_ff == 7'h33; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_6842 = _T_6840 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6843 = _T_6839 | _T_6842; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6844 = _T_6843 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6846 = _T_6844 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6856 = _T_5002 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6857 = perr_ic_index_ff == 7'h34; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_6859 = _T_6857 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6860 = _T_6856 | _T_6859; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6861 = _T_6860 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6863 = _T_6861 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6873 = _T_5003 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6874 = perr_ic_index_ff == 7'h35; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_6876 = _T_6874 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6877 = _T_6873 | _T_6876; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6878 = _T_6877 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6880 = _T_6878 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6890 = _T_5004 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6891 = perr_ic_index_ff == 7'h36; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_6893 = _T_6891 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6894 = _T_6890 | _T_6893; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6895 = _T_6894 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6897 = _T_6895 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6907 = _T_5005 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6908 = perr_ic_index_ff == 7'h37; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_6910 = _T_6908 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6911 = _T_6907 | _T_6910; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6912 = _T_6911 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6914 = _T_6912 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6924 = _T_5006 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6925 = perr_ic_index_ff == 7'h38; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_6927 = _T_6925 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6928 = _T_6924 | _T_6927; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6929 = _T_6928 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6931 = _T_6929 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6941 = _T_5007 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6942 = perr_ic_index_ff == 7'h39; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_6944 = _T_6942 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6945 = _T_6941 | _T_6944; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6946 = _T_6945 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6948 = _T_6946 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6958 = _T_5008 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6959 = perr_ic_index_ff == 7'h3a; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_6961 = _T_6959 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6962 = _T_6958 | _T_6961; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6963 = _T_6962 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6965 = _T_6963 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6975 = _T_5009 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6976 = perr_ic_index_ff == 7'h3b; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_6978 = _T_6976 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6979 = _T_6975 | _T_6978; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6980 = _T_6979 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6982 = _T_6980 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6992 = _T_5010 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6993 = perr_ic_index_ff == 7'h3c; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_6995 = _T_6993 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6996 = _T_6992 | _T_6995; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6997 = _T_6996 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6999 = _T_6997 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7009 = _T_5011 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7010 = perr_ic_index_ff == 7'h3d; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_7012 = _T_7010 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7013 = _T_7009 | _T_7012; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7014 = _T_7013 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7016 = _T_7014 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7026 = _T_5012 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7027 = perr_ic_index_ff == 7'h3e; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_7029 = _T_7027 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7030 = _T_7026 | _T_7029; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7031 = _T_7030 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7033 = _T_7031 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7043 = _T_5013 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7044 = perr_ic_index_ff == 7'h3f; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_7046 = _T_7044 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7047 = _T_7043 | _T_7046; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7048 = _T_7047 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7050 = _T_7048 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7060 = _T_4982 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7063 = _T_6517 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7064 = _T_7060 | _T_7063; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7065 = _T_7064 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7067 = _T_7065 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7077 = _T_4983 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7080 = _T_6534 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7081 = _T_7077 | _T_7080; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7082 = _T_7081 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7084 = _T_7082 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7094 = _T_4984 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7097 = _T_6551 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7098 = _T_7094 | _T_7097; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7099 = _T_7098 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7101 = _T_7099 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7111 = _T_4985 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7114 = _T_6568 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7115 = _T_7111 | _T_7114; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7116 = _T_7115 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7118 = _T_7116 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7128 = _T_4986 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7131 = _T_6585 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7132 = _T_7128 | _T_7131; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7133 = _T_7132 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7135 = _T_7133 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7145 = _T_4987 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7148 = _T_6602 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7149 = _T_7145 | _T_7148; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7150 = _T_7149 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7152 = _T_7150 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7162 = _T_4988 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7165 = _T_6619 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7166 = _T_7162 | _T_7165; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7167 = _T_7166 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7169 = _T_7167 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7179 = _T_4989 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7182 = _T_6636 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7183 = _T_7179 | _T_7182; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7184 = _T_7183 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7186 = _T_7184 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7196 = _T_4990 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7199 = _T_6653 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7200 = _T_7196 | _T_7199; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7201 = _T_7200 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7203 = _T_7201 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7213 = _T_4991 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7216 = _T_6670 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7217 = _T_7213 | _T_7216; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7218 = _T_7217 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7220 = _T_7218 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7230 = _T_4992 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7233 = _T_6687 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7234 = _T_7230 | _T_7233; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7235 = _T_7234 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7237 = _T_7235 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7247 = _T_4993 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7250 = _T_6704 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7251 = _T_7247 | _T_7250; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7252 = _T_7251 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7254 = _T_7252 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7264 = _T_4994 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7267 = _T_6721 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7268 = _T_7264 | _T_7267; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7269 = _T_7268 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7271 = _T_7269 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7281 = _T_4995 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7284 = _T_6738 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7285 = _T_7281 | _T_7284; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7286 = _T_7285 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7288 = _T_7286 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7298 = _T_4996 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7301 = _T_6755 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7302 = _T_7298 | _T_7301; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7303 = _T_7302 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7305 = _T_7303 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7315 = _T_4997 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7318 = _T_6772 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7319 = _T_7315 | _T_7318; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7320 = _T_7319 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7322 = _T_7320 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7332 = _T_4998 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7335 = _T_6789 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7336 = _T_7332 | _T_7335; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7337 = _T_7336 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7339 = _T_7337 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7349 = _T_4999 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7352 = _T_6806 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7353 = _T_7349 | _T_7352; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7354 = _T_7353 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7356 = _T_7354 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7366 = _T_5000 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7369 = _T_6823 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7370 = _T_7366 | _T_7369; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7371 = _T_7370 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7373 = _T_7371 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7383 = _T_5001 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7386 = _T_6840 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7387 = _T_7383 | _T_7386; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7388 = _T_7387 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7390 = _T_7388 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7400 = _T_5002 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7403 = _T_6857 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7404 = _T_7400 | _T_7403; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7405 = _T_7404 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7407 = _T_7405 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7417 = _T_5003 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7420 = _T_6874 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7421 = _T_7417 | _T_7420; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7422 = _T_7421 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7424 = _T_7422 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7434 = _T_5004 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7437 = _T_6891 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7438 = _T_7434 | _T_7437; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7439 = _T_7438 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7441 = _T_7439 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7451 = _T_5005 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7454 = _T_6908 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7455 = _T_7451 | _T_7454; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7456 = _T_7455 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7458 = _T_7456 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7468 = _T_5006 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7471 = _T_6925 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7472 = _T_7468 | _T_7471; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7473 = _T_7472 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7475 = _T_7473 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7485 = _T_5007 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7488 = _T_6942 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7489 = _T_7485 | _T_7488; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7490 = _T_7489 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7492 = _T_7490 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7502 = _T_5008 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7505 = _T_6959 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7506 = _T_7502 | _T_7505; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7507 = _T_7506 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7509 = _T_7507 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7519 = _T_5009 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7522 = _T_6976 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7523 = _T_7519 | _T_7522; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7524 = _T_7523 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7526 = _T_7524 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7536 = _T_5010 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7539 = _T_6993 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7540 = _T_7536 | _T_7539; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7541 = _T_7540 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7543 = _T_7541 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7553 = _T_5011 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7556 = _T_7010 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7557 = _T_7553 | _T_7556; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7558 = _T_7557 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7560 = _T_7558 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7570 = _T_5012 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7573 = _T_7027 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7574 = _T_7570 | _T_7573; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7575 = _T_7574 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7577 = _T_7575 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7587 = _T_5013 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7590 = _T_7044 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7591 = _T_7587 | _T_7590; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7592 = _T_7591 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7594 = _T_7592 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7604 = _T_5014 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7605 = perr_ic_index_ff == 7'h40; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_7607 = _T_7605 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7608 = _T_7604 | _T_7607; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7609 = _T_7608 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7611 = _T_7609 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7621 = _T_5015 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7622 = perr_ic_index_ff == 7'h41; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_7624 = _T_7622 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7625 = _T_7621 | _T_7624; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7626 = _T_7625 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7628 = _T_7626 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7638 = _T_5016 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7639 = perr_ic_index_ff == 7'h42; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_7641 = _T_7639 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7642 = _T_7638 | _T_7641; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7643 = _T_7642 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7645 = _T_7643 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7655 = _T_5017 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7656 = perr_ic_index_ff == 7'h43; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_7658 = _T_7656 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7659 = _T_7655 | _T_7658; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7660 = _T_7659 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7662 = _T_7660 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7672 = _T_5018 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7673 = perr_ic_index_ff == 7'h44; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_7675 = _T_7673 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7676 = _T_7672 | _T_7675; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7677 = _T_7676 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7679 = _T_7677 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7689 = _T_5019 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7690 = perr_ic_index_ff == 7'h45; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_7692 = _T_7690 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7693 = _T_7689 | _T_7692; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7694 = _T_7693 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7696 = _T_7694 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7706 = _T_5020 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7707 = perr_ic_index_ff == 7'h46; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_7709 = _T_7707 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7710 = _T_7706 | _T_7709; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7711 = _T_7710 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7713 = _T_7711 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7723 = _T_5021 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7724 = perr_ic_index_ff == 7'h47; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_7726 = _T_7724 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7727 = _T_7723 | _T_7726; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7728 = _T_7727 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7730 = _T_7728 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7740 = _T_5022 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7741 = perr_ic_index_ff == 7'h48; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_7743 = _T_7741 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7744 = _T_7740 | _T_7743; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7745 = _T_7744 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7747 = _T_7745 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7757 = _T_5023 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7758 = perr_ic_index_ff == 7'h49; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_7760 = _T_7758 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7761 = _T_7757 | _T_7760; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7762 = _T_7761 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7764 = _T_7762 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7774 = _T_5024 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7775 = perr_ic_index_ff == 7'h4a; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_7777 = _T_7775 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7778 = _T_7774 | _T_7777; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7779 = _T_7778 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7781 = _T_7779 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7791 = _T_5025 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7792 = perr_ic_index_ff == 7'h4b; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_7794 = _T_7792 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7795 = _T_7791 | _T_7794; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7796 = _T_7795 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7798 = _T_7796 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7808 = _T_5026 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7809 = perr_ic_index_ff == 7'h4c; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_7811 = _T_7809 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7812 = _T_7808 | _T_7811; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7813 = _T_7812 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7815 = _T_7813 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7825 = _T_5027 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7826 = perr_ic_index_ff == 7'h4d; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_7828 = _T_7826 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7829 = _T_7825 | _T_7828; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7830 = _T_7829 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7832 = _T_7830 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7842 = _T_5028 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7843 = perr_ic_index_ff == 7'h4e; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_7845 = _T_7843 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7846 = _T_7842 | _T_7845; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7847 = _T_7846 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7849 = _T_7847 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7859 = _T_5029 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7860 = perr_ic_index_ff == 7'h4f; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_7862 = _T_7860 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7863 = _T_7859 | _T_7862; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7864 = _T_7863 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7866 = _T_7864 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7876 = _T_5030 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7877 = perr_ic_index_ff == 7'h50; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_7879 = _T_7877 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7880 = _T_7876 | _T_7879; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7881 = _T_7880 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7883 = _T_7881 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7893 = _T_5031 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7894 = perr_ic_index_ff == 7'h51; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_7896 = _T_7894 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7897 = _T_7893 | _T_7896; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7898 = _T_7897 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7900 = _T_7898 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7910 = _T_5032 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7911 = perr_ic_index_ff == 7'h52; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_7913 = _T_7911 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7914 = _T_7910 | _T_7913; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7915 = _T_7914 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7917 = _T_7915 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7927 = _T_5033 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7928 = perr_ic_index_ff == 7'h53; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_7930 = _T_7928 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7931 = _T_7927 | _T_7930; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7932 = _T_7931 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7934 = _T_7932 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7944 = _T_5034 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7945 = perr_ic_index_ff == 7'h54; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_7947 = _T_7945 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7948 = _T_7944 | _T_7947; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7949 = _T_7948 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7951 = _T_7949 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7961 = _T_5035 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7962 = perr_ic_index_ff == 7'h55; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_7964 = _T_7962 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7965 = _T_7961 | _T_7964; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7966 = _T_7965 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7968 = _T_7966 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7978 = _T_5036 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7979 = perr_ic_index_ff == 7'h56; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_7981 = _T_7979 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7982 = _T_7978 | _T_7981; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7983 = _T_7982 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7985 = _T_7983 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7995 = _T_5037 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7996 = perr_ic_index_ff == 7'h57; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_7998 = _T_7996 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7999 = _T_7995 | _T_7998; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8000 = _T_7999 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8002 = _T_8000 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8012 = _T_5038 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8013 = perr_ic_index_ff == 7'h58; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_8015 = _T_8013 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8016 = _T_8012 | _T_8015; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8017 = _T_8016 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8019 = _T_8017 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8029 = _T_5039 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8030 = perr_ic_index_ff == 7'h59; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_8032 = _T_8030 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8033 = _T_8029 | _T_8032; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8034 = _T_8033 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8036 = _T_8034 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8046 = _T_5040 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8047 = perr_ic_index_ff == 7'h5a; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_8049 = _T_8047 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8050 = _T_8046 | _T_8049; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8051 = _T_8050 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8053 = _T_8051 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8063 = _T_5041 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8064 = perr_ic_index_ff == 7'h5b; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_8066 = _T_8064 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8067 = _T_8063 | _T_8066; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8068 = _T_8067 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8070 = _T_8068 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8080 = _T_5042 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8081 = perr_ic_index_ff == 7'h5c; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_8083 = _T_8081 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8084 = _T_8080 | _T_8083; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8085 = _T_8084 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8087 = _T_8085 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8097 = _T_5043 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8098 = perr_ic_index_ff == 7'h5d; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_8100 = _T_8098 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8101 = _T_8097 | _T_8100; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8102 = _T_8101 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8104 = _T_8102 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8114 = _T_5044 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8115 = perr_ic_index_ff == 7'h5e; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_8117 = _T_8115 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8118 = _T_8114 | _T_8117; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8119 = _T_8118 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8121 = _T_8119 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8131 = _T_5045 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8132 = perr_ic_index_ff == 7'h5f; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_8134 = _T_8132 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8135 = _T_8131 | _T_8134; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8136 = _T_8135 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8138 = _T_8136 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8148 = _T_5014 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8151 = _T_7605 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8152 = _T_8148 | _T_8151; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8153 = _T_8152 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8155 = _T_8153 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8165 = _T_5015 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8168 = _T_7622 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8169 = _T_8165 | _T_8168; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8170 = _T_8169 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8172 = _T_8170 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8182 = _T_5016 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8185 = _T_7639 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8186 = _T_8182 | _T_8185; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8187 = _T_8186 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8189 = _T_8187 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8199 = _T_5017 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8202 = _T_7656 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8203 = _T_8199 | _T_8202; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8204 = _T_8203 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8206 = _T_8204 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8216 = _T_5018 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8219 = _T_7673 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8220 = _T_8216 | _T_8219; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8221 = _T_8220 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8223 = _T_8221 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8233 = _T_5019 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8236 = _T_7690 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8237 = _T_8233 | _T_8236; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8238 = _T_8237 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8240 = _T_8238 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8250 = _T_5020 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8253 = _T_7707 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8254 = _T_8250 | _T_8253; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8255 = _T_8254 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8257 = _T_8255 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8267 = _T_5021 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8270 = _T_7724 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8271 = _T_8267 | _T_8270; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8272 = _T_8271 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8274 = _T_8272 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8284 = _T_5022 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8287 = _T_7741 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8288 = _T_8284 | _T_8287; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8289 = _T_8288 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8291 = _T_8289 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8301 = _T_5023 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8304 = _T_7758 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8305 = _T_8301 | _T_8304; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8306 = _T_8305 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8308 = _T_8306 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8318 = _T_5024 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8321 = _T_7775 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8322 = _T_8318 | _T_8321; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8323 = _T_8322 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8325 = _T_8323 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8335 = _T_5025 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8338 = _T_7792 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8339 = _T_8335 | _T_8338; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8340 = _T_8339 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8342 = _T_8340 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8352 = _T_5026 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8355 = _T_7809 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8356 = _T_8352 | _T_8355; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8357 = _T_8356 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8359 = _T_8357 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8369 = _T_5027 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8372 = _T_7826 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8373 = _T_8369 | _T_8372; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8374 = _T_8373 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8376 = _T_8374 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8386 = _T_5028 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8389 = _T_7843 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8390 = _T_8386 | _T_8389; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8391 = _T_8390 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8393 = _T_8391 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8403 = _T_5029 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8406 = _T_7860 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8407 = _T_8403 | _T_8406; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8408 = _T_8407 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8410 = _T_8408 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8420 = _T_5030 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8423 = _T_7877 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8424 = _T_8420 | _T_8423; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8425 = _T_8424 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8427 = _T_8425 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8437 = _T_5031 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8440 = _T_7894 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8441 = _T_8437 | _T_8440; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8442 = _T_8441 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8444 = _T_8442 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8454 = _T_5032 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8457 = _T_7911 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8458 = _T_8454 | _T_8457; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8459 = _T_8458 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8461 = _T_8459 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8471 = _T_5033 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8474 = _T_7928 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8475 = _T_8471 | _T_8474; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8476 = _T_8475 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8478 = _T_8476 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8488 = _T_5034 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8491 = _T_7945 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8492 = _T_8488 | _T_8491; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8493 = _T_8492 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8495 = _T_8493 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8505 = _T_5035 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8508 = _T_7962 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8509 = _T_8505 | _T_8508; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8510 = _T_8509 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8512 = _T_8510 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8522 = _T_5036 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8525 = _T_7979 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8526 = _T_8522 | _T_8525; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8527 = _T_8526 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8529 = _T_8527 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8539 = _T_5037 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8542 = _T_7996 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8543 = _T_8539 | _T_8542; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8544 = _T_8543 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8546 = _T_8544 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8556 = _T_5038 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8559 = _T_8013 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8560 = _T_8556 | _T_8559; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8561 = _T_8560 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8563 = _T_8561 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8573 = _T_5039 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8576 = _T_8030 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8577 = _T_8573 | _T_8576; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8578 = _T_8577 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8580 = _T_8578 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8590 = _T_5040 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8593 = _T_8047 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8594 = _T_8590 | _T_8593; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8595 = _T_8594 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8597 = _T_8595 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8607 = _T_5041 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8610 = _T_8064 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8611 = _T_8607 | _T_8610; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8612 = _T_8611 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8614 = _T_8612 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8624 = _T_5042 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8627 = _T_8081 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8628 = _T_8624 | _T_8627; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8629 = _T_8628 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8631 = _T_8629 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8641 = _T_5043 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8644 = _T_8098 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8645 = _T_8641 | _T_8644; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8646 = _T_8645 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8648 = _T_8646 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8658 = _T_5044 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8661 = _T_8115 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8662 = _T_8658 | _T_8661; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8663 = _T_8662 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8665 = _T_8663 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8675 = _T_5045 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8678 = _T_8132 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8679 = _T_8675 | _T_8678; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8680 = _T_8679 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8682 = _T_8680 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8692 = _T_5046 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8693 = perr_ic_index_ff == 7'h60; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_8695 = _T_8693 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8696 = _T_8692 | _T_8695; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8697 = _T_8696 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8699 = _T_8697 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8709 = _T_5047 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8710 = perr_ic_index_ff == 7'h61; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_8712 = _T_8710 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8713 = _T_8709 | _T_8712; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8714 = _T_8713 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8716 = _T_8714 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8726 = _T_5048 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8727 = perr_ic_index_ff == 7'h62; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_8729 = _T_8727 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8730 = _T_8726 | _T_8729; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8731 = _T_8730 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8733 = _T_8731 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8743 = _T_5049 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8744 = perr_ic_index_ff == 7'h63; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_8746 = _T_8744 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8747 = _T_8743 | _T_8746; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8748 = _T_8747 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8750 = _T_8748 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8760 = _T_5050 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8761 = perr_ic_index_ff == 7'h64; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_8763 = _T_8761 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8764 = _T_8760 | _T_8763; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8765 = _T_8764 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8767 = _T_8765 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8777 = _T_5051 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8778 = perr_ic_index_ff == 7'h65; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_8780 = _T_8778 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8781 = _T_8777 | _T_8780; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8782 = _T_8781 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8784 = _T_8782 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8794 = _T_5052 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8795 = perr_ic_index_ff == 7'h66; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_8797 = _T_8795 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8798 = _T_8794 | _T_8797; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8799 = _T_8798 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8801 = _T_8799 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8811 = _T_5053 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8812 = perr_ic_index_ff == 7'h67; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_8814 = _T_8812 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8815 = _T_8811 | _T_8814; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8816 = _T_8815 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8818 = _T_8816 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8828 = _T_5054 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8829 = perr_ic_index_ff == 7'h68; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_8831 = _T_8829 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8832 = _T_8828 | _T_8831; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8833 = _T_8832 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8835 = _T_8833 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8845 = _T_5055 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8846 = perr_ic_index_ff == 7'h69; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_8848 = _T_8846 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8849 = _T_8845 | _T_8848; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8850 = _T_8849 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8852 = _T_8850 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8862 = _T_5056 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8863 = perr_ic_index_ff == 7'h6a; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_8865 = _T_8863 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8866 = _T_8862 | _T_8865; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8867 = _T_8866 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8869 = _T_8867 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8879 = _T_5057 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8880 = perr_ic_index_ff == 7'h6b; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_8882 = _T_8880 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8883 = _T_8879 | _T_8882; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8884 = _T_8883 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8886 = _T_8884 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8896 = _T_5058 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8897 = perr_ic_index_ff == 7'h6c; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_8899 = _T_8897 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8900 = _T_8896 | _T_8899; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8901 = _T_8900 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8903 = _T_8901 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8913 = _T_5059 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8914 = perr_ic_index_ff == 7'h6d; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_8916 = _T_8914 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8917 = _T_8913 | _T_8916; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8918 = _T_8917 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8920 = _T_8918 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8930 = _T_5060 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8931 = perr_ic_index_ff == 7'h6e; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_8933 = _T_8931 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8934 = _T_8930 | _T_8933; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8935 = _T_8934 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8937 = _T_8935 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8947 = _T_5061 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8948 = perr_ic_index_ff == 7'h6f; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_8950 = _T_8948 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8951 = _T_8947 | _T_8950; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8952 = _T_8951 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8954 = _T_8952 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8964 = _T_5062 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8965 = perr_ic_index_ff == 7'h70; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_8967 = _T_8965 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8968 = _T_8964 | _T_8967; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8969 = _T_8968 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8971 = _T_8969 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8981 = _T_5063 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8982 = perr_ic_index_ff == 7'h71; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_8984 = _T_8982 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8985 = _T_8981 | _T_8984; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8986 = _T_8985 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8988 = _T_8986 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8998 = _T_5064 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8999 = perr_ic_index_ff == 7'h72; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_9001 = _T_8999 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_9002 = _T_8998 | _T_9001; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_9003 = _T_9002 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_9005 = _T_9003 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_9015 = _T_5065 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_9016 = perr_ic_index_ff == 7'h73; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_9018 = _T_9016 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_9019 = _T_9015 | _T_9018; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_9020 = _T_9019 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_9022 = _T_9020 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_9032 = _T_5066 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_9033 = perr_ic_index_ff == 7'h74; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_9035 = _T_9033 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_9036 = _T_9032 | _T_9035; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_9037 = _T_9036 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_9039 = _T_9037 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_9049 = _T_5067 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_9050 = perr_ic_index_ff == 7'h75; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_9052 = _T_9050 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_9053 = _T_9049 | _T_9052; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_9054 = _T_9053 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_9056 = _T_9054 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_9066 = _T_5068 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_9067 = perr_ic_index_ff == 7'h76; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_9069 = _T_9067 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_9070 = _T_9066 | _T_9069; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_9071 = _T_9070 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_9073 = _T_9071 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_9083 = _T_5069 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_9084 = perr_ic_index_ff == 7'h77; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_9086 = _T_9084 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_9087 = _T_9083 | _T_9086; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_9088 = _T_9087 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_9090 = _T_9088 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_9100 = _T_5070 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_9101 = perr_ic_index_ff == 7'h78; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_9103 = _T_9101 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_9104 = _T_9100 | _T_9103; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_9105 = _T_9104 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_9107 = _T_9105 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_9117 = _T_5071 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_9118 = perr_ic_index_ff == 7'h79; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_9120 = _T_9118 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_9121 = _T_9117 | _T_9120; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_9122 = _T_9121 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_9124 = _T_9122 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_9134 = _T_5072 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_9135 = perr_ic_index_ff == 7'h7a; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_9137 = _T_9135 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_9138 = _T_9134 | _T_9137; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_9139 = _T_9138 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_9141 = _T_9139 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_9151 = _T_5073 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_9152 = perr_ic_index_ff == 7'h7b; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_9154 = _T_9152 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_9155 = _T_9151 | _T_9154; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_9156 = _T_9155 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_9158 = _T_9156 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_9168 = _T_5074 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_9169 = perr_ic_index_ff == 7'h7c; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_9171 = _T_9169 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_9172 = _T_9168 | _T_9171; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_9173 = _T_9172 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_9175 = _T_9173 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_9185 = _T_5075 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_9186 = perr_ic_index_ff == 7'h7d; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_9188 = _T_9186 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_9189 = _T_9185 | _T_9188; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_9190 = _T_9189 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_9192 = _T_9190 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_9202 = _T_5076 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_9203 = perr_ic_index_ff == 7'h7e; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_9205 = _T_9203 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_9206 = _T_9202 | _T_9205; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_9207 = _T_9206 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_9209 = _T_9207 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_9219 = _T_5077 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_9220 = perr_ic_index_ff == 7'h7f; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_9222 = _T_9220 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_9223 = _T_9219 | _T_9222; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_9224 = _T_9223 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_9226 = _T_9224 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_9236 = _T_5046 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_9239 = _T_8693 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_9240 = _T_9236 | _T_9239; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_9241 = _T_9240 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_9243 = _T_9241 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_9253 = _T_5047 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_9256 = _T_8710 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_9257 = _T_9253 | _T_9256; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_9258 = _T_9257 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_9260 = _T_9258 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_9270 = _T_5048 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_9273 = _T_8727 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_9274 = _T_9270 | _T_9273; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_9275 = _T_9274 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_9277 = _T_9275 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_9287 = _T_5049 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_9290 = _T_8744 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_9291 = _T_9287 | _T_9290; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_9292 = _T_9291 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_9294 = _T_9292 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_9304 = _T_5050 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_9307 = _T_8761 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_9308 = _T_9304 | _T_9307; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_9309 = _T_9308 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_9311 = _T_9309 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_9321 = _T_5051 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_9324 = _T_8778 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_9325 = _T_9321 | _T_9324; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_9326 = _T_9325 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_9328 = _T_9326 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_9338 = _T_5052 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_9341 = _T_8795 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_9342 = _T_9338 | _T_9341; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_9343 = _T_9342 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_9345 = _T_9343 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_9355 = _T_5053 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_9358 = _T_8812 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_9359 = _T_9355 | _T_9358; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_9360 = _T_9359 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_9362 = _T_9360 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_9372 = _T_5054 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_9375 = _T_8829 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_9376 = _T_9372 | _T_9375; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_9377 = _T_9376 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_9379 = _T_9377 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_9389 = _T_5055 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_9392 = _T_8846 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_9393 = _T_9389 | _T_9392; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_9394 = _T_9393 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_9396 = _T_9394 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_9406 = _T_5056 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_9409 = _T_8863 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_9410 = _T_9406 | _T_9409; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_9411 = _T_9410 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_9413 = _T_9411 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_9423 = _T_5057 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_9426 = _T_8880 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_9427 = _T_9423 | _T_9426; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_9428 = _T_9427 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_9430 = _T_9428 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_9440 = _T_5058 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_9443 = _T_8897 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_9444 = _T_9440 | _T_9443; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_9445 = _T_9444 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_9447 = _T_9445 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_9457 = _T_5059 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_9460 = _T_8914 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_9461 = _T_9457 | _T_9460; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_9462 = _T_9461 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_9464 = _T_9462 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_9474 = _T_5060 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_9477 = _T_8931 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_9478 = _T_9474 | _T_9477; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_9479 = _T_9478 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_9481 = _T_9479 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_9491 = _T_5061 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_9494 = _T_8948 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_9495 = _T_9491 | _T_9494; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_9496 = _T_9495 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_9498 = _T_9496 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_9508 = _T_5062 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_9511 = _T_8965 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_9512 = _T_9508 | _T_9511; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_9513 = _T_9512 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_9515 = _T_9513 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_9525 = _T_5063 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_9528 = _T_8982 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_9529 = _T_9525 | _T_9528; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_9530 = _T_9529 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_9532 = _T_9530 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_9542 = _T_5064 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_9545 = _T_8999 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_9546 = _T_9542 | _T_9545; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_9547 = _T_9546 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_9549 = _T_9547 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_9559 = _T_5065 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_9562 = _T_9016 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_9563 = _T_9559 | _T_9562; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_9564 = _T_9563 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_9566 = _T_9564 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_9576 = _T_5066 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_9579 = _T_9033 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_9580 = _T_9576 | _T_9579; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_9581 = _T_9580 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_9583 = _T_9581 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_9593 = _T_5067 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_9596 = _T_9050 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_9597 = _T_9593 | _T_9596; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_9598 = _T_9597 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_9600 = _T_9598 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_9610 = _T_5068 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_9613 = _T_9067 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_9614 = _T_9610 | _T_9613; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_9615 = _T_9614 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_9617 = _T_9615 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_9627 = _T_5069 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_9630 = _T_9084 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_9631 = _T_9627 | _T_9630; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_9632 = _T_9631 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_9634 = _T_9632 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_9644 = _T_5070 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_9647 = _T_9101 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_9648 = _T_9644 | _T_9647; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_9649 = _T_9648 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_9651 = _T_9649 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_9661 = _T_5071 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_9664 = _T_9118 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_9665 = _T_9661 | _T_9664; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_9666 = _T_9665 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_9668 = _T_9666 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_9678 = _T_5072 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_9681 = _T_9135 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_9682 = _T_9678 | _T_9681; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_9683 = _T_9682 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_9685 = _T_9683 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_9695 = _T_5073 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_9698 = _T_9152 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_9699 = _T_9695 | _T_9698; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_9700 = _T_9699 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_9702 = _T_9700 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_9712 = _T_5074 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_9715 = _T_9169 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_9716 = _T_9712 | _T_9715; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_9717 = _T_9716 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_9719 = _T_9717 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_9729 = _T_5075 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_9732 = _T_9186 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_9733 = _T_9729 | _T_9732; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_9734 = _T_9733 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_9736 = _T_9734 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_9746 = _T_5076 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_9749 = _T_9203 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_9750 = _T_9746 | _T_9749; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_9751 = _T_9750 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_9753 = _T_9751 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_9763 = _T_5077 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_9766 = _T_9220 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_9767 = _T_9763 | _T_9766; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_9768 = _T_9767 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_9770 = _T_9768 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_10572 = ~fetch_uncacheable_ff; // @[el2_ifu_mem_ctl.scala 813:63]
  wire  _T_10573 = _T_10572 & ifc_fetch_req_f; // @[el2_ifu_mem_ctl.scala 813:85]
  wire [1:0] _T_10575 = _T_10573 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  reg  _T_10582; // @[el2_ifu_mem_ctl.scala 818:57]
  reg  _T_10583; // @[el2_ifu_mem_ctl.scala 819:56]
  reg  _T_10584; // @[el2_ifu_mem_ctl.scala 820:59]
  wire  _T_10585 = ~ifu_bus_arready_ff; // @[el2_ifu_mem_ctl.scala 821:80]
  wire  _T_10586 = ifu_bus_arvalid_ff & _T_10585; // @[el2_ifu_mem_ctl.scala 821:78]
  wire  _T_10587 = _T_10586 & miss_pending; // @[el2_ifu_mem_ctl.scala 821:100]
  reg  _T_10588; // @[el2_ifu_mem_ctl.scala 821:58]
  reg  _T_10589; // @[el2_ifu_mem_ctl.scala 822:58]
  wire  _T_10592 = io_dec_tlu_ic_diag_pkt_icache_dicawics[15:14] == 2'h3; // @[el2_ifu_mem_ctl.scala 829:71]
  wire  _T_10594 = io_dec_tlu_ic_diag_pkt_icache_dicawics[15:14] == 2'h2; // @[el2_ifu_mem_ctl.scala 829:124]
  wire  _T_10596 = io_dec_tlu_ic_diag_pkt_icache_dicawics[15:14] == 2'h1; // @[el2_ifu_mem_ctl.scala 830:50]
  wire  _T_10598 = io_dec_tlu_ic_diag_pkt_icache_dicawics[15:14] == 2'h0; // @[el2_ifu_mem_ctl.scala 830:103]
  wire [3:0] _T_10601 = {_T_10592,_T_10594,_T_10596,_T_10598}; // @[Cat.scala 29:58]
  wire  ic_debug_ict_array_sel_in = io_ic_debug_rd_en & io_ic_debug_tag_array; // @[el2_ifu_mem_ctl.scala 832:53]
  reg  _T_10612; // @[Reg.scala 27:20]
  assign io_ifu_miss_state_idle = miss_state == 3'h0; // @[el2_ifu_mem_ctl.scala 328:26]
  assign io_ifu_ic_mb_empty = _T_326 | _T_231; // @[el2_ifu_mem_ctl.scala 327:22]
  assign io_ic_dma_active = _T_11 | io_dec_tlu_flush_err_wb; // @[el2_ifu_mem_ctl.scala 192:20]
  assign io_ic_write_stall = write_ic_16_bytes & _T_4139; // @[el2_ifu_mem_ctl.scala 699:21]
  assign io_ifu_pmu_ic_miss = _T_10582; // @[el2_ifu_mem_ctl.scala 818:22]
  assign io_ifu_pmu_ic_hit = _T_10583; // @[el2_ifu_mem_ctl.scala 819:21]
  assign io_ifu_pmu_bus_error = _T_10584; // @[el2_ifu_mem_ctl.scala 820:24]
  assign io_ifu_pmu_bus_busy = _T_10588; // @[el2_ifu_mem_ctl.scala 821:23]
  assign io_ifu_pmu_bus_trxn = _T_10589; // @[el2_ifu_mem_ctl.scala 822:23]
  assign io_ifu_axi_awvalid = 1'h0; // @[el2_ifu_mem_ctl.scala 142:22]
  assign io_ifu_axi_awid = 3'h0; // @[el2_ifu_mem_ctl.scala 141:19]
  assign io_ifu_axi_awaddr = 32'h0; // @[el2_ifu_mem_ctl.scala 136:21]
  assign io_ifu_axi_awregion = 4'h0; // @[el2_ifu_mem_ctl.scala 140:23]
  assign io_ifu_axi_awlen = 8'h0; // @[el2_ifu_mem_ctl.scala 138:20]
  assign io_ifu_axi_awsize = 3'h0; // @[el2_ifu_mem_ctl.scala 149:21]
  assign io_ifu_axi_awburst = 2'h0; // @[el2_ifu_mem_ctl.scala 151:22]
  assign io_ifu_axi_awlock = 1'h0; // @[el2_ifu_mem_ctl.scala 146:21]
  assign io_ifu_axi_awcache = 4'h0; // @[el2_ifu_mem_ctl.scala 144:22]
  assign io_ifu_axi_awprot = 3'h0; // @[el2_ifu_mem_ctl.scala 137:21]
  assign io_ifu_axi_awqos = 4'h0; // @[el2_ifu_mem_ctl.scala 135:20]
  assign io_ifu_axi_wvalid = 1'h0; // @[el2_ifu_mem_ctl.scala 133:21]
  assign io_ifu_axi_wdata = 64'h0; // @[el2_ifu_mem_ctl.scala 134:20]
  assign io_ifu_axi_wstrb = 8'h0; // @[el2_ifu_mem_ctl.scala 143:20]
  assign io_ifu_axi_wlast = 1'h0; // @[el2_ifu_mem_ctl.scala 152:20]
  assign io_ifu_axi_bready = 1'h0; // @[el2_ifu_mem_ctl.scala 147:21]
  assign io_ifu_axi_arvalid = ifu_bus_cmd_valid; // @[el2_ifu_mem_ctl.scala 560:22]
  assign io_ifu_axi_arid = bus_rd_addr_count & _T_2572; // @[el2_ifu_mem_ctl.scala 561:19]
  assign io_ifu_axi_araddr = _T_2574 & _T_2576; // @[el2_ifu_mem_ctl.scala 562:21]
  assign io_ifu_axi_arregion = ifu_ic_req_addr_f[28:25]; // @[el2_ifu_mem_ctl.scala 565:23]
  assign io_ifu_axi_arlen = 8'h0; // @[el2_ifu_mem_ctl.scala 148:20]
  assign io_ifu_axi_arsize = 3'h3; // @[el2_ifu_mem_ctl.scala 563:21]
  assign io_ifu_axi_arburst = 2'h1; // @[el2_ifu_mem_ctl.scala 566:22]
  assign io_ifu_axi_arlock = 1'h0; // @[el2_ifu_mem_ctl.scala 139:21]
  assign io_ifu_axi_arcache = 4'hf; // @[el2_ifu_mem_ctl.scala 564:22]
  assign io_ifu_axi_arprot = 3'h0; // @[el2_ifu_mem_ctl.scala 150:21]
  assign io_ifu_axi_arqos = 4'h0; // @[el2_ifu_mem_ctl.scala 145:20]
  assign io_ifu_axi_rready = 1'h1; // @[el2_ifu_mem_ctl.scala 567:21]
  assign io_iccm_dma_ecc_error = |iccm_double_ecc_error; // @[el2_ifu_mem_ctl.scala 658:25]
  assign io_iccm_dma_rvalid = iccm_dma_rvalid_temp; // @[el2_ifu_mem_ctl.scala 656:22]
  assign io_iccm_dma_rdata = iccm_dma_rdata_temp; // @[el2_ifu_mem_ctl.scala 660:21]
  assign io_iccm_dma_rtag = iccm_dma_rtag_temp; // @[el2_ifu_mem_ctl.scala 651:20]
  assign io_iccm_ready = _T_2675 & _T_2669; // @[el2_ifu_mem_ctl.scala 630:17]
  assign io_ic_rw_addr = _T_338 | _T_339; // @[el2_ifu_mem_ctl.scala 337:17]
  assign io_ic_wr_en = bus_ic_wr_en & _T_4125; // @[el2_ifu_mem_ctl.scala 698:15]
  assign io_ic_rd_en = _T_4117 | _T_4122; // @[el2_ifu_mem_ctl.scala 689:15]
  assign io_ic_wr_data_0 = ic_wr_16bytes_data[70:0]; // @[el2_ifu_mem_ctl.scala 344:17]
  assign io_ic_wr_data_1 = ic_wr_16bytes_data[141:71]; // @[el2_ifu_mem_ctl.scala 344:17]
  assign io_ic_debug_wr_data = io_dec_tlu_ic_diag_pkt_icache_wrdata; // @[el2_ifu_mem_ctl.scala 345:23]
  assign io_ifu_ic_debug_rd_data = _T_1209; // @[el2_ifu_mem_ctl.scala 353:27]
  assign io_ic_debug_addr = io_dec_tlu_ic_diag_pkt_icache_dicawics[9:0]; // @[el2_ifu_mem_ctl.scala 825:20]
  assign io_ic_debug_rd_en = io_dec_tlu_ic_diag_pkt_icache_rd_valid; // @[el2_ifu_mem_ctl.scala 827:21]
  assign io_ic_debug_wr_en = io_dec_tlu_ic_diag_pkt_icache_wr_valid; // @[el2_ifu_mem_ctl.scala 828:21]
  assign io_ic_debug_tag_array = io_dec_tlu_ic_diag_pkt_icache_dicawics[16]; // @[el2_ifu_mem_ctl.scala 826:25]
  assign io_ic_debug_way = _T_10601[1:0]; // @[el2_ifu_mem_ctl.scala 829:19]
  assign io_ic_tag_valid = ic_tag_valid_unq & _T_10575; // @[el2_ifu_mem_ctl.scala 813:19]
  assign io_iccm_rw_addr = _T_3263 ? io_dma_mem_addr[15:1] : _T_3270; // @[el2_ifu_mem_ctl.scala 662:19]
  assign io_iccm_wren = _T_2679 | iccm_correct_ecc; // @[el2_ifu_mem_ctl.scala 632:16]
  assign io_iccm_rden = _T_2683 | _T_2684; // @[el2_ifu_mem_ctl.scala 633:16]
  assign io_iccm_wr_data = _T_3245 ? _T_3246 : _T_3253; // @[el2_ifu_mem_ctl.scala 639:19]
  assign io_iccm_wr_size = _T_2689 & io_dma_mem_sz; // @[el2_ifu_mem_ctl.scala 635:19]
  assign io_ic_hit_f = _T_263 | _T_264; // @[el2_ifu_mem_ctl.scala 289:15]
  assign io_ic_access_fault_f = _T_2457 & _T_317; // @[el2_ifu_mem_ctl.scala 385:24]
  assign io_ic_access_fault_type_f = io_iccm_rd_ecc_double_err ? 2'h1 : _T_1271; // @[el2_ifu_mem_ctl.scala 386:29]
  assign io_iccm_rd_ecc_single_err = _T_4062 & ifc_fetch_req_f; // @[el2_ifu_mem_ctl.scala 675:29]
  assign io_iccm_rd_ecc_double_err = iccm_dma_ecc_error_in & ifc_iccm_access_f; // @[el2_ifu_mem_ctl.scala 676:29]
  assign io_ic_error_start = _T_1197 | ic_rd_parity_final_err; // @[el2_ifu_mem_ctl.scala 347:21]
  assign io_ifu_async_error_start = io_iccm_rd_ecc_single_err | io_ic_error_start; // @[el2_ifu_mem_ctl.scala 191:28]
  assign io_iccm_dma_sb_error = _T_3 & dma_iccm_req_f; // @[el2_ifu_mem_ctl.scala 190:24]
  assign io_ic_fetch_val_f = {_T_1279,fetch_req_f_qual}; // @[el2_ifu_mem_ctl.scala 389:21]
  assign io_ic_data_f = io_ic_rd_data[31:0]; // @[el2_ifu_mem_ctl.scala 382:16]
  assign io_ic_premux_data = ic_premux_data_temp[63:0]; // @[el2_ifu_mem_ctl.scala 379:21]
  assign io_ic_sel_premux_data = fetch_req_iccm_f | sel_byp_data; // @[el2_ifu_mem_ctl.scala 380:25]
  assign io_ifu_ic_debug_rd_data_valid = _T_10612; // @[el2_ifu_mem_ctl.scala 836:33]
  assign io_iccm_buf_correct_ecc = iccm_correct_ecc & _T_2462; // @[el2_ifu_mem_ctl.scala 479:27]
  assign io_iccm_correction_state = _T_2490 ? 1'h0 : _GEN_60; // @[el2_ifu_mem_ctl.scala 514:28 el2_ifu_mem_ctl.scala 527:32 el2_ifu_mem_ctl.scala 534:32 el2_ifu_mem_ctl.scala 541:32]
  assign io_test = {_T_2873,_T_2870}; // @[el2_ifu_mem_ctl.scala 636:11]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  flush_final_f = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  ifc_fetch_req_f_raw = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  miss_state = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  scnd_miss_req_q = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  ifu_fetch_addr_int_f = _RAND_4[30:0];
  _RAND_5 = {1{`RANDOM}};
  ifc_iccm_access_f = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  iccm_dma_rvalid_in = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  dma_iccm_req_f = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  perr_state = _RAND_8[2:0];
  _RAND_9 = {1{`RANDOM}};
  err_stop_state = _RAND_9[1:0];
  _RAND_10 = {1{`RANDOM}};
  reset_all_tags = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  ifc_region_acc_fault_final_f = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  ifu_bus_rvalid_unq_ff = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  bus_ifu_bus_clk_en_ff = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  uncacheable_miss_ff = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  bus_data_beat_count = _RAND_15[2:0];
  _RAND_16 = {1{`RANDOM}};
  ic_miss_buff_data_valid = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  imb_ff = _RAND_17[30:0];
  _RAND_18 = {1{`RANDOM}};
  last_data_recieved_ff = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  sel_mb_addr_ff = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  way_status_mb_scnd_ff = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  ifu_ic_rw_int_addr_ff = _RAND_21[6:0];
  _RAND_22 = {1{`RANDOM}};
  way_status_out_0 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  way_status_out_1 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  way_status_out_2 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  way_status_out_3 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  way_status_out_4 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  way_status_out_5 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  way_status_out_6 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  way_status_out_7 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  way_status_out_8 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  way_status_out_9 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  way_status_out_10 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  way_status_out_11 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  way_status_out_12 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  way_status_out_13 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  way_status_out_14 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  way_status_out_15 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  way_status_out_16 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  way_status_out_17 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  way_status_out_18 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  way_status_out_19 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  way_status_out_20 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  way_status_out_21 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  way_status_out_22 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  way_status_out_23 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  way_status_out_24 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  way_status_out_25 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  way_status_out_26 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  way_status_out_27 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  way_status_out_28 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  way_status_out_29 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  way_status_out_30 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  way_status_out_31 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  way_status_out_32 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  way_status_out_33 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  way_status_out_34 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  way_status_out_35 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  way_status_out_36 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  way_status_out_37 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  way_status_out_38 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  way_status_out_39 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  way_status_out_40 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  way_status_out_41 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  way_status_out_42 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  way_status_out_43 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  way_status_out_44 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  way_status_out_45 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  way_status_out_46 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  way_status_out_47 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  way_status_out_48 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  way_status_out_49 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  way_status_out_50 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  way_status_out_51 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  way_status_out_52 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  way_status_out_53 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  way_status_out_54 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  way_status_out_55 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  way_status_out_56 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  way_status_out_57 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  way_status_out_58 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  way_status_out_59 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  way_status_out_60 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  way_status_out_61 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  way_status_out_62 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  way_status_out_63 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  way_status_out_64 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  way_status_out_65 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  way_status_out_66 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  way_status_out_67 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  way_status_out_68 = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  way_status_out_69 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  way_status_out_70 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  way_status_out_71 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  way_status_out_72 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  way_status_out_73 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  way_status_out_74 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  way_status_out_75 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  way_status_out_76 = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  way_status_out_77 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  way_status_out_78 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  way_status_out_79 = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  way_status_out_80 = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  way_status_out_81 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  way_status_out_82 = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  way_status_out_83 = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  way_status_out_84 = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  way_status_out_85 = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  way_status_out_86 = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  way_status_out_87 = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  way_status_out_88 = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  way_status_out_89 = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  way_status_out_90 = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  way_status_out_91 = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  way_status_out_92 = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  way_status_out_93 = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  way_status_out_94 = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  way_status_out_95 = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  way_status_out_96 = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  way_status_out_97 = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  way_status_out_98 = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  way_status_out_99 = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  way_status_out_100 = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  way_status_out_101 = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  way_status_out_102 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  way_status_out_103 = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  way_status_out_104 = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  way_status_out_105 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  way_status_out_106 = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  way_status_out_107 = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  way_status_out_108 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  way_status_out_109 = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  way_status_out_110 = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  way_status_out_111 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  way_status_out_112 = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  way_status_out_113 = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  way_status_out_114 = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  way_status_out_115 = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  way_status_out_116 = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  way_status_out_117 = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  way_status_out_118 = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  way_status_out_119 = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  way_status_out_120 = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  way_status_out_121 = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  way_status_out_122 = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  way_status_out_123 = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  way_status_out_124 = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  way_status_out_125 = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  way_status_out_126 = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  way_status_out_127 = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  tagv_mb_scnd_ff = _RAND_150[1:0];
  _RAND_151 = {1{`RANDOM}};
  uncacheable_miss_scnd_ff = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  imb_scnd_ff = _RAND_152[30:0];
  _RAND_153 = {1{`RANDOM}};
  ifu_bus_rid_ff = _RAND_153[2:0];
  _RAND_154 = {1{`RANDOM}};
  ifu_bus_rresp_ff = _RAND_154[1:0];
  _RAND_155 = {1{`RANDOM}};
  ifu_wr_data_comb_err_ff = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  way_status_mb_ff = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  tagv_mb_ff = _RAND_157[1:0];
  _RAND_158 = {1{`RANDOM}};
  reset_ic_ff = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  fetch_uncacheable_ff = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  miss_addr = _RAND_160[25:0];
  _RAND_161 = {1{`RANDOM}};
  ifc_region_acc_fault_f = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  bus_rd_addr_count = _RAND_162[2:0];
  _RAND_163 = {1{`RANDOM}};
  ic_act_miss_f_delayed = _RAND_163[0:0];
  _RAND_164 = {2{`RANDOM}};
  ifu_bus_rdata_ff = _RAND_164[63:0];
  _RAND_165 = {1{`RANDOM}};
  ic_miss_buff_data_0 = _RAND_165[31:0];
  _RAND_166 = {1{`RANDOM}};
  ic_miss_buff_data_1 = _RAND_166[31:0];
  _RAND_167 = {1{`RANDOM}};
  ic_miss_buff_data_2 = _RAND_167[31:0];
  _RAND_168 = {1{`RANDOM}};
  ic_miss_buff_data_3 = _RAND_168[31:0];
  _RAND_169 = {1{`RANDOM}};
  ic_miss_buff_data_4 = _RAND_169[31:0];
  _RAND_170 = {1{`RANDOM}};
  ic_miss_buff_data_5 = _RAND_170[31:0];
  _RAND_171 = {1{`RANDOM}};
  ic_miss_buff_data_6 = _RAND_171[31:0];
  _RAND_172 = {1{`RANDOM}};
  ic_miss_buff_data_7 = _RAND_172[31:0];
  _RAND_173 = {1{`RANDOM}};
  ic_miss_buff_data_8 = _RAND_173[31:0];
  _RAND_174 = {1{`RANDOM}};
  ic_miss_buff_data_9 = _RAND_174[31:0];
  _RAND_175 = {1{`RANDOM}};
  ic_miss_buff_data_10 = _RAND_175[31:0];
  _RAND_176 = {1{`RANDOM}};
  ic_miss_buff_data_11 = _RAND_176[31:0];
  _RAND_177 = {1{`RANDOM}};
  ic_miss_buff_data_12 = _RAND_177[31:0];
  _RAND_178 = {1{`RANDOM}};
  ic_miss_buff_data_13 = _RAND_178[31:0];
  _RAND_179 = {1{`RANDOM}};
  ic_miss_buff_data_14 = _RAND_179[31:0];
  _RAND_180 = {1{`RANDOM}};
  ic_miss_buff_data_15 = _RAND_180[31:0];
  _RAND_181 = {1{`RANDOM}};
  ic_crit_wd_rdy_new_ff = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  ic_miss_buff_data_error = _RAND_182[7:0];
  _RAND_183 = {1{`RANDOM}};
  ic_debug_ict_array_sel_ff = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  ic_tag_valid_out_1_0 = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  ic_tag_valid_out_1_1 = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  ic_tag_valid_out_1_2 = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  ic_tag_valid_out_1_3 = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  ic_tag_valid_out_1_4 = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  ic_tag_valid_out_1_5 = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  ic_tag_valid_out_1_6 = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  ic_tag_valid_out_1_7 = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  ic_tag_valid_out_1_8 = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  ic_tag_valid_out_1_9 = _RAND_193[0:0];
  _RAND_194 = {1{`RANDOM}};
  ic_tag_valid_out_1_10 = _RAND_194[0:0];
  _RAND_195 = {1{`RANDOM}};
  ic_tag_valid_out_1_11 = _RAND_195[0:0];
  _RAND_196 = {1{`RANDOM}};
  ic_tag_valid_out_1_12 = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  ic_tag_valid_out_1_13 = _RAND_197[0:0];
  _RAND_198 = {1{`RANDOM}};
  ic_tag_valid_out_1_14 = _RAND_198[0:0];
  _RAND_199 = {1{`RANDOM}};
  ic_tag_valid_out_1_15 = _RAND_199[0:0];
  _RAND_200 = {1{`RANDOM}};
  ic_tag_valid_out_1_16 = _RAND_200[0:0];
  _RAND_201 = {1{`RANDOM}};
  ic_tag_valid_out_1_17 = _RAND_201[0:0];
  _RAND_202 = {1{`RANDOM}};
  ic_tag_valid_out_1_18 = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  ic_tag_valid_out_1_19 = _RAND_203[0:0];
  _RAND_204 = {1{`RANDOM}};
  ic_tag_valid_out_1_20 = _RAND_204[0:0];
  _RAND_205 = {1{`RANDOM}};
  ic_tag_valid_out_1_21 = _RAND_205[0:0];
  _RAND_206 = {1{`RANDOM}};
  ic_tag_valid_out_1_22 = _RAND_206[0:0];
  _RAND_207 = {1{`RANDOM}};
  ic_tag_valid_out_1_23 = _RAND_207[0:0];
  _RAND_208 = {1{`RANDOM}};
  ic_tag_valid_out_1_24 = _RAND_208[0:0];
  _RAND_209 = {1{`RANDOM}};
  ic_tag_valid_out_1_25 = _RAND_209[0:0];
  _RAND_210 = {1{`RANDOM}};
  ic_tag_valid_out_1_26 = _RAND_210[0:0];
  _RAND_211 = {1{`RANDOM}};
  ic_tag_valid_out_1_27 = _RAND_211[0:0];
  _RAND_212 = {1{`RANDOM}};
  ic_tag_valid_out_1_28 = _RAND_212[0:0];
  _RAND_213 = {1{`RANDOM}};
  ic_tag_valid_out_1_29 = _RAND_213[0:0];
  _RAND_214 = {1{`RANDOM}};
  ic_tag_valid_out_1_30 = _RAND_214[0:0];
  _RAND_215 = {1{`RANDOM}};
  ic_tag_valid_out_1_31 = _RAND_215[0:0];
  _RAND_216 = {1{`RANDOM}};
  ic_tag_valid_out_1_32 = _RAND_216[0:0];
  _RAND_217 = {1{`RANDOM}};
  ic_tag_valid_out_1_33 = _RAND_217[0:0];
  _RAND_218 = {1{`RANDOM}};
  ic_tag_valid_out_1_34 = _RAND_218[0:0];
  _RAND_219 = {1{`RANDOM}};
  ic_tag_valid_out_1_35 = _RAND_219[0:0];
  _RAND_220 = {1{`RANDOM}};
  ic_tag_valid_out_1_36 = _RAND_220[0:0];
  _RAND_221 = {1{`RANDOM}};
  ic_tag_valid_out_1_37 = _RAND_221[0:0];
  _RAND_222 = {1{`RANDOM}};
  ic_tag_valid_out_1_38 = _RAND_222[0:0];
  _RAND_223 = {1{`RANDOM}};
  ic_tag_valid_out_1_39 = _RAND_223[0:0];
  _RAND_224 = {1{`RANDOM}};
  ic_tag_valid_out_1_40 = _RAND_224[0:0];
  _RAND_225 = {1{`RANDOM}};
  ic_tag_valid_out_1_41 = _RAND_225[0:0];
  _RAND_226 = {1{`RANDOM}};
  ic_tag_valid_out_1_42 = _RAND_226[0:0];
  _RAND_227 = {1{`RANDOM}};
  ic_tag_valid_out_1_43 = _RAND_227[0:0];
  _RAND_228 = {1{`RANDOM}};
  ic_tag_valid_out_1_44 = _RAND_228[0:0];
  _RAND_229 = {1{`RANDOM}};
  ic_tag_valid_out_1_45 = _RAND_229[0:0];
  _RAND_230 = {1{`RANDOM}};
  ic_tag_valid_out_1_46 = _RAND_230[0:0];
  _RAND_231 = {1{`RANDOM}};
  ic_tag_valid_out_1_47 = _RAND_231[0:0];
  _RAND_232 = {1{`RANDOM}};
  ic_tag_valid_out_1_48 = _RAND_232[0:0];
  _RAND_233 = {1{`RANDOM}};
  ic_tag_valid_out_1_49 = _RAND_233[0:0];
  _RAND_234 = {1{`RANDOM}};
  ic_tag_valid_out_1_50 = _RAND_234[0:0];
  _RAND_235 = {1{`RANDOM}};
  ic_tag_valid_out_1_51 = _RAND_235[0:0];
  _RAND_236 = {1{`RANDOM}};
  ic_tag_valid_out_1_52 = _RAND_236[0:0];
  _RAND_237 = {1{`RANDOM}};
  ic_tag_valid_out_1_53 = _RAND_237[0:0];
  _RAND_238 = {1{`RANDOM}};
  ic_tag_valid_out_1_54 = _RAND_238[0:0];
  _RAND_239 = {1{`RANDOM}};
  ic_tag_valid_out_1_55 = _RAND_239[0:0];
  _RAND_240 = {1{`RANDOM}};
  ic_tag_valid_out_1_56 = _RAND_240[0:0];
  _RAND_241 = {1{`RANDOM}};
  ic_tag_valid_out_1_57 = _RAND_241[0:0];
  _RAND_242 = {1{`RANDOM}};
  ic_tag_valid_out_1_58 = _RAND_242[0:0];
  _RAND_243 = {1{`RANDOM}};
  ic_tag_valid_out_1_59 = _RAND_243[0:0];
  _RAND_244 = {1{`RANDOM}};
  ic_tag_valid_out_1_60 = _RAND_244[0:0];
  _RAND_245 = {1{`RANDOM}};
  ic_tag_valid_out_1_61 = _RAND_245[0:0];
  _RAND_246 = {1{`RANDOM}};
  ic_tag_valid_out_1_62 = _RAND_246[0:0];
  _RAND_247 = {1{`RANDOM}};
  ic_tag_valid_out_1_63 = _RAND_247[0:0];
  _RAND_248 = {1{`RANDOM}};
  ic_tag_valid_out_1_64 = _RAND_248[0:0];
  _RAND_249 = {1{`RANDOM}};
  ic_tag_valid_out_1_65 = _RAND_249[0:0];
  _RAND_250 = {1{`RANDOM}};
  ic_tag_valid_out_1_66 = _RAND_250[0:0];
  _RAND_251 = {1{`RANDOM}};
  ic_tag_valid_out_1_67 = _RAND_251[0:0];
  _RAND_252 = {1{`RANDOM}};
  ic_tag_valid_out_1_68 = _RAND_252[0:0];
  _RAND_253 = {1{`RANDOM}};
  ic_tag_valid_out_1_69 = _RAND_253[0:0];
  _RAND_254 = {1{`RANDOM}};
  ic_tag_valid_out_1_70 = _RAND_254[0:0];
  _RAND_255 = {1{`RANDOM}};
  ic_tag_valid_out_1_71 = _RAND_255[0:0];
  _RAND_256 = {1{`RANDOM}};
  ic_tag_valid_out_1_72 = _RAND_256[0:0];
  _RAND_257 = {1{`RANDOM}};
  ic_tag_valid_out_1_73 = _RAND_257[0:0];
  _RAND_258 = {1{`RANDOM}};
  ic_tag_valid_out_1_74 = _RAND_258[0:0];
  _RAND_259 = {1{`RANDOM}};
  ic_tag_valid_out_1_75 = _RAND_259[0:0];
  _RAND_260 = {1{`RANDOM}};
  ic_tag_valid_out_1_76 = _RAND_260[0:0];
  _RAND_261 = {1{`RANDOM}};
  ic_tag_valid_out_1_77 = _RAND_261[0:0];
  _RAND_262 = {1{`RANDOM}};
  ic_tag_valid_out_1_78 = _RAND_262[0:0];
  _RAND_263 = {1{`RANDOM}};
  ic_tag_valid_out_1_79 = _RAND_263[0:0];
  _RAND_264 = {1{`RANDOM}};
  ic_tag_valid_out_1_80 = _RAND_264[0:0];
  _RAND_265 = {1{`RANDOM}};
  ic_tag_valid_out_1_81 = _RAND_265[0:0];
  _RAND_266 = {1{`RANDOM}};
  ic_tag_valid_out_1_82 = _RAND_266[0:0];
  _RAND_267 = {1{`RANDOM}};
  ic_tag_valid_out_1_83 = _RAND_267[0:0];
  _RAND_268 = {1{`RANDOM}};
  ic_tag_valid_out_1_84 = _RAND_268[0:0];
  _RAND_269 = {1{`RANDOM}};
  ic_tag_valid_out_1_85 = _RAND_269[0:0];
  _RAND_270 = {1{`RANDOM}};
  ic_tag_valid_out_1_86 = _RAND_270[0:0];
  _RAND_271 = {1{`RANDOM}};
  ic_tag_valid_out_1_87 = _RAND_271[0:0];
  _RAND_272 = {1{`RANDOM}};
  ic_tag_valid_out_1_88 = _RAND_272[0:0];
  _RAND_273 = {1{`RANDOM}};
  ic_tag_valid_out_1_89 = _RAND_273[0:0];
  _RAND_274 = {1{`RANDOM}};
  ic_tag_valid_out_1_90 = _RAND_274[0:0];
  _RAND_275 = {1{`RANDOM}};
  ic_tag_valid_out_1_91 = _RAND_275[0:0];
  _RAND_276 = {1{`RANDOM}};
  ic_tag_valid_out_1_92 = _RAND_276[0:0];
  _RAND_277 = {1{`RANDOM}};
  ic_tag_valid_out_1_93 = _RAND_277[0:0];
  _RAND_278 = {1{`RANDOM}};
  ic_tag_valid_out_1_94 = _RAND_278[0:0];
  _RAND_279 = {1{`RANDOM}};
  ic_tag_valid_out_1_95 = _RAND_279[0:0];
  _RAND_280 = {1{`RANDOM}};
  ic_tag_valid_out_1_96 = _RAND_280[0:0];
  _RAND_281 = {1{`RANDOM}};
  ic_tag_valid_out_1_97 = _RAND_281[0:0];
  _RAND_282 = {1{`RANDOM}};
  ic_tag_valid_out_1_98 = _RAND_282[0:0];
  _RAND_283 = {1{`RANDOM}};
  ic_tag_valid_out_1_99 = _RAND_283[0:0];
  _RAND_284 = {1{`RANDOM}};
  ic_tag_valid_out_1_100 = _RAND_284[0:0];
  _RAND_285 = {1{`RANDOM}};
  ic_tag_valid_out_1_101 = _RAND_285[0:0];
  _RAND_286 = {1{`RANDOM}};
  ic_tag_valid_out_1_102 = _RAND_286[0:0];
  _RAND_287 = {1{`RANDOM}};
  ic_tag_valid_out_1_103 = _RAND_287[0:0];
  _RAND_288 = {1{`RANDOM}};
  ic_tag_valid_out_1_104 = _RAND_288[0:0];
  _RAND_289 = {1{`RANDOM}};
  ic_tag_valid_out_1_105 = _RAND_289[0:0];
  _RAND_290 = {1{`RANDOM}};
  ic_tag_valid_out_1_106 = _RAND_290[0:0];
  _RAND_291 = {1{`RANDOM}};
  ic_tag_valid_out_1_107 = _RAND_291[0:0];
  _RAND_292 = {1{`RANDOM}};
  ic_tag_valid_out_1_108 = _RAND_292[0:0];
  _RAND_293 = {1{`RANDOM}};
  ic_tag_valid_out_1_109 = _RAND_293[0:0];
  _RAND_294 = {1{`RANDOM}};
  ic_tag_valid_out_1_110 = _RAND_294[0:0];
  _RAND_295 = {1{`RANDOM}};
  ic_tag_valid_out_1_111 = _RAND_295[0:0];
  _RAND_296 = {1{`RANDOM}};
  ic_tag_valid_out_1_112 = _RAND_296[0:0];
  _RAND_297 = {1{`RANDOM}};
  ic_tag_valid_out_1_113 = _RAND_297[0:0];
  _RAND_298 = {1{`RANDOM}};
  ic_tag_valid_out_1_114 = _RAND_298[0:0];
  _RAND_299 = {1{`RANDOM}};
  ic_tag_valid_out_1_115 = _RAND_299[0:0];
  _RAND_300 = {1{`RANDOM}};
  ic_tag_valid_out_1_116 = _RAND_300[0:0];
  _RAND_301 = {1{`RANDOM}};
  ic_tag_valid_out_1_117 = _RAND_301[0:0];
  _RAND_302 = {1{`RANDOM}};
  ic_tag_valid_out_1_118 = _RAND_302[0:0];
  _RAND_303 = {1{`RANDOM}};
  ic_tag_valid_out_1_119 = _RAND_303[0:0];
  _RAND_304 = {1{`RANDOM}};
  ic_tag_valid_out_1_120 = _RAND_304[0:0];
  _RAND_305 = {1{`RANDOM}};
  ic_tag_valid_out_1_121 = _RAND_305[0:0];
  _RAND_306 = {1{`RANDOM}};
  ic_tag_valid_out_1_122 = _RAND_306[0:0];
  _RAND_307 = {1{`RANDOM}};
  ic_tag_valid_out_1_123 = _RAND_307[0:0];
  _RAND_308 = {1{`RANDOM}};
  ic_tag_valid_out_1_124 = _RAND_308[0:0];
  _RAND_309 = {1{`RANDOM}};
  ic_tag_valid_out_1_125 = _RAND_309[0:0];
  _RAND_310 = {1{`RANDOM}};
  ic_tag_valid_out_1_126 = _RAND_310[0:0];
  _RAND_311 = {1{`RANDOM}};
  ic_tag_valid_out_1_127 = _RAND_311[0:0];
  _RAND_312 = {1{`RANDOM}};
  ic_tag_valid_out_0_0 = _RAND_312[0:0];
  _RAND_313 = {1{`RANDOM}};
  ic_tag_valid_out_0_1 = _RAND_313[0:0];
  _RAND_314 = {1{`RANDOM}};
  ic_tag_valid_out_0_2 = _RAND_314[0:0];
  _RAND_315 = {1{`RANDOM}};
  ic_tag_valid_out_0_3 = _RAND_315[0:0];
  _RAND_316 = {1{`RANDOM}};
  ic_tag_valid_out_0_4 = _RAND_316[0:0];
  _RAND_317 = {1{`RANDOM}};
  ic_tag_valid_out_0_5 = _RAND_317[0:0];
  _RAND_318 = {1{`RANDOM}};
  ic_tag_valid_out_0_6 = _RAND_318[0:0];
  _RAND_319 = {1{`RANDOM}};
  ic_tag_valid_out_0_7 = _RAND_319[0:0];
  _RAND_320 = {1{`RANDOM}};
  ic_tag_valid_out_0_8 = _RAND_320[0:0];
  _RAND_321 = {1{`RANDOM}};
  ic_tag_valid_out_0_9 = _RAND_321[0:0];
  _RAND_322 = {1{`RANDOM}};
  ic_tag_valid_out_0_10 = _RAND_322[0:0];
  _RAND_323 = {1{`RANDOM}};
  ic_tag_valid_out_0_11 = _RAND_323[0:0];
  _RAND_324 = {1{`RANDOM}};
  ic_tag_valid_out_0_12 = _RAND_324[0:0];
  _RAND_325 = {1{`RANDOM}};
  ic_tag_valid_out_0_13 = _RAND_325[0:0];
  _RAND_326 = {1{`RANDOM}};
  ic_tag_valid_out_0_14 = _RAND_326[0:0];
  _RAND_327 = {1{`RANDOM}};
  ic_tag_valid_out_0_15 = _RAND_327[0:0];
  _RAND_328 = {1{`RANDOM}};
  ic_tag_valid_out_0_16 = _RAND_328[0:0];
  _RAND_329 = {1{`RANDOM}};
  ic_tag_valid_out_0_17 = _RAND_329[0:0];
  _RAND_330 = {1{`RANDOM}};
  ic_tag_valid_out_0_18 = _RAND_330[0:0];
  _RAND_331 = {1{`RANDOM}};
  ic_tag_valid_out_0_19 = _RAND_331[0:0];
  _RAND_332 = {1{`RANDOM}};
  ic_tag_valid_out_0_20 = _RAND_332[0:0];
  _RAND_333 = {1{`RANDOM}};
  ic_tag_valid_out_0_21 = _RAND_333[0:0];
  _RAND_334 = {1{`RANDOM}};
  ic_tag_valid_out_0_22 = _RAND_334[0:0];
  _RAND_335 = {1{`RANDOM}};
  ic_tag_valid_out_0_23 = _RAND_335[0:0];
  _RAND_336 = {1{`RANDOM}};
  ic_tag_valid_out_0_24 = _RAND_336[0:0];
  _RAND_337 = {1{`RANDOM}};
  ic_tag_valid_out_0_25 = _RAND_337[0:0];
  _RAND_338 = {1{`RANDOM}};
  ic_tag_valid_out_0_26 = _RAND_338[0:0];
  _RAND_339 = {1{`RANDOM}};
  ic_tag_valid_out_0_27 = _RAND_339[0:0];
  _RAND_340 = {1{`RANDOM}};
  ic_tag_valid_out_0_28 = _RAND_340[0:0];
  _RAND_341 = {1{`RANDOM}};
  ic_tag_valid_out_0_29 = _RAND_341[0:0];
  _RAND_342 = {1{`RANDOM}};
  ic_tag_valid_out_0_30 = _RAND_342[0:0];
  _RAND_343 = {1{`RANDOM}};
  ic_tag_valid_out_0_31 = _RAND_343[0:0];
  _RAND_344 = {1{`RANDOM}};
  ic_tag_valid_out_0_32 = _RAND_344[0:0];
  _RAND_345 = {1{`RANDOM}};
  ic_tag_valid_out_0_33 = _RAND_345[0:0];
  _RAND_346 = {1{`RANDOM}};
  ic_tag_valid_out_0_34 = _RAND_346[0:0];
  _RAND_347 = {1{`RANDOM}};
  ic_tag_valid_out_0_35 = _RAND_347[0:0];
  _RAND_348 = {1{`RANDOM}};
  ic_tag_valid_out_0_36 = _RAND_348[0:0];
  _RAND_349 = {1{`RANDOM}};
  ic_tag_valid_out_0_37 = _RAND_349[0:0];
  _RAND_350 = {1{`RANDOM}};
  ic_tag_valid_out_0_38 = _RAND_350[0:0];
  _RAND_351 = {1{`RANDOM}};
  ic_tag_valid_out_0_39 = _RAND_351[0:0];
  _RAND_352 = {1{`RANDOM}};
  ic_tag_valid_out_0_40 = _RAND_352[0:0];
  _RAND_353 = {1{`RANDOM}};
  ic_tag_valid_out_0_41 = _RAND_353[0:0];
  _RAND_354 = {1{`RANDOM}};
  ic_tag_valid_out_0_42 = _RAND_354[0:0];
  _RAND_355 = {1{`RANDOM}};
  ic_tag_valid_out_0_43 = _RAND_355[0:0];
  _RAND_356 = {1{`RANDOM}};
  ic_tag_valid_out_0_44 = _RAND_356[0:0];
  _RAND_357 = {1{`RANDOM}};
  ic_tag_valid_out_0_45 = _RAND_357[0:0];
  _RAND_358 = {1{`RANDOM}};
  ic_tag_valid_out_0_46 = _RAND_358[0:0];
  _RAND_359 = {1{`RANDOM}};
  ic_tag_valid_out_0_47 = _RAND_359[0:0];
  _RAND_360 = {1{`RANDOM}};
  ic_tag_valid_out_0_48 = _RAND_360[0:0];
  _RAND_361 = {1{`RANDOM}};
  ic_tag_valid_out_0_49 = _RAND_361[0:0];
  _RAND_362 = {1{`RANDOM}};
  ic_tag_valid_out_0_50 = _RAND_362[0:0];
  _RAND_363 = {1{`RANDOM}};
  ic_tag_valid_out_0_51 = _RAND_363[0:0];
  _RAND_364 = {1{`RANDOM}};
  ic_tag_valid_out_0_52 = _RAND_364[0:0];
  _RAND_365 = {1{`RANDOM}};
  ic_tag_valid_out_0_53 = _RAND_365[0:0];
  _RAND_366 = {1{`RANDOM}};
  ic_tag_valid_out_0_54 = _RAND_366[0:0];
  _RAND_367 = {1{`RANDOM}};
  ic_tag_valid_out_0_55 = _RAND_367[0:0];
  _RAND_368 = {1{`RANDOM}};
  ic_tag_valid_out_0_56 = _RAND_368[0:0];
  _RAND_369 = {1{`RANDOM}};
  ic_tag_valid_out_0_57 = _RAND_369[0:0];
  _RAND_370 = {1{`RANDOM}};
  ic_tag_valid_out_0_58 = _RAND_370[0:0];
  _RAND_371 = {1{`RANDOM}};
  ic_tag_valid_out_0_59 = _RAND_371[0:0];
  _RAND_372 = {1{`RANDOM}};
  ic_tag_valid_out_0_60 = _RAND_372[0:0];
  _RAND_373 = {1{`RANDOM}};
  ic_tag_valid_out_0_61 = _RAND_373[0:0];
  _RAND_374 = {1{`RANDOM}};
  ic_tag_valid_out_0_62 = _RAND_374[0:0];
  _RAND_375 = {1{`RANDOM}};
  ic_tag_valid_out_0_63 = _RAND_375[0:0];
  _RAND_376 = {1{`RANDOM}};
  ic_tag_valid_out_0_64 = _RAND_376[0:0];
  _RAND_377 = {1{`RANDOM}};
  ic_tag_valid_out_0_65 = _RAND_377[0:0];
  _RAND_378 = {1{`RANDOM}};
  ic_tag_valid_out_0_66 = _RAND_378[0:0];
  _RAND_379 = {1{`RANDOM}};
  ic_tag_valid_out_0_67 = _RAND_379[0:0];
  _RAND_380 = {1{`RANDOM}};
  ic_tag_valid_out_0_68 = _RAND_380[0:0];
  _RAND_381 = {1{`RANDOM}};
  ic_tag_valid_out_0_69 = _RAND_381[0:0];
  _RAND_382 = {1{`RANDOM}};
  ic_tag_valid_out_0_70 = _RAND_382[0:0];
  _RAND_383 = {1{`RANDOM}};
  ic_tag_valid_out_0_71 = _RAND_383[0:0];
  _RAND_384 = {1{`RANDOM}};
  ic_tag_valid_out_0_72 = _RAND_384[0:0];
  _RAND_385 = {1{`RANDOM}};
  ic_tag_valid_out_0_73 = _RAND_385[0:0];
  _RAND_386 = {1{`RANDOM}};
  ic_tag_valid_out_0_74 = _RAND_386[0:0];
  _RAND_387 = {1{`RANDOM}};
  ic_tag_valid_out_0_75 = _RAND_387[0:0];
  _RAND_388 = {1{`RANDOM}};
  ic_tag_valid_out_0_76 = _RAND_388[0:0];
  _RAND_389 = {1{`RANDOM}};
  ic_tag_valid_out_0_77 = _RAND_389[0:0];
  _RAND_390 = {1{`RANDOM}};
  ic_tag_valid_out_0_78 = _RAND_390[0:0];
  _RAND_391 = {1{`RANDOM}};
  ic_tag_valid_out_0_79 = _RAND_391[0:0];
  _RAND_392 = {1{`RANDOM}};
  ic_tag_valid_out_0_80 = _RAND_392[0:0];
  _RAND_393 = {1{`RANDOM}};
  ic_tag_valid_out_0_81 = _RAND_393[0:0];
  _RAND_394 = {1{`RANDOM}};
  ic_tag_valid_out_0_82 = _RAND_394[0:0];
  _RAND_395 = {1{`RANDOM}};
  ic_tag_valid_out_0_83 = _RAND_395[0:0];
  _RAND_396 = {1{`RANDOM}};
  ic_tag_valid_out_0_84 = _RAND_396[0:0];
  _RAND_397 = {1{`RANDOM}};
  ic_tag_valid_out_0_85 = _RAND_397[0:0];
  _RAND_398 = {1{`RANDOM}};
  ic_tag_valid_out_0_86 = _RAND_398[0:0];
  _RAND_399 = {1{`RANDOM}};
  ic_tag_valid_out_0_87 = _RAND_399[0:0];
  _RAND_400 = {1{`RANDOM}};
  ic_tag_valid_out_0_88 = _RAND_400[0:0];
  _RAND_401 = {1{`RANDOM}};
  ic_tag_valid_out_0_89 = _RAND_401[0:0];
  _RAND_402 = {1{`RANDOM}};
  ic_tag_valid_out_0_90 = _RAND_402[0:0];
  _RAND_403 = {1{`RANDOM}};
  ic_tag_valid_out_0_91 = _RAND_403[0:0];
  _RAND_404 = {1{`RANDOM}};
  ic_tag_valid_out_0_92 = _RAND_404[0:0];
  _RAND_405 = {1{`RANDOM}};
  ic_tag_valid_out_0_93 = _RAND_405[0:0];
  _RAND_406 = {1{`RANDOM}};
  ic_tag_valid_out_0_94 = _RAND_406[0:0];
  _RAND_407 = {1{`RANDOM}};
  ic_tag_valid_out_0_95 = _RAND_407[0:0];
  _RAND_408 = {1{`RANDOM}};
  ic_tag_valid_out_0_96 = _RAND_408[0:0];
  _RAND_409 = {1{`RANDOM}};
  ic_tag_valid_out_0_97 = _RAND_409[0:0];
  _RAND_410 = {1{`RANDOM}};
  ic_tag_valid_out_0_98 = _RAND_410[0:0];
  _RAND_411 = {1{`RANDOM}};
  ic_tag_valid_out_0_99 = _RAND_411[0:0];
  _RAND_412 = {1{`RANDOM}};
  ic_tag_valid_out_0_100 = _RAND_412[0:0];
  _RAND_413 = {1{`RANDOM}};
  ic_tag_valid_out_0_101 = _RAND_413[0:0];
  _RAND_414 = {1{`RANDOM}};
  ic_tag_valid_out_0_102 = _RAND_414[0:0];
  _RAND_415 = {1{`RANDOM}};
  ic_tag_valid_out_0_103 = _RAND_415[0:0];
  _RAND_416 = {1{`RANDOM}};
  ic_tag_valid_out_0_104 = _RAND_416[0:0];
  _RAND_417 = {1{`RANDOM}};
  ic_tag_valid_out_0_105 = _RAND_417[0:0];
  _RAND_418 = {1{`RANDOM}};
  ic_tag_valid_out_0_106 = _RAND_418[0:0];
  _RAND_419 = {1{`RANDOM}};
  ic_tag_valid_out_0_107 = _RAND_419[0:0];
  _RAND_420 = {1{`RANDOM}};
  ic_tag_valid_out_0_108 = _RAND_420[0:0];
  _RAND_421 = {1{`RANDOM}};
  ic_tag_valid_out_0_109 = _RAND_421[0:0];
  _RAND_422 = {1{`RANDOM}};
  ic_tag_valid_out_0_110 = _RAND_422[0:0];
  _RAND_423 = {1{`RANDOM}};
  ic_tag_valid_out_0_111 = _RAND_423[0:0];
  _RAND_424 = {1{`RANDOM}};
  ic_tag_valid_out_0_112 = _RAND_424[0:0];
  _RAND_425 = {1{`RANDOM}};
  ic_tag_valid_out_0_113 = _RAND_425[0:0];
  _RAND_426 = {1{`RANDOM}};
  ic_tag_valid_out_0_114 = _RAND_426[0:0];
  _RAND_427 = {1{`RANDOM}};
  ic_tag_valid_out_0_115 = _RAND_427[0:0];
  _RAND_428 = {1{`RANDOM}};
  ic_tag_valid_out_0_116 = _RAND_428[0:0];
  _RAND_429 = {1{`RANDOM}};
  ic_tag_valid_out_0_117 = _RAND_429[0:0];
  _RAND_430 = {1{`RANDOM}};
  ic_tag_valid_out_0_118 = _RAND_430[0:0];
  _RAND_431 = {1{`RANDOM}};
  ic_tag_valid_out_0_119 = _RAND_431[0:0];
  _RAND_432 = {1{`RANDOM}};
  ic_tag_valid_out_0_120 = _RAND_432[0:0];
  _RAND_433 = {1{`RANDOM}};
  ic_tag_valid_out_0_121 = _RAND_433[0:0];
  _RAND_434 = {1{`RANDOM}};
  ic_tag_valid_out_0_122 = _RAND_434[0:0];
  _RAND_435 = {1{`RANDOM}};
  ic_tag_valid_out_0_123 = _RAND_435[0:0];
  _RAND_436 = {1{`RANDOM}};
  ic_tag_valid_out_0_124 = _RAND_436[0:0];
  _RAND_437 = {1{`RANDOM}};
  ic_tag_valid_out_0_125 = _RAND_437[0:0];
  _RAND_438 = {1{`RANDOM}};
  ic_tag_valid_out_0_126 = _RAND_438[0:0];
  _RAND_439 = {1{`RANDOM}};
  ic_tag_valid_out_0_127 = _RAND_439[0:0];
  _RAND_440 = {1{`RANDOM}};
  ic_debug_way_ff = _RAND_440[1:0];
  _RAND_441 = {1{`RANDOM}};
  ic_debug_rd_en_ff = _RAND_441[0:0];
  _RAND_442 = {3{`RANDOM}};
  _T_1209 = _RAND_442[70:0];
  _RAND_443 = {1{`RANDOM}};
  perr_ic_index_ff = _RAND_443[6:0];
  _RAND_444 = {1{`RANDOM}};
  dma_sb_err_state_ff = _RAND_444[0:0];
  _RAND_445 = {1{`RANDOM}};
  ifu_bus_cmd_valid = _RAND_445[0:0];
  _RAND_446 = {1{`RANDOM}};
  bus_cmd_beat_count = _RAND_446[2:0];
  _RAND_447 = {1{`RANDOM}};
  ifu_bus_arready_unq_ff = _RAND_447[0:0];
  _RAND_448 = {1{`RANDOM}};
  ifu_bus_arvalid_ff = _RAND_448[0:0];
  _RAND_449 = {1{`RANDOM}};
  ifc_dma_access_ok_prev = _RAND_449[0:0];
  _RAND_450 = {2{`RANDOM}};
  iccm_ecc_corr_data_ff = _RAND_450[38:0];
  _RAND_451 = {1{`RANDOM}};
  dma_mem_addr_ff = _RAND_451[1:0];
  _RAND_452 = {1{`RANDOM}};
  dma_mem_tag_ff = _RAND_452[2:0];
  _RAND_453 = {1{`RANDOM}};
  iccm_dma_rtag_temp = _RAND_453[2:0];
  _RAND_454 = {1{`RANDOM}};
  iccm_dma_rvalid_temp = _RAND_454[0:0];
  _RAND_455 = {2{`RANDOM}};
  iccm_dma_rdata_temp = _RAND_455[63:0];
  _RAND_456 = {1{`RANDOM}};
  iccm_ecc_corr_index_ff = _RAND_456[13:0];
  _RAND_457 = {1{`RANDOM}};
  iccm_rd_ecc_single_err_ff = _RAND_457[0:0];
  _RAND_458 = {1{`RANDOM}};
  iccm_rw_addr_f = _RAND_458[13:0];
  _RAND_459 = {1{`RANDOM}};
  ifu_status_wr_addr_ff = _RAND_459[6:0];
  _RAND_460 = {1{`RANDOM}};
  way_status_wr_en_ff = _RAND_460[0:0];
  _RAND_461 = {1{`RANDOM}};
  way_status_new_ff = _RAND_461[0:0];
  _RAND_462 = {1{`RANDOM}};
  ifu_tag_wren_ff = _RAND_462[1:0];
  _RAND_463 = {1{`RANDOM}};
  ic_valid_ff = _RAND_463[0:0];
  _RAND_464 = {1{`RANDOM}};
  _T_10582 = _RAND_464[0:0];
  _RAND_465 = {1{`RANDOM}};
  _T_10583 = _RAND_465[0:0];
  _RAND_466 = {1{`RANDOM}};
  _T_10584 = _RAND_466[0:0];
  _RAND_467 = {1{`RANDOM}};
  _T_10588 = _RAND_467[0:0];
  _RAND_468 = {1{`RANDOM}};
  _T_10589 = _RAND_468[0:0];
  _RAND_469 = {1{`RANDOM}};
  _T_10612 = _RAND_469[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      flush_final_f <= 1'h0;
    end else begin
      flush_final_f <= io_exu_flush_final;
    end
    if (reset) begin
      ifc_fetch_req_f_raw <= 1'h0;
    end else begin
      ifc_fetch_req_f_raw <= ifc_fetch_req_qual_bf;
    end
    if (reset) begin
      miss_state <= 3'h0;
    end else if (miss_state_en) begin
      if (_T_24) begin
        if (_T_26) begin
          miss_state <= 3'h1;
        end else begin
          miss_state <= 3'h2;
        end
      end else if (_T_31) begin
        if (_T_36) begin
          miss_state <= 3'h0;
        end else if (_T_40) begin
          miss_state <= 3'h3;
        end else if (_T_47) begin
          miss_state <= 3'h4;
        end else if (_T_51) begin
          miss_state <= 3'h0;
        end else if (_T_61) begin
          miss_state <= 3'h6;
        end else if (_T_71) begin
          miss_state <= 3'h6;
        end else if (_T_79) begin
          miss_state <= 3'h0;
        end else if (_T_84) begin
          miss_state <= 3'h2;
        end else begin
          miss_state <= 3'h0;
        end
      end else if (_T_102) begin
        miss_state <= 3'h0;
      end else if (_T_106) begin
        if (_T_113) begin
          miss_state <= 3'h2;
        end else begin
          miss_state <= 3'h0;
        end
      end else if (_T_121) begin
        if (_T_126) begin
          miss_state <= 3'h2;
        end else begin
          miss_state <= 3'h0;
        end
      end else if (_T_132) begin
        if (_T_137) begin
          miss_state <= 3'h5;
        end else if (_T_143) begin
          miss_state <= 3'h7;
        end else begin
          miss_state <= 3'h0;
        end
      end else if (_T_151) begin
        if (io_dec_tlu_force_halt) begin
          miss_state <= 3'h0;
        end else if (io_exu_flush_final) begin
          if (_T_32) begin
            miss_state <= 3'h0;
          end else begin
            miss_state <= 3'h2;
          end
        end else begin
          miss_state <= 3'h1;
        end
      end else if (_T_160) begin
        if (io_dec_tlu_force_halt) begin
          miss_state <= 3'h0;
        end else if (io_exu_flush_final) begin
          if (_T_32) begin
            miss_state <= 3'h0;
          end else begin
            miss_state <= 3'h2;
          end
        end else begin
          miss_state <= 3'h0;
        end
      end else begin
        miss_state <= 3'h0;
      end
    end
    if (reset) begin
      ifu_fetch_addr_int_f <= 31'h0;
    end else begin
      ifu_fetch_addr_int_f <= io_ifc_fetch_addr_bf;
    end
    if (reset) begin
      ifc_iccm_access_f <= 1'h0;
    end else begin
      ifc_iccm_access_f <= io_ifc_iccm_access_bf;
    end
    if (reset) begin
      ifc_region_acc_fault_final_f <= 1'h0;
    end else begin
      ifc_region_acc_fault_final_f <= io_ifc_region_acc_fault_bf;
    end
    if (reset) begin
      ifu_bus_rvalid_unq_ff <= 1'h0;
    end else if (io_ifu_bus_clk_en) begin
      ifu_bus_rvalid_unq_ff <= io_ifu_axi_rvalid;
    end
    if (reset) begin
      uncacheable_miss_ff <= 1'h0;
    end else if (scnd_miss_req) begin
      uncacheable_miss_ff <= uncacheable_miss_scnd_ff;
    end else if (!(sel_hold_imb)) begin
      uncacheable_miss_ff <= io_ifc_fetch_uncacheable_bf;
    end
    if (scnd_miss_req) begin
      imb_ff <= imb_scnd_ff;
    end else if (!(sel_hold_imb)) begin
      imb_ff <= io_ifc_fetch_addr_bf;
    end
    if (reset) begin
      way_status_mb_scnd_ff <= 1'h0;
    end else if (!(_T_19)) begin
      way_status_mb_scnd_ff <= way_status;
    end
    if (reset) begin
      way_status_out_0 <= 1'h0;
    end else if (_T_4173) begin
      way_status_out_0 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_1 <= 1'h0;
    end else if (_T_4178) begin
      way_status_out_1 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_2 <= 1'h0;
    end else if (_T_4183) begin
      way_status_out_2 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_3 <= 1'h0;
    end else if (_T_4188) begin
      way_status_out_3 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_4 <= 1'h0;
    end else if (_T_4193) begin
      way_status_out_4 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_5 <= 1'h0;
    end else if (_T_4198) begin
      way_status_out_5 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_6 <= 1'h0;
    end else if (_T_4203) begin
      way_status_out_6 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_7 <= 1'h0;
    end else if (_T_4208) begin
      way_status_out_7 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_8 <= 1'h0;
    end else if (_T_4213) begin
      way_status_out_8 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_9 <= 1'h0;
    end else if (_T_4218) begin
      way_status_out_9 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_10 <= 1'h0;
    end else if (_T_4223) begin
      way_status_out_10 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_11 <= 1'h0;
    end else if (_T_4228) begin
      way_status_out_11 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_12 <= 1'h0;
    end else if (_T_4233) begin
      way_status_out_12 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_13 <= 1'h0;
    end else if (_T_4238) begin
      way_status_out_13 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_14 <= 1'h0;
    end else if (_T_4243) begin
      way_status_out_14 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_15 <= 1'h0;
    end else if (_T_4248) begin
      way_status_out_15 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_16 <= 1'h0;
    end else if (_T_4253) begin
      way_status_out_16 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_17 <= 1'h0;
    end else if (_T_4258) begin
      way_status_out_17 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_18 <= 1'h0;
    end else if (_T_4263) begin
      way_status_out_18 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_19 <= 1'h0;
    end else if (_T_4268) begin
      way_status_out_19 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_20 <= 1'h0;
    end else if (_T_4273) begin
      way_status_out_20 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_21 <= 1'h0;
    end else if (_T_4278) begin
      way_status_out_21 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_22 <= 1'h0;
    end else if (_T_4283) begin
      way_status_out_22 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_23 <= 1'h0;
    end else if (_T_4288) begin
      way_status_out_23 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_24 <= 1'h0;
    end else if (_T_4293) begin
      way_status_out_24 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_25 <= 1'h0;
    end else if (_T_4298) begin
      way_status_out_25 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_26 <= 1'h0;
    end else if (_T_4303) begin
      way_status_out_26 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_27 <= 1'h0;
    end else if (_T_4308) begin
      way_status_out_27 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_28 <= 1'h0;
    end else if (_T_4313) begin
      way_status_out_28 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_29 <= 1'h0;
    end else if (_T_4318) begin
      way_status_out_29 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_30 <= 1'h0;
    end else if (_T_4323) begin
      way_status_out_30 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_31 <= 1'h0;
    end else if (_T_4328) begin
      way_status_out_31 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_32 <= 1'h0;
    end else if (_T_4333) begin
      way_status_out_32 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_33 <= 1'h0;
    end else if (_T_4338) begin
      way_status_out_33 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_34 <= 1'h0;
    end else if (_T_4343) begin
      way_status_out_34 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_35 <= 1'h0;
    end else if (_T_4348) begin
      way_status_out_35 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_36 <= 1'h0;
    end else if (_T_4353) begin
      way_status_out_36 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_37 <= 1'h0;
    end else if (_T_4358) begin
      way_status_out_37 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_38 <= 1'h0;
    end else if (_T_4363) begin
      way_status_out_38 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_39 <= 1'h0;
    end else if (_T_4368) begin
      way_status_out_39 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_40 <= 1'h0;
    end else if (_T_4373) begin
      way_status_out_40 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_41 <= 1'h0;
    end else if (_T_4378) begin
      way_status_out_41 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_42 <= 1'h0;
    end else if (_T_4383) begin
      way_status_out_42 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_43 <= 1'h0;
    end else if (_T_4388) begin
      way_status_out_43 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_44 <= 1'h0;
    end else if (_T_4393) begin
      way_status_out_44 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_45 <= 1'h0;
    end else if (_T_4398) begin
      way_status_out_45 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_46 <= 1'h0;
    end else if (_T_4403) begin
      way_status_out_46 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_47 <= 1'h0;
    end else if (_T_4408) begin
      way_status_out_47 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_48 <= 1'h0;
    end else if (_T_4413) begin
      way_status_out_48 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_49 <= 1'h0;
    end else if (_T_4418) begin
      way_status_out_49 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_50 <= 1'h0;
    end else if (_T_4423) begin
      way_status_out_50 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_51 <= 1'h0;
    end else if (_T_4428) begin
      way_status_out_51 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_52 <= 1'h0;
    end else if (_T_4433) begin
      way_status_out_52 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_53 <= 1'h0;
    end else if (_T_4438) begin
      way_status_out_53 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_54 <= 1'h0;
    end else if (_T_4443) begin
      way_status_out_54 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_55 <= 1'h0;
    end else if (_T_4448) begin
      way_status_out_55 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_56 <= 1'h0;
    end else if (_T_4453) begin
      way_status_out_56 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_57 <= 1'h0;
    end else if (_T_4458) begin
      way_status_out_57 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_58 <= 1'h0;
    end else if (_T_4463) begin
      way_status_out_58 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_59 <= 1'h0;
    end else if (_T_4468) begin
      way_status_out_59 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_60 <= 1'h0;
    end else if (_T_4473) begin
      way_status_out_60 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_61 <= 1'h0;
    end else if (_T_4478) begin
      way_status_out_61 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_62 <= 1'h0;
    end else if (_T_4483) begin
      way_status_out_62 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_63 <= 1'h0;
    end else if (_T_4488) begin
      way_status_out_63 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_64 <= 1'h0;
    end else if (_T_4493) begin
      way_status_out_64 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_65 <= 1'h0;
    end else if (_T_4498) begin
      way_status_out_65 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_66 <= 1'h0;
    end else if (_T_4503) begin
      way_status_out_66 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_67 <= 1'h0;
    end else if (_T_4508) begin
      way_status_out_67 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_68 <= 1'h0;
    end else if (_T_4513) begin
      way_status_out_68 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_69 <= 1'h0;
    end else if (_T_4518) begin
      way_status_out_69 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_70 <= 1'h0;
    end else if (_T_4523) begin
      way_status_out_70 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_71 <= 1'h0;
    end else if (_T_4528) begin
      way_status_out_71 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_72 <= 1'h0;
    end else if (_T_4533) begin
      way_status_out_72 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_73 <= 1'h0;
    end else if (_T_4538) begin
      way_status_out_73 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_74 <= 1'h0;
    end else if (_T_4543) begin
      way_status_out_74 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_75 <= 1'h0;
    end else if (_T_4548) begin
      way_status_out_75 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_76 <= 1'h0;
    end else if (_T_4553) begin
      way_status_out_76 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_77 <= 1'h0;
    end else if (_T_4558) begin
      way_status_out_77 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_78 <= 1'h0;
    end else if (_T_4563) begin
      way_status_out_78 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_79 <= 1'h0;
    end else if (_T_4568) begin
      way_status_out_79 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_80 <= 1'h0;
    end else if (_T_4573) begin
      way_status_out_80 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_81 <= 1'h0;
    end else if (_T_4578) begin
      way_status_out_81 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_82 <= 1'h0;
    end else if (_T_4583) begin
      way_status_out_82 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_83 <= 1'h0;
    end else if (_T_4588) begin
      way_status_out_83 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_84 <= 1'h0;
    end else if (_T_4593) begin
      way_status_out_84 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_85 <= 1'h0;
    end else if (_T_4598) begin
      way_status_out_85 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_86 <= 1'h0;
    end else if (_T_4603) begin
      way_status_out_86 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_87 <= 1'h0;
    end else if (_T_4608) begin
      way_status_out_87 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_88 <= 1'h0;
    end else if (_T_4613) begin
      way_status_out_88 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_89 <= 1'h0;
    end else if (_T_4618) begin
      way_status_out_89 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_90 <= 1'h0;
    end else if (_T_4623) begin
      way_status_out_90 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_91 <= 1'h0;
    end else if (_T_4628) begin
      way_status_out_91 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_92 <= 1'h0;
    end else if (_T_4633) begin
      way_status_out_92 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_93 <= 1'h0;
    end else if (_T_4638) begin
      way_status_out_93 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_94 <= 1'h0;
    end else if (_T_4643) begin
      way_status_out_94 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_95 <= 1'h0;
    end else if (_T_4648) begin
      way_status_out_95 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_96 <= 1'h0;
    end else if (_T_4653) begin
      way_status_out_96 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_97 <= 1'h0;
    end else if (_T_4658) begin
      way_status_out_97 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_98 <= 1'h0;
    end else if (_T_4663) begin
      way_status_out_98 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_99 <= 1'h0;
    end else if (_T_4668) begin
      way_status_out_99 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_100 <= 1'h0;
    end else if (_T_4673) begin
      way_status_out_100 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_101 <= 1'h0;
    end else if (_T_4678) begin
      way_status_out_101 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_102 <= 1'h0;
    end else if (_T_4683) begin
      way_status_out_102 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_103 <= 1'h0;
    end else if (_T_4688) begin
      way_status_out_103 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_104 <= 1'h0;
    end else if (_T_4693) begin
      way_status_out_104 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_105 <= 1'h0;
    end else if (_T_4698) begin
      way_status_out_105 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_106 <= 1'h0;
    end else if (_T_4703) begin
      way_status_out_106 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_107 <= 1'h0;
    end else if (_T_4708) begin
      way_status_out_107 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_108 <= 1'h0;
    end else if (_T_4713) begin
      way_status_out_108 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_109 <= 1'h0;
    end else if (_T_4718) begin
      way_status_out_109 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_110 <= 1'h0;
    end else if (_T_4723) begin
      way_status_out_110 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_111 <= 1'h0;
    end else if (_T_4728) begin
      way_status_out_111 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_112 <= 1'h0;
    end else if (_T_4733) begin
      way_status_out_112 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_113 <= 1'h0;
    end else if (_T_4738) begin
      way_status_out_113 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_114 <= 1'h0;
    end else if (_T_4743) begin
      way_status_out_114 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_115 <= 1'h0;
    end else if (_T_4748) begin
      way_status_out_115 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_116 <= 1'h0;
    end else if (_T_4753) begin
      way_status_out_116 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_117 <= 1'h0;
    end else if (_T_4758) begin
      way_status_out_117 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_118 <= 1'h0;
    end else if (_T_4763) begin
      way_status_out_118 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_119 <= 1'h0;
    end else if (_T_4768) begin
      way_status_out_119 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_120 <= 1'h0;
    end else if (_T_4773) begin
      way_status_out_120 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_121 <= 1'h0;
    end else if (_T_4778) begin
      way_status_out_121 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_122 <= 1'h0;
    end else if (_T_4783) begin
      way_status_out_122 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_123 <= 1'h0;
    end else if (_T_4788) begin
      way_status_out_123 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_124 <= 1'h0;
    end else if (_T_4793) begin
      way_status_out_124 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_125 <= 1'h0;
    end else if (_T_4798) begin
      way_status_out_125 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_126 <= 1'h0;
    end else if (_T_4803) begin
      way_status_out_126 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_127 <= 1'h0;
    end else if (_T_4808) begin
      way_status_out_127 <= way_status_new_ff;
    end
    if (reset) begin
      tagv_mb_scnd_ff <= 2'h0;
    end else if (!(_T_19)) begin
      tagv_mb_scnd_ff <= _T_198;
    end
    if (reset) begin
      uncacheable_miss_scnd_ff <= 1'h0;
    end else if (!(sel_hold_imb_scnd)) begin
      uncacheable_miss_scnd_ff <= io_ifc_fetch_uncacheable_bf;
    end
    if (reset) begin
      imb_scnd_ff <= 31'h0;
    end else if (!(sel_hold_imb_scnd)) begin
      imb_scnd_ff <= io_ifc_fetch_addr_bf;
    end
    if (reset) begin
      ifu_bus_rid_ff <= 3'h0;
    end else if (io_ifu_bus_clk_en) begin
      ifu_bus_rid_ff <= io_ifu_axi_rid;
    end
    if (reset) begin
      ifu_bus_rresp_ff <= 2'h0;
    end else if (io_ifu_bus_clk_en) begin
      ifu_bus_rresp_ff <= io_ifu_axi_rresp;
    end
    if (reset) begin
      way_status_mb_ff <= 1'h0;
    end else if (_T_278) begin
      way_status_mb_ff <= way_status_mb_scnd_ff;
    end else if (_T_280) begin
      way_status_mb_ff <= replace_way_mb_any_0;
    end else if (!(miss_pending)) begin
      way_status_mb_ff <= way_status;
    end
    if (reset) begin
      tagv_mb_ff <= 2'h0;
    end else if (scnd_miss_req) begin
      tagv_mb_ff <= _T_290;
    end else if (!(miss_pending)) begin
      tagv_mb_ff <= _T_295;
    end
    reset_ic_ff <= _T_298 & _T_299;
    if (reset) begin
      fetch_uncacheable_ff <= 1'h0;
    end else begin
      fetch_uncacheable_ff <= io_ifc_fetch_uncacheable_bf;
    end
    if (reset) begin
      miss_addr <= 26'h0;
    end else if (_T_231) begin
      miss_addr <= imb_ff[30:5];
    end else if (scnd_miss_req_q) begin
      miss_addr <= imb_scnd_ff[30:5];
    end
    if (reset) begin
      ifc_region_acc_fault_f <= 1'h0;
    end else begin
      ifc_region_acc_fault_f <= io_ifc_region_acc_fault_bf;
    end
    if (reset) begin
      bus_rd_addr_count <= 3'h0;
    end else if (_T_2615) begin
      if (_T_231) begin
        bus_rd_addr_count <= imb_ff[4:2];
      end else if (scnd_miss_req_q) begin
        bus_rd_addr_count <= imb_scnd_ff[4:2];
      end else if (bus_cmd_sent) begin
        bus_rd_addr_count <= _T_2611;
      end
    end
    if (reset) begin
      ifu_bus_rdata_ff <= 64'h0;
    end else if (io_ifu_bus_clk_en) begin
      ifu_bus_rdata_ff <= io_ifu_axi_rdata;
    end
    if (reset) begin
      ic_miss_buff_data_0 <= 32'h0;
    end else if (write_fill_data_0) begin
      ic_miss_buff_data_0 <= io_ifu_axi_rdata[31:0];
    end
    if (reset) begin
      ic_miss_buff_data_1 <= 32'h0;
    end else if (write_fill_data_0) begin
      ic_miss_buff_data_1 <= io_ifu_axi_rdata[63:32];
    end
    if (reset) begin
      ic_miss_buff_data_2 <= 32'h0;
    end else if (write_fill_data_1) begin
      ic_miss_buff_data_2 <= io_ifu_axi_rdata[31:0];
    end
    if (reset) begin
      ic_miss_buff_data_3 <= 32'h0;
    end else if (write_fill_data_1) begin
      ic_miss_buff_data_3 <= io_ifu_axi_rdata[63:32];
    end
    if (reset) begin
      ic_miss_buff_data_4 <= 32'h0;
    end else if (write_fill_data_2) begin
      ic_miss_buff_data_4 <= io_ifu_axi_rdata[31:0];
    end
    if (reset) begin
      ic_miss_buff_data_5 <= 32'h0;
    end else if (write_fill_data_2) begin
      ic_miss_buff_data_5 <= io_ifu_axi_rdata[63:32];
    end
    if (reset) begin
      ic_miss_buff_data_6 <= 32'h0;
    end else if (write_fill_data_3) begin
      ic_miss_buff_data_6 <= io_ifu_axi_rdata[31:0];
    end
    if (reset) begin
      ic_miss_buff_data_7 <= 32'h0;
    end else if (write_fill_data_3) begin
      ic_miss_buff_data_7 <= io_ifu_axi_rdata[63:32];
    end
    if (reset) begin
      ic_miss_buff_data_8 <= 32'h0;
    end else if (write_fill_data_4) begin
      ic_miss_buff_data_8 <= io_ifu_axi_rdata[31:0];
    end
    if (reset) begin
      ic_miss_buff_data_9 <= 32'h0;
    end else if (write_fill_data_4) begin
      ic_miss_buff_data_9 <= io_ifu_axi_rdata[63:32];
    end
    if (reset) begin
      ic_miss_buff_data_10 <= 32'h0;
    end else if (write_fill_data_5) begin
      ic_miss_buff_data_10 <= io_ifu_axi_rdata[31:0];
    end
    if (reset) begin
      ic_miss_buff_data_11 <= 32'h0;
    end else if (write_fill_data_5) begin
      ic_miss_buff_data_11 <= io_ifu_axi_rdata[63:32];
    end
    if (reset) begin
      ic_miss_buff_data_12 <= 32'h0;
    end else if (write_fill_data_6) begin
      ic_miss_buff_data_12 <= io_ifu_axi_rdata[31:0];
    end
    if (reset) begin
      ic_miss_buff_data_13 <= 32'h0;
    end else if (write_fill_data_6) begin
      ic_miss_buff_data_13 <= io_ifu_axi_rdata[63:32];
    end
    if (reset) begin
      ic_miss_buff_data_14 <= 32'h0;
    end else if (write_fill_data_7) begin
      ic_miss_buff_data_14 <= io_ifu_axi_rdata[31:0];
    end
    if (reset) begin
      ic_miss_buff_data_15 <= 32'h0;
    end else if (write_fill_data_7) begin
      ic_miss_buff_data_15 <= io_ifu_axi_rdata[63:32];
    end
    if (reset) begin
      ic_debug_ict_array_sel_ff <= 1'h0;
    end else if (debug_c1_clken) begin
      ic_debug_ict_array_sel_ff <= ic_debug_ict_array_sel_in;
    end
    if (reset) begin
      ic_tag_valid_out_1_0 <= 1'h0;
    end else if (_T_5979) begin
      ic_tag_valid_out_1_0 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_1 <= 1'h0;
    end else if (_T_5996) begin
      ic_tag_valid_out_1_1 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_2 <= 1'h0;
    end else if (_T_6013) begin
      ic_tag_valid_out_1_2 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_3 <= 1'h0;
    end else if (_T_6030) begin
      ic_tag_valid_out_1_3 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_4 <= 1'h0;
    end else if (_T_6047) begin
      ic_tag_valid_out_1_4 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_5 <= 1'h0;
    end else if (_T_6064) begin
      ic_tag_valid_out_1_5 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_6 <= 1'h0;
    end else if (_T_6081) begin
      ic_tag_valid_out_1_6 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_7 <= 1'h0;
    end else if (_T_6098) begin
      ic_tag_valid_out_1_7 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_8 <= 1'h0;
    end else if (_T_6115) begin
      ic_tag_valid_out_1_8 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_9 <= 1'h0;
    end else if (_T_6132) begin
      ic_tag_valid_out_1_9 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_10 <= 1'h0;
    end else if (_T_6149) begin
      ic_tag_valid_out_1_10 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_11 <= 1'h0;
    end else if (_T_6166) begin
      ic_tag_valid_out_1_11 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_12 <= 1'h0;
    end else if (_T_6183) begin
      ic_tag_valid_out_1_12 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_13 <= 1'h0;
    end else if (_T_6200) begin
      ic_tag_valid_out_1_13 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_14 <= 1'h0;
    end else if (_T_6217) begin
      ic_tag_valid_out_1_14 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_15 <= 1'h0;
    end else if (_T_6234) begin
      ic_tag_valid_out_1_15 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_16 <= 1'h0;
    end else if (_T_6251) begin
      ic_tag_valid_out_1_16 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_17 <= 1'h0;
    end else if (_T_6268) begin
      ic_tag_valid_out_1_17 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_18 <= 1'h0;
    end else if (_T_6285) begin
      ic_tag_valid_out_1_18 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_19 <= 1'h0;
    end else if (_T_6302) begin
      ic_tag_valid_out_1_19 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_20 <= 1'h0;
    end else if (_T_6319) begin
      ic_tag_valid_out_1_20 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_21 <= 1'h0;
    end else if (_T_6336) begin
      ic_tag_valid_out_1_21 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_22 <= 1'h0;
    end else if (_T_6353) begin
      ic_tag_valid_out_1_22 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_23 <= 1'h0;
    end else if (_T_6370) begin
      ic_tag_valid_out_1_23 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_24 <= 1'h0;
    end else if (_T_6387) begin
      ic_tag_valid_out_1_24 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_25 <= 1'h0;
    end else if (_T_6404) begin
      ic_tag_valid_out_1_25 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_26 <= 1'h0;
    end else if (_T_6421) begin
      ic_tag_valid_out_1_26 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_27 <= 1'h0;
    end else if (_T_6438) begin
      ic_tag_valid_out_1_27 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_28 <= 1'h0;
    end else if (_T_6455) begin
      ic_tag_valid_out_1_28 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_29 <= 1'h0;
    end else if (_T_6472) begin
      ic_tag_valid_out_1_29 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_30 <= 1'h0;
    end else if (_T_6489) begin
      ic_tag_valid_out_1_30 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_31 <= 1'h0;
    end else if (_T_6506) begin
      ic_tag_valid_out_1_31 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_32 <= 1'h0;
    end else if (_T_7067) begin
      ic_tag_valid_out_1_32 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_33 <= 1'h0;
    end else if (_T_7084) begin
      ic_tag_valid_out_1_33 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_34 <= 1'h0;
    end else if (_T_7101) begin
      ic_tag_valid_out_1_34 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_35 <= 1'h0;
    end else if (_T_7118) begin
      ic_tag_valid_out_1_35 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_36 <= 1'h0;
    end else if (_T_7135) begin
      ic_tag_valid_out_1_36 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_37 <= 1'h0;
    end else if (_T_7152) begin
      ic_tag_valid_out_1_37 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_38 <= 1'h0;
    end else if (_T_7169) begin
      ic_tag_valid_out_1_38 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_39 <= 1'h0;
    end else if (_T_7186) begin
      ic_tag_valid_out_1_39 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_40 <= 1'h0;
    end else if (_T_7203) begin
      ic_tag_valid_out_1_40 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_41 <= 1'h0;
    end else if (_T_7220) begin
      ic_tag_valid_out_1_41 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_42 <= 1'h0;
    end else if (_T_7237) begin
      ic_tag_valid_out_1_42 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_43 <= 1'h0;
    end else if (_T_7254) begin
      ic_tag_valid_out_1_43 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_44 <= 1'h0;
    end else if (_T_7271) begin
      ic_tag_valid_out_1_44 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_45 <= 1'h0;
    end else if (_T_7288) begin
      ic_tag_valid_out_1_45 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_46 <= 1'h0;
    end else if (_T_7305) begin
      ic_tag_valid_out_1_46 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_47 <= 1'h0;
    end else if (_T_7322) begin
      ic_tag_valid_out_1_47 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_48 <= 1'h0;
    end else if (_T_7339) begin
      ic_tag_valid_out_1_48 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_49 <= 1'h0;
    end else if (_T_7356) begin
      ic_tag_valid_out_1_49 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_50 <= 1'h0;
    end else if (_T_7373) begin
      ic_tag_valid_out_1_50 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_51 <= 1'h0;
    end else if (_T_7390) begin
      ic_tag_valid_out_1_51 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_52 <= 1'h0;
    end else if (_T_7407) begin
      ic_tag_valid_out_1_52 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_53 <= 1'h0;
    end else if (_T_7424) begin
      ic_tag_valid_out_1_53 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_54 <= 1'h0;
    end else if (_T_7441) begin
      ic_tag_valid_out_1_54 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_55 <= 1'h0;
    end else if (_T_7458) begin
      ic_tag_valid_out_1_55 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_56 <= 1'h0;
    end else if (_T_7475) begin
      ic_tag_valid_out_1_56 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_57 <= 1'h0;
    end else if (_T_7492) begin
      ic_tag_valid_out_1_57 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_58 <= 1'h0;
    end else if (_T_7509) begin
      ic_tag_valid_out_1_58 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_59 <= 1'h0;
    end else if (_T_7526) begin
      ic_tag_valid_out_1_59 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_60 <= 1'h0;
    end else if (_T_7543) begin
      ic_tag_valid_out_1_60 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_61 <= 1'h0;
    end else if (_T_7560) begin
      ic_tag_valid_out_1_61 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_62 <= 1'h0;
    end else if (_T_7577) begin
      ic_tag_valid_out_1_62 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_63 <= 1'h0;
    end else if (_T_7594) begin
      ic_tag_valid_out_1_63 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_64 <= 1'h0;
    end else if (_T_8155) begin
      ic_tag_valid_out_1_64 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_65 <= 1'h0;
    end else if (_T_8172) begin
      ic_tag_valid_out_1_65 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_66 <= 1'h0;
    end else if (_T_8189) begin
      ic_tag_valid_out_1_66 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_67 <= 1'h0;
    end else if (_T_8206) begin
      ic_tag_valid_out_1_67 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_68 <= 1'h0;
    end else if (_T_8223) begin
      ic_tag_valid_out_1_68 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_69 <= 1'h0;
    end else if (_T_8240) begin
      ic_tag_valid_out_1_69 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_70 <= 1'h0;
    end else if (_T_8257) begin
      ic_tag_valid_out_1_70 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_71 <= 1'h0;
    end else if (_T_8274) begin
      ic_tag_valid_out_1_71 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_72 <= 1'h0;
    end else if (_T_8291) begin
      ic_tag_valid_out_1_72 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_73 <= 1'h0;
    end else if (_T_8308) begin
      ic_tag_valid_out_1_73 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_74 <= 1'h0;
    end else if (_T_8325) begin
      ic_tag_valid_out_1_74 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_75 <= 1'h0;
    end else if (_T_8342) begin
      ic_tag_valid_out_1_75 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_76 <= 1'h0;
    end else if (_T_8359) begin
      ic_tag_valid_out_1_76 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_77 <= 1'h0;
    end else if (_T_8376) begin
      ic_tag_valid_out_1_77 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_78 <= 1'h0;
    end else if (_T_8393) begin
      ic_tag_valid_out_1_78 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_79 <= 1'h0;
    end else if (_T_8410) begin
      ic_tag_valid_out_1_79 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_80 <= 1'h0;
    end else if (_T_8427) begin
      ic_tag_valid_out_1_80 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_81 <= 1'h0;
    end else if (_T_8444) begin
      ic_tag_valid_out_1_81 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_82 <= 1'h0;
    end else if (_T_8461) begin
      ic_tag_valid_out_1_82 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_83 <= 1'h0;
    end else if (_T_8478) begin
      ic_tag_valid_out_1_83 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_84 <= 1'h0;
    end else if (_T_8495) begin
      ic_tag_valid_out_1_84 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_85 <= 1'h0;
    end else if (_T_8512) begin
      ic_tag_valid_out_1_85 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_86 <= 1'h0;
    end else if (_T_8529) begin
      ic_tag_valid_out_1_86 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_87 <= 1'h0;
    end else if (_T_8546) begin
      ic_tag_valid_out_1_87 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_88 <= 1'h0;
    end else if (_T_8563) begin
      ic_tag_valid_out_1_88 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_89 <= 1'h0;
    end else if (_T_8580) begin
      ic_tag_valid_out_1_89 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_90 <= 1'h0;
    end else if (_T_8597) begin
      ic_tag_valid_out_1_90 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_91 <= 1'h0;
    end else if (_T_8614) begin
      ic_tag_valid_out_1_91 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_92 <= 1'h0;
    end else if (_T_8631) begin
      ic_tag_valid_out_1_92 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_93 <= 1'h0;
    end else if (_T_8648) begin
      ic_tag_valid_out_1_93 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_94 <= 1'h0;
    end else if (_T_8665) begin
      ic_tag_valid_out_1_94 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_95 <= 1'h0;
    end else if (_T_8682) begin
      ic_tag_valid_out_1_95 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_96 <= 1'h0;
    end else if (_T_9243) begin
      ic_tag_valid_out_1_96 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_97 <= 1'h0;
    end else if (_T_9260) begin
      ic_tag_valid_out_1_97 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_98 <= 1'h0;
    end else if (_T_9277) begin
      ic_tag_valid_out_1_98 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_99 <= 1'h0;
    end else if (_T_9294) begin
      ic_tag_valid_out_1_99 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_100 <= 1'h0;
    end else if (_T_9311) begin
      ic_tag_valid_out_1_100 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_101 <= 1'h0;
    end else if (_T_9328) begin
      ic_tag_valid_out_1_101 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_102 <= 1'h0;
    end else if (_T_9345) begin
      ic_tag_valid_out_1_102 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_103 <= 1'h0;
    end else if (_T_9362) begin
      ic_tag_valid_out_1_103 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_104 <= 1'h0;
    end else if (_T_9379) begin
      ic_tag_valid_out_1_104 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_105 <= 1'h0;
    end else if (_T_9396) begin
      ic_tag_valid_out_1_105 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_106 <= 1'h0;
    end else if (_T_9413) begin
      ic_tag_valid_out_1_106 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_107 <= 1'h0;
    end else if (_T_9430) begin
      ic_tag_valid_out_1_107 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_108 <= 1'h0;
    end else if (_T_9447) begin
      ic_tag_valid_out_1_108 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_109 <= 1'h0;
    end else if (_T_9464) begin
      ic_tag_valid_out_1_109 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_110 <= 1'h0;
    end else if (_T_9481) begin
      ic_tag_valid_out_1_110 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_111 <= 1'h0;
    end else if (_T_9498) begin
      ic_tag_valid_out_1_111 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_112 <= 1'h0;
    end else if (_T_9515) begin
      ic_tag_valid_out_1_112 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_113 <= 1'h0;
    end else if (_T_9532) begin
      ic_tag_valid_out_1_113 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_114 <= 1'h0;
    end else if (_T_9549) begin
      ic_tag_valid_out_1_114 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_115 <= 1'h0;
    end else if (_T_9566) begin
      ic_tag_valid_out_1_115 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_116 <= 1'h0;
    end else if (_T_9583) begin
      ic_tag_valid_out_1_116 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_117 <= 1'h0;
    end else if (_T_9600) begin
      ic_tag_valid_out_1_117 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_118 <= 1'h0;
    end else if (_T_9617) begin
      ic_tag_valid_out_1_118 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_119 <= 1'h0;
    end else if (_T_9634) begin
      ic_tag_valid_out_1_119 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_120 <= 1'h0;
    end else if (_T_9651) begin
      ic_tag_valid_out_1_120 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_121 <= 1'h0;
    end else if (_T_9668) begin
      ic_tag_valid_out_1_121 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_122 <= 1'h0;
    end else if (_T_9685) begin
      ic_tag_valid_out_1_122 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_123 <= 1'h0;
    end else if (_T_9702) begin
      ic_tag_valid_out_1_123 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_124 <= 1'h0;
    end else if (_T_9719) begin
      ic_tag_valid_out_1_124 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_125 <= 1'h0;
    end else if (_T_9736) begin
      ic_tag_valid_out_1_125 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_126 <= 1'h0;
    end else if (_T_9753) begin
      ic_tag_valid_out_1_126 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_1_127 <= 1'h0;
    end else if (_T_9770) begin
      ic_tag_valid_out_1_127 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_0 <= 1'h0;
    end else if (_T_5435) begin
      ic_tag_valid_out_0_0 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_1 <= 1'h0;
    end else if (_T_5452) begin
      ic_tag_valid_out_0_1 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_2 <= 1'h0;
    end else if (_T_5469) begin
      ic_tag_valid_out_0_2 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_3 <= 1'h0;
    end else if (_T_5486) begin
      ic_tag_valid_out_0_3 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_4 <= 1'h0;
    end else if (_T_5503) begin
      ic_tag_valid_out_0_4 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_5 <= 1'h0;
    end else if (_T_5520) begin
      ic_tag_valid_out_0_5 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_6 <= 1'h0;
    end else if (_T_5537) begin
      ic_tag_valid_out_0_6 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_7 <= 1'h0;
    end else if (_T_5554) begin
      ic_tag_valid_out_0_7 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_8 <= 1'h0;
    end else if (_T_5571) begin
      ic_tag_valid_out_0_8 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_9 <= 1'h0;
    end else if (_T_5588) begin
      ic_tag_valid_out_0_9 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_10 <= 1'h0;
    end else if (_T_5605) begin
      ic_tag_valid_out_0_10 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_11 <= 1'h0;
    end else if (_T_5622) begin
      ic_tag_valid_out_0_11 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_12 <= 1'h0;
    end else if (_T_5639) begin
      ic_tag_valid_out_0_12 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_13 <= 1'h0;
    end else if (_T_5656) begin
      ic_tag_valid_out_0_13 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_14 <= 1'h0;
    end else if (_T_5673) begin
      ic_tag_valid_out_0_14 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_15 <= 1'h0;
    end else if (_T_5690) begin
      ic_tag_valid_out_0_15 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_16 <= 1'h0;
    end else if (_T_5707) begin
      ic_tag_valid_out_0_16 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_17 <= 1'h0;
    end else if (_T_5724) begin
      ic_tag_valid_out_0_17 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_18 <= 1'h0;
    end else if (_T_5741) begin
      ic_tag_valid_out_0_18 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_19 <= 1'h0;
    end else if (_T_5758) begin
      ic_tag_valid_out_0_19 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_20 <= 1'h0;
    end else if (_T_5775) begin
      ic_tag_valid_out_0_20 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_21 <= 1'h0;
    end else if (_T_5792) begin
      ic_tag_valid_out_0_21 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_22 <= 1'h0;
    end else if (_T_5809) begin
      ic_tag_valid_out_0_22 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_23 <= 1'h0;
    end else if (_T_5826) begin
      ic_tag_valid_out_0_23 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_24 <= 1'h0;
    end else if (_T_5843) begin
      ic_tag_valid_out_0_24 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_25 <= 1'h0;
    end else if (_T_5860) begin
      ic_tag_valid_out_0_25 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_26 <= 1'h0;
    end else if (_T_5877) begin
      ic_tag_valid_out_0_26 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_27 <= 1'h0;
    end else if (_T_5894) begin
      ic_tag_valid_out_0_27 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_28 <= 1'h0;
    end else if (_T_5911) begin
      ic_tag_valid_out_0_28 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_29 <= 1'h0;
    end else if (_T_5928) begin
      ic_tag_valid_out_0_29 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_30 <= 1'h0;
    end else if (_T_5945) begin
      ic_tag_valid_out_0_30 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_31 <= 1'h0;
    end else if (_T_5962) begin
      ic_tag_valid_out_0_31 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_32 <= 1'h0;
    end else if (_T_6523) begin
      ic_tag_valid_out_0_32 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_33 <= 1'h0;
    end else if (_T_6540) begin
      ic_tag_valid_out_0_33 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_34 <= 1'h0;
    end else if (_T_6557) begin
      ic_tag_valid_out_0_34 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_35 <= 1'h0;
    end else if (_T_6574) begin
      ic_tag_valid_out_0_35 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_36 <= 1'h0;
    end else if (_T_6591) begin
      ic_tag_valid_out_0_36 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_37 <= 1'h0;
    end else if (_T_6608) begin
      ic_tag_valid_out_0_37 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_38 <= 1'h0;
    end else if (_T_6625) begin
      ic_tag_valid_out_0_38 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_39 <= 1'h0;
    end else if (_T_6642) begin
      ic_tag_valid_out_0_39 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_40 <= 1'h0;
    end else if (_T_6659) begin
      ic_tag_valid_out_0_40 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_41 <= 1'h0;
    end else if (_T_6676) begin
      ic_tag_valid_out_0_41 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_42 <= 1'h0;
    end else if (_T_6693) begin
      ic_tag_valid_out_0_42 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_43 <= 1'h0;
    end else if (_T_6710) begin
      ic_tag_valid_out_0_43 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_44 <= 1'h0;
    end else if (_T_6727) begin
      ic_tag_valid_out_0_44 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_45 <= 1'h0;
    end else if (_T_6744) begin
      ic_tag_valid_out_0_45 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_46 <= 1'h0;
    end else if (_T_6761) begin
      ic_tag_valid_out_0_46 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_47 <= 1'h0;
    end else if (_T_6778) begin
      ic_tag_valid_out_0_47 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_48 <= 1'h0;
    end else if (_T_6795) begin
      ic_tag_valid_out_0_48 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_49 <= 1'h0;
    end else if (_T_6812) begin
      ic_tag_valid_out_0_49 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_50 <= 1'h0;
    end else if (_T_6829) begin
      ic_tag_valid_out_0_50 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_51 <= 1'h0;
    end else if (_T_6846) begin
      ic_tag_valid_out_0_51 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_52 <= 1'h0;
    end else if (_T_6863) begin
      ic_tag_valid_out_0_52 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_53 <= 1'h0;
    end else if (_T_6880) begin
      ic_tag_valid_out_0_53 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_54 <= 1'h0;
    end else if (_T_6897) begin
      ic_tag_valid_out_0_54 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_55 <= 1'h0;
    end else if (_T_6914) begin
      ic_tag_valid_out_0_55 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_56 <= 1'h0;
    end else if (_T_6931) begin
      ic_tag_valid_out_0_56 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_57 <= 1'h0;
    end else if (_T_6948) begin
      ic_tag_valid_out_0_57 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_58 <= 1'h0;
    end else if (_T_6965) begin
      ic_tag_valid_out_0_58 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_59 <= 1'h0;
    end else if (_T_6982) begin
      ic_tag_valid_out_0_59 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_60 <= 1'h0;
    end else if (_T_6999) begin
      ic_tag_valid_out_0_60 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_61 <= 1'h0;
    end else if (_T_7016) begin
      ic_tag_valid_out_0_61 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_62 <= 1'h0;
    end else if (_T_7033) begin
      ic_tag_valid_out_0_62 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_63 <= 1'h0;
    end else if (_T_7050) begin
      ic_tag_valid_out_0_63 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_64 <= 1'h0;
    end else if (_T_7611) begin
      ic_tag_valid_out_0_64 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_65 <= 1'h0;
    end else if (_T_7628) begin
      ic_tag_valid_out_0_65 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_66 <= 1'h0;
    end else if (_T_7645) begin
      ic_tag_valid_out_0_66 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_67 <= 1'h0;
    end else if (_T_7662) begin
      ic_tag_valid_out_0_67 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_68 <= 1'h0;
    end else if (_T_7679) begin
      ic_tag_valid_out_0_68 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_69 <= 1'h0;
    end else if (_T_7696) begin
      ic_tag_valid_out_0_69 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_70 <= 1'h0;
    end else if (_T_7713) begin
      ic_tag_valid_out_0_70 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_71 <= 1'h0;
    end else if (_T_7730) begin
      ic_tag_valid_out_0_71 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_72 <= 1'h0;
    end else if (_T_7747) begin
      ic_tag_valid_out_0_72 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_73 <= 1'h0;
    end else if (_T_7764) begin
      ic_tag_valid_out_0_73 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_74 <= 1'h0;
    end else if (_T_7781) begin
      ic_tag_valid_out_0_74 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_75 <= 1'h0;
    end else if (_T_7798) begin
      ic_tag_valid_out_0_75 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_76 <= 1'h0;
    end else if (_T_7815) begin
      ic_tag_valid_out_0_76 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_77 <= 1'h0;
    end else if (_T_7832) begin
      ic_tag_valid_out_0_77 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_78 <= 1'h0;
    end else if (_T_7849) begin
      ic_tag_valid_out_0_78 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_79 <= 1'h0;
    end else if (_T_7866) begin
      ic_tag_valid_out_0_79 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_80 <= 1'h0;
    end else if (_T_7883) begin
      ic_tag_valid_out_0_80 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_81 <= 1'h0;
    end else if (_T_7900) begin
      ic_tag_valid_out_0_81 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_82 <= 1'h0;
    end else if (_T_7917) begin
      ic_tag_valid_out_0_82 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_83 <= 1'h0;
    end else if (_T_7934) begin
      ic_tag_valid_out_0_83 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_84 <= 1'h0;
    end else if (_T_7951) begin
      ic_tag_valid_out_0_84 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_85 <= 1'h0;
    end else if (_T_7968) begin
      ic_tag_valid_out_0_85 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_86 <= 1'h0;
    end else if (_T_7985) begin
      ic_tag_valid_out_0_86 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_87 <= 1'h0;
    end else if (_T_8002) begin
      ic_tag_valid_out_0_87 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_88 <= 1'h0;
    end else if (_T_8019) begin
      ic_tag_valid_out_0_88 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_89 <= 1'h0;
    end else if (_T_8036) begin
      ic_tag_valid_out_0_89 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_90 <= 1'h0;
    end else if (_T_8053) begin
      ic_tag_valid_out_0_90 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_91 <= 1'h0;
    end else if (_T_8070) begin
      ic_tag_valid_out_0_91 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_92 <= 1'h0;
    end else if (_T_8087) begin
      ic_tag_valid_out_0_92 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_93 <= 1'h0;
    end else if (_T_8104) begin
      ic_tag_valid_out_0_93 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_94 <= 1'h0;
    end else if (_T_8121) begin
      ic_tag_valid_out_0_94 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_95 <= 1'h0;
    end else if (_T_8138) begin
      ic_tag_valid_out_0_95 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_96 <= 1'h0;
    end else if (_T_8699) begin
      ic_tag_valid_out_0_96 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_97 <= 1'h0;
    end else if (_T_8716) begin
      ic_tag_valid_out_0_97 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_98 <= 1'h0;
    end else if (_T_8733) begin
      ic_tag_valid_out_0_98 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_99 <= 1'h0;
    end else if (_T_8750) begin
      ic_tag_valid_out_0_99 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_100 <= 1'h0;
    end else if (_T_8767) begin
      ic_tag_valid_out_0_100 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_101 <= 1'h0;
    end else if (_T_8784) begin
      ic_tag_valid_out_0_101 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_102 <= 1'h0;
    end else if (_T_8801) begin
      ic_tag_valid_out_0_102 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_103 <= 1'h0;
    end else if (_T_8818) begin
      ic_tag_valid_out_0_103 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_104 <= 1'h0;
    end else if (_T_8835) begin
      ic_tag_valid_out_0_104 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_105 <= 1'h0;
    end else if (_T_8852) begin
      ic_tag_valid_out_0_105 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_106 <= 1'h0;
    end else if (_T_8869) begin
      ic_tag_valid_out_0_106 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_107 <= 1'h0;
    end else if (_T_8886) begin
      ic_tag_valid_out_0_107 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_108 <= 1'h0;
    end else if (_T_8903) begin
      ic_tag_valid_out_0_108 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_109 <= 1'h0;
    end else if (_T_8920) begin
      ic_tag_valid_out_0_109 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_110 <= 1'h0;
    end else if (_T_8937) begin
      ic_tag_valid_out_0_110 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_111 <= 1'h0;
    end else if (_T_8954) begin
      ic_tag_valid_out_0_111 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_112 <= 1'h0;
    end else if (_T_8971) begin
      ic_tag_valid_out_0_112 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_113 <= 1'h0;
    end else if (_T_8988) begin
      ic_tag_valid_out_0_113 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_114 <= 1'h0;
    end else if (_T_9005) begin
      ic_tag_valid_out_0_114 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_115 <= 1'h0;
    end else if (_T_9022) begin
      ic_tag_valid_out_0_115 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_116 <= 1'h0;
    end else if (_T_9039) begin
      ic_tag_valid_out_0_116 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_117 <= 1'h0;
    end else if (_T_9056) begin
      ic_tag_valid_out_0_117 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_118 <= 1'h0;
    end else if (_T_9073) begin
      ic_tag_valid_out_0_118 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_119 <= 1'h0;
    end else if (_T_9090) begin
      ic_tag_valid_out_0_119 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_120 <= 1'h0;
    end else if (_T_9107) begin
      ic_tag_valid_out_0_120 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_121 <= 1'h0;
    end else if (_T_9124) begin
      ic_tag_valid_out_0_121 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_122 <= 1'h0;
    end else if (_T_9141) begin
      ic_tag_valid_out_0_122 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_123 <= 1'h0;
    end else if (_T_9158) begin
      ic_tag_valid_out_0_123 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_124 <= 1'h0;
    end else if (_T_9175) begin
      ic_tag_valid_out_0_124 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_125 <= 1'h0;
    end else if (_T_9192) begin
      ic_tag_valid_out_0_125 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_126 <= 1'h0;
    end else if (_T_9209) begin
      ic_tag_valid_out_0_126 <= _T_5425;
    end
    if (reset) begin
      ic_tag_valid_out_0_127 <= 1'h0;
    end else if (_T_9226) begin
      ic_tag_valid_out_0_127 <= _T_5425;
    end
    if (reset) begin
      ic_debug_way_ff <= 2'h0;
    end else if (debug_c1_clken) begin
      ic_debug_way_ff <= io_ic_debug_way;
    end
    if (reset) begin
      _T_1209 <= 71'h0;
    end else if (ic_debug_rd_en_ff) begin
      if (ic_debug_ict_array_sel_ff) begin
        _T_1209 <= {{5'd0}, _T_1208};
      end else begin
        _T_1209 <= io_ic_debug_rd_data;
      end
    end
    if (reset) begin
      ifu_bus_cmd_valid <= 1'h0;
    end else if (_T_2564) begin
      ifu_bus_cmd_valid <= ifc_bus_ic_req_ff_in;
    end
    if (reset) begin
      bus_cmd_beat_count <= 3'h0;
    end else if (_T_2639) begin
      bus_cmd_beat_count <= bus_new_cmd_beat_count;
    end
    if (reset) begin
      ifu_bus_arready_unq_ff <= 1'h0;
    end else if (io_ifu_bus_clk_en) begin
      ifu_bus_arready_unq_ff <= io_ifu_axi_arready;
    end
    if (reset) begin
      ifu_bus_arvalid_ff <= 1'h0;
    end else if (io_ifu_bus_clk_en) begin
      ifu_bus_arvalid_ff <= io_ifu_axi_arvalid;
    end
  end
  always @(posedge io_free_clk) begin
    if (reset) begin
      scnd_miss_req_q <= 1'h0;
    end else begin
      scnd_miss_req_q <= scnd_miss_req_in;
    end
    if (reset) begin
      iccm_dma_rvalid_in <= 1'h0;
    end else begin
      iccm_dma_rvalid_in <= _T_2683;
    end
    if (reset) begin
      dma_iccm_req_f <= 1'h0;
    end else begin
      dma_iccm_req_f <= io_dma_iccm_req;
    end
    if (reset) begin
      perr_state <= 3'h0;
    end else if (perr_state_en) begin
      if (_T_2465) begin
        if (io_iccm_dma_sb_error) begin
          perr_state <= 3'h4;
        end else if (_T_2467) begin
          perr_state <= 3'h1;
        end else begin
          perr_state <= 3'h2;
        end
      end else if (_T_2477) begin
        perr_state <= 3'h0;
      end else if (_T_2480) begin
        if (_T_2482) begin
          perr_state <= 3'h0;
        end else begin
          perr_state <= 3'h3;
        end
      end else if (_T_2486) begin
        if (io_dec_tlu_force_halt) begin
          perr_state <= 3'h0;
        end else begin
          perr_state <= 3'h3;
        end
      end else begin
        perr_state <= 3'h0;
      end
    end
    if (reset) begin
      err_stop_state <= 2'h0;
    end else if (err_stop_state_en) begin
      if (_T_2490) begin
        err_stop_state <= 2'h1;
      end else if (_T_2495) begin
        if (_T_2497) begin
          err_stop_state <= 2'h0;
        end else if (_T_2518) begin
          err_stop_state <= 2'h3;
        end else if (io_ifu_fetch_val[0]) begin
          err_stop_state <= 2'h2;
        end else begin
          err_stop_state <= 2'h1;
        end
      end else if (_T_2522) begin
        if (_T_2497) begin
          err_stop_state <= 2'h0;
        end else if (io_ifu_fetch_val[0]) begin
          err_stop_state <= 2'h3;
        end else begin
          err_stop_state <= 2'h2;
        end
      end else if (_T_2539) begin
        if (_T_2543) begin
          err_stop_state <= 2'h0;
        end else if (io_dec_tlu_flush_err_wb) begin
          err_stop_state <= 2'h1;
        end else begin
          err_stop_state <= 2'h3;
        end
      end else begin
        err_stop_state <= 2'h0;
      end
    end
    if (reset) begin
      bus_ifu_bus_clk_en_ff <= 1'h0;
    end else begin
      bus_ifu_bus_clk_en_ff <= io_ifu_bus_clk_en;
    end
    if (reset) begin
      bus_data_beat_count <= 3'h0;
    end else begin
      bus_data_beat_count <= bus_new_data_beat_count;
    end
    if (reset) begin
      ic_miss_buff_data_valid <= 8'h0;
    end else begin
      ic_miss_buff_data_valid <= _T_1368;
    end
    if (reset) begin
      last_data_recieved_ff <= 1'h0;
    end else begin
      last_data_recieved_ff <= last_data_recieved_in;
    end
    if (reset) begin
      sel_mb_addr_ff <= 1'h0;
    end else begin
      sel_mb_addr_ff <= sel_mb_addr;
    end
    if (reset) begin
      ifu_ic_rw_int_addr_ff <= 7'h0;
    end else if (_T_4148) begin
      ifu_ic_rw_int_addr_ff <= io_ic_debug_addr[9:3];
    end else begin
      ifu_ic_rw_int_addr_ff <= ifu_ic_rw_int_addr[11:5];
    end
    if (reset) begin
      ifu_wr_data_comb_err_ff <= 1'h0;
    end else begin
      ifu_wr_data_comb_err_ff <= ifu_wr_cumulative_err;
    end
    if (reset) begin
      ic_act_miss_f_delayed <= 1'h0;
    end else begin
      ic_act_miss_f_delayed <= ic_act_miss_f;
    end
    if (reset) begin
      ic_crit_wd_rdy_new_ff <= 1'h0;
    end else begin
      ic_crit_wd_rdy_new_ff <= ic_crit_wd_rdy_new_in;
    end
    if (reset) begin
      ic_miss_buff_data_error <= 8'h0;
    end else begin
      ic_miss_buff_data_error <= _T_1408;
    end
    if (reset) begin
      ic_debug_rd_en_ff <= 1'h0;
    end else begin
      ic_debug_rd_en_ff <= io_ic_debug_rd_en;
    end
    if (reset) begin
      ifc_dma_access_ok_prev <= 1'h0;
    end else begin
      ifc_dma_access_ok_prev <= ifc_dma_access_ok_d;
    end
    if (reset) begin
      iccm_ecc_corr_data_ff <= 39'h0;
    end else if (iccm_ecc_write_status) begin
      iccm_ecc_corr_data_ff <= _T_4083;
    end
    if (reset) begin
      dma_mem_addr_ff <= 2'h0;
    end else begin
      dma_mem_addr_ff <= io_dma_mem_addr[3:2];
    end
    if (reset) begin
      dma_mem_tag_ff <= 3'h0;
    end else begin
      dma_mem_tag_ff <= io_dma_mem_tag;
    end
    if (reset) begin
      iccm_dma_rtag_temp <= 3'h0;
    end else begin
      iccm_dma_rtag_temp <= dma_mem_tag_ff;
    end
    if (reset) begin
      iccm_dma_rvalid_temp <= 1'h0;
    end else begin
      iccm_dma_rvalid_temp <= iccm_dma_rvalid_in;
    end
    if (reset) begin
      iccm_dma_rdata_temp <= 64'h0;
    end else if (iccm_dma_ecc_error_in) begin
      iccm_dma_rdata_temp <= _T_3257;
    end else begin
      iccm_dma_rdata_temp <= _T_3258;
    end
    if (reset) begin
      iccm_ecc_corr_index_ff <= 14'h0;
    end else if (iccm_ecc_write_status) begin
      if (iccm_single_ecc_error[0]) begin
        iccm_ecc_corr_index_ff <= iccm_rw_addr_f;
      end else begin
        iccm_ecc_corr_index_ff <= _T_4079;
      end
    end
    if (reset) begin
      iccm_rd_ecc_single_err_ff <= 1'h0;
    end else begin
      iccm_rd_ecc_single_err_ff <= iccm_rd_ecc_single_err_hold_in;
    end
    if (reset) begin
      iccm_rw_addr_f <= 14'h0;
    end else begin
      iccm_rw_addr_f <= io_iccm_rw_addr[14:1];
    end
    if (reset) begin
      ifu_status_wr_addr_ff <= 7'h0;
    end else if (_T_4148) begin
      ifu_status_wr_addr_ff <= io_ic_debug_addr[9:3];
    end else begin
      ifu_status_wr_addr_ff <= ifu_status_wr_addr[11:5];
    end
    if (reset) begin
      way_status_wr_en_ff <= 1'h0;
    end else begin
      way_status_wr_en_ff <= way_status_wr_en_w_debug;
    end
    if (reset) begin
      way_status_new_ff <= 1'h0;
    end else if (_T_4151) begin
      way_status_new_ff <= io_ic_debug_wr_data[4];
    end else if (_T_10560) begin
      way_status_new_ff <= replace_way_mb_any_0;
    end else begin
      way_status_new_ff <= way_status_hit_new;
    end
    if (reset) begin
      ifu_tag_wren_ff <= 2'h0;
    end else begin
      ifu_tag_wren_ff <= ifu_tag_wren_w_debug;
    end
    if (reset) begin
      ic_valid_ff <= 1'h0;
    end else if (_T_4151) begin
      ic_valid_ff <= io_ic_debug_wr_data[0];
    end else begin
      ic_valid_ff <= ic_valid;
    end
    if (reset) begin
      _T_10612 <= 1'h0;
    end else if (ic_debug_rd_en_ff) begin
      _T_10612 <= ic_debug_rd_en_ff;
    end
  end
  always @(posedge io_active_clk) begin
    if (reset) begin
      reset_all_tags <= 1'h0;
    end else begin
      reset_all_tags <= io_dec_tlu_fence_i_wb;
    end
    if (reset) begin
      perr_ic_index_ff <= 7'h0;
    end else if (perr_sb_write_status) begin
      perr_ic_index_ff <= ifu_ic_rw_int_addr_ff;
    end
    if (reset) begin
      dma_sb_err_state_ff <= 1'h0;
    end else begin
      dma_sb_err_state_ff <= _T_7;
    end
    if (reset) begin
      _T_10582 <= 1'h0;
    end else begin
      _T_10582 <= ic_act_miss_f;
    end
    if (reset) begin
      _T_10583 <= 1'h0;
    end else begin
      _T_10583 <= ic_act_hit_f;
    end
    if (reset) begin
      _T_10584 <= 1'h0;
    end else begin
      _T_10584 <= ifc_bus_acc_fault_f;
    end
    if (reset) begin
      _T_10588 <= 1'h0;
    end else begin
      _T_10588 <= _T_10587;
    end
    if (reset) begin
      _T_10589 <= 1'h0;
    end else begin
      _T_10589 <= bus_cmd_sent;
    end
  end
endmodule
