module lsu_trigger(
  input         clock,
  input         reset,
  input         io_trigger_pkt_any_0_select,
  input         io_trigger_pkt_any_0_match_pkt,
  input         io_trigger_pkt_any_0_store,
  input         io_trigger_pkt_any_0_load,
  input         io_trigger_pkt_any_0_execute,
  input         io_trigger_pkt_any_0_m,
  input  [31:0] io_trigger_pkt_any_0_tdata2,
  input         io_trigger_pkt_any_1_select,
  input         io_trigger_pkt_any_1_match_pkt,
  input         io_trigger_pkt_any_1_store,
  input         io_trigger_pkt_any_1_load,
  input         io_trigger_pkt_any_1_execute,
  input         io_trigger_pkt_any_1_m,
  input  [31:0] io_trigger_pkt_any_1_tdata2,
  input         io_trigger_pkt_any_2_select,
  input         io_trigger_pkt_any_2_match_pkt,
  input         io_trigger_pkt_any_2_store,
  input         io_trigger_pkt_any_2_load,
  input         io_trigger_pkt_any_2_execute,
  input         io_trigger_pkt_any_2_m,
  input  [31:0] io_trigger_pkt_any_2_tdata2,
  input         io_trigger_pkt_any_3_select,
  input         io_trigger_pkt_any_3_match_pkt,
  input         io_trigger_pkt_any_3_store,
  input         io_trigger_pkt_any_3_load,
  input         io_trigger_pkt_any_3_execute,
  input         io_trigger_pkt_any_3_m,
  input  [31:0] io_trigger_pkt_any_3_tdata2,
  input         io_lsu_pkt_m_valid,
  input         io_lsu_pkt_m_bits_fast_int,
  input         io_lsu_pkt_m_bits_by,
  input         io_lsu_pkt_m_bits_half,
  input         io_lsu_pkt_m_bits_word,
  input         io_lsu_pkt_m_bits_dword,
  input         io_lsu_pkt_m_bits_load,
  input         io_lsu_pkt_m_bits_store,
  input         io_lsu_pkt_m_bits_unsign,
  input         io_lsu_pkt_m_bits_dma,
  input         io_lsu_pkt_m_bits_store_data_bypass_d,
  input         io_lsu_pkt_m_bits_load_ldst_bypass_d,
  input         io_lsu_pkt_m_bits_store_data_bypass_m,
  input  [31:0] io_lsu_addr_m,
  input  [31:0] io_store_data_m,
  output [3:0]  io_lsu_trigger_match_m
);
  wire  _T = io_trigger_pkt_any_0_m | io_trigger_pkt_any_1_m; // @[lsu_trigger.scala 16:73]
  wire  _T_1 = _T | io_trigger_pkt_any_2_m; // @[lsu_trigger.scala 16:73]
  wire  trigger_enable = _T_1 | io_trigger_pkt_any_3_m; // @[lsu_trigger.scala 16:73]
  wire [15:0] _T_4 = io_lsu_pkt_m_bits_word ? 16'hffff : 16'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _T_6 = _T_4 & io_store_data_m[31:16]; // @[lsu_trigger.scala 17:66]
  wire  _T_7 = io_lsu_pkt_m_bits_half | io_lsu_pkt_m_bits_word; // @[lsu_trigger.scala 17:124]
  wire [7:0] _T_9 = _T_7 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_11 = _T_9 & io_store_data_m[15:8]; // @[lsu_trigger.scala 17:151]
  wire [31:0] store_data_trigger_m = {_T_6,_T_11,io_store_data_m[7:0]}; // @[Cat.scala 29:58]
  wire [31:0] _T_15 = trigger_enable ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] ldst_addr_trigger_m = io_lsu_addr_m & _T_15; // @[lsu_trigger.scala 18:43]
  wire  _T_17 = ~io_trigger_pkt_any_0_select; // @[lsu_trigger.scala 19:53]
  wire  _T_18 = io_trigger_pkt_any_0_select & io_trigger_pkt_any_0_store; // @[lsu_trigger.scala 19:143]
  wire [31:0] _T_20 = _T_17 ? ldst_addr_trigger_m : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_21 = _T_18 ? store_data_trigger_m : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] lsu_match_data_0 = _T_20 | _T_21; // @[Mux.scala 27:72]
  wire  _T_24 = ~io_trigger_pkt_any_1_select; // @[lsu_trigger.scala 19:53]
  wire  _T_25 = io_trigger_pkt_any_1_select & io_trigger_pkt_any_1_store; // @[lsu_trigger.scala 19:143]
  wire [31:0] _T_27 = _T_24 ? ldst_addr_trigger_m : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_28 = _T_25 ? store_data_trigger_m : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] lsu_match_data_1 = _T_27 | _T_28; // @[Mux.scala 27:72]
  wire  _T_31 = ~io_trigger_pkt_any_2_select; // @[lsu_trigger.scala 19:53]
  wire  _T_32 = io_trigger_pkt_any_2_select & io_trigger_pkt_any_2_store; // @[lsu_trigger.scala 19:143]
  wire [31:0] _T_34 = _T_31 ? ldst_addr_trigger_m : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_35 = _T_32 ? store_data_trigger_m : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] lsu_match_data_2 = _T_34 | _T_35; // @[Mux.scala 27:72]
  wire  _T_38 = ~io_trigger_pkt_any_3_select; // @[lsu_trigger.scala 19:53]
  wire  _T_39 = io_trigger_pkt_any_3_select & io_trigger_pkt_any_3_store; // @[lsu_trigger.scala 19:143]
  wire [31:0] _T_41 = _T_38 ? ldst_addr_trigger_m : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_42 = _T_39 ? store_data_trigger_m : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] lsu_match_data_3 = _T_41 | _T_42; // @[Mux.scala 27:72]
  wire  _T_44 = ~io_lsu_pkt_m_bits_dma; // @[lsu_trigger.scala 20:70]
  wire  _T_45 = io_lsu_pkt_m_valid & _T_44; // @[lsu_trigger.scala 20:68]
  wire  _T_46 = _T_45 & trigger_enable; // @[lsu_trigger.scala 20:93]
  wire  _T_47 = io_trigger_pkt_any_0_store & io_lsu_pkt_m_bits_store; // @[lsu_trigger.scala 20:142]
  wire  _T_48 = io_trigger_pkt_any_0_load & io_lsu_pkt_m_bits_load; // @[lsu_trigger.scala 21:33]
  wire  _T_50 = _T_48 & _T_17; // @[lsu_trigger.scala 21:58]
  wire  _T_51 = _T_47 | _T_50; // @[lsu_trigger.scala 20:168]
  wire  _T_52 = _T_46 & _T_51; // @[lsu_trigger.scala 20:110]
  wire  _T_55 = &io_trigger_pkt_any_0_tdata2; // @[lib.scala 101:45]
  wire  _T_56 = ~_T_55; // @[lib.scala 101:39]
  wire  _T_57 = io_trigger_pkt_any_0_match_pkt & _T_56; // @[lib.scala 101:37]
  wire  _T_60 = io_trigger_pkt_any_0_tdata2[0] == lsu_match_data_0[0]; // @[lib.scala 102:52]
  wire  _T_61 = _T_57 | _T_60; // @[lib.scala 102:41]
  wire  _T_63 = &io_trigger_pkt_any_0_tdata2[0]; // @[lib.scala 104:36]
  wire  _T_64 = _T_63 & _T_57; // @[lib.scala 104:41]
  wire  _T_67 = io_trigger_pkt_any_0_tdata2[1] == lsu_match_data_0[1]; // @[lib.scala 104:78]
  wire  _T_68 = _T_64 | _T_67; // @[lib.scala 104:23]
  wire  _T_70 = &io_trigger_pkt_any_0_tdata2[1:0]; // @[lib.scala 104:36]
  wire  _T_71 = _T_70 & _T_57; // @[lib.scala 104:41]
  wire  _T_74 = io_trigger_pkt_any_0_tdata2[2] == lsu_match_data_0[2]; // @[lib.scala 104:78]
  wire  _T_75 = _T_71 | _T_74; // @[lib.scala 104:23]
  wire  _T_77 = &io_trigger_pkt_any_0_tdata2[2:0]; // @[lib.scala 104:36]
  wire  _T_78 = _T_77 & _T_57; // @[lib.scala 104:41]
  wire  _T_81 = io_trigger_pkt_any_0_tdata2[3] == lsu_match_data_0[3]; // @[lib.scala 104:78]
  wire  _T_82 = _T_78 | _T_81; // @[lib.scala 104:23]
  wire  _T_84 = &io_trigger_pkt_any_0_tdata2[3:0]; // @[lib.scala 104:36]
  wire  _T_85 = _T_84 & _T_57; // @[lib.scala 104:41]
  wire  _T_88 = io_trigger_pkt_any_0_tdata2[4] == lsu_match_data_0[4]; // @[lib.scala 104:78]
  wire  _T_89 = _T_85 | _T_88; // @[lib.scala 104:23]
  wire  _T_91 = &io_trigger_pkt_any_0_tdata2[4:0]; // @[lib.scala 104:36]
  wire  _T_92 = _T_91 & _T_57; // @[lib.scala 104:41]
  wire  _T_95 = io_trigger_pkt_any_0_tdata2[5] == lsu_match_data_0[5]; // @[lib.scala 104:78]
  wire  _T_96 = _T_92 | _T_95; // @[lib.scala 104:23]
  wire  _T_98 = &io_trigger_pkt_any_0_tdata2[5:0]; // @[lib.scala 104:36]
  wire  _T_99 = _T_98 & _T_57; // @[lib.scala 104:41]
  wire  _T_102 = io_trigger_pkt_any_0_tdata2[6] == lsu_match_data_0[6]; // @[lib.scala 104:78]
  wire  _T_103 = _T_99 | _T_102; // @[lib.scala 104:23]
  wire  _T_105 = &io_trigger_pkt_any_0_tdata2[6:0]; // @[lib.scala 104:36]
  wire  _T_106 = _T_105 & _T_57; // @[lib.scala 104:41]
  wire  _T_109 = io_trigger_pkt_any_0_tdata2[7] == lsu_match_data_0[7]; // @[lib.scala 104:78]
  wire  _T_110 = _T_106 | _T_109; // @[lib.scala 104:23]
  wire  _T_112 = &io_trigger_pkt_any_0_tdata2[7:0]; // @[lib.scala 104:36]
  wire  _T_113 = _T_112 & _T_57; // @[lib.scala 104:41]
  wire  _T_116 = io_trigger_pkt_any_0_tdata2[8] == lsu_match_data_0[8]; // @[lib.scala 104:78]
  wire  _T_117 = _T_113 | _T_116; // @[lib.scala 104:23]
  wire  _T_119 = &io_trigger_pkt_any_0_tdata2[8:0]; // @[lib.scala 104:36]
  wire  _T_120 = _T_119 & _T_57; // @[lib.scala 104:41]
  wire  _T_123 = io_trigger_pkt_any_0_tdata2[9] == lsu_match_data_0[9]; // @[lib.scala 104:78]
  wire  _T_124 = _T_120 | _T_123; // @[lib.scala 104:23]
  wire  _T_126 = &io_trigger_pkt_any_0_tdata2[9:0]; // @[lib.scala 104:36]
  wire  _T_127 = _T_126 & _T_57; // @[lib.scala 104:41]
  wire  _T_130 = io_trigger_pkt_any_0_tdata2[10] == lsu_match_data_0[10]; // @[lib.scala 104:78]
  wire  _T_131 = _T_127 | _T_130; // @[lib.scala 104:23]
  wire  _T_133 = &io_trigger_pkt_any_0_tdata2[10:0]; // @[lib.scala 104:36]
  wire  _T_134 = _T_133 & _T_57; // @[lib.scala 104:41]
  wire  _T_137 = io_trigger_pkt_any_0_tdata2[11] == lsu_match_data_0[11]; // @[lib.scala 104:78]
  wire  _T_138 = _T_134 | _T_137; // @[lib.scala 104:23]
  wire  _T_140 = &io_trigger_pkt_any_0_tdata2[11:0]; // @[lib.scala 104:36]
  wire  _T_141 = _T_140 & _T_57; // @[lib.scala 104:41]
  wire  _T_144 = io_trigger_pkt_any_0_tdata2[12] == lsu_match_data_0[12]; // @[lib.scala 104:78]
  wire  _T_145 = _T_141 | _T_144; // @[lib.scala 104:23]
  wire  _T_147 = &io_trigger_pkt_any_0_tdata2[12:0]; // @[lib.scala 104:36]
  wire  _T_148 = _T_147 & _T_57; // @[lib.scala 104:41]
  wire  _T_151 = io_trigger_pkt_any_0_tdata2[13] == lsu_match_data_0[13]; // @[lib.scala 104:78]
  wire  _T_152 = _T_148 | _T_151; // @[lib.scala 104:23]
  wire  _T_154 = &io_trigger_pkt_any_0_tdata2[13:0]; // @[lib.scala 104:36]
  wire  _T_155 = _T_154 & _T_57; // @[lib.scala 104:41]
  wire  _T_158 = io_trigger_pkt_any_0_tdata2[14] == lsu_match_data_0[14]; // @[lib.scala 104:78]
  wire  _T_159 = _T_155 | _T_158; // @[lib.scala 104:23]
  wire  _T_161 = &io_trigger_pkt_any_0_tdata2[14:0]; // @[lib.scala 104:36]
  wire  _T_162 = _T_161 & _T_57; // @[lib.scala 104:41]
  wire  _T_165 = io_trigger_pkt_any_0_tdata2[15] == lsu_match_data_0[15]; // @[lib.scala 104:78]
  wire  _T_166 = _T_162 | _T_165; // @[lib.scala 104:23]
  wire  _T_168 = &io_trigger_pkt_any_0_tdata2[15:0]; // @[lib.scala 104:36]
  wire  _T_169 = _T_168 & _T_57; // @[lib.scala 104:41]
  wire  _T_172 = io_trigger_pkt_any_0_tdata2[16] == lsu_match_data_0[16]; // @[lib.scala 104:78]
  wire  _T_173 = _T_169 | _T_172; // @[lib.scala 104:23]
  wire  _T_175 = &io_trigger_pkt_any_0_tdata2[16:0]; // @[lib.scala 104:36]
  wire  _T_176 = _T_175 & _T_57; // @[lib.scala 104:41]
  wire  _T_179 = io_trigger_pkt_any_0_tdata2[17] == lsu_match_data_0[17]; // @[lib.scala 104:78]
  wire  _T_180 = _T_176 | _T_179; // @[lib.scala 104:23]
  wire  _T_182 = &io_trigger_pkt_any_0_tdata2[17:0]; // @[lib.scala 104:36]
  wire  _T_183 = _T_182 & _T_57; // @[lib.scala 104:41]
  wire  _T_186 = io_trigger_pkt_any_0_tdata2[18] == lsu_match_data_0[18]; // @[lib.scala 104:78]
  wire  _T_187 = _T_183 | _T_186; // @[lib.scala 104:23]
  wire  _T_189 = &io_trigger_pkt_any_0_tdata2[18:0]; // @[lib.scala 104:36]
  wire  _T_190 = _T_189 & _T_57; // @[lib.scala 104:41]
  wire  _T_193 = io_trigger_pkt_any_0_tdata2[19] == lsu_match_data_0[19]; // @[lib.scala 104:78]
  wire  _T_194 = _T_190 | _T_193; // @[lib.scala 104:23]
  wire  _T_196 = &io_trigger_pkt_any_0_tdata2[19:0]; // @[lib.scala 104:36]
  wire  _T_197 = _T_196 & _T_57; // @[lib.scala 104:41]
  wire  _T_200 = io_trigger_pkt_any_0_tdata2[20] == lsu_match_data_0[20]; // @[lib.scala 104:78]
  wire  _T_201 = _T_197 | _T_200; // @[lib.scala 104:23]
  wire  _T_203 = &io_trigger_pkt_any_0_tdata2[20:0]; // @[lib.scala 104:36]
  wire  _T_204 = _T_203 & _T_57; // @[lib.scala 104:41]
  wire  _T_207 = io_trigger_pkt_any_0_tdata2[21] == lsu_match_data_0[21]; // @[lib.scala 104:78]
  wire  _T_208 = _T_204 | _T_207; // @[lib.scala 104:23]
  wire  _T_210 = &io_trigger_pkt_any_0_tdata2[21:0]; // @[lib.scala 104:36]
  wire  _T_211 = _T_210 & _T_57; // @[lib.scala 104:41]
  wire  _T_214 = io_trigger_pkt_any_0_tdata2[22] == lsu_match_data_0[22]; // @[lib.scala 104:78]
  wire  _T_215 = _T_211 | _T_214; // @[lib.scala 104:23]
  wire  _T_217 = &io_trigger_pkt_any_0_tdata2[22:0]; // @[lib.scala 104:36]
  wire  _T_218 = _T_217 & _T_57; // @[lib.scala 104:41]
  wire  _T_221 = io_trigger_pkt_any_0_tdata2[23] == lsu_match_data_0[23]; // @[lib.scala 104:78]
  wire  _T_222 = _T_218 | _T_221; // @[lib.scala 104:23]
  wire  _T_224 = &io_trigger_pkt_any_0_tdata2[23:0]; // @[lib.scala 104:36]
  wire  _T_225 = _T_224 & _T_57; // @[lib.scala 104:41]
  wire  _T_228 = io_trigger_pkt_any_0_tdata2[24] == lsu_match_data_0[24]; // @[lib.scala 104:78]
  wire  _T_229 = _T_225 | _T_228; // @[lib.scala 104:23]
  wire  _T_231 = &io_trigger_pkt_any_0_tdata2[24:0]; // @[lib.scala 104:36]
  wire  _T_232 = _T_231 & _T_57; // @[lib.scala 104:41]
  wire  _T_235 = io_trigger_pkt_any_0_tdata2[25] == lsu_match_data_0[25]; // @[lib.scala 104:78]
  wire  _T_236 = _T_232 | _T_235; // @[lib.scala 104:23]
  wire  _T_238 = &io_trigger_pkt_any_0_tdata2[25:0]; // @[lib.scala 104:36]
  wire  _T_239 = _T_238 & _T_57; // @[lib.scala 104:41]
  wire  _T_242 = io_trigger_pkt_any_0_tdata2[26] == lsu_match_data_0[26]; // @[lib.scala 104:78]
  wire  _T_243 = _T_239 | _T_242; // @[lib.scala 104:23]
  wire  _T_245 = &io_trigger_pkt_any_0_tdata2[26:0]; // @[lib.scala 104:36]
  wire  _T_246 = _T_245 & _T_57; // @[lib.scala 104:41]
  wire  _T_249 = io_trigger_pkt_any_0_tdata2[27] == lsu_match_data_0[27]; // @[lib.scala 104:78]
  wire  _T_250 = _T_246 | _T_249; // @[lib.scala 104:23]
  wire  _T_252 = &io_trigger_pkt_any_0_tdata2[27:0]; // @[lib.scala 104:36]
  wire  _T_253 = _T_252 & _T_57; // @[lib.scala 104:41]
  wire  _T_256 = io_trigger_pkt_any_0_tdata2[28] == lsu_match_data_0[28]; // @[lib.scala 104:78]
  wire  _T_257 = _T_253 | _T_256; // @[lib.scala 104:23]
  wire  _T_259 = &io_trigger_pkt_any_0_tdata2[28:0]; // @[lib.scala 104:36]
  wire  _T_260 = _T_259 & _T_57; // @[lib.scala 104:41]
  wire  _T_263 = io_trigger_pkt_any_0_tdata2[29] == lsu_match_data_0[29]; // @[lib.scala 104:78]
  wire  _T_264 = _T_260 | _T_263; // @[lib.scala 104:23]
  wire  _T_266 = &io_trigger_pkt_any_0_tdata2[29:0]; // @[lib.scala 104:36]
  wire  _T_267 = _T_266 & _T_57; // @[lib.scala 104:41]
  wire  _T_270 = io_trigger_pkt_any_0_tdata2[30] == lsu_match_data_0[30]; // @[lib.scala 104:78]
  wire  _T_271 = _T_267 | _T_270; // @[lib.scala 104:23]
  wire  _T_273 = &io_trigger_pkt_any_0_tdata2[30:0]; // @[lib.scala 104:36]
  wire  _T_274 = _T_273 & _T_57; // @[lib.scala 104:41]
  wire  _T_277 = io_trigger_pkt_any_0_tdata2[31] == lsu_match_data_0[31]; // @[lib.scala 104:78]
  wire  _T_278 = _T_274 | _T_277; // @[lib.scala 104:23]
  wire [7:0] _T_285 = {_T_110,_T_103,_T_96,_T_89,_T_82,_T_75,_T_68,_T_61}; // @[lib.scala 105:14]
  wire [15:0] _T_293 = {_T_166,_T_159,_T_152,_T_145,_T_138,_T_131,_T_124,_T_117,_T_285}; // @[lib.scala 105:14]
  wire [7:0] _T_300 = {_T_222,_T_215,_T_208,_T_201,_T_194,_T_187,_T_180,_T_173}; // @[lib.scala 105:14]
  wire [31:0] _T_309 = {_T_278,_T_271,_T_264,_T_257,_T_250,_T_243,_T_236,_T_229,_T_300,_T_293}; // @[lib.scala 105:14]
  wire  _T_310 = &_T_309; // @[lib.scala 105:25]
  wire  _T_311 = _T_52 & _T_310; // @[lsu_trigger.scala 21:92]
  wire  _T_315 = io_trigger_pkt_any_1_store & io_lsu_pkt_m_bits_store; // @[lsu_trigger.scala 20:142]
  wire  _T_316 = io_trigger_pkt_any_1_load & io_lsu_pkt_m_bits_load; // @[lsu_trigger.scala 21:33]
  wire  _T_318 = _T_316 & _T_24; // @[lsu_trigger.scala 21:58]
  wire  _T_319 = _T_315 | _T_318; // @[lsu_trigger.scala 20:168]
  wire  _T_320 = _T_46 & _T_319; // @[lsu_trigger.scala 20:110]
  wire  _T_323 = &io_trigger_pkt_any_1_tdata2; // @[lib.scala 101:45]
  wire  _T_324 = ~_T_323; // @[lib.scala 101:39]
  wire  _T_325 = io_trigger_pkt_any_1_match_pkt & _T_324; // @[lib.scala 101:37]
  wire  _T_328 = io_trigger_pkt_any_1_tdata2[0] == lsu_match_data_1[0]; // @[lib.scala 102:52]
  wire  _T_329 = _T_325 | _T_328; // @[lib.scala 102:41]
  wire  _T_331 = &io_trigger_pkt_any_1_tdata2[0]; // @[lib.scala 104:36]
  wire  _T_332 = _T_331 & _T_325; // @[lib.scala 104:41]
  wire  _T_335 = io_trigger_pkt_any_1_tdata2[1] == lsu_match_data_1[1]; // @[lib.scala 104:78]
  wire  _T_336 = _T_332 | _T_335; // @[lib.scala 104:23]
  wire  _T_338 = &io_trigger_pkt_any_1_tdata2[1:0]; // @[lib.scala 104:36]
  wire  _T_339 = _T_338 & _T_325; // @[lib.scala 104:41]
  wire  _T_342 = io_trigger_pkt_any_1_tdata2[2] == lsu_match_data_1[2]; // @[lib.scala 104:78]
  wire  _T_343 = _T_339 | _T_342; // @[lib.scala 104:23]
  wire  _T_345 = &io_trigger_pkt_any_1_tdata2[2:0]; // @[lib.scala 104:36]
  wire  _T_346 = _T_345 & _T_325; // @[lib.scala 104:41]
  wire  _T_349 = io_trigger_pkt_any_1_tdata2[3] == lsu_match_data_1[3]; // @[lib.scala 104:78]
  wire  _T_350 = _T_346 | _T_349; // @[lib.scala 104:23]
  wire  _T_352 = &io_trigger_pkt_any_1_tdata2[3:0]; // @[lib.scala 104:36]
  wire  _T_353 = _T_352 & _T_325; // @[lib.scala 104:41]
  wire  _T_356 = io_trigger_pkt_any_1_tdata2[4] == lsu_match_data_1[4]; // @[lib.scala 104:78]
  wire  _T_357 = _T_353 | _T_356; // @[lib.scala 104:23]
  wire  _T_359 = &io_trigger_pkt_any_1_tdata2[4:0]; // @[lib.scala 104:36]
  wire  _T_360 = _T_359 & _T_325; // @[lib.scala 104:41]
  wire  _T_363 = io_trigger_pkt_any_1_tdata2[5] == lsu_match_data_1[5]; // @[lib.scala 104:78]
  wire  _T_364 = _T_360 | _T_363; // @[lib.scala 104:23]
  wire  _T_366 = &io_trigger_pkt_any_1_tdata2[5:0]; // @[lib.scala 104:36]
  wire  _T_367 = _T_366 & _T_325; // @[lib.scala 104:41]
  wire  _T_370 = io_trigger_pkt_any_1_tdata2[6] == lsu_match_data_1[6]; // @[lib.scala 104:78]
  wire  _T_371 = _T_367 | _T_370; // @[lib.scala 104:23]
  wire  _T_373 = &io_trigger_pkt_any_1_tdata2[6:0]; // @[lib.scala 104:36]
  wire  _T_374 = _T_373 & _T_325; // @[lib.scala 104:41]
  wire  _T_377 = io_trigger_pkt_any_1_tdata2[7] == lsu_match_data_1[7]; // @[lib.scala 104:78]
  wire  _T_378 = _T_374 | _T_377; // @[lib.scala 104:23]
  wire  _T_380 = &io_trigger_pkt_any_1_tdata2[7:0]; // @[lib.scala 104:36]
  wire  _T_381 = _T_380 & _T_325; // @[lib.scala 104:41]
  wire  _T_384 = io_trigger_pkt_any_1_tdata2[8] == lsu_match_data_1[8]; // @[lib.scala 104:78]
  wire  _T_385 = _T_381 | _T_384; // @[lib.scala 104:23]
  wire  _T_387 = &io_trigger_pkt_any_1_tdata2[8:0]; // @[lib.scala 104:36]
  wire  _T_388 = _T_387 & _T_325; // @[lib.scala 104:41]
  wire  _T_391 = io_trigger_pkt_any_1_tdata2[9] == lsu_match_data_1[9]; // @[lib.scala 104:78]
  wire  _T_392 = _T_388 | _T_391; // @[lib.scala 104:23]
  wire  _T_394 = &io_trigger_pkt_any_1_tdata2[9:0]; // @[lib.scala 104:36]
  wire  _T_395 = _T_394 & _T_325; // @[lib.scala 104:41]
  wire  _T_398 = io_trigger_pkt_any_1_tdata2[10] == lsu_match_data_1[10]; // @[lib.scala 104:78]
  wire  _T_399 = _T_395 | _T_398; // @[lib.scala 104:23]
  wire  _T_401 = &io_trigger_pkt_any_1_tdata2[10:0]; // @[lib.scala 104:36]
  wire  _T_402 = _T_401 & _T_325; // @[lib.scala 104:41]
  wire  _T_405 = io_trigger_pkt_any_1_tdata2[11] == lsu_match_data_1[11]; // @[lib.scala 104:78]
  wire  _T_406 = _T_402 | _T_405; // @[lib.scala 104:23]
  wire  _T_408 = &io_trigger_pkt_any_1_tdata2[11:0]; // @[lib.scala 104:36]
  wire  _T_409 = _T_408 & _T_325; // @[lib.scala 104:41]
  wire  _T_412 = io_trigger_pkt_any_1_tdata2[12] == lsu_match_data_1[12]; // @[lib.scala 104:78]
  wire  _T_413 = _T_409 | _T_412; // @[lib.scala 104:23]
  wire  _T_415 = &io_trigger_pkt_any_1_tdata2[12:0]; // @[lib.scala 104:36]
  wire  _T_416 = _T_415 & _T_325; // @[lib.scala 104:41]
  wire  _T_419 = io_trigger_pkt_any_1_tdata2[13] == lsu_match_data_1[13]; // @[lib.scala 104:78]
  wire  _T_420 = _T_416 | _T_419; // @[lib.scala 104:23]
  wire  _T_422 = &io_trigger_pkt_any_1_tdata2[13:0]; // @[lib.scala 104:36]
  wire  _T_423 = _T_422 & _T_325; // @[lib.scala 104:41]
  wire  _T_426 = io_trigger_pkt_any_1_tdata2[14] == lsu_match_data_1[14]; // @[lib.scala 104:78]
  wire  _T_427 = _T_423 | _T_426; // @[lib.scala 104:23]
  wire  _T_429 = &io_trigger_pkt_any_1_tdata2[14:0]; // @[lib.scala 104:36]
  wire  _T_430 = _T_429 & _T_325; // @[lib.scala 104:41]
  wire  _T_433 = io_trigger_pkt_any_1_tdata2[15] == lsu_match_data_1[15]; // @[lib.scala 104:78]
  wire  _T_434 = _T_430 | _T_433; // @[lib.scala 104:23]
  wire  _T_436 = &io_trigger_pkt_any_1_tdata2[15:0]; // @[lib.scala 104:36]
  wire  _T_437 = _T_436 & _T_325; // @[lib.scala 104:41]
  wire  _T_440 = io_trigger_pkt_any_1_tdata2[16] == lsu_match_data_1[16]; // @[lib.scala 104:78]
  wire  _T_441 = _T_437 | _T_440; // @[lib.scala 104:23]
  wire  _T_443 = &io_trigger_pkt_any_1_tdata2[16:0]; // @[lib.scala 104:36]
  wire  _T_444 = _T_443 & _T_325; // @[lib.scala 104:41]
  wire  _T_447 = io_trigger_pkt_any_1_tdata2[17] == lsu_match_data_1[17]; // @[lib.scala 104:78]
  wire  _T_448 = _T_444 | _T_447; // @[lib.scala 104:23]
  wire  _T_450 = &io_trigger_pkt_any_1_tdata2[17:0]; // @[lib.scala 104:36]
  wire  _T_451 = _T_450 & _T_325; // @[lib.scala 104:41]
  wire  _T_454 = io_trigger_pkt_any_1_tdata2[18] == lsu_match_data_1[18]; // @[lib.scala 104:78]
  wire  _T_455 = _T_451 | _T_454; // @[lib.scala 104:23]
  wire  _T_457 = &io_trigger_pkt_any_1_tdata2[18:0]; // @[lib.scala 104:36]
  wire  _T_458 = _T_457 & _T_325; // @[lib.scala 104:41]
  wire  _T_461 = io_trigger_pkt_any_1_tdata2[19] == lsu_match_data_1[19]; // @[lib.scala 104:78]
  wire  _T_462 = _T_458 | _T_461; // @[lib.scala 104:23]
  wire  _T_464 = &io_trigger_pkt_any_1_tdata2[19:0]; // @[lib.scala 104:36]
  wire  _T_465 = _T_464 & _T_325; // @[lib.scala 104:41]
  wire  _T_468 = io_trigger_pkt_any_1_tdata2[20] == lsu_match_data_1[20]; // @[lib.scala 104:78]
  wire  _T_469 = _T_465 | _T_468; // @[lib.scala 104:23]
  wire  _T_471 = &io_trigger_pkt_any_1_tdata2[20:0]; // @[lib.scala 104:36]
  wire  _T_472 = _T_471 & _T_325; // @[lib.scala 104:41]
  wire  _T_475 = io_trigger_pkt_any_1_tdata2[21] == lsu_match_data_1[21]; // @[lib.scala 104:78]
  wire  _T_476 = _T_472 | _T_475; // @[lib.scala 104:23]
  wire  _T_478 = &io_trigger_pkt_any_1_tdata2[21:0]; // @[lib.scala 104:36]
  wire  _T_479 = _T_478 & _T_325; // @[lib.scala 104:41]
  wire  _T_482 = io_trigger_pkt_any_1_tdata2[22] == lsu_match_data_1[22]; // @[lib.scala 104:78]
  wire  _T_483 = _T_479 | _T_482; // @[lib.scala 104:23]
  wire  _T_485 = &io_trigger_pkt_any_1_tdata2[22:0]; // @[lib.scala 104:36]
  wire  _T_486 = _T_485 & _T_325; // @[lib.scala 104:41]
  wire  _T_489 = io_trigger_pkt_any_1_tdata2[23] == lsu_match_data_1[23]; // @[lib.scala 104:78]
  wire  _T_490 = _T_486 | _T_489; // @[lib.scala 104:23]
  wire  _T_492 = &io_trigger_pkt_any_1_tdata2[23:0]; // @[lib.scala 104:36]
  wire  _T_493 = _T_492 & _T_325; // @[lib.scala 104:41]
  wire  _T_496 = io_trigger_pkt_any_1_tdata2[24] == lsu_match_data_1[24]; // @[lib.scala 104:78]
  wire  _T_497 = _T_493 | _T_496; // @[lib.scala 104:23]
  wire  _T_499 = &io_trigger_pkt_any_1_tdata2[24:0]; // @[lib.scala 104:36]
  wire  _T_500 = _T_499 & _T_325; // @[lib.scala 104:41]
  wire  _T_503 = io_trigger_pkt_any_1_tdata2[25] == lsu_match_data_1[25]; // @[lib.scala 104:78]
  wire  _T_504 = _T_500 | _T_503; // @[lib.scala 104:23]
  wire  _T_506 = &io_trigger_pkt_any_1_tdata2[25:0]; // @[lib.scala 104:36]
  wire  _T_507 = _T_506 & _T_325; // @[lib.scala 104:41]
  wire  _T_510 = io_trigger_pkt_any_1_tdata2[26] == lsu_match_data_1[26]; // @[lib.scala 104:78]
  wire  _T_511 = _T_507 | _T_510; // @[lib.scala 104:23]
  wire  _T_513 = &io_trigger_pkt_any_1_tdata2[26:0]; // @[lib.scala 104:36]
  wire  _T_514 = _T_513 & _T_325; // @[lib.scala 104:41]
  wire  _T_517 = io_trigger_pkt_any_1_tdata2[27] == lsu_match_data_1[27]; // @[lib.scala 104:78]
  wire  _T_518 = _T_514 | _T_517; // @[lib.scala 104:23]
  wire  _T_520 = &io_trigger_pkt_any_1_tdata2[27:0]; // @[lib.scala 104:36]
  wire  _T_521 = _T_520 & _T_325; // @[lib.scala 104:41]
  wire  _T_524 = io_trigger_pkt_any_1_tdata2[28] == lsu_match_data_1[28]; // @[lib.scala 104:78]
  wire  _T_525 = _T_521 | _T_524; // @[lib.scala 104:23]
  wire  _T_527 = &io_trigger_pkt_any_1_tdata2[28:0]; // @[lib.scala 104:36]
  wire  _T_528 = _T_527 & _T_325; // @[lib.scala 104:41]
  wire  _T_531 = io_trigger_pkt_any_1_tdata2[29] == lsu_match_data_1[29]; // @[lib.scala 104:78]
  wire  _T_532 = _T_528 | _T_531; // @[lib.scala 104:23]
  wire  _T_534 = &io_trigger_pkt_any_1_tdata2[29:0]; // @[lib.scala 104:36]
  wire  _T_535 = _T_534 & _T_325; // @[lib.scala 104:41]
  wire  _T_538 = io_trigger_pkt_any_1_tdata2[30] == lsu_match_data_1[30]; // @[lib.scala 104:78]
  wire  _T_539 = _T_535 | _T_538; // @[lib.scala 104:23]
  wire  _T_541 = &io_trigger_pkt_any_1_tdata2[30:0]; // @[lib.scala 104:36]
  wire  _T_542 = _T_541 & _T_325; // @[lib.scala 104:41]
  wire  _T_545 = io_trigger_pkt_any_1_tdata2[31] == lsu_match_data_1[31]; // @[lib.scala 104:78]
  wire  _T_546 = _T_542 | _T_545; // @[lib.scala 104:23]
  wire [7:0] _T_553 = {_T_378,_T_371,_T_364,_T_357,_T_350,_T_343,_T_336,_T_329}; // @[lib.scala 105:14]
  wire [15:0] _T_561 = {_T_434,_T_427,_T_420,_T_413,_T_406,_T_399,_T_392,_T_385,_T_553}; // @[lib.scala 105:14]
  wire [7:0] _T_568 = {_T_490,_T_483,_T_476,_T_469,_T_462,_T_455,_T_448,_T_441}; // @[lib.scala 105:14]
  wire [31:0] _T_577 = {_T_546,_T_539,_T_532,_T_525,_T_518,_T_511,_T_504,_T_497,_T_568,_T_561}; // @[lib.scala 105:14]
  wire  _T_578 = &_T_577; // @[lib.scala 105:25]
  wire  _T_579 = _T_320 & _T_578; // @[lsu_trigger.scala 21:92]
  wire  _T_583 = io_trigger_pkt_any_2_store & io_lsu_pkt_m_bits_store; // @[lsu_trigger.scala 20:142]
  wire  _T_584 = io_trigger_pkt_any_2_load & io_lsu_pkt_m_bits_load; // @[lsu_trigger.scala 21:33]
  wire  _T_586 = _T_584 & _T_31; // @[lsu_trigger.scala 21:58]
  wire  _T_587 = _T_583 | _T_586; // @[lsu_trigger.scala 20:168]
  wire  _T_588 = _T_46 & _T_587; // @[lsu_trigger.scala 20:110]
  wire  _T_591 = &io_trigger_pkt_any_2_tdata2; // @[lib.scala 101:45]
  wire  _T_592 = ~_T_591; // @[lib.scala 101:39]
  wire  _T_593 = io_trigger_pkt_any_2_match_pkt & _T_592; // @[lib.scala 101:37]
  wire  _T_596 = io_trigger_pkt_any_2_tdata2[0] == lsu_match_data_2[0]; // @[lib.scala 102:52]
  wire  _T_597 = _T_593 | _T_596; // @[lib.scala 102:41]
  wire  _T_599 = &io_trigger_pkt_any_2_tdata2[0]; // @[lib.scala 104:36]
  wire  _T_600 = _T_599 & _T_593; // @[lib.scala 104:41]
  wire  _T_603 = io_trigger_pkt_any_2_tdata2[1] == lsu_match_data_2[1]; // @[lib.scala 104:78]
  wire  _T_604 = _T_600 | _T_603; // @[lib.scala 104:23]
  wire  _T_606 = &io_trigger_pkt_any_2_tdata2[1:0]; // @[lib.scala 104:36]
  wire  _T_607 = _T_606 & _T_593; // @[lib.scala 104:41]
  wire  _T_610 = io_trigger_pkt_any_2_tdata2[2] == lsu_match_data_2[2]; // @[lib.scala 104:78]
  wire  _T_611 = _T_607 | _T_610; // @[lib.scala 104:23]
  wire  _T_613 = &io_trigger_pkt_any_2_tdata2[2:0]; // @[lib.scala 104:36]
  wire  _T_614 = _T_613 & _T_593; // @[lib.scala 104:41]
  wire  _T_617 = io_trigger_pkt_any_2_tdata2[3] == lsu_match_data_2[3]; // @[lib.scala 104:78]
  wire  _T_618 = _T_614 | _T_617; // @[lib.scala 104:23]
  wire  _T_620 = &io_trigger_pkt_any_2_tdata2[3:0]; // @[lib.scala 104:36]
  wire  _T_621 = _T_620 & _T_593; // @[lib.scala 104:41]
  wire  _T_624 = io_trigger_pkt_any_2_tdata2[4] == lsu_match_data_2[4]; // @[lib.scala 104:78]
  wire  _T_625 = _T_621 | _T_624; // @[lib.scala 104:23]
  wire  _T_627 = &io_trigger_pkt_any_2_tdata2[4:0]; // @[lib.scala 104:36]
  wire  _T_628 = _T_627 & _T_593; // @[lib.scala 104:41]
  wire  _T_631 = io_trigger_pkt_any_2_tdata2[5] == lsu_match_data_2[5]; // @[lib.scala 104:78]
  wire  _T_632 = _T_628 | _T_631; // @[lib.scala 104:23]
  wire  _T_634 = &io_trigger_pkt_any_2_tdata2[5:0]; // @[lib.scala 104:36]
  wire  _T_635 = _T_634 & _T_593; // @[lib.scala 104:41]
  wire  _T_638 = io_trigger_pkt_any_2_tdata2[6] == lsu_match_data_2[6]; // @[lib.scala 104:78]
  wire  _T_639 = _T_635 | _T_638; // @[lib.scala 104:23]
  wire  _T_641 = &io_trigger_pkt_any_2_tdata2[6:0]; // @[lib.scala 104:36]
  wire  _T_642 = _T_641 & _T_593; // @[lib.scala 104:41]
  wire  _T_645 = io_trigger_pkt_any_2_tdata2[7] == lsu_match_data_2[7]; // @[lib.scala 104:78]
  wire  _T_646 = _T_642 | _T_645; // @[lib.scala 104:23]
  wire  _T_648 = &io_trigger_pkt_any_2_tdata2[7:0]; // @[lib.scala 104:36]
  wire  _T_649 = _T_648 & _T_593; // @[lib.scala 104:41]
  wire  _T_652 = io_trigger_pkt_any_2_tdata2[8] == lsu_match_data_2[8]; // @[lib.scala 104:78]
  wire  _T_653 = _T_649 | _T_652; // @[lib.scala 104:23]
  wire  _T_655 = &io_trigger_pkt_any_2_tdata2[8:0]; // @[lib.scala 104:36]
  wire  _T_656 = _T_655 & _T_593; // @[lib.scala 104:41]
  wire  _T_659 = io_trigger_pkt_any_2_tdata2[9] == lsu_match_data_2[9]; // @[lib.scala 104:78]
  wire  _T_660 = _T_656 | _T_659; // @[lib.scala 104:23]
  wire  _T_662 = &io_trigger_pkt_any_2_tdata2[9:0]; // @[lib.scala 104:36]
  wire  _T_663 = _T_662 & _T_593; // @[lib.scala 104:41]
  wire  _T_666 = io_trigger_pkt_any_2_tdata2[10] == lsu_match_data_2[10]; // @[lib.scala 104:78]
  wire  _T_667 = _T_663 | _T_666; // @[lib.scala 104:23]
  wire  _T_669 = &io_trigger_pkt_any_2_tdata2[10:0]; // @[lib.scala 104:36]
  wire  _T_670 = _T_669 & _T_593; // @[lib.scala 104:41]
  wire  _T_673 = io_trigger_pkt_any_2_tdata2[11] == lsu_match_data_2[11]; // @[lib.scala 104:78]
  wire  _T_674 = _T_670 | _T_673; // @[lib.scala 104:23]
  wire  _T_676 = &io_trigger_pkt_any_2_tdata2[11:0]; // @[lib.scala 104:36]
  wire  _T_677 = _T_676 & _T_593; // @[lib.scala 104:41]
  wire  _T_680 = io_trigger_pkt_any_2_tdata2[12] == lsu_match_data_2[12]; // @[lib.scala 104:78]
  wire  _T_681 = _T_677 | _T_680; // @[lib.scala 104:23]
  wire  _T_683 = &io_trigger_pkt_any_2_tdata2[12:0]; // @[lib.scala 104:36]
  wire  _T_684 = _T_683 & _T_593; // @[lib.scala 104:41]
  wire  _T_687 = io_trigger_pkt_any_2_tdata2[13] == lsu_match_data_2[13]; // @[lib.scala 104:78]
  wire  _T_688 = _T_684 | _T_687; // @[lib.scala 104:23]
  wire  _T_690 = &io_trigger_pkt_any_2_tdata2[13:0]; // @[lib.scala 104:36]
  wire  _T_691 = _T_690 & _T_593; // @[lib.scala 104:41]
  wire  _T_694 = io_trigger_pkt_any_2_tdata2[14] == lsu_match_data_2[14]; // @[lib.scala 104:78]
  wire  _T_695 = _T_691 | _T_694; // @[lib.scala 104:23]
  wire  _T_697 = &io_trigger_pkt_any_2_tdata2[14:0]; // @[lib.scala 104:36]
  wire  _T_698 = _T_697 & _T_593; // @[lib.scala 104:41]
  wire  _T_701 = io_trigger_pkt_any_2_tdata2[15] == lsu_match_data_2[15]; // @[lib.scala 104:78]
  wire  _T_702 = _T_698 | _T_701; // @[lib.scala 104:23]
  wire  _T_704 = &io_trigger_pkt_any_2_tdata2[15:0]; // @[lib.scala 104:36]
  wire  _T_705 = _T_704 & _T_593; // @[lib.scala 104:41]
  wire  _T_708 = io_trigger_pkt_any_2_tdata2[16] == lsu_match_data_2[16]; // @[lib.scala 104:78]
  wire  _T_709 = _T_705 | _T_708; // @[lib.scala 104:23]
  wire  _T_711 = &io_trigger_pkt_any_2_tdata2[16:0]; // @[lib.scala 104:36]
  wire  _T_712 = _T_711 & _T_593; // @[lib.scala 104:41]
  wire  _T_715 = io_trigger_pkt_any_2_tdata2[17] == lsu_match_data_2[17]; // @[lib.scala 104:78]
  wire  _T_716 = _T_712 | _T_715; // @[lib.scala 104:23]
  wire  _T_718 = &io_trigger_pkt_any_2_tdata2[17:0]; // @[lib.scala 104:36]
  wire  _T_719 = _T_718 & _T_593; // @[lib.scala 104:41]
  wire  _T_722 = io_trigger_pkt_any_2_tdata2[18] == lsu_match_data_2[18]; // @[lib.scala 104:78]
  wire  _T_723 = _T_719 | _T_722; // @[lib.scala 104:23]
  wire  _T_725 = &io_trigger_pkt_any_2_tdata2[18:0]; // @[lib.scala 104:36]
  wire  _T_726 = _T_725 & _T_593; // @[lib.scala 104:41]
  wire  _T_729 = io_trigger_pkt_any_2_tdata2[19] == lsu_match_data_2[19]; // @[lib.scala 104:78]
  wire  _T_730 = _T_726 | _T_729; // @[lib.scala 104:23]
  wire  _T_732 = &io_trigger_pkt_any_2_tdata2[19:0]; // @[lib.scala 104:36]
  wire  _T_733 = _T_732 & _T_593; // @[lib.scala 104:41]
  wire  _T_736 = io_trigger_pkt_any_2_tdata2[20] == lsu_match_data_2[20]; // @[lib.scala 104:78]
  wire  _T_737 = _T_733 | _T_736; // @[lib.scala 104:23]
  wire  _T_739 = &io_trigger_pkt_any_2_tdata2[20:0]; // @[lib.scala 104:36]
  wire  _T_740 = _T_739 & _T_593; // @[lib.scala 104:41]
  wire  _T_743 = io_trigger_pkt_any_2_tdata2[21] == lsu_match_data_2[21]; // @[lib.scala 104:78]
  wire  _T_744 = _T_740 | _T_743; // @[lib.scala 104:23]
  wire  _T_746 = &io_trigger_pkt_any_2_tdata2[21:0]; // @[lib.scala 104:36]
  wire  _T_747 = _T_746 & _T_593; // @[lib.scala 104:41]
  wire  _T_750 = io_trigger_pkt_any_2_tdata2[22] == lsu_match_data_2[22]; // @[lib.scala 104:78]
  wire  _T_751 = _T_747 | _T_750; // @[lib.scala 104:23]
  wire  _T_753 = &io_trigger_pkt_any_2_tdata2[22:0]; // @[lib.scala 104:36]
  wire  _T_754 = _T_753 & _T_593; // @[lib.scala 104:41]
  wire  _T_757 = io_trigger_pkt_any_2_tdata2[23] == lsu_match_data_2[23]; // @[lib.scala 104:78]
  wire  _T_758 = _T_754 | _T_757; // @[lib.scala 104:23]
  wire  _T_760 = &io_trigger_pkt_any_2_tdata2[23:0]; // @[lib.scala 104:36]
  wire  _T_761 = _T_760 & _T_593; // @[lib.scala 104:41]
  wire  _T_764 = io_trigger_pkt_any_2_tdata2[24] == lsu_match_data_2[24]; // @[lib.scala 104:78]
  wire  _T_765 = _T_761 | _T_764; // @[lib.scala 104:23]
  wire  _T_767 = &io_trigger_pkt_any_2_tdata2[24:0]; // @[lib.scala 104:36]
  wire  _T_768 = _T_767 & _T_593; // @[lib.scala 104:41]
  wire  _T_771 = io_trigger_pkt_any_2_tdata2[25] == lsu_match_data_2[25]; // @[lib.scala 104:78]
  wire  _T_772 = _T_768 | _T_771; // @[lib.scala 104:23]
  wire  _T_774 = &io_trigger_pkt_any_2_tdata2[25:0]; // @[lib.scala 104:36]
  wire  _T_775 = _T_774 & _T_593; // @[lib.scala 104:41]
  wire  _T_778 = io_trigger_pkt_any_2_tdata2[26] == lsu_match_data_2[26]; // @[lib.scala 104:78]
  wire  _T_779 = _T_775 | _T_778; // @[lib.scala 104:23]
  wire  _T_781 = &io_trigger_pkt_any_2_tdata2[26:0]; // @[lib.scala 104:36]
  wire  _T_782 = _T_781 & _T_593; // @[lib.scala 104:41]
  wire  _T_785 = io_trigger_pkt_any_2_tdata2[27] == lsu_match_data_2[27]; // @[lib.scala 104:78]
  wire  _T_786 = _T_782 | _T_785; // @[lib.scala 104:23]
  wire  _T_788 = &io_trigger_pkt_any_2_tdata2[27:0]; // @[lib.scala 104:36]
  wire  _T_789 = _T_788 & _T_593; // @[lib.scala 104:41]
  wire  _T_792 = io_trigger_pkt_any_2_tdata2[28] == lsu_match_data_2[28]; // @[lib.scala 104:78]
  wire  _T_793 = _T_789 | _T_792; // @[lib.scala 104:23]
  wire  _T_795 = &io_trigger_pkt_any_2_tdata2[28:0]; // @[lib.scala 104:36]
  wire  _T_796 = _T_795 & _T_593; // @[lib.scala 104:41]
  wire  _T_799 = io_trigger_pkt_any_2_tdata2[29] == lsu_match_data_2[29]; // @[lib.scala 104:78]
  wire  _T_800 = _T_796 | _T_799; // @[lib.scala 104:23]
  wire  _T_802 = &io_trigger_pkt_any_2_tdata2[29:0]; // @[lib.scala 104:36]
  wire  _T_803 = _T_802 & _T_593; // @[lib.scala 104:41]
  wire  _T_806 = io_trigger_pkt_any_2_tdata2[30] == lsu_match_data_2[30]; // @[lib.scala 104:78]
  wire  _T_807 = _T_803 | _T_806; // @[lib.scala 104:23]
  wire  _T_809 = &io_trigger_pkt_any_2_tdata2[30:0]; // @[lib.scala 104:36]
  wire  _T_810 = _T_809 & _T_593; // @[lib.scala 104:41]
  wire  _T_813 = io_trigger_pkt_any_2_tdata2[31] == lsu_match_data_2[31]; // @[lib.scala 104:78]
  wire  _T_814 = _T_810 | _T_813; // @[lib.scala 104:23]
  wire [7:0] _T_821 = {_T_646,_T_639,_T_632,_T_625,_T_618,_T_611,_T_604,_T_597}; // @[lib.scala 105:14]
  wire [15:0] _T_829 = {_T_702,_T_695,_T_688,_T_681,_T_674,_T_667,_T_660,_T_653,_T_821}; // @[lib.scala 105:14]
  wire [7:0] _T_836 = {_T_758,_T_751,_T_744,_T_737,_T_730,_T_723,_T_716,_T_709}; // @[lib.scala 105:14]
  wire [31:0] _T_845 = {_T_814,_T_807,_T_800,_T_793,_T_786,_T_779,_T_772,_T_765,_T_836,_T_829}; // @[lib.scala 105:14]
  wire  _T_846 = &_T_845; // @[lib.scala 105:25]
  wire  _T_847 = _T_588 & _T_846; // @[lsu_trigger.scala 21:92]
  wire  _T_851 = io_trigger_pkt_any_3_store & io_lsu_pkt_m_bits_store; // @[lsu_trigger.scala 20:142]
  wire  _T_852 = io_trigger_pkt_any_3_load & io_lsu_pkt_m_bits_load; // @[lsu_trigger.scala 21:33]
  wire  _T_854 = _T_852 & _T_38; // @[lsu_trigger.scala 21:58]
  wire  _T_855 = _T_851 | _T_854; // @[lsu_trigger.scala 20:168]
  wire  _T_856 = _T_46 & _T_855; // @[lsu_trigger.scala 20:110]
  wire  _T_859 = &io_trigger_pkt_any_3_tdata2; // @[lib.scala 101:45]
  wire  _T_860 = ~_T_859; // @[lib.scala 101:39]
  wire  _T_861 = io_trigger_pkt_any_3_match_pkt & _T_860; // @[lib.scala 101:37]
  wire  _T_864 = io_trigger_pkt_any_3_tdata2[0] == lsu_match_data_3[0]; // @[lib.scala 102:52]
  wire  _T_865 = _T_861 | _T_864; // @[lib.scala 102:41]
  wire  _T_867 = &io_trigger_pkt_any_3_tdata2[0]; // @[lib.scala 104:36]
  wire  _T_868 = _T_867 & _T_861; // @[lib.scala 104:41]
  wire  _T_871 = io_trigger_pkt_any_3_tdata2[1] == lsu_match_data_3[1]; // @[lib.scala 104:78]
  wire  _T_872 = _T_868 | _T_871; // @[lib.scala 104:23]
  wire  _T_874 = &io_trigger_pkt_any_3_tdata2[1:0]; // @[lib.scala 104:36]
  wire  _T_875 = _T_874 & _T_861; // @[lib.scala 104:41]
  wire  _T_878 = io_trigger_pkt_any_3_tdata2[2] == lsu_match_data_3[2]; // @[lib.scala 104:78]
  wire  _T_879 = _T_875 | _T_878; // @[lib.scala 104:23]
  wire  _T_881 = &io_trigger_pkt_any_3_tdata2[2:0]; // @[lib.scala 104:36]
  wire  _T_882 = _T_881 & _T_861; // @[lib.scala 104:41]
  wire  _T_885 = io_trigger_pkt_any_3_tdata2[3] == lsu_match_data_3[3]; // @[lib.scala 104:78]
  wire  _T_886 = _T_882 | _T_885; // @[lib.scala 104:23]
  wire  _T_888 = &io_trigger_pkt_any_3_tdata2[3:0]; // @[lib.scala 104:36]
  wire  _T_889 = _T_888 & _T_861; // @[lib.scala 104:41]
  wire  _T_892 = io_trigger_pkt_any_3_tdata2[4] == lsu_match_data_3[4]; // @[lib.scala 104:78]
  wire  _T_893 = _T_889 | _T_892; // @[lib.scala 104:23]
  wire  _T_895 = &io_trigger_pkt_any_3_tdata2[4:0]; // @[lib.scala 104:36]
  wire  _T_896 = _T_895 & _T_861; // @[lib.scala 104:41]
  wire  _T_899 = io_trigger_pkt_any_3_tdata2[5] == lsu_match_data_3[5]; // @[lib.scala 104:78]
  wire  _T_900 = _T_896 | _T_899; // @[lib.scala 104:23]
  wire  _T_902 = &io_trigger_pkt_any_3_tdata2[5:0]; // @[lib.scala 104:36]
  wire  _T_903 = _T_902 & _T_861; // @[lib.scala 104:41]
  wire  _T_906 = io_trigger_pkt_any_3_tdata2[6] == lsu_match_data_3[6]; // @[lib.scala 104:78]
  wire  _T_907 = _T_903 | _T_906; // @[lib.scala 104:23]
  wire  _T_909 = &io_trigger_pkt_any_3_tdata2[6:0]; // @[lib.scala 104:36]
  wire  _T_910 = _T_909 & _T_861; // @[lib.scala 104:41]
  wire  _T_913 = io_trigger_pkt_any_3_tdata2[7] == lsu_match_data_3[7]; // @[lib.scala 104:78]
  wire  _T_914 = _T_910 | _T_913; // @[lib.scala 104:23]
  wire  _T_916 = &io_trigger_pkt_any_3_tdata2[7:0]; // @[lib.scala 104:36]
  wire  _T_917 = _T_916 & _T_861; // @[lib.scala 104:41]
  wire  _T_920 = io_trigger_pkt_any_3_tdata2[8] == lsu_match_data_3[8]; // @[lib.scala 104:78]
  wire  _T_921 = _T_917 | _T_920; // @[lib.scala 104:23]
  wire  _T_923 = &io_trigger_pkt_any_3_tdata2[8:0]; // @[lib.scala 104:36]
  wire  _T_924 = _T_923 & _T_861; // @[lib.scala 104:41]
  wire  _T_927 = io_trigger_pkt_any_3_tdata2[9] == lsu_match_data_3[9]; // @[lib.scala 104:78]
  wire  _T_928 = _T_924 | _T_927; // @[lib.scala 104:23]
  wire  _T_930 = &io_trigger_pkt_any_3_tdata2[9:0]; // @[lib.scala 104:36]
  wire  _T_931 = _T_930 & _T_861; // @[lib.scala 104:41]
  wire  _T_934 = io_trigger_pkt_any_3_tdata2[10] == lsu_match_data_3[10]; // @[lib.scala 104:78]
  wire  _T_935 = _T_931 | _T_934; // @[lib.scala 104:23]
  wire  _T_937 = &io_trigger_pkt_any_3_tdata2[10:0]; // @[lib.scala 104:36]
  wire  _T_938 = _T_937 & _T_861; // @[lib.scala 104:41]
  wire  _T_941 = io_trigger_pkt_any_3_tdata2[11] == lsu_match_data_3[11]; // @[lib.scala 104:78]
  wire  _T_942 = _T_938 | _T_941; // @[lib.scala 104:23]
  wire  _T_944 = &io_trigger_pkt_any_3_tdata2[11:0]; // @[lib.scala 104:36]
  wire  _T_945 = _T_944 & _T_861; // @[lib.scala 104:41]
  wire  _T_948 = io_trigger_pkt_any_3_tdata2[12] == lsu_match_data_3[12]; // @[lib.scala 104:78]
  wire  _T_949 = _T_945 | _T_948; // @[lib.scala 104:23]
  wire  _T_951 = &io_trigger_pkt_any_3_tdata2[12:0]; // @[lib.scala 104:36]
  wire  _T_952 = _T_951 & _T_861; // @[lib.scala 104:41]
  wire  _T_955 = io_trigger_pkt_any_3_tdata2[13] == lsu_match_data_3[13]; // @[lib.scala 104:78]
  wire  _T_956 = _T_952 | _T_955; // @[lib.scala 104:23]
  wire  _T_958 = &io_trigger_pkt_any_3_tdata2[13:0]; // @[lib.scala 104:36]
  wire  _T_959 = _T_958 & _T_861; // @[lib.scala 104:41]
  wire  _T_962 = io_trigger_pkt_any_3_tdata2[14] == lsu_match_data_3[14]; // @[lib.scala 104:78]
  wire  _T_963 = _T_959 | _T_962; // @[lib.scala 104:23]
  wire  _T_965 = &io_trigger_pkt_any_3_tdata2[14:0]; // @[lib.scala 104:36]
  wire  _T_966 = _T_965 & _T_861; // @[lib.scala 104:41]
  wire  _T_969 = io_trigger_pkt_any_3_tdata2[15] == lsu_match_data_3[15]; // @[lib.scala 104:78]
  wire  _T_970 = _T_966 | _T_969; // @[lib.scala 104:23]
  wire  _T_972 = &io_trigger_pkt_any_3_tdata2[15:0]; // @[lib.scala 104:36]
  wire  _T_973 = _T_972 & _T_861; // @[lib.scala 104:41]
  wire  _T_976 = io_trigger_pkt_any_3_tdata2[16] == lsu_match_data_3[16]; // @[lib.scala 104:78]
  wire  _T_977 = _T_973 | _T_976; // @[lib.scala 104:23]
  wire  _T_979 = &io_trigger_pkt_any_3_tdata2[16:0]; // @[lib.scala 104:36]
  wire  _T_980 = _T_979 & _T_861; // @[lib.scala 104:41]
  wire  _T_983 = io_trigger_pkt_any_3_tdata2[17] == lsu_match_data_3[17]; // @[lib.scala 104:78]
  wire  _T_984 = _T_980 | _T_983; // @[lib.scala 104:23]
  wire  _T_986 = &io_trigger_pkt_any_3_tdata2[17:0]; // @[lib.scala 104:36]
  wire  _T_987 = _T_986 & _T_861; // @[lib.scala 104:41]
  wire  _T_990 = io_trigger_pkt_any_3_tdata2[18] == lsu_match_data_3[18]; // @[lib.scala 104:78]
  wire  _T_991 = _T_987 | _T_990; // @[lib.scala 104:23]
  wire  _T_993 = &io_trigger_pkt_any_3_tdata2[18:0]; // @[lib.scala 104:36]
  wire  _T_994 = _T_993 & _T_861; // @[lib.scala 104:41]
  wire  _T_997 = io_trigger_pkt_any_3_tdata2[19] == lsu_match_data_3[19]; // @[lib.scala 104:78]
  wire  _T_998 = _T_994 | _T_997; // @[lib.scala 104:23]
  wire  _T_1000 = &io_trigger_pkt_any_3_tdata2[19:0]; // @[lib.scala 104:36]
  wire  _T_1001 = _T_1000 & _T_861; // @[lib.scala 104:41]
  wire  _T_1004 = io_trigger_pkt_any_3_tdata2[20] == lsu_match_data_3[20]; // @[lib.scala 104:78]
  wire  _T_1005 = _T_1001 | _T_1004; // @[lib.scala 104:23]
  wire  _T_1007 = &io_trigger_pkt_any_3_tdata2[20:0]; // @[lib.scala 104:36]
  wire  _T_1008 = _T_1007 & _T_861; // @[lib.scala 104:41]
  wire  _T_1011 = io_trigger_pkt_any_3_tdata2[21] == lsu_match_data_3[21]; // @[lib.scala 104:78]
  wire  _T_1012 = _T_1008 | _T_1011; // @[lib.scala 104:23]
  wire  _T_1014 = &io_trigger_pkt_any_3_tdata2[21:0]; // @[lib.scala 104:36]
  wire  _T_1015 = _T_1014 & _T_861; // @[lib.scala 104:41]
  wire  _T_1018 = io_trigger_pkt_any_3_tdata2[22] == lsu_match_data_3[22]; // @[lib.scala 104:78]
  wire  _T_1019 = _T_1015 | _T_1018; // @[lib.scala 104:23]
  wire  _T_1021 = &io_trigger_pkt_any_3_tdata2[22:0]; // @[lib.scala 104:36]
  wire  _T_1022 = _T_1021 & _T_861; // @[lib.scala 104:41]
  wire  _T_1025 = io_trigger_pkt_any_3_tdata2[23] == lsu_match_data_3[23]; // @[lib.scala 104:78]
  wire  _T_1026 = _T_1022 | _T_1025; // @[lib.scala 104:23]
  wire  _T_1028 = &io_trigger_pkt_any_3_tdata2[23:0]; // @[lib.scala 104:36]
  wire  _T_1029 = _T_1028 & _T_861; // @[lib.scala 104:41]
  wire  _T_1032 = io_trigger_pkt_any_3_tdata2[24] == lsu_match_data_3[24]; // @[lib.scala 104:78]
  wire  _T_1033 = _T_1029 | _T_1032; // @[lib.scala 104:23]
  wire  _T_1035 = &io_trigger_pkt_any_3_tdata2[24:0]; // @[lib.scala 104:36]
  wire  _T_1036 = _T_1035 & _T_861; // @[lib.scala 104:41]
  wire  _T_1039 = io_trigger_pkt_any_3_tdata2[25] == lsu_match_data_3[25]; // @[lib.scala 104:78]
  wire  _T_1040 = _T_1036 | _T_1039; // @[lib.scala 104:23]
  wire  _T_1042 = &io_trigger_pkt_any_3_tdata2[25:0]; // @[lib.scala 104:36]
  wire  _T_1043 = _T_1042 & _T_861; // @[lib.scala 104:41]
  wire  _T_1046 = io_trigger_pkt_any_3_tdata2[26] == lsu_match_data_3[26]; // @[lib.scala 104:78]
  wire  _T_1047 = _T_1043 | _T_1046; // @[lib.scala 104:23]
  wire  _T_1049 = &io_trigger_pkt_any_3_tdata2[26:0]; // @[lib.scala 104:36]
  wire  _T_1050 = _T_1049 & _T_861; // @[lib.scala 104:41]
  wire  _T_1053 = io_trigger_pkt_any_3_tdata2[27] == lsu_match_data_3[27]; // @[lib.scala 104:78]
  wire  _T_1054 = _T_1050 | _T_1053; // @[lib.scala 104:23]
  wire  _T_1056 = &io_trigger_pkt_any_3_tdata2[27:0]; // @[lib.scala 104:36]
  wire  _T_1057 = _T_1056 & _T_861; // @[lib.scala 104:41]
  wire  _T_1060 = io_trigger_pkt_any_3_tdata2[28] == lsu_match_data_3[28]; // @[lib.scala 104:78]
  wire  _T_1061 = _T_1057 | _T_1060; // @[lib.scala 104:23]
  wire  _T_1063 = &io_trigger_pkt_any_3_tdata2[28:0]; // @[lib.scala 104:36]
  wire  _T_1064 = _T_1063 & _T_861; // @[lib.scala 104:41]
  wire  _T_1067 = io_trigger_pkt_any_3_tdata2[29] == lsu_match_data_3[29]; // @[lib.scala 104:78]
  wire  _T_1068 = _T_1064 | _T_1067; // @[lib.scala 104:23]
  wire  _T_1070 = &io_trigger_pkt_any_3_tdata2[29:0]; // @[lib.scala 104:36]
  wire  _T_1071 = _T_1070 & _T_861; // @[lib.scala 104:41]
  wire  _T_1074 = io_trigger_pkt_any_3_tdata2[30] == lsu_match_data_3[30]; // @[lib.scala 104:78]
  wire  _T_1075 = _T_1071 | _T_1074; // @[lib.scala 104:23]
  wire  _T_1077 = &io_trigger_pkt_any_3_tdata2[30:0]; // @[lib.scala 104:36]
  wire  _T_1078 = _T_1077 & _T_861; // @[lib.scala 104:41]
  wire  _T_1081 = io_trigger_pkt_any_3_tdata2[31] == lsu_match_data_3[31]; // @[lib.scala 104:78]
  wire  _T_1082 = _T_1078 | _T_1081; // @[lib.scala 104:23]
  wire [7:0] _T_1089 = {_T_914,_T_907,_T_900,_T_893,_T_886,_T_879,_T_872,_T_865}; // @[lib.scala 105:14]
  wire [15:0] _T_1097 = {_T_970,_T_963,_T_956,_T_949,_T_942,_T_935,_T_928,_T_921,_T_1089}; // @[lib.scala 105:14]
  wire [7:0] _T_1104 = {_T_1026,_T_1019,_T_1012,_T_1005,_T_998,_T_991,_T_984,_T_977}; // @[lib.scala 105:14]
  wire [31:0] _T_1113 = {_T_1082,_T_1075,_T_1068,_T_1061,_T_1054,_T_1047,_T_1040,_T_1033,_T_1104,_T_1097}; // @[lib.scala 105:14]
  wire  _T_1114 = &_T_1113; // @[lib.scala 105:25]
  wire  _T_1115 = _T_856 & _T_1114; // @[lsu_trigger.scala 21:92]
  wire [2:0] _T_1117 = {_T_1115,_T_847,_T_579}; // @[Cat.scala 29:58]
  assign io_lsu_trigger_match_m = {_T_1117,_T_311}; // @[lsu_trigger.scala 20:25]
endmodule
