module el2_ifu_mem_ctl(
  input         clock,
  input         reset,
  input         io_free_clk,
  input         io_active_clk,
  input         io_exu_flush_final,
  input         io_dec_tlu_flush_lower_wb,
  input         io_dec_tlu_flush_err_wb,
  input         io_dec_tlu_i0_commit_cmt,
  input         io_dec_tlu_force_halt,
  input  [30:0] io_ifc_fetch_addr_bf,
  input         io_ifc_fetch_uncacheable_bf,
  input         io_ifc_fetch_req_bf,
  input         io_ifc_fetch_req_bf_raw,
  input         io_ifc_iccm_access_bf,
  input         io_ifc_region_acc_fault_bf,
  input         io_ifc_dma_access_ok,
  input         io_dec_tlu_fence_i_wb,
  input         io_ifu_bp_hit_taken_f,
  input         io_ifu_bp_inst_mask_f,
  input         io_ifu_axi_arready,
  input         io_ifu_axi_rvalid,
  input  [2:0]  io_ifu_axi_rid,
  input  [63:0] io_ifu_axi_rdata,
  input  [1:0]  io_ifu_axi_rresp,
  input         io_ifu_bus_clk_en,
  input         io_dma_iccm_req,
  input  [31:0] io_dma_mem_addr,
  input  [2:0]  io_dma_mem_sz,
  input         io_dma_mem_write,
  input  [63:0] io_dma_mem_wdata,
  input  [2:0]  io_dma_mem_tag,
  input  [63:0] io_ic_rd_data,
  input  [70:0] io_ic_debug_rd_data,
  input  [25:0] io_ictag_debug_rd_data,
  input  [1:0]  io_ic_eccerr,
  input  [1:0]  io_ic_parerr,
  input  [1:0]  io_ic_rd_hit,
  input         io_ic_tag_perr,
  input  [63:0] io_iccm_rd_data,
  input  [77:0] io_iccm_rd_data_ecc,
  input  [1:0]  io_ifu_fetch_val,
  input  [70:0] io_dec_tlu_ic_diag_pkt_icache_wrdata,
  input  [16:0] io_dec_tlu_ic_diag_pkt_icache_dicawics,
  input         io_dec_tlu_ic_diag_pkt_icache_rd_valid,
  input         io_dec_tlu_ic_diag_pkt_icache_wr_valid,
  output        io_ifu_miss_state_idle,
  output        io_ifu_ic_mb_empty,
  output        io_ic_dma_active,
  output        io_ic_write_stall,
  output        io_ifu_pmu_ic_miss,
  output        io_ifu_pmu_ic_hit,
  output        io_ifu_pmu_bus_error,
  output        io_ifu_pmu_bus_busy,
  output        io_ifu_pmu_bus_trxn,
  output        io_ifu_axi_awvalid,
  output [2:0]  io_ifu_axi_awid,
  output [31:0] io_ifu_axi_awaddr,
  output [3:0]  io_ifu_axi_awregion,
  output [7:0]  io_ifu_axi_awlen,
  output [2:0]  io_ifu_axi_awsize,
  output [1:0]  io_ifu_axi_awburst,
  output        io_ifu_axi_awlock,
  output [3:0]  io_ifu_axi_awcache,
  output [2:0]  io_ifu_axi_awprot,
  output [3:0]  io_ifu_axi_awqos,
  output        io_ifu_axi_wvalid,
  output [63:0] io_ifu_axi_wdata,
  output [7:0]  io_ifu_axi_wstrb,
  output        io_ifu_axi_wlast,
  output        io_ifu_axi_bready,
  output        io_ifu_axi_arvalid,
  output [2:0]  io_ifu_axi_arid,
  output [31:0] io_ifu_axi_araddr,
  output [3:0]  io_ifu_axi_arregion,
  output [7:0]  io_ifu_axi_arlen,
  output [2:0]  io_ifu_axi_arsize,
  output [1:0]  io_ifu_axi_arburst,
  output        io_ifu_axi_arlock,
  output [3:0]  io_ifu_axi_arcache,
  output [2:0]  io_ifu_axi_arprot,
  output [3:0]  io_ifu_axi_arqos,
  output        io_ifu_axi_rready,
  output        io_iccm_dma_ecc_error,
  output        io_iccm_dma_rvalid,
  output [63:0] io_iccm_dma_rdata,
  output [2:0]  io_iccm_dma_rtag,
  output        io_iccm_ready,
  output [30:0] io_ic_rw_addr,
  output [1:0]  io_ic_wr_en,
  output        io_ic_rd_en,
  output [70:0] io_ic_wr_data_0,
  output [70:0] io_ic_wr_data_1,
  output [70:0] io_ic_debug_wr_data,
  output [70:0] io_ifu_ic_debug_rd_data,
  output [9:0]  io_ic_debug_addr,
  output        io_ic_debug_rd_en,
  output        io_ic_debug_wr_en,
  output        io_ic_debug_tag_array,
  output [1:0]  io_ic_debug_way,
  output [1:0]  io_ic_tag_valid,
  output [14:0] io_iccm_rw_addr,
  output        io_iccm_wren,
  output        io_iccm_rden,
  output [77:0] io_iccm_wr_data,
  output [2:0]  io_iccm_wr_size,
  output        io_ic_hit_f,
  output        io_ic_access_fault_f,
  output [1:0]  io_ic_access_fault_type_f,
  output        io_iccm_rd_ecc_single_err,
  output        io_iccm_rd_ecc_double_err,
  output        io_ic_error_start,
  output        io_ifu_async_error_start,
  output        io_iccm_dma_sb_error,
  output [1:0]  io_ic_fetch_val_f,
  output [31:0] io_ic_data_f,
  output [63:0] io_ic_premux_data,
  output        io_ic_sel_premux_data,
  input         io_dec_tlu_core_ecc_disable,
  output        io_ifu_ic_debug_rd_data_valid,
  output        io_iccm_buf_correct_ecc,
  output        io_iccm_correction_state,
  input         io_scan_mode,
  output [6:0]  io_ic_miss_buff_ecc,
  output [6:0]  io_ic_wr_ecc
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [63:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [95:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [63:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [63:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
`endif // RANDOMIZE_REG_INIT
  reg  flush_final_f; // @[el2_ifu_mem_ctl.scala 185:30]
  reg  ifc_fetch_req_f_raw; // @[el2_ifu_mem_ctl.scala 321:36]
  wire  _T_317 = ~io_exu_flush_final; // @[el2_ifu_mem_ctl.scala 322:44]
  wire  ifc_fetch_req_f = ifc_fetch_req_f_raw & _T_317; // @[el2_ifu_mem_ctl.scala 322:42]
  reg [2:0] miss_state; // @[Reg.scala 27:20]
  wire  miss_pending = miss_state != 3'h0; // @[el2_ifu_mem_ctl.scala 254:30]
  reg  scnd_miss_req_q; // @[el2_ifu_mem_ctl.scala 550:52]
  wire  scnd_miss_req = scnd_miss_req_q & _T_317; // @[el2_ifu_mem_ctl.scala 552:36]
  wire  debug_c1_clken = io_ic_debug_rd_en | io_ic_debug_wr_en; // @[el2_ifu_mem_ctl.scala 187:42]
  wire [3:0] ic_fetch_val_int_f = {2'h0,io_ic_fetch_val_f}; // @[Cat.scala 29:58]
  reg [30:0] ifu_fetch_addr_int_f; // @[el2_ifu_mem_ctl.scala 309:34]
  wire [4:0] _GEN_463 = {{1'd0}, ic_fetch_val_int_f}; // @[el2_ifu_mem_ctl.scala 667:53]
  wire [4:0] ic_fetch_val_shift_right = _GEN_463 << ifu_fetch_addr_int_f[0]; // @[el2_ifu_mem_ctl.scala 667:53]
  wire [1:0] _GEN_464 = {{1'd0}, _T_317}; // @[el2_ifu_mem_ctl.scala 670:91]
  wire [1:0] _T_3083 = ic_fetch_val_shift_right[3:2] & _GEN_464; // @[el2_ifu_mem_ctl.scala 670:91]
  reg  ifc_iccm_access_f; // @[el2_ifu_mem_ctl.scala 323:31]
  wire  fetch_req_iccm_f = ifc_fetch_req_f & ifc_iccm_access_f; // @[el2_ifu_mem_ctl.scala 276:46]
  wire [1:0] _GEN_465 = {{1'd0}, fetch_req_iccm_f}; // @[el2_ifu_mem_ctl.scala 670:113]
  wire [1:0] _T_3084 = _T_3083 & _GEN_465; // @[el2_ifu_mem_ctl.scala 670:113]
  reg  iccm_dma_rvalid_in; // @[el2_ifu_mem_ctl.scala 656:59]
  wire [1:0] _GEN_466 = {{1'd0}, iccm_dma_rvalid_in}; // @[el2_ifu_mem_ctl.scala 670:130]
  wire [1:0] _T_3085 = _T_3084 | _GEN_466; // @[el2_ifu_mem_ctl.scala 670:130]
  wire  _T_3086 = ~io_dec_tlu_core_ecc_disable; // @[el2_ifu_mem_ctl.scala 670:154]
  wire [1:0] _GEN_467 = {{1'd0}, _T_3086}; // @[el2_ifu_mem_ctl.scala 670:152]
  wire [1:0] _T_3087 = _T_3085 & _GEN_467; // @[el2_ifu_mem_ctl.scala 670:152]
  wire [1:0] _T_3076 = ic_fetch_val_shift_right[1:0] & _GEN_464; // @[el2_ifu_mem_ctl.scala 670:91]
  wire [1:0] _T_3077 = _T_3076 & _GEN_465; // @[el2_ifu_mem_ctl.scala 670:113]
  wire [1:0] _T_3078 = _T_3077 | _GEN_466; // @[el2_ifu_mem_ctl.scala 670:130]
  wire [1:0] _T_3080 = _T_3078 & _GEN_467; // @[el2_ifu_mem_ctl.scala 670:152]
  wire [3:0] iccm_ecc_word_enable = {_T_3087,_T_3080}; // @[Cat.scala 29:58]
  wire  _T_3187 = ^io_iccm_rd_data_ecc[31:0]; // @[el2_lib.scala 301:30]
  wire  _T_3188 = ^io_iccm_rd_data_ecc[38:32]; // @[el2_lib.scala 301:44]
  wire  _T_3189 = _T_3187 ^ _T_3188; // @[el2_lib.scala 301:35]
  wire [5:0] _T_3197 = {io_iccm_rd_data_ecc[31],io_iccm_rd_data_ecc[30],io_iccm_rd_data_ecc[29],io_iccm_rd_data_ecc[28],io_iccm_rd_data_ecc[27],io_iccm_rd_data_ecc[26]}; // @[el2_lib.scala 301:76]
  wire  _T_3198 = ^_T_3197; // @[el2_lib.scala 301:83]
  wire  _T_3199 = io_iccm_rd_data_ecc[37] ^ _T_3198; // @[el2_lib.scala 301:71]
  wire [6:0] _T_3206 = {io_iccm_rd_data_ecc[17],io_iccm_rd_data_ecc[16],io_iccm_rd_data_ecc[15],io_iccm_rd_data_ecc[14],io_iccm_rd_data_ecc[13],io_iccm_rd_data_ecc[12],io_iccm_rd_data_ecc[11]}; // @[el2_lib.scala 301:103]
  wire [14:0] _T_3214 = {io_iccm_rd_data_ecc[25],io_iccm_rd_data_ecc[24],io_iccm_rd_data_ecc[23],io_iccm_rd_data_ecc[22],io_iccm_rd_data_ecc[21],io_iccm_rd_data_ecc[20],io_iccm_rd_data_ecc[19],io_iccm_rd_data_ecc[18],_T_3206}; // @[el2_lib.scala 301:103]
  wire  _T_3215 = ^_T_3214; // @[el2_lib.scala 301:110]
  wire  _T_3216 = io_iccm_rd_data_ecc[36] ^ _T_3215; // @[el2_lib.scala 301:98]
  wire [6:0] _T_3223 = {io_iccm_rd_data_ecc[10],io_iccm_rd_data_ecc[9],io_iccm_rd_data_ecc[8],io_iccm_rd_data_ecc[7],io_iccm_rd_data_ecc[6],io_iccm_rd_data_ecc[5],io_iccm_rd_data_ecc[4]}; // @[el2_lib.scala 301:130]
  wire [14:0] _T_3231 = {io_iccm_rd_data_ecc[25],io_iccm_rd_data_ecc[24],io_iccm_rd_data_ecc[23],io_iccm_rd_data_ecc[22],io_iccm_rd_data_ecc[21],io_iccm_rd_data_ecc[20],io_iccm_rd_data_ecc[19],io_iccm_rd_data_ecc[18],_T_3223}; // @[el2_lib.scala 301:130]
  wire  _T_3232 = ^_T_3231; // @[el2_lib.scala 301:137]
  wire  _T_3233 = io_iccm_rd_data_ecc[35] ^ _T_3232; // @[el2_lib.scala 301:125]
  wire [8:0] _T_3242 = {io_iccm_rd_data_ecc[15],io_iccm_rd_data_ecc[14],io_iccm_rd_data_ecc[10],io_iccm_rd_data_ecc[9],io_iccm_rd_data_ecc[8],io_iccm_rd_data_ecc[7],io_iccm_rd_data_ecc[3],io_iccm_rd_data_ecc[2],io_iccm_rd_data_ecc[1]}; // @[el2_lib.scala 301:157]
  wire [17:0] _T_3251 = {io_iccm_rd_data_ecc[31],io_iccm_rd_data_ecc[30],io_iccm_rd_data_ecc[29],io_iccm_rd_data_ecc[25],io_iccm_rd_data_ecc[24],io_iccm_rd_data_ecc[23],io_iccm_rd_data_ecc[22],io_iccm_rd_data_ecc[17],io_iccm_rd_data_ecc[16],_T_3242}; // @[el2_lib.scala 301:157]
  wire  _T_3252 = ^_T_3251; // @[el2_lib.scala 301:164]
  wire  _T_3253 = io_iccm_rd_data_ecc[34] ^ _T_3252; // @[el2_lib.scala 301:152]
  wire [8:0] _T_3262 = {io_iccm_rd_data_ecc[13],io_iccm_rd_data_ecc[12],io_iccm_rd_data_ecc[10],io_iccm_rd_data_ecc[9],io_iccm_rd_data_ecc[6],io_iccm_rd_data_ecc[5],io_iccm_rd_data_ecc[3],io_iccm_rd_data_ecc[2],io_iccm_rd_data_ecc[0]}; // @[el2_lib.scala 301:184]
  wire [17:0] _T_3271 = {io_iccm_rd_data_ecc[31],io_iccm_rd_data_ecc[28],io_iccm_rd_data_ecc[27],io_iccm_rd_data_ecc[25],io_iccm_rd_data_ecc[24],io_iccm_rd_data_ecc[21],io_iccm_rd_data_ecc[20],io_iccm_rd_data_ecc[17],io_iccm_rd_data_ecc[16],_T_3262}; // @[el2_lib.scala 301:184]
  wire  _T_3272 = ^_T_3271; // @[el2_lib.scala 301:191]
  wire  _T_3273 = io_iccm_rd_data_ecc[33] ^ _T_3272; // @[el2_lib.scala 301:179]
  wire [8:0] _T_3282 = {io_iccm_rd_data_ecc[13],io_iccm_rd_data_ecc[11],io_iccm_rd_data_ecc[10],io_iccm_rd_data_ecc[8],io_iccm_rd_data_ecc[6],io_iccm_rd_data_ecc[4],io_iccm_rd_data_ecc[3],io_iccm_rd_data_ecc[1],io_iccm_rd_data_ecc[0]}; // @[el2_lib.scala 301:211]
  wire [17:0] _T_3291 = {io_iccm_rd_data_ecc[30],io_iccm_rd_data_ecc[28],io_iccm_rd_data_ecc[26],io_iccm_rd_data_ecc[25],io_iccm_rd_data_ecc[23],io_iccm_rd_data_ecc[21],io_iccm_rd_data_ecc[19],io_iccm_rd_data_ecc[17],io_iccm_rd_data_ecc[15],_T_3282}; // @[el2_lib.scala 301:211]
  wire  _T_3292 = ^_T_3291; // @[el2_lib.scala 301:218]
  wire  _T_3293 = io_iccm_rd_data_ecc[32] ^ _T_3292; // @[el2_lib.scala 301:206]
  wire [6:0] _T_3299 = {_T_3189,_T_3199,_T_3216,_T_3233,_T_3253,_T_3273,_T_3293}; // @[Cat.scala 29:58]
  wire  _T_3300 = _T_3299 != 7'h0; // @[el2_lib.scala 302:44]
  wire  _T_3301 = iccm_ecc_word_enable[0] & _T_3300; // @[el2_lib.scala 302:32]
  wire  _T_3303 = _T_3301 & _T_3299[6]; // @[el2_lib.scala 302:53]
  wire  _T_3572 = ^io_iccm_rd_data_ecc[70:39]; // @[el2_lib.scala 301:30]
  wire  _T_3573 = ^io_iccm_rd_data_ecc[77:71]; // @[el2_lib.scala 301:44]
  wire  _T_3574 = _T_3572 ^ _T_3573; // @[el2_lib.scala 301:35]
  wire [5:0] _T_3582 = {io_iccm_rd_data_ecc[70],io_iccm_rd_data_ecc[69],io_iccm_rd_data_ecc[68],io_iccm_rd_data_ecc[67],io_iccm_rd_data_ecc[66],io_iccm_rd_data_ecc[65]}; // @[el2_lib.scala 301:76]
  wire  _T_3583 = ^_T_3582; // @[el2_lib.scala 301:83]
  wire  _T_3584 = io_iccm_rd_data_ecc[76] ^ _T_3583; // @[el2_lib.scala 301:71]
  wire [6:0] _T_3591 = {io_iccm_rd_data_ecc[56],io_iccm_rd_data_ecc[55],io_iccm_rd_data_ecc[54],io_iccm_rd_data_ecc[53],io_iccm_rd_data_ecc[52],io_iccm_rd_data_ecc[51],io_iccm_rd_data_ecc[50]}; // @[el2_lib.scala 301:103]
  wire [14:0] _T_3599 = {io_iccm_rd_data_ecc[64],io_iccm_rd_data_ecc[63],io_iccm_rd_data_ecc[62],io_iccm_rd_data_ecc[61],io_iccm_rd_data_ecc[60],io_iccm_rd_data_ecc[59],io_iccm_rd_data_ecc[58],io_iccm_rd_data_ecc[57],_T_3591}; // @[el2_lib.scala 301:103]
  wire  _T_3600 = ^_T_3599; // @[el2_lib.scala 301:110]
  wire  _T_3601 = io_iccm_rd_data_ecc[75] ^ _T_3600; // @[el2_lib.scala 301:98]
  wire [6:0] _T_3608 = {io_iccm_rd_data_ecc[49],io_iccm_rd_data_ecc[48],io_iccm_rd_data_ecc[47],io_iccm_rd_data_ecc[46],io_iccm_rd_data_ecc[45],io_iccm_rd_data_ecc[44],io_iccm_rd_data_ecc[43]}; // @[el2_lib.scala 301:130]
  wire [14:0] _T_3616 = {io_iccm_rd_data_ecc[64],io_iccm_rd_data_ecc[63],io_iccm_rd_data_ecc[62],io_iccm_rd_data_ecc[61],io_iccm_rd_data_ecc[60],io_iccm_rd_data_ecc[59],io_iccm_rd_data_ecc[58],io_iccm_rd_data_ecc[57],_T_3608}; // @[el2_lib.scala 301:130]
  wire  _T_3617 = ^_T_3616; // @[el2_lib.scala 301:137]
  wire  _T_3618 = io_iccm_rd_data_ecc[74] ^ _T_3617; // @[el2_lib.scala 301:125]
  wire [8:0] _T_3627 = {io_iccm_rd_data_ecc[54],io_iccm_rd_data_ecc[53],io_iccm_rd_data_ecc[49],io_iccm_rd_data_ecc[48],io_iccm_rd_data_ecc[47],io_iccm_rd_data_ecc[46],io_iccm_rd_data_ecc[42],io_iccm_rd_data_ecc[41],io_iccm_rd_data_ecc[40]}; // @[el2_lib.scala 301:157]
  wire [17:0] _T_3636 = {io_iccm_rd_data_ecc[70],io_iccm_rd_data_ecc[69],io_iccm_rd_data_ecc[68],io_iccm_rd_data_ecc[64],io_iccm_rd_data_ecc[63],io_iccm_rd_data_ecc[62],io_iccm_rd_data_ecc[61],io_iccm_rd_data_ecc[56],io_iccm_rd_data_ecc[55],_T_3627}; // @[el2_lib.scala 301:157]
  wire  _T_3637 = ^_T_3636; // @[el2_lib.scala 301:164]
  wire  _T_3638 = io_iccm_rd_data_ecc[73] ^ _T_3637; // @[el2_lib.scala 301:152]
  wire [8:0] _T_3647 = {io_iccm_rd_data_ecc[52],io_iccm_rd_data_ecc[51],io_iccm_rd_data_ecc[49],io_iccm_rd_data_ecc[48],io_iccm_rd_data_ecc[45],io_iccm_rd_data_ecc[44],io_iccm_rd_data_ecc[42],io_iccm_rd_data_ecc[41],io_iccm_rd_data_ecc[39]}; // @[el2_lib.scala 301:184]
  wire [17:0] _T_3656 = {io_iccm_rd_data_ecc[70],io_iccm_rd_data_ecc[67],io_iccm_rd_data_ecc[66],io_iccm_rd_data_ecc[64],io_iccm_rd_data_ecc[63],io_iccm_rd_data_ecc[60],io_iccm_rd_data_ecc[59],io_iccm_rd_data_ecc[56],io_iccm_rd_data_ecc[55],_T_3647}; // @[el2_lib.scala 301:184]
  wire  _T_3657 = ^_T_3656; // @[el2_lib.scala 301:191]
  wire  _T_3658 = io_iccm_rd_data_ecc[72] ^ _T_3657; // @[el2_lib.scala 301:179]
  wire [8:0] _T_3667 = {io_iccm_rd_data_ecc[52],io_iccm_rd_data_ecc[50],io_iccm_rd_data_ecc[49],io_iccm_rd_data_ecc[47],io_iccm_rd_data_ecc[45],io_iccm_rd_data_ecc[43],io_iccm_rd_data_ecc[42],io_iccm_rd_data_ecc[40],io_iccm_rd_data_ecc[39]}; // @[el2_lib.scala 301:211]
  wire [17:0] _T_3676 = {io_iccm_rd_data_ecc[69],io_iccm_rd_data_ecc[67],io_iccm_rd_data_ecc[65],io_iccm_rd_data_ecc[64],io_iccm_rd_data_ecc[62],io_iccm_rd_data_ecc[60],io_iccm_rd_data_ecc[58],io_iccm_rd_data_ecc[56],io_iccm_rd_data_ecc[54],_T_3667}; // @[el2_lib.scala 301:211]
  wire  _T_3677 = ^_T_3676; // @[el2_lib.scala 301:218]
  wire  _T_3678 = io_iccm_rd_data_ecc[71] ^ _T_3677; // @[el2_lib.scala 301:206]
  wire [6:0] _T_3684 = {_T_3574,_T_3584,_T_3601,_T_3618,_T_3638,_T_3658,_T_3678}; // @[Cat.scala 29:58]
  wire  _T_3685 = _T_3684 != 7'h0; // @[el2_lib.scala 302:44]
  wire  _T_3686 = iccm_ecc_word_enable[1] & _T_3685; // @[el2_lib.scala 302:32]
  wire  _T_3688 = _T_3686 & _T_3684[6]; // @[el2_lib.scala 302:53]
  wire [1:0] iccm_single_ecc_error = {_T_3303,_T_3688}; // @[Cat.scala 29:58]
  wire  _T_3 = |iccm_single_ecc_error; // @[el2_ifu_mem_ctl.scala 190:52]
  reg  dma_iccm_req_f; // @[el2_ifu_mem_ctl.scala 634:51]
  wire  _T_6 = io_iccm_rd_ecc_single_err | io_ic_error_start; // @[el2_ifu_mem_ctl.scala 191:57]
  reg [2:0] perr_state; // @[Reg.scala 27:20]
  wire  _T_7 = perr_state == 3'h4; // @[el2_ifu_mem_ctl.scala 192:54]
  wire  iccm_correct_ecc = perr_state == 3'h3; // @[el2_ifu_mem_ctl.scala 479:34]
  wire  _T_8 = iccm_correct_ecc | _T_7; // @[el2_ifu_mem_ctl.scala 192:40]
  reg [1:0] err_stop_state; // @[Reg.scala 27:20]
  wire  _T_9 = err_stop_state == 2'h3; // @[el2_ifu_mem_ctl.scala 192:90]
  wire  _T_10 = _T_8 | _T_9; // @[el2_ifu_mem_ctl.scala 192:72]
  wire  _T_2452 = 2'h0 == err_stop_state; // @[Conditional.scala 37:30]
  wire  _T_2457 = 2'h1 == err_stop_state; // @[Conditional.scala 37:30]
  wire  _T_2477 = io_ifu_fetch_val == 2'h3; // @[el2_ifu_mem_ctl.scala 529:48]
  wire  two_byte_instr = io_ic_data_f[1:0] != 2'h3; // @[el2_ifu_mem_ctl.scala 395:42]
  wire  _T_2479 = io_ifu_fetch_val[0] & two_byte_instr; // @[el2_ifu_mem_ctl.scala 529:79]
  wire  _T_2480 = _T_2477 | _T_2479; // @[el2_ifu_mem_ctl.scala 529:56]
  wire  _T_2481 = io_exu_flush_final | io_dec_tlu_i0_commit_cmt; // @[el2_ifu_mem_ctl.scala 529:122]
  wire  _T_2482 = ~_T_2481; // @[el2_ifu_mem_ctl.scala 529:101]
  wire  _T_2483 = _T_2480 & _T_2482; // @[el2_ifu_mem_ctl.scala 529:99]
  wire  _T_2484 = 2'h2 == err_stop_state; // @[Conditional.scala 37:30]
  wire  _T_2498 = io_ifu_fetch_val[0] & _T_317; // @[el2_ifu_mem_ctl.scala 536:45]
  wire  _T_2499 = ~io_dec_tlu_i0_commit_cmt; // @[el2_ifu_mem_ctl.scala 536:69]
  wire  _T_2500 = _T_2498 & _T_2499; // @[el2_ifu_mem_ctl.scala 536:67]
  wire  _T_2501 = 2'h3 == err_stop_state; // @[Conditional.scala 37:30]
  wire  _GEN_54 = _T_2484 ? _T_2500 : _T_2501; // @[Conditional.scala 39:67]
  wire  _GEN_58 = _T_2457 ? _T_2483 : _GEN_54; // @[Conditional.scala 39:67]
  wire  err_stop_fetch = _T_2452 ? 1'h0 : _GEN_58; // @[Conditional.scala 40:58]
  wire  _T_11 = _T_10 | err_stop_fetch; // @[el2_ifu_mem_ctl.scala 192:112]
  wire  _T_13 = io_ifu_axi_rvalid & io_ifu_bus_clk_en; // @[el2_ifu_mem_ctl.scala 194:44]
  wire  _T_14 = _T_13 & io_ifu_axi_rready; // @[el2_ifu_mem_ctl.scala 194:65]
  wire  _T_227 = |io_ic_rd_hit; // @[el2_ifu_mem_ctl.scala 284:37]
  wire  _T_228 = ~_T_227; // @[el2_ifu_mem_ctl.scala 284:23]
  reg  reset_all_tags; // @[el2_ifu_mem_ctl.scala 702:53]
  wire  _T_229 = _T_228 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 284:41]
  wire  _T_207 = ~ifc_iccm_access_f; // @[el2_ifu_mem_ctl.scala 275:48]
  wire  _T_208 = ifc_fetch_req_f & _T_207; // @[el2_ifu_mem_ctl.scala 275:46]
  reg  ifc_region_acc_fault_final_f; // @[el2_ifu_mem_ctl.scala 325:42]
  wire  _T_209 = ~ifc_region_acc_fault_final_f; // @[el2_ifu_mem_ctl.scala 275:69]
  wire  fetch_req_icache_f = _T_208 & _T_209; // @[el2_ifu_mem_ctl.scala 275:67]
  wire  _T_230 = _T_229 & fetch_req_icache_f; // @[el2_ifu_mem_ctl.scala 284:59]
  wire  _T_231 = ~miss_pending; // @[el2_ifu_mem_ctl.scala 284:82]
  wire  _T_232 = _T_230 & _T_231; // @[el2_ifu_mem_ctl.scala 284:80]
  wire  _T_233 = _T_232 | scnd_miss_req; // @[el2_ifu_mem_ctl.scala 284:97]
  wire  ic_act_miss_f = _T_233 & _T_209; // @[el2_ifu_mem_ctl.scala 284:114]
  reg  ifu_bus_rvalid_unq_ff; // @[Reg.scala 27:20]
  reg  bus_ifu_bus_clk_en_ff; // @[el2_ifu_mem_ctl.scala 549:61]
  wire  ifu_bus_rvalid_ff = ifu_bus_rvalid_unq_ff & bus_ifu_bus_clk_en_ff; // @[el2_ifu_mem_ctl.scala 591:49]
  wire  bus_ifu_wr_en_ff = ifu_bus_rvalid_ff & miss_pending; // @[el2_ifu_mem_ctl.scala 618:41]
  reg  uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 311:33]
  reg [2:0] bus_data_beat_count; // @[el2_ifu_mem_ctl.scala 599:56]
  wire  _T_2603 = bus_data_beat_count == 3'h1; // @[el2_ifu_mem_ctl.scala 616:69]
  wire  _T_2604 = &bus_data_beat_count; // @[el2_ifu_mem_ctl.scala 616:101]
  wire  bus_last_data_beat = uncacheable_miss_ff ? _T_2603 : _T_2604; // @[el2_ifu_mem_ctl.scala 616:28]
  wire  _T_2550 = bus_ifu_wr_en_ff & bus_last_data_beat; // @[el2_ifu_mem_ctl.scala 595:68]
  wire  _T_2551 = ic_act_miss_f | _T_2550; // @[el2_ifu_mem_ctl.scala 595:48]
  wire  bus_reset_data_beat_cnt = _T_2551 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 595:91]
  wire  _T_2547 = ~bus_last_data_beat; // @[el2_ifu_mem_ctl.scala 594:50]
  wire  _T_2548 = bus_ifu_wr_en_ff & _T_2547; // @[el2_ifu_mem_ctl.scala 594:48]
  wire  _T_2549 = ~io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 594:72]
  wire  bus_inc_data_beat_cnt = _T_2548 & _T_2549; // @[el2_ifu_mem_ctl.scala 594:70]
  wire [2:0] _T_2555 = bus_data_beat_count + 3'h1; // @[el2_ifu_mem_ctl.scala 598:115]
  wire [2:0] _T_2557 = bus_inc_data_beat_cnt ? _T_2555 : 3'h0; // @[Mux.scala 27:72]
  wire  _T_2552 = ~bus_inc_data_beat_cnt; // @[el2_ifu_mem_ctl.scala 596:32]
  wire  _T_2553 = ~bus_reset_data_beat_cnt; // @[el2_ifu_mem_ctl.scala 596:57]
  wire  bus_hold_data_beat_cnt = _T_2552 & _T_2553; // @[el2_ifu_mem_ctl.scala 596:55]
  wire [2:0] _T_2558 = bus_hold_data_beat_cnt ? bus_data_beat_count : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] bus_new_data_beat_count = _T_2557 | _T_2558; // @[Mux.scala 27:72]
  wire  _T_15 = &bus_new_data_beat_count; // @[el2_ifu_mem_ctl.scala 194:112]
  wire  _T_16 = _T_14 & _T_15; // @[el2_ifu_mem_ctl.scala 194:85]
  wire  _T_17 = ~uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 195:5]
  wire  _T_18 = _T_16 & _T_17; // @[el2_ifu_mem_ctl.scala 194:118]
  wire  _T_19 = miss_state == 3'h5; // @[el2_ifu_mem_ctl.scala 195:41]
  wire  _T_24 = 3'h0 == miss_state; // @[Conditional.scala 37:30]
  wire  _T_26 = ic_act_miss_f & _T_317; // @[el2_ifu_mem_ctl.scala 201:43]
  wire [2:0] _T_28 = _T_26 ? 3'h1 : 3'h2; // @[el2_ifu_mem_ctl.scala 201:27]
  wire  _T_31 = 3'h1 == miss_state; // @[Conditional.scala 37:30]
  wire [4:0] byp_fetch_index = ifu_fetch_addr_int_f[4:0]; // @[el2_ifu_mem_ctl.scala 431:45]
  wire  _T_2122 = byp_fetch_index[4:2] == 3'h0; // @[el2_ifu_mem_ctl.scala 452:127]
  reg [7:0] ic_miss_buff_data_valid; // @[el2_ifu_mem_ctl.scala 408:60]
  wire  _T_2153 = _T_2122 & ic_miss_buff_data_valid[0]; // @[Mux.scala 27:72]
  wire  _T_2126 = byp_fetch_index[4:2] == 3'h1; // @[el2_ifu_mem_ctl.scala 452:127]
  wire  _T_2154 = _T_2126 & ic_miss_buff_data_valid[1]; // @[Mux.scala 27:72]
  wire  _T_2161 = _T_2153 | _T_2154; // @[Mux.scala 27:72]
  wire  _T_2130 = byp_fetch_index[4:2] == 3'h2; // @[el2_ifu_mem_ctl.scala 452:127]
  wire  _T_2155 = _T_2130 & ic_miss_buff_data_valid[2]; // @[Mux.scala 27:72]
  wire  _T_2162 = _T_2161 | _T_2155; // @[Mux.scala 27:72]
  wire  _T_2134 = byp_fetch_index[4:2] == 3'h3; // @[el2_ifu_mem_ctl.scala 452:127]
  wire  _T_2156 = _T_2134 & ic_miss_buff_data_valid[3]; // @[Mux.scala 27:72]
  wire  _T_2163 = _T_2162 | _T_2156; // @[Mux.scala 27:72]
  wire  _T_2138 = byp_fetch_index[4:2] == 3'h4; // @[el2_ifu_mem_ctl.scala 452:127]
  wire  _T_2157 = _T_2138 & ic_miss_buff_data_valid[4]; // @[Mux.scala 27:72]
  wire  _T_2164 = _T_2163 | _T_2157; // @[Mux.scala 27:72]
  wire  _T_2142 = byp_fetch_index[4:2] == 3'h5; // @[el2_ifu_mem_ctl.scala 452:127]
  wire  _T_2158 = _T_2142 & ic_miss_buff_data_valid[5]; // @[Mux.scala 27:72]
  wire  _T_2165 = _T_2164 | _T_2158; // @[Mux.scala 27:72]
  wire  _T_2146 = byp_fetch_index[4:2] == 3'h6; // @[el2_ifu_mem_ctl.scala 452:127]
  wire  _T_2159 = _T_2146 & ic_miss_buff_data_valid[6]; // @[Mux.scala 27:72]
  wire  _T_2166 = _T_2165 | _T_2159; // @[Mux.scala 27:72]
  wire  _T_2150 = byp_fetch_index[4:2] == 3'h7; // @[el2_ifu_mem_ctl.scala 452:127]
  wire  _T_2160 = _T_2150 & ic_miss_buff_data_valid[7]; // @[Mux.scala 27:72]
  wire  ic_miss_buff_data_valid_bypass_index = _T_2166 | _T_2160; // @[Mux.scala 27:72]
  wire  _T_2208 = ~byp_fetch_index[1]; // @[el2_ifu_mem_ctl.scala 454:69]
  wire  _T_2209 = ic_miss_buff_data_valid_bypass_index & _T_2208; // @[el2_ifu_mem_ctl.scala 454:67]
  wire  _T_2211 = ~byp_fetch_index[0]; // @[el2_ifu_mem_ctl.scala 454:91]
  wire  _T_2212 = _T_2209 & _T_2211; // @[el2_ifu_mem_ctl.scala 454:89]
  wire  _T_2217 = _T_2209 & byp_fetch_index[0]; // @[el2_ifu_mem_ctl.scala 455:65]
  wire  _T_2218 = _T_2212 | _T_2217; // @[el2_ifu_mem_ctl.scala 454:112]
  wire  _T_2220 = ic_miss_buff_data_valid_bypass_index & byp_fetch_index[1]; // @[el2_ifu_mem_ctl.scala 456:43]
  wire  _T_2223 = _T_2220 & _T_2211; // @[el2_ifu_mem_ctl.scala 456:65]
  wire  _T_2224 = _T_2218 | _T_2223; // @[el2_ifu_mem_ctl.scala 455:88]
  wire  _T_2228 = _T_2220 & byp_fetch_index[0]; // @[el2_ifu_mem_ctl.scala 457:65]
  wire [2:0] byp_fetch_index_inc = ifu_fetch_addr_int_f[4:2] + 3'h1; // @[el2_ifu_mem_ctl.scala 434:75]
  wire  _T_2168 = byp_fetch_index_inc == 3'h0; // @[el2_ifu_mem_ctl.scala 453:110]
  wire  _T_2192 = _T_2168 & ic_miss_buff_data_valid[0]; // @[Mux.scala 27:72]
  wire  _T_2171 = byp_fetch_index_inc == 3'h1; // @[el2_ifu_mem_ctl.scala 453:110]
  wire  _T_2193 = _T_2171 & ic_miss_buff_data_valid[1]; // @[Mux.scala 27:72]
  wire  _T_2200 = _T_2192 | _T_2193; // @[Mux.scala 27:72]
  wire  _T_2174 = byp_fetch_index_inc == 3'h2; // @[el2_ifu_mem_ctl.scala 453:110]
  wire  _T_2194 = _T_2174 & ic_miss_buff_data_valid[2]; // @[Mux.scala 27:72]
  wire  _T_2201 = _T_2200 | _T_2194; // @[Mux.scala 27:72]
  wire  _T_2177 = byp_fetch_index_inc == 3'h3; // @[el2_ifu_mem_ctl.scala 453:110]
  wire  _T_2195 = _T_2177 & ic_miss_buff_data_valid[3]; // @[Mux.scala 27:72]
  wire  _T_2202 = _T_2201 | _T_2195; // @[Mux.scala 27:72]
  wire  _T_2180 = byp_fetch_index_inc == 3'h4; // @[el2_ifu_mem_ctl.scala 453:110]
  wire  _T_2196 = _T_2180 & ic_miss_buff_data_valid[4]; // @[Mux.scala 27:72]
  wire  _T_2203 = _T_2202 | _T_2196; // @[Mux.scala 27:72]
  wire  _T_2183 = byp_fetch_index_inc == 3'h5; // @[el2_ifu_mem_ctl.scala 453:110]
  wire  _T_2197 = _T_2183 & ic_miss_buff_data_valid[5]; // @[Mux.scala 27:72]
  wire  _T_2204 = _T_2203 | _T_2197; // @[Mux.scala 27:72]
  wire  _T_2186 = byp_fetch_index_inc == 3'h6; // @[el2_ifu_mem_ctl.scala 453:110]
  wire  _T_2198 = _T_2186 & ic_miss_buff_data_valid[6]; // @[Mux.scala 27:72]
  wire  _T_2205 = _T_2204 | _T_2198; // @[Mux.scala 27:72]
  wire  _T_2189 = byp_fetch_index_inc == 3'h7; // @[el2_ifu_mem_ctl.scala 453:110]
  wire  _T_2199 = _T_2189 & ic_miss_buff_data_valid[7]; // @[Mux.scala 27:72]
  wire  ic_miss_buff_data_valid_inc_bypass_index = _T_2205 | _T_2199; // @[Mux.scala 27:72]
  wire  _T_2229 = _T_2228 & ic_miss_buff_data_valid_inc_bypass_index; // @[el2_ifu_mem_ctl.scala 457:87]
  wire  _T_2230 = _T_2224 | _T_2229; // @[el2_ifu_mem_ctl.scala 456:88]
  wire  _T_2234 = ic_miss_buff_data_valid_bypass_index & _T_2150; // @[el2_ifu_mem_ctl.scala 458:43]
  wire  miss_buff_hit_unq_f = _T_2230 | _T_2234; // @[el2_ifu_mem_ctl.scala 457:131]
  wire  _T_2250 = miss_state == 3'h4; // @[el2_ifu_mem_ctl.scala 463:55]
  wire  _T_2251 = miss_state == 3'h1; // @[el2_ifu_mem_ctl.scala 463:87]
  wire  _T_2252 = _T_2250 | _T_2251; // @[el2_ifu_mem_ctl.scala 463:74]
  wire  crit_byp_hit_f = miss_buff_hit_unq_f & _T_2252; // @[el2_ifu_mem_ctl.scala 463:41]
  wire  _T_2235 = miss_state == 3'h6; // @[el2_ifu_mem_ctl.scala 460:30]
  reg [30:0] imb_ff; // @[el2_ifu_mem_ctl.scala 312:20]
  wire  miss_wrap_f = imb_ff[5] != ifu_fetch_addr_int_f[6]; // @[el2_ifu_mem_ctl.scala 451:51]
  wire  _T_2236 = ~miss_wrap_f; // @[el2_ifu_mem_ctl.scala 460:68]
  wire  _T_2237 = miss_buff_hit_unq_f & _T_2236; // @[el2_ifu_mem_ctl.scala 460:66]
  wire  stream_hit_f = _T_2235 & _T_2237; // @[el2_ifu_mem_ctl.scala 460:43]
  wire  _T_215 = crit_byp_hit_f | stream_hit_f; // @[el2_ifu_mem_ctl.scala 279:35]
  wire  _T_216 = _T_215 & fetch_req_icache_f; // @[el2_ifu_mem_ctl.scala 279:52]
  wire  ic_byp_hit_f = _T_216 & miss_pending; // @[el2_ifu_mem_ctl.scala 279:73]
  reg  last_data_recieved_ff; // @[el2_ifu_mem_ctl.scala 601:58]
  wire  last_beat = bus_last_data_beat & bus_ifu_wr_en_ff; // @[el2_ifu_mem_ctl.scala 628:35]
  wire  _T_32 = bus_ifu_wr_en_ff & last_beat; // @[el2_ifu_mem_ctl.scala 205:113]
  wire  _T_33 = last_data_recieved_ff | _T_32; // @[el2_ifu_mem_ctl.scala 205:93]
  wire  _T_34 = ic_byp_hit_f & _T_33; // @[el2_ifu_mem_ctl.scala 205:67]
  wire  _T_35 = _T_34 & uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 205:127]
  wire  _T_36 = io_dec_tlu_force_halt | _T_35; // @[el2_ifu_mem_ctl.scala 205:51]
  wire  _T_38 = ~last_data_recieved_ff; // @[el2_ifu_mem_ctl.scala 206:30]
  wire  _T_39 = ic_byp_hit_f & _T_38; // @[el2_ifu_mem_ctl.scala 206:27]
  wire  _T_40 = _T_39 & uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 206:53]
  wire  _T_42 = ~ic_byp_hit_f; // @[el2_ifu_mem_ctl.scala 207:16]
  wire  _T_44 = _T_42 & _T_317; // @[el2_ifu_mem_ctl.scala 207:30]
  wire  _T_46 = _T_44 & _T_32; // @[el2_ifu_mem_ctl.scala 207:52]
  wire  _T_47 = _T_46 & uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 207:85]
  wire  _T_51 = _T_32 & _T_17; // @[el2_ifu_mem_ctl.scala 208:49]
  wire  _T_54 = ic_byp_hit_f & _T_317; // @[el2_ifu_mem_ctl.scala 209:33]
  wire  _T_56 = ~_T_32; // @[el2_ifu_mem_ctl.scala 209:57]
  wire  _T_57 = _T_54 & _T_56; // @[el2_ifu_mem_ctl.scala 209:55]
  wire  ifu_bp_hit_taken_q_f = io_ifu_bp_hit_taken_f & io_ic_hit_f; // @[el2_ifu_mem_ctl.scala 197:52]
  wire  _T_58 = ~ifu_bp_hit_taken_q_f; // @[el2_ifu_mem_ctl.scala 209:91]
  wire  _T_59 = _T_57 & _T_58; // @[el2_ifu_mem_ctl.scala 209:89]
  wire  _T_61 = _T_59 & _T_17; // @[el2_ifu_mem_ctl.scala 209:113]
  wire  _T_64 = bus_ifu_wr_en_ff & _T_317; // @[el2_ifu_mem_ctl.scala 210:39]
  wire  _T_67 = _T_64 & _T_56; // @[el2_ifu_mem_ctl.scala 210:61]
  wire  _T_69 = _T_67 & _T_58; // @[el2_ifu_mem_ctl.scala 210:95]
  wire  _T_71 = _T_69 & _T_17; // @[el2_ifu_mem_ctl.scala 210:119]
  wire  _T_79 = _T_46 & _T_17; // @[el2_ifu_mem_ctl.scala 211:100]
  wire  _T_81 = io_exu_flush_final | ifu_bp_hit_taken_q_f; // @[el2_ifu_mem_ctl.scala 212:44]
  wire  _T_84 = _T_81 & _T_56; // @[el2_ifu_mem_ctl.scala 212:68]
  wire [2:0] _T_86 = _T_84 ? 3'h2 : 3'h0; // @[el2_ifu_mem_ctl.scala 212:22]
  wire [2:0] _T_87 = _T_79 ? 3'h0 : _T_86; // @[el2_ifu_mem_ctl.scala 211:20]
  wire [2:0] _T_88 = _T_71 ? 3'h6 : _T_87; // @[el2_ifu_mem_ctl.scala 210:20]
  wire [2:0] _T_89 = _T_61 ? 3'h6 : _T_88; // @[el2_ifu_mem_ctl.scala 209:18]
  wire [2:0] _T_90 = _T_51 ? 3'h0 : _T_89; // @[el2_ifu_mem_ctl.scala 208:16]
  wire [2:0] _T_91 = _T_47 ? 3'h4 : _T_90; // @[el2_ifu_mem_ctl.scala 207:14]
  wire [2:0] _T_92 = _T_40 ? 3'h3 : _T_91; // @[el2_ifu_mem_ctl.scala 206:12]
  wire [2:0] _T_93 = _T_36 ? 3'h0 : _T_92; // @[el2_ifu_mem_ctl.scala 205:27]
  wire  _T_102 = 3'h4 == miss_state; // @[Conditional.scala 37:30]
  wire  _T_106 = 3'h6 == miss_state; // @[Conditional.scala 37:30]
  wire  _T_2247 = byp_fetch_index[4:1] == 4'h7; // @[el2_ifu_mem_ctl.scala 462:60]
  wire  _T_2248 = _T_2247 & ifc_fetch_req_f; // @[el2_ifu_mem_ctl.scala 462:92]
  wire  stream_eol_f = _T_2248 & stream_hit_f; // @[el2_ifu_mem_ctl.scala 462:110]
  wire  _T_108 = _T_81 | stream_eol_f; // @[el2_ifu_mem_ctl.scala 220:72]
  wire  _T_111 = _T_108 & _T_56; // @[el2_ifu_mem_ctl.scala 220:87]
  wire  _T_113 = _T_111 & _T_2549; // @[el2_ifu_mem_ctl.scala 220:122]
  wire [2:0] _T_115 = _T_113 ? 3'h2 : 3'h0; // @[el2_ifu_mem_ctl.scala 220:27]
  wire  _T_121 = 3'h3 == miss_state; // @[Conditional.scala 37:30]
  wire  _T_124 = io_exu_flush_final & _T_56; // @[el2_ifu_mem_ctl.scala 224:48]
  wire  _T_126 = _T_124 & _T_2549; // @[el2_ifu_mem_ctl.scala 224:82]
  wire [2:0] _T_128 = _T_126 ? 3'h2 : 3'h0; // @[el2_ifu_mem_ctl.scala 224:27]
  wire  _T_132 = 3'h2 == miss_state; // @[Conditional.scala 37:30]
  wire  _T_236 = io_ic_rd_hit == 2'h0; // @[el2_ifu_mem_ctl.scala 285:28]
  wire  _T_237 = _T_236 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 285:42]
  wire  _T_238 = _T_237 & fetch_req_icache_f; // @[el2_ifu_mem_ctl.scala 285:60]
  wire  _T_239 = miss_state == 3'h2; // @[el2_ifu_mem_ctl.scala 285:94]
  wire  _T_240 = _T_238 & _T_239; // @[el2_ifu_mem_ctl.scala 285:81]
  wire  _T_243 = imb_ff[30:5] != ifu_fetch_addr_int_f[30:5]; // @[el2_ifu_mem_ctl.scala 286:39]
  wire  _T_244 = _T_240 & _T_243; // @[el2_ifu_mem_ctl.scala 285:111]
  wire  _T_246 = _T_244 & _T_17; // @[el2_ifu_mem_ctl.scala 286:91]
  reg  sel_mb_addr_ff; // @[el2_ifu_mem_ctl.scala 339:51]
  wire  _T_247 = ~sel_mb_addr_ff; // @[el2_ifu_mem_ctl.scala 286:116]
  wire  _T_248 = _T_246 & _T_247; // @[el2_ifu_mem_ctl.scala 286:114]
  wire  ic_miss_under_miss_f = _T_248 & _T_209; // @[el2_ifu_mem_ctl.scala 286:132]
  wire  _T_135 = ic_miss_under_miss_f & _T_56; // @[el2_ifu_mem_ctl.scala 228:50]
  wire  _T_137 = _T_135 & _T_2549; // @[el2_ifu_mem_ctl.scala 228:84]
  wire  _T_256 = _T_230 & _T_239; // @[el2_ifu_mem_ctl.scala 287:85]
  wire  _T_259 = imb_ff[30:5] == ifu_fetch_addr_int_f[30:5]; // @[el2_ifu_mem_ctl.scala 288:39]
  wire  _T_260 = _T_259 | uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 288:91]
  wire  ic_ignore_2nd_miss_f = _T_256 & _T_260; // @[el2_ifu_mem_ctl.scala 287:117]
  wire  _T_141 = ic_ignore_2nd_miss_f & _T_56; // @[el2_ifu_mem_ctl.scala 229:35]
  wire  _T_143 = _T_141 & _T_2549; // @[el2_ifu_mem_ctl.scala 229:69]
  wire [2:0] _T_145 = _T_143 ? 3'h7 : 3'h0; // @[el2_ifu_mem_ctl.scala 229:12]
  wire [2:0] _T_146 = _T_137 ? 3'h5 : _T_145; // @[el2_ifu_mem_ctl.scala 228:27]
  wire  _T_151 = 3'h5 == miss_state; // @[Conditional.scala 37:30]
  wire [2:0] _T_154 = _T_32 ? 3'h0 : 3'h2; // @[el2_ifu_mem_ctl.scala 234:12]
  wire [2:0] _T_155 = io_exu_flush_final ? _T_154 : 3'h1; // @[el2_ifu_mem_ctl.scala 233:62]
  wire [2:0] _T_156 = io_dec_tlu_force_halt ? 3'h0 : _T_155; // @[el2_ifu_mem_ctl.scala 233:27]
  wire  _T_160 = 3'h7 == miss_state; // @[Conditional.scala 37:30]
  wire [2:0] _T_164 = io_exu_flush_final ? _T_154 : 3'h0; // @[el2_ifu_mem_ctl.scala 238:62]
  wire [2:0] _T_165 = io_dec_tlu_force_halt ? 3'h0 : _T_164; // @[el2_ifu_mem_ctl.scala 238:27]
  wire [2:0] _GEN_0 = _T_160 ? _T_165 : 3'h0; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_2 = _T_151 ? _T_156 : _GEN_0; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_4 = _T_132 ? _T_146 : _GEN_2; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_6 = _T_121 ? _T_128 : _GEN_4; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_8 = _T_106 ? _T_115 : _GEN_6; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_10 = _T_102 ? 3'h0 : _GEN_8; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_12 = _T_31 ? _T_93 : _GEN_10; // @[Conditional.scala 39:67]
  wire [2:0] miss_nxtstate = _T_24 ? _T_28 : _GEN_12; // @[Conditional.scala 40:58]
  wire  _T_20 = miss_nxtstate == 3'h5; // @[el2_ifu_mem_ctl.scala 195:73]
  wire  _T_21 = _T_19 | _T_20; // @[el2_ifu_mem_ctl.scala 195:57]
  wire  _T_22 = _T_18 & _T_21; // @[el2_ifu_mem_ctl.scala 195:26]
  wire  scnd_miss_req_in = _T_22 & _T_317; // @[el2_ifu_mem_ctl.scala 195:91]
  wire  _T_30 = ic_act_miss_f & _T_2549; // @[el2_ifu_mem_ctl.scala 202:38]
  wire  _T_94 = io_dec_tlu_force_halt | io_exu_flush_final; // @[el2_ifu_mem_ctl.scala 213:46]
  wire  _T_95 = _T_94 | ic_byp_hit_f; // @[el2_ifu_mem_ctl.scala 213:67]
  wire  _T_96 = _T_95 | ifu_bp_hit_taken_q_f; // @[el2_ifu_mem_ctl.scala 213:82]
  wire  _T_98 = _T_96 | _T_32; // @[el2_ifu_mem_ctl.scala 213:105]
  wire  _T_100 = bus_ifu_wr_en_ff & _T_17; // @[el2_ifu_mem_ctl.scala 213:158]
  wire  _T_101 = _T_98 | _T_100; // @[el2_ifu_mem_ctl.scala 213:138]
  wire  _T_103 = io_exu_flush_final | flush_final_f; // @[el2_ifu_mem_ctl.scala 217:43]
  wire  _T_104 = _T_103 | ic_byp_hit_f; // @[el2_ifu_mem_ctl.scala 217:59]
  wire  _T_105 = _T_104 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 217:74]
  wire  _T_119 = _T_108 | _T_32; // @[el2_ifu_mem_ctl.scala 221:84]
  wire  _T_120 = _T_119 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 221:118]
  wire  _T_130 = io_exu_flush_final | _T_32; // @[el2_ifu_mem_ctl.scala 225:43]
  wire  _T_131 = _T_130 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 225:76]
  wire  _T_148 = _T_32 | ic_miss_under_miss_f; // @[el2_ifu_mem_ctl.scala 230:55]
  wire  _T_149 = _T_148 | ic_ignore_2nd_miss_f; // @[el2_ifu_mem_ctl.scala 230:78]
  wire  _T_150 = _T_149 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 230:101]
  wire  _T_158 = _T_32 | io_exu_flush_final; // @[el2_ifu_mem_ctl.scala 235:55]
  wire  _T_159 = _T_158 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 235:76]
  wire  _GEN_1 = _T_160 & _T_159; // @[Conditional.scala 39:67]
  wire  _GEN_3 = _T_151 ? _T_159 : _GEN_1; // @[Conditional.scala 39:67]
  wire  _GEN_5 = _T_132 ? _T_150 : _GEN_3; // @[Conditional.scala 39:67]
  wire  _GEN_7 = _T_121 ? _T_131 : _GEN_5; // @[Conditional.scala 39:67]
  wire  _GEN_9 = _T_106 ? _T_120 : _GEN_7; // @[Conditional.scala 39:67]
  wire  _GEN_11 = _T_102 ? _T_105 : _GEN_9; // @[Conditional.scala 39:67]
  wire  _GEN_13 = _T_31 ? _T_101 : _GEN_11; // @[Conditional.scala 39:67]
  wire  miss_state_en = _T_24 ? _T_30 : _GEN_13; // @[Conditional.scala 40:58]
  wire  _T_174 = ~flush_final_f; // @[el2_ifu_mem_ctl.scala 255:95]
  wire  _T_175 = _T_2250 & _T_174; // @[el2_ifu_mem_ctl.scala 255:93]
  wire  crit_wd_byp_ok_ff = _T_2251 | _T_175; // @[el2_ifu_mem_ctl.scala 255:58]
  wire  _T_178 = miss_pending & _T_56; // @[el2_ifu_mem_ctl.scala 256:36]
  wire  _T_180 = _T_2250 & io_exu_flush_final; // @[el2_ifu_mem_ctl.scala 256:106]
  wire  _T_181 = ~_T_180; // @[el2_ifu_mem_ctl.scala 256:72]
  wire  _T_182 = _T_178 & _T_181; // @[el2_ifu_mem_ctl.scala 256:70]
  wire  _T_184 = _T_2250 & crit_byp_hit_f; // @[el2_ifu_mem_ctl.scala 257:57]
  wire  _T_185 = ~_T_184; // @[el2_ifu_mem_ctl.scala 257:23]
  wire  _T_186 = _T_182 & _T_185; // @[el2_ifu_mem_ctl.scala 256:128]
  wire  _T_187 = _T_186 | ic_act_miss_f; // @[el2_ifu_mem_ctl.scala 257:77]
  wire  _T_188 = miss_nxtstate == 3'h4; // @[el2_ifu_mem_ctl.scala 258:36]
  wire  _T_189 = miss_pending & _T_188; // @[el2_ifu_mem_ctl.scala 258:19]
  wire  sel_hold_imb = _T_187 | _T_189; // @[el2_ifu_mem_ctl.scala 257:93]
  wire  _T_191 = _T_19 | ic_miss_under_miss_f; // @[el2_ifu_mem_ctl.scala 260:57]
  wire  sel_hold_imb_scnd = _T_191 & _T_174; // @[el2_ifu_mem_ctl.scala 260:81]
  reg  way_status_mb_scnd_ff; // @[el2_ifu_mem_ctl.scala 268:35]
  reg [6:0] _T_5128; // @[el2_ifu_mem_ctl.scala 730:14]
  wire [5:0] ifu_ic_rw_int_addr_ff = _T_5128[5:0]; // @[el2_ifu_mem_ctl.scala 729:27]
  wire [6:0] _GEN_472 = {{1'd0}, ifu_ic_rw_int_addr_ff}; // @[el2_ifu_mem_ctl.scala 726:121]
  wire  _T_4993 = _GEN_472 == 7'h7f; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4995 = _T_4993 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4484; // @[Reg.scala 27:20]
  wire  way_status_out_127 = _T_4484[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_473 = {{5'd0}, way_status_out_127}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4996 = _T_4995 & _GEN_473; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4989 = _GEN_472 == 7'h7e; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4991 = _T_4989 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4480; // @[Reg.scala 27:20]
  wire  way_status_out_126 = _T_4480[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_475 = {{5'd0}, way_status_out_126}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4992 = _T_4991 & _GEN_475; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4985 = _GEN_472 == 7'h7d; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4987 = _T_4985 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4476; // @[Reg.scala 27:20]
  wire  way_status_out_125 = _T_4476[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_477 = {{5'd0}, way_status_out_125}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4988 = _T_4987 & _GEN_477; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4981 = _GEN_472 == 7'h7c; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4983 = _T_4981 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4472; // @[Reg.scala 27:20]
  wire  way_status_out_124 = _T_4472[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_479 = {{5'd0}, way_status_out_124}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4984 = _T_4983 & _GEN_479; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4977 = _GEN_472 == 7'h7b; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4979 = _T_4977 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4468; // @[Reg.scala 27:20]
  wire  way_status_out_123 = _T_4468[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_481 = {{5'd0}, way_status_out_123}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4980 = _T_4979 & _GEN_481; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4973 = _GEN_472 == 7'h7a; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4975 = _T_4973 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4464; // @[Reg.scala 27:20]
  wire  way_status_out_122 = _T_4464[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_483 = {{5'd0}, way_status_out_122}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4976 = _T_4975 & _GEN_483; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4969 = _GEN_472 == 7'h79; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4971 = _T_4969 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4460; // @[Reg.scala 27:20]
  wire  way_status_out_121 = _T_4460[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_485 = {{5'd0}, way_status_out_121}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4972 = _T_4971 & _GEN_485; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4965 = _GEN_472 == 7'h78; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4967 = _T_4965 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4456; // @[Reg.scala 27:20]
  wire  way_status_out_120 = _T_4456[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_487 = {{5'd0}, way_status_out_120}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4968 = _T_4967 & _GEN_487; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4961 = _GEN_472 == 7'h77; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4963 = _T_4961 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4452; // @[Reg.scala 27:20]
  wire  way_status_out_119 = _T_4452[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_489 = {{5'd0}, way_status_out_119}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4964 = _T_4963 & _GEN_489; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4957 = _GEN_472 == 7'h76; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4959 = _T_4957 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4448; // @[Reg.scala 27:20]
  wire  way_status_out_118 = _T_4448[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_491 = {{5'd0}, way_status_out_118}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4960 = _T_4959 & _GEN_491; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [59:0] _T_5005 = {_T_4996,_T_4992,_T_4988,_T_4984,_T_4980,_T_4976,_T_4972,_T_4968,_T_4964,_T_4960}; // @[Cat.scala 29:58]
  wire  _T_4953 = _GEN_472 == 7'h75; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4955 = _T_4953 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4444; // @[Reg.scala 27:20]
  wire  way_status_out_117 = _T_4444[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_493 = {{5'd0}, way_status_out_117}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4956 = _T_4955 & _GEN_493; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4949 = _GEN_472 == 7'h74; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4951 = _T_4949 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4440; // @[Reg.scala 27:20]
  wire  way_status_out_116 = _T_4440[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_495 = {{5'd0}, way_status_out_116}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4952 = _T_4951 & _GEN_495; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4945 = _GEN_472 == 7'h73; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4947 = _T_4945 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4436; // @[Reg.scala 27:20]
  wire  way_status_out_115 = _T_4436[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_497 = {{5'd0}, way_status_out_115}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4948 = _T_4947 & _GEN_497; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4941 = _GEN_472 == 7'h72; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4943 = _T_4941 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4432; // @[Reg.scala 27:20]
  wire  way_status_out_114 = _T_4432[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_499 = {{5'd0}, way_status_out_114}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4944 = _T_4943 & _GEN_499; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4937 = _GEN_472 == 7'h71; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4939 = _T_4937 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4428; // @[Reg.scala 27:20]
  wire  way_status_out_113 = _T_4428[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_501 = {{5'd0}, way_status_out_113}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4940 = _T_4939 & _GEN_501; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4933 = _GEN_472 == 7'h70; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4935 = _T_4933 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4424; // @[Reg.scala 27:20]
  wire  way_status_out_112 = _T_4424[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_503 = {{5'd0}, way_status_out_112}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4936 = _T_4935 & _GEN_503; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4929 = _GEN_472 == 7'h6f; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4931 = _T_4929 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4420; // @[Reg.scala 27:20]
  wire  way_status_out_111 = _T_4420[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_505 = {{5'd0}, way_status_out_111}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4932 = _T_4931 & _GEN_505; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4925 = _GEN_472 == 7'h6e; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4927 = _T_4925 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4416; // @[Reg.scala 27:20]
  wire  way_status_out_110 = _T_4416[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_507 = {{5'd0}, way_status_out_110}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4928 = _T_4927 & _GEN_507; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4921 = _GEN_472 == 7'h6d; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4923 = _T_4921 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4412; // @[Reg.scala 27:20]
  wire  way_status_out_109 = _T_4412[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_509 = {{5'd0}, way_status_out_109}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4924 = _T_4923 & _GEN_509; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [113:0] _T_5014 = {_T_5005,_T_4956,_T_4952,_T_4948,_T_4944,_T_4940,_T_4936,_T_4932,_T_4928,_T_4924}; // @[Cat.scala 29:58]
  wire  _T_4917 = _GEN_472 == 7'h6c; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4919 = _T_4917 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4408; // @[Reg.scala 27:20]
  wire  way_status_out_108 = _T_4408[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_511 = {{5'd0}, way_status_out_108}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4920 = _T_4919 & _GEN_511; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4913 = _GEN_472 == 7'h6b; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4915 = _T_4913 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4404; // @[Reg.scala 27:20]
  wire  way_status_out_107 = _T_4404[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_513 = {{5'd0}, way_status_out_107}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4916 = _T_4915 & _GEN_513; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4909 = _GEN_472 == 7'h6a; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4911 = _T_4909 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4400; // @[Reg.scala 27:20]
  wire  way_status_out_106 = _T_4400[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_515 = {{5'd0}, way_status_out_106}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4912 = _T_4911 & _GEN_515; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4905 = _GEN_472 == 7'h69; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4907 = _T_4905 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4396; // @[Reg.scala 27:20]
  wire  way_status_out_105 = _T_4396[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_517 = {{5'd0}, way_status_out_105}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4908 = _T_4907 & _GEN_517; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4901 = _GEN_472 == 7'h68; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4903 = _T_4901 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4392; // @[Reg.scala 27:20]
  wire  way_status_out_104 = _T_4392[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_519 = {{5'd0}, way_status_out_104}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4904 = _T_4903 & _GEN_519; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4897 = _GEN_472 == 7'h67; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4899 = _T_4897 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4388; // @[Reg.scala 27:20]
  wire  way_status_out_103 = _T_4388[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_521 = {{5'd0}, way_status_out_103}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4900 = _T_4899 & _GEN_521; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4893 = _GEN_472 == 7'h66; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4895 = _T_4893 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4384; // @[Reg.scala 27:20]
  wire  way_status_out_102 = _T_4384[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_523 = {{5'd0}, way_status_out_102}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4896 = _T_4895 & _GEN_523; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4889 = _GEN_472 == 7'h65; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4891 = _T_4889 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4380; // @[Reg.scala 27:20]
  wire  way_status_out_101 = _T_4380[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_525 = {{5'd0}, way_status_out_101}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4892 = _T_4891 & _GEN_525; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4885 = _GEN_472 == 7'h64; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4887 = _T_4885 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4376; // @[Reg.scala 27:20]
  wire  way_status_out_100 = _T_4376[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_527 = {{5'd0}, way_status_out_100}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4888 = _T_4887 & _GEN_527; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [167:0] _T_5023 = {_T_5014,_T_4920,_T_4916,_T_4912,_T_4908,_T_4904,_T_4900,_T_4896,_T_4892,_T_4888}; // @[Cat.scala 29:58]
  wire  _T_4881 = _GEN_472 == 7'h63; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4883 = _T_4881 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4372; // @[Reg.scala 27:20]
  wire  way_status_out_99 = _T_4372[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_529 = {{5'd0}, way_status_out_99}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4884 = _T_4883 & _GEN_529; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4877 = _GEN_472 == 7'h62; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4879 = _T_4877 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4368; // @[Reg.scala 27:20]
  wire  way_status_out_98 = _T_4368[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_531 = {{5'd0}, way_status_out_98}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4880 = _T_4879 & _GEN_531; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4873 = _GEN_472 == 7'h61; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4875 = _T_4873 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4364; // @[Reg.scala 27:20]
  wire  way_status_out_97 = _T_4364[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_533 = {{5'd0}, way_status_out_97}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4876 = _T_4875 & _GEN_533; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4869 = _GEN_472 == 7'h60; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4871 = _T_4869 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4360; // @[Reg.scala 27:20]
  wire  way_status_out_96 = _T_4360[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_535 = {{5'd0}, way_status_out_96}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4872 = _T_4871 & _GEN_535; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4865 = _GEN_472 == 7'h5f; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4867 = _T_4865 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4356; // @[Reg.scala 27:20]
  wire  way_status_out_95 = _T_4356[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_537 = {{5'd0}, way_status_out_95}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4868 = _T_4867 & _GEN_537; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4861 = _GEN_472 == 7'h5e; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4863 = _T_4861 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4352; // @[Reg.scala 27:20]
  wire  way_status_out_94 = _T_4352[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_539 = {{5'd0}, way_status_out_94}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4864 = _T_4863 & _GEN_539; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4857 = _GEN_472 == 7'h5d; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4859 = _T_4857 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4348; // @[Reg.scala 27:20]
  wire  way_status_out_93 = _T_4348[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_541 = {{5'd0}, way_status_out_93}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4860 = _T_4859 & _GEN_541; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4853 = _GEN_472 == 7'h5c; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4855 = _T_4853 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4344; // @[Reg.scala 27:20]
  wire  way_status_out_92 = _T_4344[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_543 = {{5'd0}, way_status_out_92}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4856 = _T_4855 & _GEN_543; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4849 = _GEN_472 == 7'h5b; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4851 = _T_4849 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4340; // @[Reg.scala 27:20]
  wire  way_status_out_91 = _T_4340[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_545 = {{5'd0}, way_status_out_91}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4852 = _T_4851 & _GEN_545; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [221:0] _T_5032 = {_T_5023,_T_4884,_T_4880,_T_4876,_T_4872,_T_4868,_T_4864,_T_4860,_T_4856,_T_4852}; // @[Cat.scala 29:58]
  wire  _T_4845 = _GEN_472 == 7'h5a; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4847 = _T_4845 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4336; // @[Reg.scala 27:20]
  wire  way_status_out_90 = _T_4336[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_547 = {{5'd0}, way_status_out_90}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4848 = _T_4847 & _GEN_547; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4841 = _GEN_472 == 7'h59; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4843 = _T_4841 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4332; // @[Reg.scala 27:20]
  wire  way_status_out_89 = _T_4332[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_549 = {{5'd0}, way_status_out_89}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4844 = _T_4843 & _GEN_549; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4837 = _GEN_472 == 7'h58; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4839 = _T_4837 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4328; // @[Reg.scala 27:20]
  wire  way_status_out_88 = _T_4328[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_551 = {{5'd0}, way_status_out_88}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4840 = _T_4839 & _GEN_551; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4833 = _GEN_472 == 7'h57; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4835 = _T_4833 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4324; // @[Reg.scala 27:20]
  wire  way_status_out_87 = _T_4324[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_553 = {{5'd0}, way_status_out_87}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4836 = _T_4835 & _GEN_553; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4829 = _GEN_472 == 7'h56; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4831 = _T_4829 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4320; // @[Reg.scala 27:20]
  wire  way_status_out_86 = _T_4320[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_555 = {{5'd0}, way_status_out_86}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4832 = _T_4831 & _GEN_555; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4825 = _GEN_472 == 7'h55; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4827 = _T_4825 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4316; // @[Reg.scala 27:20]
  wire  way_status_out_85 = _T_4316[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_557 = {{5'd0}, way_status_out_85}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4828 = _T_4827 & _GEN_557; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4821 = _GEN_472 == 7'h54; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4823 = _T_4821 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4312; // @[Reg.scala 27:20]
  wire  way_status_out_84 = _T_4312[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_559 = {{5'd0}, way_status_out_84}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4824 = _T_4823 & _GEN_559; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4817 = _GEN_472 == 7'h53; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4819 = _T_4817 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4308; // @[Reg.scala 27:20]
  wire  way_status_out_83 = _T_4308[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_561 = {{5'd0}, way_status_out_83}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4820 = _T_4819 & _GEN_561; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4813 = _GEN_472 == 7'h52; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4815 = _T_4813 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4304; // @[Reg.scala 27:20]
  wire  way_status_out_82 = _T_4304[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_563 = {{5'd0}, way_status_out_82}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4816 = _T_4815 & _GEN_563; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [275:0] _T_5041 = {_T_5032,_T_4848,_T_4844,_T_4840,_T_4836,_T_4832,_T_4828,_T_4824,_T_4820,_T_4816}; // @[Cat.scala 29:58]
  wire  _T_4809 = _GEN_472 == 7'h51; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4811 = _T_4809 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4300; // @[Reg.scala 27:20]
  wire  way_status_out_81 = _T_4300[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_565 = {{5'd0}, way_status_out_81}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4812 = _T_4811 & _GEN_565; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4805 = _GEN_472 == 7'h50; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4807 = _T_4805 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4296; // @[Reg.scala 27:20]
  wire  way_status_out_80 = _T_4296[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_567 = {{5'd0}, way_status_out_80}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4808 = _T_4807 & _GEN_567; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4801 = _GEN_472 == 7'h4f; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4803 = _T_4801 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4292; // @[Reg.scala 27:20]
  wire  way_status_out_79 = _T_4292[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_569 = {{5'd0}, way_status_out_79}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4804 = _T_4803 & _GEN_569; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4797 = _GEN_472 == 7'h4e; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4799 = _T_4797 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4288; // @[Reg.scala 27:20]
  wire  way_status_out_78 = _T_4288[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_571 = {{5'd0}, way_status_out_78}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4800 = _T_4799 & _GEN_571; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4793 = _GEN_472 == 7'h4d; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4795 = _T_4793 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4284; // @[Reg.scala 27:20]
  wire  way_status_out_77 = _T_4284[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_573 = {{5'd0}, way_status_out_77}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4796 = _T_4795 & _GEN_573; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4789 = _GEN_472 == 7'h4c; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4791 = _T_4789 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4280; // @[Reg.scala 27:20]
  wire  way_status_out_76 = _T_4280[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_575 = {{5'd0}, way_status_out_76}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4792 = _T_4791 & _GEN_575; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4785 = _GEN_472 == 7'h4b; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4787 = _T_4785 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4276; // @[Reg.scala 27:20]
  wire  way_status_out_75 = _T_4276[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_577 = {{5'd0}, way_status_out_75}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4788 = _T_4787 & _GEN_577; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4781 = _GEN_472 == 7'h4a; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4783 = _T_4781 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4272; // @[Reg.scala 27:20]
  wire  way_status_out_74 = _T_4272[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_579 = {{5'd0}, way_status_out_74}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4784 = _T_4783 & _GEN_579; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4777 = _GEN_472 == 7'h49; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4779 = _T_4777 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4268; // @[Reg.scala 27:20]
  wire  way_status_out_73 = _T_4268[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_581 = {{5'd0}, way_status_out_73}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4780 = _T_4779 & _GEN_581; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [329:0] _T_5050 = {_T_5041,_T_4812,_T_4808,_T_4804,_T_4800,_T_4796,_T_4792,_T_4788,_T_4784,_T_4780}; // @[Cat.scala 29:58]
  wire  _T_4773 = _GEN_472 == 7'h48; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4775 = _T_4773 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4264; // @[Reg.scala 27:20]
  wire  way_status_out_72 = _T_4264[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_583 = {{5'd0}, way_status_out_72}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4776 = _T_4775 & _GEN_583; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4769 = _GEN_472 == 7'h47; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4771 = _T_4769 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4260; // @[Reg.scala 27:20]
  wire  way_status_out_71 = _T_4260[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_585 = {{5'd0}, way_status_out_71}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4772 = _T_4771 & _GEN_585; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4765 = _GEN_472 == 7'h46; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4767 = _T_4765 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4256; // @[Reg.scala 27:20]
  wire  way_status_out_70 = _T_4256[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_587 = {{5'd0}, way_status_out_70}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4768 = _T_4767 & _GEN_587; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4761 = _GEN_472 == 7'h45; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4763 = _T_4761 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4252; // @[Reg.scala 27:20]
  wire  way_status_out_69 = _T_4252[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_589 = {{5'd0}, way_status_out_69}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4764 = _T_4763 & _GEN_589; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4757 = _GEN_472 == 7'h44; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4759 = _T_4757 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4248; // @[Reg.scala 27:20]
  wire  way_status_out_68 = _T_4248[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_591 = {{5'd0}, way_status_out_68}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4760 = _T_4759 & _GEN_591; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4753 = _GEN_472 == 7'h43; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4755 = _T_4753 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4244; // @[Reg.scala 27:20]
  wire  way_status_out_67 = _T_4244[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_593 = {{5'd0}, way_status_out_67}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4756 = _T_4755 & _GEN_593; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4749 = _GEN_472 == 7'h42; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4751 = _T_4749 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4240; // @[Reg.scala 27:20]
  wire  way_status_out_66 = _T_4240[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_595 = {{5'd0}, way_status_out_66}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4752 = _T_4751 & _GEN_595; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4745 = _GEN_472 == 7'h41; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4747 = _T_4745 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4236; // @[Reg.scala 27:20]
  wire  way_status_out_65 = _T_4236[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_597 = {{5'd0}, way_status_out_65}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4748 = _T_4747 & _GEN_597; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4741 = _GEN_472 == 7'h40; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4743 = _T_4741 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4232; // @[Reg.scala 27:20]
  wire  way_status_out_64 = _T_4232[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_599 = {{5'd0}, way_status_out_64}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4744 = _T_4743 & _GEN_599; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [383:0] _T_5059 = {_T_5050,_T_4776,_T_4772,_T_4768,_T_4764,_T_4760,_T_4756,_T_4752,_T_4748,_T_4744}; // @[Cat.scala 29:58]
  wire  _T_4737 = ifu_ic_rw_int_addr_ff == 6'h3f; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4739 = _T_4737 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4228; // @[Reg.scala 27:20]
  wire  way_status_out_63 = _T_4228[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_600 = {{5'd0}, way_status_out_63}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4740 = _T_4739 & _GEN_600; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4733 = ifu_ic_rw_int_addr_ff == 6'h3e; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4735 = _T_4733 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4224; // @[Reg.scala 27:20]
  wire  way_status_out_62 = _T_4224[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_601 = {{5'd0}, way_status_out_62}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4736 = _T_4735 & _GEN_601; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4729 = ifu_ic_rw_int_addr_ff == 6'h3d; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4731 = _T_4729 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4220; // @[Reg.scala 27:20]
  wire  way_status_out_61 = _T_4220[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_602 = {{5'd0}, way_status_out_61}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4732 = _T_4731 & _GEN_602; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4725 = ifu_ic_rw_int_addr_ff == 6'h3c; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4727 = _T_4725 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4216; // @[Reg.scala 27:20]
  wire  way_status_out_60 = _T_4216[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_603 = {{5'd0}, way_status_out_60}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4728 = _T_4727 & _GEN_603; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4721 = ifu_ic_rw_int_addr_ff == 6'h3b; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4723 = _T_4721 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4212; // @[Reg.scala 27:20]
  wire  way_status_out_59 = _T_4212[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_604 = {{5'd0}, way_status_out_59}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4724 = _T_4723 & _GEN_604; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4717 = ifu_ic_rw_int_addr_ff == 6'h3a; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4719 = _T_4717 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4208; // @[Reg.scala 27:20]
  wire  way_status_out_58 = _T_4208[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_605 = {{5'd0}, way_status_out_58}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4720 = _T_4719 & _GEN_605; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4713 = ifu_ic_rw_int_addr_ff == 6'h39; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4715 = _T_4713 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4204; // @[Reg.scala 27:20]
  wire  way_status_out_57 = _T_4204[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_606 = {{5'd0}, way_status_out_57}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4716 = _T_4715 & _GEN_606; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4709 = ifu_ic_rw_int_addr_ff == 6'h38; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4711 = _T_4709 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4200; // @[Reg.scala 27:20]
  wire  way_status_out_56 = _T_4200[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_607 = {{5'd0}, way_status_out_56}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4712 = _T_4711 & _GEN_607; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4705 = ifu_ic_rw_int_addr_ff == 6'h37; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4707 = _T_4705 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4196; // @[Reg.scala 27:20]
  wire  way_status_out_55 = _T_4196[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_608 = {{5'd0}, way_status_out_55}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4708 = _T_4707 & _GEN_608; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [437:0] _T_5068 = {_T_5059,_T_4740,_T_4736,_T_4732,_T_4728,_T_4724,_T_4720,_T_4716,_T_4712,_T_4708}; // @[Cat.scala 29:58]
  wire  _T_4701 = ifu_ic_rw_int_addr_ff == 6'h36; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4703 = _T_4701 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4192; // @[Reg.scala 27:20]
  wire  way_status_out_54 = _T_4192[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_609 = {{5'd0}, way_status_out_54}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4704 = _T_4703 & _GEN_609; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4697 = ifu_ic_rw_int_addr_ff == 6'h35; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4699 = _T_4697 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4188; // @[Reg.scala 27:20]
  wire  way_status_out_53 = _T_4188[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_610 = {{5'd0}, way_status_out_53}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4700 = _T_4699 & _GEN_610; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4693 = ifu_ic_rw_int_addr_ff == 6'h34; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4695 = _T_4693 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4184; // @[Reg.scala 27:20]
  wire  way_status_out_52 = _T_4184[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_611 = {{5'd0}, way_status_out_52}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4696 = _T_4695 & _GEN_611; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4689 = ifu_ic_rw_int_addr_ff == 6'h33; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4691 = _T_4689 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4180; // @[Reg.scala 27:20]
  wire  way_status_out_51 = _T_4180[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_612 = {{5'd0}, way_status_out_51}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4692 = _T_4691 & _GEN_612; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4685 = ifu_ic_rw_int_addr_ff == 6'h32; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4687 = _T_4685 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4176; // @[Reg.scala 27:20]
  wire  way_status_out_50 = _T_4176[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_613 = {{5'd0}, way_status_out_50}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4688 = _T_4687 & _GEN_613; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4681 = ifu_ic_rw_int_addr_ff == 6'h31; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4683 = _T_4681 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4172; // @[Reg.scala 27:20]
  wire  way_status_out_49 = _T_4172[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_614 = {{5'd0}, way_status_out_49}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4684 = _T_4683 & _GEN_614; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4677 = ifu_ic_rw_int_addr_ff == 6'h30; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4679 = _T_4677 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4168; // @[Reg.scala 27:20]
  wire  way_status_out_48 = _T_4168[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_615 = {{5'd0}, way_status_out_48}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4680 = _T_4679 & _GEN_615; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4673 = ifu_ic_rw_int_addr_ff == 6'h2f; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4675 = _T_4673 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4164; // @[Reg.scala 27:20]
  wire  way_status_out_47 = _T_4164[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_616 = {{5'd0}, way_status_out_47}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4676 = _T_4675 & _GEN_616; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4669 = ifu_ic_rw_int_addr_ff == 6'h2e; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4671 = _T_4669 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4160; // @[Reg.scala 27:20]
  wire  way_status_out_46 = _T_4160[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_617 = {{5'd0}, way_status_out_46}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4672 = _T_4671 & _GEN_617; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [491:0] _T_5077 = {_T_5068,_T_4704,_T_4700,_T_4696,_T_4692,_T_4688,_T_4684,_T_4680,_T_4676,_T_4672}; // @[Cat.scala 29:58]
  wire  _T_4665 = ifu_ic_rw_int_addr_ff == 6'h2d; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4667 = _T_4665 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4156; // @[Reg.scala 27:20]
  wire  way_status_out_45 = _T_4156[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_618 = {{5'd0}, way_status_out_45}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4668 = _T_4667 & _GEN_618; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4661 = ifu_ic_rw_int_addr_ff == 6'h2c; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4663 = _T_4661 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4152; // @[Reg.scala 27:20]
  wire  way_status_out_44 = _T_4152[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_619 = {{5'd0}, way_status_out_44}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4664 = _T_4663 & _GEN_619; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4657 = ifu_ic_rw_int_addr_ff == 6'h2b; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4659 = _T_4657 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4148; // @[Reg.scala 27:20]
  wire  way_status_out_43 = _T_4148[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_620 = {{5'd0}, way_status_out_43}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4660 = _T_4659 & _GEN_620; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4653 = ifu_ic_rw_int_addr_ff == 6'h2a; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4655 = _T_4653 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4144; // @[Reg.scala 27:20]
  wire  way_status_out_42 = _T_4144[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_621 = {{5'd0}, way_status_out_42}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4656 = _T_4655 & _GEN_621; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4649 = ifu_ic_rw_int_addr_ff == 6'h29; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4651 = _T_4649 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4140; // @[Reg.scala 27:20]
  wire  way_status_out_41 = _T_4140[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_622 = {{5'd0}, way_status_out_41}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4652 = _T_4651 & _GEN_622; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4645 = ifu_ic_rw_int_addr_ff == 6'h28; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4647 = _T_4645 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4136; // @[Reg.scala 27:20]
  wire  way_status_out_40 = _T_4136[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_623 = {{5'd0}, way_status_out_40}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4648 = _T_4647 & _GEN_623; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4641 = ifu_ic_rw_int_addr_ff == 6'h27; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4643 = _T_4641 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4132; // @[Reg.scala 27:20]
  wire  way_status_out_39 = _T_4132[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_624 = {{5'd0}, way_status_out_39}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4644 = _T_4643 & _GEN_624; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4637 = ifu_ic_rw_int_addr_ff == 6'h26; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4639 = _T_4637 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4128; // @[Reg.scala 27:20]
  wire  way_status_out_38 = _T_4128[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_625 = {{5'd0}, way_status_out_38}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4640 = _T_4639 & _GEN_625; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4633 = ifu_ic_rw_int_addr_ff == 6'h25; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4635 = _T_4633 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4124; // @[Reg.scala 27:20]
  wire  way_status_out_37 = _T_4124[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_626 = {{5'd0}, way_status_out_37}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4636 = _T_4635 & _GEN_626; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [545:0] _T_5086 = {_T_5077,_T_4668,_T_4664,_T_4660,_T_4656,_T_4652,_T_4648,_T_4644,_T_4640,_T_4636}; // @[Cat.scala 29:58]
  wire  _T_4629 = ifu_ic_rw_int_addr_ff == 6'h24; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4631 = _T_4629 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4120; // @[Reg.scala 27:20]
  wire  way_status_out_36 = _T_4120[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_627 = {{5'd0}, way_status_out_36}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4632 = _T_4631 & _GEN_627; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4625 = ifu_ic_rw_int_addr_ff == 6'h23; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4627 = _T_4625 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4116; // @[Reg.scala 27:20]
  wire  way_status_out_35 = _T_4116[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_628 = {{5'd0}, way_status_out_35}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4628 = _T_4627 & _GEN_628; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4621 = ifu_ic_rw_int_addr_ff == 6'h22; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4623 = _T_4621 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4112; // @[Reg.scala 27:20]
  wire  way_status_out_34 = _T_4112[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_629 = {{5'd0}, way_status_out_34}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4624 = _T_4623 & _GEN_629; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4617 = ifu_ic_rw_int_addr_ff == 6'h21; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4619 = _T_4617 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4108; // @[Reg.scala 27:20]
  wire  way_status_out_33 = _T_4108[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_630 = {{5'd0}, way_status_out_33}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4620 = _T_4619 & _GEN_630; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4613 = ifu_ic_rw_int_addr_ff == 6'h20; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4615 = _T_4613 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4104; // @[Reg.scala 27:20]
  wire  way_status_out_32 = _T_4104[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_631 = {{5'd0}, way_status_out_32}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4616 = _T_4615 & _GEN_631; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4609 = ifu_ic_rw_int_addr_ff == 6'h1f; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4611 = _T_4609 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4100; // @[Reg.scala 27:20]
  wire  way_status_out_31 = _T_4100[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_632 = {{5'd0}, way_status_out_31}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4612 = _T_4611 & _GEN_632; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4605 = ifu_ic_rw_int_addr_ff == 6'h1e; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4607 = _T_4605 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4096; // @[Reg.scala 27:20]
  wire  way_status_out_30 = _T_4096[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_633 = {{5'd0}, way_status_out_30}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4608 = _T_4607 & _GEN_633; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4601 = ifu_ic_rw_int_addr_ff == 6'h1d; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4603 = _T_4601 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4092; // @[Reg.scala 27:20]
  wire  way_status_out_29 = _T_4092[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_634 = {{5'd0}, way_status_out_29}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4604 = _T_4603 & _GEN_634; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4597 = ifu_ic_rw_int_addr_ff == 6'h1c; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4599 = _T_4597 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4088; // @[Reg.scala 27:20]
  wire  way_status_out_28 = _T_4088[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_635 = {{5'd0}, way_status_out_28}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4600 = _T_4599 & _GEN_635; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [599:0] _T_5095 = {_T_5086,_T_4632,_T_4628,_T_4624,_T_4620,_T_4616,_T_4612,_T_4608,_T_4604,_T_4600}; // @[Cat.scala 29:58]
  wire  _T_4593 = ifu_ic_rw_int_addr_ff == 6'h1b; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4595 = _T_4593 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4084; // @[Reg.scala 27:20]
  wire  way_status_out_27 = _T_4084[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_636 = {{5'd0}, way_status_out_27}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4596 = _T_4595 & _GEN_636; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4589 = ifu_ic_rw_int_addr_ff == 6'h1a; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4591 = _T_4589 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4080; // @[Reg.scala 27:20]
  wire  way_status_out_26 = _T_4080[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_637 = {{5'd0}, way_status_out_26}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4592 = _T_4591 & _GEN_637; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4585 = ifu_ic_rw_int_addr_ff == 6'h19; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4587 = _T_4585 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4076; // @[Reg.scala 27:20]
  wire  way_status_out_25 = _T_4076[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_638 = {{5'd0}, way_status_out_25}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4588 = _T_4587 & _GEN_638; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4581 = ifu_ic_rw_int_addr_ff == 6'h18; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4583 = _T_4581 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4072; // @[Reg.scala 27:20]
  wire  way_status_out_24 = _T_4072[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_639 = {{5'd0}, way_status_out_24}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4584 = _T_4583 & _GEN_639; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4577 = ifu_ic_rw_int_addr_ff == 6'h17; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4579 = _T_4577 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4068; // @[Reg.scala 27:20]
  wire  way_status_out_23 = _T_4068[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_640 = {{5'd0}, way_status_out_23}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4580 = _T_4579 & _GEN_640; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4573 = ifu_ic_rw_int_addr_ff == 6'h16; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4575 = _T_4573 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4064; // @[Reg.scala 27:20]
  wire  way_status_out_22 = _T_4064[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_641 = {{5'd0}, way_status_out_22}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4576 = _T_4575 & _GEN_641; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4569 = ifu_ic_rw_int_addr_ff == 6'h15; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4571 = _T_4569 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4060; // @[Reg.scala 27:20]
  wire  way_status_out_21 = _T_4060[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_642 = {{5'd0}, way_status_out_21}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4572 = _T_4571 & _GEN_642; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4565 = ifu_ic_rw_int_addr_ff == 6'h14; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4567 = _T_4565 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4056; // @[Reg.scala 27:20]
  wire  way_status_out_20 = _T_4056[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_643 = {{5'd0}, way_status_out_20}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4568 = _T_4567 & _GEN_643; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4561 = ifu_ic_rw_int_addr_ff == 6'h13; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4563 = _T_4561 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4052; // @[Reg.scala 27:20]
  wire  way_status_out_19 = _T_4052[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_644 = {{5'd0}, way_status_out_19}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4564 = _T_4563 & _GEN_644; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [653:0] _T_5104 = {_T_5095,_T_4596,_T_4592,_T_4588,_T_4584,_T_4580,_T_4576,_T_4572,_T_4568,_T_4564}; // @[Cat.scala 29:58]
  wire  _T_4557 = ifu_ic_rw_int_addr_ff == 6'h12; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4559 = _T_4557 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4048; // @[Reg.scala 27:20]
  wire  way_status_out_18 = _T_4048[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_645 = {{5'd0}, way_status_out_18}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4560 = _T_4559 & _GEN_645; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4553 = ifu_ic_rw_int_addr_ff == 6'h11; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4555 = _T_4553 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4044; // @[Reg.scala 27:20]
  wire  way_status_out_17 = _T_4044[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_646 = {{5'd0}, way_status_out_17}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4556 = _T_4555 & _GEN_646; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4549 = ifu_ic_rw_int_addr_ff == 6'h10; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4551 = _T_4549 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4040; // @[Reg.scala 27:20]
  wire  way_status_out_16 = _T_4040[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_647 = {{5'd0}, way_status_out_16}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4552 = _T_4551 & _GEN_647; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4545 = ifu_ic_rw_int_addr_ff == 6'hf; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4547 = _T_4545 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4036; // @[Reg.scala 27:20]
  wire  way_status_out_15 = _T_4036[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_648 = {{5'd0}, way_status_out_15}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4548 = _T_4547 & _GEN_648; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4541 = ifu_ic_rw_int_addr_ff == 6'he; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4543 = _T_4541 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4032; // @[Reg.scala 27:20]
  wire  way_status_out_14 = _T_4032[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_649 = {{5'd0}, way_status_out_14}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4544 = _T_4543 & _GEN_649; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4537 = ifu_ic_rw_int_addr_ff == 6'hd; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4539 = _T_4537 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4028; // @[Reg.scala 27:20]
  wire  way_status_out_13 = _T_4028[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_650 = {{5'd0}, way_status_out_13}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4540 = _T_4539 & _GEN_650; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4533 = ifu_ic_rw_int_addr_ff == 6'hc; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4535 = _T_4533 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4024; // @[Reg.scala 27:20]
  wire  way_status_out_12 = _T_4024[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_651 = {{5'd0}, way_status_out_12}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4536 = _T_4535 & _GEN_651; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4529 = ifu_ic_rw_int_addr_ff == 6'hb; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4531 = _T_4529 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4020; // @[Reg.scala 27:20]
  wire  way_status_out_11 = _T_4020[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_652 = {{5'd0}, way_status_out_11}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4532 = _T_4531 & _GEN_652; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4525 = ifu_ic_rw_int_addr_ff == 6'ha; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4527 = _T_4525 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4016; // @[Reg.scala 27:20]
  wire  way_status_out_10 = _T_4016[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_653 = {{5'd0}, way_status_out_10}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4528 = _T_4527 & _GEN_653; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [707:0] _T_5113 = {_T_5104,_T_4560,_T_4556,_T_4552,_T_4548,_T_4544,_T_4540,_T_4536,_T_4532,_T_4528}; // @[Cat.scala 29:58]
  wire  _T_4521 = ifu_ic_rw_int_addr_ff == 6'h9; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4523 = _T_4521 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4012; // @[Reg.scala 27:20]
  wire  way_status_out_9 = _T_4012[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_654 = {{5'd0}, way_status_out_9}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4524 = _T_4523 & _GEN_654; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4517 = ifu_ic_rw_int_addr_ff == 6'h8; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4519 = _T_4517 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4008; // @[Reg.scala 27:20]
  wire  way_status_out_8 = _T_4008[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_655 = {{5'd0}, way_status_out_8}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4520 = _T_4519 & _GEN_655; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4513 = ifu_ic_rw_int_addr_ff == 6'h7; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4515 = _T_4513 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4004; // @[Reg.scala 27:20]
  wire  way_status_out_7 = _T_4004[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_656 = {{5'd0}, way_status_out_7}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4516 = _T_4515 & _GEN_656; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4509 = ifu_ic_rw_int_addr_ff == 6'h6; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4511 = _T_4509 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4000; // @[Reg.scala 27:20]
  wire  way_status_out_6 = _T_4000[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_657 = {{5'd0}, way_status_out_6}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4512 = _T_4511 & _GEN_657; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4505 = ifu_ic_rw_int_addr_ff == 6'h5; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4507 = _T_4505 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3996; // @[Reg.scala 27:20]
  wire  way_status_out_5 = _T_3996[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_658 = {{5'd0}, way_status_out_5}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4508 = _T_4507 & _GEN_658; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4501 = ifu_ic_rw_int_addr_ff == 6'h4; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4503 = _T_4501 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3992; // @[Reg.scala 27:20]
  wire  way_status_out_4 = _T_3992[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_659 = {{5'd0}, way_status_out_4}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4504 = _T_4503 & _GEN_659; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4497 = ifu_ic_rw_int_addr_ff == 6'h3; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4499 = _T_4497 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3988; // @[Reg.scala 27:20]
  wire  way_status_out_3 = _T_3988[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_660 = {{5'd0}, way_status_out_3}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4500 = _T_4499 & _GEN_660; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4493 = ifu_ic_rw_int_addr_ff == 6'h2; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4495 = _T_4493 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3984; // @[Reg.scala 27:20]
  wire  way_status_out_2 = _T_3984[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_661 = {{5'd0}, way_status_out_2}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4496 = _T_4495 & _GEN_661; // @[el2_ifu_mem_ctl.scala 726:130]
  wire  _T_4489 = ifu_ic_rw_int_addr_ff == 6'h1; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4491 = _T_4489 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3980; // @[Reg.scala 27:20]
  wire  way_status_out_1 = _T_3980[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_662 = {{5'd0}, way_status_out_1}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4492 = _T_4491 & _GEN_662; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [761:0] _T_5122 = {_T_5113,_T_4524,_T_4520,_T_4516,_T_4512,_T_4508,_T_4504,_T_4500,_T_4496,_T_4492}; // @[Cat.scala 29:58]
  wire  _T_4485 = ifu_ic_rw_int_addr_ff == 6'h0; // @[el2_ifu_mem_ctl.scala 726:121]
  wire [5:0] _T_4487 = _T_4485 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3976; // @[Reg.scala 27:20]
  wire  way_status_out_0 = _T_3976[0]; // @[el2_ifu_mem_ctl.scala 723:30 el2_ifu_mem_ctl.scala 725:33]
  wire [5:0] _GEN_663 = {{5'd0}, way_status_out_0}; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [5:0] _T_4488 = _T_4487 & _GEN_663; // @[el2_ifu_mem_ctl.scala 726:130]
  wire [767:0] _T_5123 = {_T_5122,_T_4488}; // @[Cat.scala 29:58]
  wire  way_status = _T_5123[0]; // @[el2_ifu_mem_ctl.scala 726:16]
  wire  _T_195 = ~reset_all_tags; // @[el2_ifu_mem_ctl.scala 263:96]
  reg  uncacheable_miss_scnd_ff; // @[el2_ifu_mem_ctl.scala 265:38]
  reg [30:0] imb_scnd_ff; // @[el2_ifu_mem_ctl.scala 267:25]
  wire [2:0] _T_206 = bus_ifu_wr_en_ff ? 3'h7 : 3'h0; // @[Bitwise.scala 72:12]
  reg [2:0] ifu_bus_rid_ff; // @[Reg.scala 27:20]
  wire [2:0] ic_wr_addr_bits_hi_3 = ifu_bus_rid_ff & _T_206; // @[el2_ifu_mem_ctl.scala 272:45]
  wire  _T_212 = _T_231 | _T_239; // @[el2_ifu_mem_ctl.scala 277:59]
  wire  _T_214 = _T_212 | _T_2235; // @[el2_ifu_mem_ctl.scala 277:91]
  wire  ic_iccm_hit_f = fetch_req_iccm_f & _T_214; // @[el2_ifu_mem_ctl.scala 277:41]
  wire  _T_219 = _T_227 & fetch_req_icache_f; // @[el2_ifu_mem_ctl.scala 283:39]
  wire  _T_221 = _T_219 & _T_195; // @[el2_ifu_mem_ctl.scala 283:60]
  wire  _T_225 = _T_221 & _T_212; // @[el2_ifu_mem_ctl.scala 283:78]
  wire  ic_act_hit_f = _T_225 & _T_247; // @[el2_ifu_mem_ctl.scala 283:126]
  wire  _T_262 = ic_act_hit_f | ic_byp_hit_f; // @[el2_ifu_mem_ctl.scala 290:31]
  wire  _T_263 = _T_262 | ic_iccm_hit_f; // @[el2_ifu_mem_ctl.scala 290:46]
  wire  _T_264 = ifc_region_acc_fault_final_f & ifc_fetch_req_f; // @[el2_ifu_mem_ctl.scala 290:94]
  wire  _T_268 = sel_hold_imb ? uncacheable_miss_ff : io_ifc_fetch_uncacheable_bf; // @[el2_ifu_mem_ctl.scala 291:84]
  wire  uncacheable_miss_in = scnd_miss_req ? uncacheable_miss_scnd_ff : _T_268; // @[el2_ifu_mem_ctl.scala 291:32]
  wire  _T_274 = imb_ff[12:6] == imb_scnd_ff[12:6]; // @[el2_ifu_mem_ctl.scala 294:75]
  wire  _T_275 = _T_274 & scnd_miss_req; // @[el2_ifu_mem_ctl.scala 294:127]
  reg [1:0] ifu_bus_rresp_ff; // @[Reg.scala 27:20]
  wire  _T_2624 = |ifu_bus_rresp_ff; // @[el2_ifu_mem_ctl.scala 624:48]
  wire  _T_2625 = _T_2624 & ifu_bus_rvalid_ff; // @[el2_ifu_mem_ctl.scala 624:52]
  wire  bus_ifu_wr_data_error_ff = _T_2625 & miss_pending; // @[el2_ifu_mem_ctl.scala 624:73]
  reg  ifu_wr_data_comb_err_ff; // @[el2_ifu_mem_ctl.scala 370:61]
  wire  ifu_wr_cumulative_err_data = bus_ifu_wr_data_error_ff | ifu_wr_data_comb_err_ff; // @[el2_ifu_mem_ctl.scala 369:55]
  wire  _T_276 = ~ifu_wr_cumulative_err_data; // @[el2_ifu_mem_ctl.scala 294:145]
  wire  scnd_miss_index_match = _T_275 & _T_276; // @[el2_ifu_mem_ctl.scala 294:143]
  wire  _T_277 = ~scnd_miss_index_match; // @[el2_ifu_mem_ctl.scala 297:47]
  wire  _T_278 = scnd_miss_req & _T_277; // @[el2_ifu_mem_ctl.scala 297:45]
  wire  _T_280 = scnd_miss_req & scnd_miss_index_match; // @[el2_ifu_mem_ctl.scala 298:26]
  reg  way_status_mb_ff; // @[el2_ifu_mem_ctl.scala 317:30]
  wire  _T_10073 = ~way_status_mb_ff; // @[el2_ifu_mem_ctl.scala 779:33]
  reg [1:0] tagv_mb_ff; // @[el2_ifu_mem_ctl.scala 318:24]
  wire  _T_10075 = _T_10073 & tagv_mb_ff[0]; // @[el2_ifu_mem_ctl.scala 779:51]
  wire  _T_10077 = _T_10075 & tagv_mb_ff[1]; // @[el2_ifu_mem_ctl.scala 779:67]
  wire  _T_10079 = ~tagv_mb_ff[0]; // @[el2_ifu_mem_ctl.scala 779:86]
  wire  replace_way_mb_any_0 = _T_10077 | _T_10079; // @[el2_ifu_mem_ctl.scala 779:84]
  wire [1:0] _T_287 = scnd_miss_index_match ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire  _T_10082 = way_status_mb_ff & tagv_mb_ff[0]; // @[el2_ifu_mem_ctl.scala 780:50]
  wire  _T_10084 = _T_10082 & tagv_mb_ff[1]; // @[el2_ifu_mem_ctl.scala 780:66]
  wire  _T_10086 = ~tagv_mb_ff[1]; // @[el2_ifu_mem_ctl.scala 780:85]
  wire  _T_10088 = _T_10086 & tagv_mb_ff[0]; // @[el2_ifu_mem_ctl.scala 780:100]
  wire  replace_way_mb_any_1 = _T_10084 | _T_10088; // @[el2_ifu_mem_ctl.scala 780:83]
  wire [1:0] _T_288 = {replace_way_mb_any_1,replace_way_mb_any_0}; // @[Cat.scala 29:58]
  wire [1:0] _T_289 = _T_287 & _T_288; // @[el2_ifu_mem_ctl.scala 302:110]
  wire  _T_297 = ~scnd_miss_req_q; // @[el2_ifu_mem_ctl.scala 306:36]
  wire  _T_298 = miss_pending & _T_297; // @[el2_ifu_mem_ctl.scala 306:34]
  reg  reset_ic_ff; // @[el2_ifu_mem_ctl.scala 307:25]
  wire  _T_299 = reset_all_tags | reset_ic_ff; // @[el2_ifu_mem_ctl.scala 306:72]
  wire  reset_ic_in = _T_298 & _T_299; // @[el2_ifu_mem_ctl.scala 306:53]
  reg  fetch_uncacheable_ff; // @[el2_ifu_mem_ctl.scala 308:37]
  reg [25:0] miss_addr; // @[el2_ifu_mem_ctl.scala 316:23]
  wire  _T_313 = _T_2250 & flush_final_f; // @[el2_ifu_mem_ctl.scala 320:87]
  wire  _T_314 = ~_T_313; // @[el2_ifu_mem_ctl.scala 320:55]
  wire  _T_315 = io_ifc_fetch_req_bf & _T_314; // @[el2_ifu_mem_ctl.scala 320:53]
  wire  _T_2242 = ~_T_2237; // @[el2_ifu_mem_ctl.scala 461:46]
  wire  _T_2243 = _T_2235 & _T_2242; // @[el2_ifu_mem_ctl.scala 461:44]
  wire  stream_miss_f = _T_2243 & ifc_fetch_req_f; // @[el2_ifu_mem_ctl.scala 461:84]
  wire  _T_316 = ~stream_miss_f; // @[el2_ifu_mem_ctl.scala 320:106]
  wire  ifc_fetch_req_qual_bf = _T_315 & _T_316; // @[el2_ifu_mem_ctl.scala 320:104]
  reg  ifc_region_acc_fault_f; // @[el2_ifu_mem_ctl.scala 326:39]
  reg [2:0] bus_rd_addr_count; // @[Reg.scala 27:20]
  wire [28:0] ifu_ic_req_addr_f = {miss_addr,bus_rd_addr_count}; // @[Cat.scala 29:58]
  wire  _T_323 = _T_239 | _T_2235; // @[el2_ifu_mem_ctl.scala 328:55]
  wire  _T_326 = _T_323 & _T_56; // @[el2_ifu_mem_ctl.scala 328:82]
  wire  _T_2256 = ~ifu_bus_rid_ff[0]; // @[el2_ifu_mem_ctl.scala 466:55]
  wire [2:0] other_tag = {ifu_bus_rid_ff[2:1],_T_2256}; // @[Cat.scala 29:58]
  wire  _T_2257 = other_tag == 3'h0; // @[el2_ifu_mem_ctl.scala 467:81]
  wire  _T_2281 = _T_2257 & ic_miss_buff_data_valid[0]; // @[Mux.scala 27:72]
  wire  _T_2260 = other_tag == 3'h1; // @[el2_ifu_mem_ctl.scala 467:81]
  wire  _T_2282 = _T_2260 & ic_miss_buff_data_valid[1]; // @[Mux.scala 27:72]
  wire  _T_2289 = _T_2281 | _T_2282; // @[Mux.scala 27:72]
  wire  _T_2263 = other_tag == 3'h2; // @[el2_ifu_mem_ctl.scala 467:81]
  wire  _T_2283 = _T_2263 & ic_miss_buff_data_valid[2]; // @[Mux.scala 27:72]
  wire  _T_2290 = _T_2289 | _T_2283; // @[Mux.scala 27:72]
  wire  _T_2266 = other_tag == 3'h3; // @[el2_ifu_mem_ctl.scala 467:81]
  wire  _T_2284 = _T_2266 & ic_miss_buff_data_valid[3]; // @[Mux.scala 27:72]
  wire  _T_2291 = _T_2290 | _T_2284; // @[Mux.scala 27:72]
  wire  _T_2269 = other_tag == 3'h4; // @[el2_ifu_mem_ctl.scala 467:81]
  wire  _T_2285 = _T_2269 & ic_miss_buff_data_valid[4]; // @[Mux.scala 27:72]
  wire  _T_2292 = _T_2291 | _T_2285; // @[Mux.scala 27:72]
  wire  _T_2272 = other_tag == 3'h5; // @[el2_ifu_mem_ctl.scala 467:81]
  wire  _T_2286 = _T_2272 & ic_miss_buff_data_valid[5]; // @[Mux.scala 27:72]
  wire  _T_2293 = _T_2292 | _T_2286; // @[Mux.scala 27:72]
  wire  _T_2275 = other_tag == 3'h6; // @[el2_ifu_mem_ctl.scala 467:81]
  wire  _T_2287 = _T_2275 & ic_miss_buff_data_valid[6]; // @[Mux.scala 27:72]
  wire  _T_2294 = _T_2293 | _T_2287; // @[Mux.scala 27:72]
  wire  _T_2278 = other_tag == 3'h7; // @[el2_ifu_mem_ctl.scala 467:81]
  wire  _T_2288 = _T_2278 & ic_miss_buff_data_valid[7]; // @[Mux.scala 27:72]
  wire  second_half_available = _T_2294 | _T_2288; // @[Mux.scala 27:72]
  wire  write_ic_16_bytes = second_half_available & bus_ifu_wr_en_ff; // @[el2_ifu_mem_ctl.scala 468:46]
  wire  _T_330 = miss_pending & write_ic_16_bytes; // @[el2_ifu_mem_ctl.scala 332:35]
  wire  _T_332 = _T_330 & _T_17; // @[el2_ifu_mem_ctl.scala 332:55]
  reg  ic_act_miss_f_delayed; // @[el2_ifu_mem_ctl.scala 621:61]
  wire  _T_2618 = ic_act_miss_f_delayed & _T_2251; // @[el2_ifu_mem_ctl.scala 622:53]
  wire  reset_tag_valid_for_miss = _T_2618 & _T_17; // @[el2_ifu_mem_ctl.scala 622:84]
  wire  sel_mb_addr = _T_332 | reset_tag_valid_for_miss; // @[el2_ifu_mem_ctl.scala 332:79]
  wire [30:0] _T_336 = {imb_ff[30:5],ic_wr_addr_bits_hi_3,imb_ff[1:0]}; // @[Cat.scala 29:58]
  wire  _T_337 = ~sel_mb_addr; // @[el2_ifu_mem_ctl.scala 334:37]
  wire [30:0] _T_338 = sel_mb_addr ? _T_336 : 31'h0; // @[Mux.scala 27:72]
  wire [30:0] _T_339 = _T_337 ? io_ifc_fetch_addr_bf : 31'h0; // @[Mux.scala 27:72]
  wire [30:0] ifu_ic_rw_int_addr = _T_338 | _T_339; // @[Mux.scala 27:72]
  wire  _T_344 = _T_332 & last_beat; // @[el2_ifu_mem_ctl.scala 336:84]
  wire  _T_2612 = ~_T_2624; // @[el2_ifu_mem_ctl.scala 619:84]
  wire  _T_2613 = _T_100 & _T_2612; // @[el2_ifu_mem_ctl.scala 619:82]
  wire  bus_ifu_wr_en_ff_q = _T_2613 & write_ic_16_bytes; // @[el2_ifu_mem_ctl.scala 619:108]
  wire  sel_mb_status_addr = _T_344 & bus_ifu_wr_en_ff_q; // @[el2_ifu_mem_ctl.scala 336:96]
  wire [30:0] ifu_status_wr_addr = sel_mb_status_addr ? _T_336 : ifu_fetch_addr_int_f; // @[el2_ifu_mem_ctl.scala 337:31]
  reg [63:0] ifu_bus_rdata_ff; // @[Reg.scala 27:20]
  wire [7:0] _T_568 = {ifu_bus_rdata_ff[11],ifu_bus_rdata_ff[10],ifu_bus_rdata_ff[8],ifu_bus_rdata_ff[6],ifu_bus_rdata_ff[4],ifu_bus_rdata_ff[3],ifu_bus_rdata_ff[1],ifu_bus_rdata_ff[0]}; // @[el2_lib.scala 347:27]
  wire [16:0] _T_577 = {ifu_bus_rdata_ff[28],ifu_bus_rdata_ff[26],ifu_bus_rdata_ff[25],ifu_bus_rdata_ff[23],ifu_bus_rdata_ff[21],ifu_bus_rdata_ff[19],ifu_bus_rdata_ff[17],ifu_bus_rdata_ff[15],ifu_bus_rdata_ff[13],_T_568}; // @[el2_lib.scala 347:27]
  wire [8:0] _T_585 = {ifu_bus_rdata_ff[46],ifu_bus_rdata_ff[44],ifu_bus_rdata_ff[42],ifu_bus_rdata_ff[40],ifu_bus_rdata_ff[38],ifu_bus_rdata_ff[36],ifu_bus_rdata_ff[34],ifu_bus_rdata_ff[32],ifu_bus_rdata_ff[30]}; // @[el2_lib.scala 347:27]
  wire [17:0] _T_594 = {ifu_bus_rdata_ff[63],ifu_bus_rdata_ff[61],ifu_bus_rdata_ff[59],ifu_bus_rdata_ff[57],ifu_bus_rdata_ff[56],ifu_bus_rdata_ff[54],ifu_bus_rdata_ff[52],ifu_bus_rdata_ff[50],ifu_bus_rdata_ff[48],_T_585}; // @[el2_lib.scala 347:27]
  wire [34:0] _T_595 = {_T_594,_T_577}; // @[el2_lib.scala 347:27]
  wire  _T_596 = ^_T_595; // @[el2_lib.scala 347:34]
  wire [7:0] _T_603 = {ifu_bus_rdata_ff[12],ifu_bus_rdata_ff[10],ifu_bus_rdata_ff[9],ifu_bus_rdata_ff[6],ifu_bus_rdata_ff[5],ifu_bus_rdata_ff[3],ifu_bus_rdata_ff[2],ifu_bus_rdata_ff[0]}; // @[el2_lib.scala 347:44]
  wire [16:0] _T_612 = {ifu_bus_rdata_ff[28],ifu_bus_rdata_ff[27],ifu_bus_rdata_ff[25],ifu_bus_rdata_ff[24],ifu_bus_rdata_ff[21],ifu_bus_rdata_ff[20],ifu_bus_rdata_ff[17],ifu_bus_rdata_ff[16],ifu_bus_rdata_ff[13],_T_603}; // @[el2_lib.scala 347:44]
  wire [8:0] _T_620 = {ifu_bus_rdata_ff[47],ifu_bus_rdata_ff[44],ifu_bus_rdata_ff[43],ifu_bus_rdata_ff[40],ifu_bus_rdata_ff[39],ifu_bus_rdata_ff[36],ifu_bus_rdata_ff[35],ifu_bus_rdata_ff[32],ifu_bus_rdata_ff[31]}; // @[el2_lib.scala 347:44]
  wire [17:0] _T_629 = {ifu_bus_rdata_ff[63],ifu_bus_rdata_ff[62],ifu_bus_rdata_ff[59],ifu_bus_rdata_ff[58],ifu_bus_rdata_ff[56],ifu_bus_rdata_ff[55],ifu_bus_rdata_ff[52],ifu_bus_rdata_ff[51],ifu_bus_rdata_ff[48],_T_620}; // @[el2_lib.scala 347:44]
  wire [34:0] _T_630 = {_T_629,_T_612}; // @[el2_lib.scala 347:44]
  wire  _T_631 = ^_T_630; // @[el2_lib.scala 347:51]
  wire [7:0] _T_638 = {ifu_bus_rdata_ff[14],ifu_bus_rdata_ff[10],ifu_bus_rdata_ff[9],ifu_bus_rdata_ff[8],ifu_bus_rdata_ff[7],ifu_bus_rdata_ff[3],ifu_bus_rdata_ff[2],ifu_bus_rdata_ff[1]}; // @[el2_lib.scala 347:61]
  wire [16:0] _T_647 = {ifu_bus_rdata_ff[30],ifu_bus_rdata_ff[29],ifu_bus_rdata_ff[25],ifu_bus_rdata_ff[24],ifu_bus_rdata_ff[23],ifu_bus_rdata_ff[22],ifu_bus_rdata_ff[17],ifu_bus_rdata_ff[16],ifu_bus_rdata_ff[15],_T_638}; // @[el2_lib.scala 347:61]
  wire [8:0] _T_655 = {ifu_bus_rdata_ff[47],ifu_bus_rdata_ff[46],ifu_bus_rdata_ff[45],ifu_bus_rdata_ff[40],ifu_bus_rdata_ff[39],ifu_bus_rdata_ff[38],ifu_bus_rdata_ff[37],ifu_bus_rdata_ff[32],ifu_bus_rdata_ff[31]}; // @[el2_lib.scala 347:61]
  wire [17:0] _T_664 = {ifu_bus_rdata_ff[63],ifu_bus_rdata_ff[62],ifu_bus_rdata_ff[61],ifu_bus_rdata_ff[60],ifu_bus_rdata_ff[56],ifu_bus_rdata_ff[55],ifu_bus_rdata_ff[54],ifu_bus_rdata_ff[53],ifu_bus_rdata_ff[48],_T_655}; // @[el2_lib.scala 347:61]
  wire [34:0] _T_665 = {_T_664,_T_647}; // @[el2_lib.scala 347:61]
  wire  _T_666 = ^_T_665; // @[el2_lib.scala 347:68]
  wire [6:0] _T_672 = {ifu_bus_rdata_ff[10],ifu_bus_rdata_ff[9],ifu_bus_rdata_ff[8],ifu_bus_rdata_ff[7],ifu_bus_rdata_ff[6],ifu_bus_rdata_ff[5],ifu_bus_rdata_ff[4]}; // @[el2_lib.scala 347:78]
  wire [14:0] _T_680 = {ifu_bus_rdata_ff[25],ifu_bus_rdata_ff[24],ifu_bus_rdata_ff[23],ifu_bus_rdata_ff[22],ifu_bus_rdata_ff[21],ifu_bus_rdata_ff[20],ifu_bus_rdata_ff[19],ifu_bus_rdata_ff[18],_T_672}; // @[el2_lib.scala 347:78]
  wire [7:0] _T_687 = {ifu_bus_rdata_ff[40],ifu_bus_rdata_ff[39],ifu_bus_rdata_ff[38],ifu_bus_rdata_ff[37],ifu_bus_rdata_ff[36],ifu_bus_rdata_ff[35],ifu_bus_rdata_ff[34],ifu_bus_rdata_ff[33]}; // @[el2_lib.scala 347:78]
  wire [30:0] _T_696 = {ifu_bus_rdata_ff[56],ifu_bus_rdata_ff[55],ifu_bus_rdata_ff[54],ifu_bus_rdata_ff[53],ifu_bus_rdata_ff[52],ifu_bus_rdata_ff[51],ifu_bus_rdata_ff[50],ifu_bus_rdata_ff[49],_T_687,_T_680}; // @[el2_lib.scala 347:78]
  wire  _T_697 = ^_T_696; // @[el2_lib.scala 347:85]
  wire [6:0] _T_703 = {ifu_bus_rdata_ff[17],ifu_bus_rdata_ff[16],ifu_bus_rdata_ff[15],ifu_bus_rdata_ff[14],ifu_bus_rdata_ff[13],ifu_bus_rdata_ff[12],ifu_bus_rdata_ff[11]}; // @[el2_lib.scala 347:95]
  wire [14:0] _T_711 = {ifu_bus_rdata_ff[25],ifu_bus_rdata_ff[24],ifu_bus_rdata_ff[23],ifu_bus_rdata_ff[22],ifu_bus_rdata_ff[21],ifu_bus_rdata_ff[20],ifu_bus_rdata_ff[19],ifu_bus_rdata_ff[18],_T_703}; // @[el2_lib.scala 347:95]
  wire [7:0] _T_718 = {ifu_bus_rdata_ff[48],ifu_bus_rdata_ff[47],ifu_bus_rdata_ff[46],ifu_bus_rdata_ff[45],ifu_bus_rdata_ff[44],ifu_bus_rdata_ff[43],ifu_bus_rdata_ff[42],ifu_bus_rdata_ff[41]}; // @[el2_lib.scala 347:95]
  wire [30:0] _T_727 = {ifu_bus_rdata_ff[56],ifu_bus_rdata_ff[55],ifu_bus_rdata_ff[54],ifu_bus_rdata_ff[53],ifu_bus_rdata_ff[52],ifu_bus_rdata_ff[51],ifu_bus_rdata_ff[50],ifu_bus_rdata_ff[49],_T_718,_T_711}; // @[el2_lib.scala 347:95]
  wire  _T_728 = ^_T_727; // @[el2_lib.scala 347:102]
  wire [6:0] _T_734 = {ifu_bus_rdata_ff[32],ifu_bus_rdata_ff[31],ifu_bus_rdata_ff[30],ifu_bus_rdata_ff[29],ifu_bus_rdata_ff[28],ifu_bus_rdata_ff[27],ifu_bus_rdata_ff[26]}; // @[el2_lib.scala 347:112]
  wire [14:0] _T_742 = {ifu_bus_rdata_ff[40],ifu_bus_rdata_ff[39],ifu_bus_rdata_ff[38],ifu_bus_rdata_ff[37],ifu_bus_rdata_ff[36],ifu_bus_rdata_ff[35],ifu_bus_rdata_ff[34],ifu_bus_rdata_ff[33],_T_734}; // @[el2_lib.scala 347:112]
  wire [30:0] _T_758 = {ifu_bus_rdata_ff[56],ifu_bus_rdata_ff[55],ifu_bus_rdata_ff[54],ifu_bus_rdata_ff[53],ifu_bus_rdata_ff[52],ifu_bus_rdata_ff[51],ifu_bus_rdata_ff[50],ifu_bus_rdata_ff[49],_T_718,_T_742}; // @[el2_lib.scala 347:112]
  wire  _T_759 = ^_T_758; // @[el2_lib.scala 347:119]
  wire [6:0] _T_765 = {ifu_bus_rdata_ff[63],ifu_bus_rdata_ff[62],ifu_bus_rdata_ff[61],ifu_bus_rdata_ff[60],ifu_bus_rdata_ff[59],ifu_bus_rdata_ff[58],ifu_bus_rdata_ff[57]}; // @[el2_lib.scala 347:129]
  wire  _T_766 = ^_T_765; // @[el2_lib.scala 347:136]
  wire [2:0] _T_768 = {_T_728,_T_759,_T_766}; // @[Cat.scala 29:58]
  wire [3:0] _T_771 = {_T_596,_T_631,_T_666,_T_697}; // @[Cat.scala 29:58]
  wire [3:0] _T_2297 = {ifu_bus_rid_ff[2:1],_T_2256,1'h1}; // @[Cat.scala 29:58]
  wire  _T_2298 = _T_2297 == 4'h0; // @[el2_ifu_mem_ctl.scala 469:89]
  reg [31:0] ic_miss_buff_data_0; // @[Reg.scala 27:20]
  wire [31:0] _T_2345 = _T_2298 ? ic_miss_buff_data_0 : 32'h0; // @[Mux.scala 27:72]
  wire  _T_2301 = _T_2297 == 4'h1; // @[el2_ifu_mem_ctl.scala 469:89]
  reg [31:0] ic_miss_buff_data_1; // @[Reg.scala 27:20]
  wire [31:0] _T_2346 = _T_2301 ? ic_miss_buff_data_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2361 = _T_2345 | _T_2346; // @[Mux.scala 27:72]
  wire  _T_2304 = _T_2297 == 4'h2; // @[el2_ifu_mem_ctl.scala 469:89]
  reg [31:0] ic_miss_buff_data_2; // @[Reg.scala 27:20]
  wire [31:0] _T_2347 = _T_2304 ? ic_miss_buff_data_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2362 = _T_2361 | _T_2347; // @[Mux.scala 27:72]
  wire  _T_2307 = _T_2297 == 4'h3; // @[el2_ifu_mem_ctl.scala 469:89]
  reg [31:0] ic_miss_buff_data_3; // @[Reg.scala 27:20]
  wire [31:0] _T_2348 = _T_2307 ? ic_miss_buff_data_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2363 = _T_2362 | _T_2348; // @[Mux.scala 27:72]
  wire  _T_2310 = _T_2297 == 4'h4; // @[el2_ifu_mem_ctl.scala 469:89]
  reg [31:0] ic_miss_buff_data_4; // @[Reg.scala 27:20]
  wire [31:0] _T_2349 = _T_2310 ? ic_miss_buff_data_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2364 = _T_2363 | _T_2349; // @[Mux.scala 27:72]
  wire  _T_2313 = _T_2297 == 4'h5; // @[el2_ifu_mem_ctl.scala 469:89]
  reg [31:0] ic_miss_buff_data_5; // @[Reg.scala 27:20]
  wire [31:0] _T_2350 = _T_2313 ? ic_miss_buff_data_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2365 = _T_2364 | _T_2350; // @[Mux.scala 27:72]
  wire  _T_2316 = _T_2297 == 4'h6; // @[el2_ifu_mem_ctl.scala 469:89]
  reg [31:0] ic_miss_buff_data_6; // @[Reg.scala 27:20]
  wire [31:0] _T_2351 = _T_2316 ? ic_miss_buff_data_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2366 = _T_2365 | _T_2351; // @[Mux.scala 27:72]
  wire  _T_2319 = _T_2297 == 4'h7; // @[el2_ifu_mem_ctl.scala 469:89]
  reg [31:0] ic_miss_buff_data_7; // @[Reg.scala 27:20]
  wire [31:0] _T_2352 = _T_2319 ? ic_miss_buff_data_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2367 = _T_2366 | _T_2352; // @[Mux.scala 27:72]
  wire  _T_2322 = _T_2297 == 4'h8; // @[el2_ifu_mem_ctl.scala 469:89]
  reg [31:0] ic_miss_buff_data_8; // @[Reg.scala 27:20]
  wire [31:0] _T_2353 = _T_2322 ? ic_miss_buff_data_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2368 = _T_2367 | _T_2353; // @[Mux.scala 27:72]
  wire  _T_2325 = _T_2297 == 4'h9; // @[el2_ifu_mem_ctl.scala 469:89]
  reg [31:0] ic_miss_buff_data_9; // @[Reg.scala 27:20]
  wire [31:0] _T_2354 = _T_2325 ? ic_miss_buff_data_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2369 = _T_2368 | _T_2354; // @[Mux.scala 27:72]
  wire  _T_2328 = _T_2297 == 4'ha; // @[el2_ifu_mem_ctl.scala 469:89]
  reg [31:0] ic_miss_buff_data_10; // @[Reg.scala 27:20]
  wire [31:0] _T_2355 = _T_2328 ? ic_miss_buff_data_10 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2370 = _T_2369 | _T_2355; // @[Mux.scala 27:72]
  wire  _T_2331 = _T_2297 == 4'hb; // @[el2_ifu_mem_ctl.scala 469:89]
  reg [31:0] ic_miss_buff_data_11; // @[Reg.scala 27:20]
  wire [31:0] _T_2356 = _T_2331 ? ic_miss_buff_data_11 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2371 = _T_2370 | _T_2356; // @[Mux.scala 27:72]
  wire  _T_2334 = _T_2297 == 4'hc; // @[el2_ifu_mem_ctl.scala 469:89]
  reg [31:0] ic_miss_buff_data_12; // @[Reg.scala 27:20]
  wire [31:0] _T_2357 = _T_2334 ? ic_miss_buff_data_12 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2372 = _T_2371 | _T_2357; // @[Mux.scala 27:72]
  wire  _T_2337 = _T_2297 == 4'hd; // @[el2_ifu_mem_ctl.scala 469:89]
  reg [31:0] ic_miss_buff_data_13; // @[Reg.scala 27:20]
  wire [31:0] _T_2358 = _T_2337 ? ic_miss_buff_data_13 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2373 = _T_2372 | _T_2358; // @[Mux.scala 27:72]
  wire  _T_2340 = _T_2297 == 4'he; // @[el2_ifu_mem_ctl.scala 469:89]
  reg [31:0] ic_miss_buff_data_14; // @[Reg.scala 27:20]
  wire [31:0] _T_2359 = _T_2340 ? ic_miss_buff_data_14 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2374 = _T_2373 | _T_2359; // @[Mux.scala 27:72]
  wire  _T_2343 = _T_2297 == 4'hf; // @[el2_ifu_mem_ctl.scala 469:89]
  reg [31:0] ic_miss_buff_data_15; // @[Reg.scala 27:20]
  wire [31:0] _T_2360 = _T_2343 ? ic_miss_buff_data_15 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2375 = _T_2374 | _T_2360; // @[Mux.scala 27:72]
  wire [3:0] _T_2377 = {ifu_bus_rid_ff[2:1],_T_2256,1'h0}; // @[Cat.scala 29:58]
  wire  _T_2378 = _T_2377 == 4'h0; // @[el2_ifu_mem_ctl.scala 470:64]
  wire [31:0] _T_2401 = _T_2378 ? ic_miss_buff_data_0 : 32'h0; // @[Mux.scala 27:72]
  wire  _T_2381 = _T_2377 == 4'h1; // @[el2_ifu_mem_ctl.scala 470:64]
  wire [31:0] _T_2402 = _T_2381 ? ic_miss_buff_data_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2409 = _T_2401 | _T_2402; // @[Mux.scala 27:72]
  wire  _T_2384 = _T_2377 == 4'h2; // @[el2_ifu_mem_ctl.scala 470:64]
  wire [31:0] _T_2403 = _T_2384 ? ic_miss_buff_data_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2410 = _T_2409 | _T_2403; // @[Mux.scala 27:72]
  wire  _T_2387 = _T_2377 == 4'h3; // @[el2_ifu_mem_ctl.scala 470:64]
  wire [31:0] _T_2404 = _T_2387 ? ic_miss_buff_data_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2411 = _T_2410 | _T_2404; // @[Mux.scala 27:72]
  wire  _T_2390 = _T_2377 == 4'h4; // @[el2_ifu_mem_ctl.scala 470:64]
  wire [31:0] _T_2405 = _T_2390 ? ic_miss_buff_data_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2412 = _T_2411 | _T_2405; // @[Mux.scala 27:72]
  wire  _T_2393 = _T_2377 == 4'h5; // @[el2_ifu_mem_ctl.scala 470:64]
  wire [31:0] _T_2406 = _T_2393 ? ic_miss_buff_data_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2413 = _T_2412 | _T_2406; // @[Mux.scala 27:72]
  wire  _T_2396 = _T_2377 == 4'h6; // @[el2_ifu_mem_ctl.scala 470:64]
  wire [31:0] _T_2407 = _T_2396 ? ic_miss_buff_data_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2414 = _T_2413 | _T_2407; // @[Mux.scala 27:72]
  wire  _T_2399 = _T_2377 == 4'h7; // @[el2_ifu_mem_ctl.scala 470:64]
  wire [31:0] _T_2408 = _T_2399 ? ic_miss_buff_data_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2415 = _T_2414 | _T_2408; // @[Mux.scala 27:72]
  wire [63:0] ic_miss_buff_half = {_T_2375,_T_2415}; // @[Cat.scala 29:58]
  wire [7:0] _T_990 = {ic_miss_buff_half[11],ic_miss_buff_half[10],ic_miss_buff_half[8],ic_miss_buff_half[6],ic_miss_buff_half[4],ic_miss_buff_half[3],ic_miss_buff_half[1],ic_miss_buff_half[0]}; // @[el2_lib.scala 347:27]
  wire [16:0] _T_999 = {ic_miss_buff_half[28],ic_miss_buff_half[26],ic_miss_buff_half[25],ic_miss_buff_half[23],ic_miss_buff_half[21],ic_miss_buff_half[19],ic_miss_buff_half[17],ic_miss_buff_half[15],ic_miss_buff_half[13],_T_990}; // @[el2_lib.scala 347:27]
  wire [8:0] _T_1007 = {ic_miss_buff_half[46],ic_miss_buff_half[44],ic_miss_buff_half[42],ic_miss_buff_half[40],ic_miss_buff_half[38],ic_miss_buff_half[36],ic_miss_buff_half[34],ic_miss_buff_half[32],ic_miss_buff_half[30]}; // @[el2_lib.scala 347:27]
  wire [17:0] _T_1016 = {ic_miss_buff_half[63],ic_miss_buff_half[61],ic_miss_buff_half[59],ic_miss_buff_half[57],ic_miss_buff_half[56],ic_miss_buff_half[54],ic_miss_buff_half[52],ic_miss_buff_half[50],ic_miss_buff_half[48],_T_1007}; // @[el2_lib.scala 347:27]
  wire [34:0] _T_1017 = {_T_1016,_T_999}; // @[el2_lib.scala 347:27]
  wire  _T_1018 = ^_T_1017; // @[el2_lib.scala 347:34]
  wire [7:0] _T_1025 = {ic_miss_buff_half[12],ic_miss_buff_half[10],ic_miss_buff_half[9],ic_miss_buff_half[6],ic_miss_buff_half[5],ic_miss_buff_half[3],ic_miss_buff_half[2],ic_miss_buff_half[0]}; // @[el2_lib.scala 347:44]
  wire [16:0] _T_1034 = {ic_miss_buff_half[28],ic_miss_buff_half[27],ic_miss_buff_half[25],ic_miss_buff_half[24],ic_miss_buff_half[21],ic_miss_buff_half[20],ic_miss_buff_half[17],ic_miss_buff_half[16],ic_miss_buff_half[13],_T_1025}; // @[el2_lib.scala 347:44]
  wire [8:0] _T_1042 = {ic_miss_buff_half[47],ic_miss_buff_half[44],ic_miss_buff_half[43],ic_miss_buff_half[40],ic_miss_buff_half[39],ic_miss_buff_half[36],ic_miss_buff_half[35],ic_miss_buff_half[32],ic_miss_buff_half[31]}; // @[el2_lib.scala 347:44]
  wire [17:0] _T_1051 = {ic_miss_buff_half[63],ic_miss_buff_half[62],ic_miss_buff_half[59],ic_miss_buff_half[58],ic_miss_buff_half[56],ic_miss_buff_half[55],ic_miss_buff_half[52],ic_miss_buff_half[51],ic_miss_buff_half[48],_T_1042}; // @[el2_lib.scala 347:44]
  wire [34:0] _T_1052 = {_T_1051,_T_1034}; // @[el2_lib.scala 347:44]
  wire  _T_1053 = ^_T_1052; // @[el2_lib.scala 347:51]
  wire [7:0] _T_1060 = {ic_miss_buff_half[14],ic_miss_buff_half[10],ic_miss_buff_half[9],ic_miss_buff_half[8],ic_miss_buff_half[7],ic_miss_buff_half[3],ic_miss_buff_half[2],ic_miss_buff_half[1]}; // @[el2_lib.scala 347:61]
  wire [16:0] _T_1069 = {ic_miss_buff_half[30],ic_miss_buff_half[29],ic_miss_buff_half[25],ic_miss_buff_half[24],ic_miss_buff_half[23],ic_miss_buff_half[22],ic_miss_buff_half[17],ic_miss_buff_half[16],ic_miss_buff_half[15],_T_1060}; // @[el2_lib.scala 347:61]
  wire [8:0] _T_1077 = {ic_miss_buff_half[47],ic_miss_buff_half[46],ic_miss_buff_half[45],ic_miss_buff_half[40],ic_miss_buff_half[39],ic_miss_buff_half[38],ic_miss_buff_half[37],ic_miss_buff_half[32],ic_miss_buff_half[31]}; // @[el2_lib.scala 347:61]
  wire [17:0] _T_1086 = {ic_miss_buff_half[63],ic_miss_buff_half[62],ic_miss_buff_half[61],ic_miss_buff_half[60],ic_miss_buff_half[56],ic_miss_buff_half[55],ic_miss_buff_half[54],ic_miss_buff_half[53],ic_miss_buff_half[48],_T_1077}; // @[el2_lib.scala 347:61]
  wire [34:0] _T_1087 = {_T_1086,_T_1069}; // @[el2_lib.scala 347:61]
  wire  _T_1088 = ^_T_1087; // @[el2_lib.scala 347:68]
  wire [6:0] _T_1094 = {ic_miss_buff_half[10],ic_miss_buff_half[9],ic_miss_buff_half[8],ic_miss_buff_half[7],ic_miss_buff_half[6],ic_miss_buff_half[5],ic_miss_buff_half[4]}; // @[el2_lib.scala 347:78]
  wire [14:0] _T_1102 = {ic_miss_buff_half[25],ic_miss_buff_half[24],ic_miss_buff_half[23],ic_miss_buff_half[22],ic_miss_buff_half[21],ic_miss_buff_half[20],ic_miss_buff_half[19],ic_miss_buff_half[18],_T_1094}; // @[el2_lib.scala 347:78]
  wire [7:0] _T_1109 = {ic_miss_buff_half[40],ic_miss_buff_half[39],ic_miss_buff_half[38],ic_miss_buff_half[37],ic_miss_buff_half[36],ic_miss_buff_half[35],ic_miss_buff_half[34],ic_miss_buff_half[33]}; // @[el2_lib.scala 347:78]
  wire [30:0] _T_1118 = {ic_miss_buff_half[56],ic_miss_buff_half[55],ic_miss_buff_half[54],ic_miss_buff_half[53],ic_miss_buff_half[52],ic_miss_buff_half[51],ic_miss_buff_half[50],ic_miss_buff_half[49],_T_1109,_T_1102}; // @[el2_lib.scala 347:78]
  wire  _T_1119 = ^_T_1118; // @[el2_lib.scala 347:85]
  wire [6:0] _T_1125 = {ic_miss_buff_half[17],ic_miss_buff_half[16],ic_miss_buff_half[15],ic_miss_buff_half[14],ic_miss_buff_half[13],ic_miss_buff_half[12],ic_miss_buff_half[11]}; // @[el2_lib.scala 347:95]
  wire [14:0] _T_1133 = {ic_miss_buff_half[25],ic_miss_buff_half[24],ic_miss_buff_half[23],ic_miss_buff_half[22],ic_miss_buff_half[21],ic_miss_buff_half[20],ic_miss_buff_half[19],ic_miss_buff_half[18],_T_1125}; // @[el2_lib.scala 347:95]
  wire [7:0] _T_1140 = {ic_miss_buff_half[48],ic_miss_buff_half[47],ic_miss_buff_half[46],ic_miss_buff_half[45],ic_miss_buff_half[44],ic_miss_buff_half[43],ic_miss_buff_half[42],ic_miss_buff_half[41]}; // @[el2_lib.scala 347:95]
  wire [30:0] _T_1149 = {ic_miss_buff_half[56],ic_miss_buff_half[55],ic_miss_buff_half[54],ic_miss_buff_half[53],ic_miss_buff_half[52],ic_miss_buff_half[51],ic_miss_buff_half[50],ic_miss_buff_half[49],_T_1140,_T_1133}; // @[el2_lib.scala 347:95]
  wire  _T_1150 = ^_T_1149; // @[el2_lib.scala 347:102]
  wire [6:0] _T_1156 = {ic_miss_buff_half[32],ic_miss_buff_half[31],ic_miss_buff_half[30],ic_miss_buff_half[29],ic_miss_buff_half[28],ic_miss_buff_half[27],ic_miss_buff_half[26]}; // @[el2_lib.scala 347:112]
  wire [14:0] _T_1164 = {ic_miss_buff_half[40],ic_miss_buff_half[39],ic_miss_buff_half[38],ic_miss_buff_half[37],ic_miss_buff_half[36],ic_miss_buff_half[35],ic_miss_buff_half[34],ic_miss_buff_half[33],_T_1156}; // @[el2_lib.scala 347:112]
  wire [30:0] _T_1180 = {ic_miss_buff_half[56],ic_miss_buff_half[55],ic_miss_buff_half[54],ic_miss_buff_half[53],ic_miss_buff_half[52],ic_miss_buff_half[51],ic_miss_buff_half[50],ic_miss_buff_half[49],_T_1140,_T_1164}; // @[el2_lib.scala 347:112]
  wire  _T_1181 = ^_T_1180; // @[el2_lib.scala 347:119]
  wire [6:0] _T_1187 = {ic_miss_buff_half[63],ic_miss_buff_half[62],ic_miss_buff_half[61],ic_miss_buff_half[60],ic_miss_buff_half[59],ic_miss_buff_half[58],ic_miss_buff_half[57]}; // @[el2_lib.scala 347:129]
  wire  _T_1188 = ^_T_1187; // @[el2_lib.scala 347:136]
  wire [2:0] _T_1190 = {_T_1150,_T_1181,_T_1188}; // @[Cat.scala 29:58]
  wire [3:0] _T_1193 = {_T_1018,_T_1053,_T_1088,_T_1119}; // @[Cat.scala 29:58]
  wire [70:0] _T_1235 = {_T_596,_T_631,_T_666,_T_697,_T_728,_T_759,_T_766,ifu_bus_rdata_ff}; // @[Cat.scala 29:58]
  wire [70:0] _T_1234 = {_T_1018,_T_1053,_T_1088,_T_1119,_T_1150,_T_1181,_T_1188,_T_2375,_T_2415}; // @[Cat.scala 29:58]
  wire [141:0] _T_1236 = {_T_596,_T_631,_T_666,_T_697,_T_728,_T_759,_T_766,ifu_bus_rdata_ff,_T_1234}; // @[Cat.scala 29:58]
  wire [141:0] _T_1239 = {_T_1018,_T_1053,_T_1088,_T_1119,_T_1150,_T_1181,_T_1188,_T_2375,_T_2415,_T_1235}; // @[Cat.scala 29:58]
  wire [141:0] ic_wr_16bytes_data = ifu_bus_rid_ff[0] ? _T_1236 : _T_1239; // @[el2_ifu_mem_ctl.scala 360:28]
  wire  _T_1196 = |io_ic_eccerr; // @[el2_ifu_mem_ctl.scala 350:56]
  wire  _T_1197 = _T_1196 & ic_act_hit_f; // @[el2_ifu_mem_ctl.scala 350:83]
  wire [4:0] bypass_index = imb_ff[4:0]; // @[el2_ifu_mem_ctl.scala 416:28]
  wire  _T_1415 = bypass_index[4:2] == 3'h0; // @[el2_ifu_mem_ctl.scala 418:114]
  wire  bus_ifu_wr_en = _T_13 & miss_pending; // @[el2_ifu_mem_ctl.scala 617:35]
  wire  _T_1284 = io_ifu_axi_rid == 3'h0; // @[el2_ifu_mem_ctl.scala 401:91]
  wire  write_fill_data_0 = bus_ifu_wr_en & _T_1284; // @[el2_ifu_mem_ctl.scala 401:73]
  wire  _T_1341 = ~ic_act_miss_f; // @[el2_ifu_mem_ctl.scala 407:118]
  wire  _T_1342 = ic_miss_buff_data_valid[0] & _T_1341; // @[el2_ifu_mem_ctl.scala 407:116]
  wire  ic_miss_buff_data_valid_in_0 = write_fill_data_0 | _T_1342; // @[el2_ifu_mem_ctl.scala 407:88]
  wire  _T_1438 = _T_1415 & ic_miss_buff_data_valid_in_0; // @[Mux.scala 27:72]
  wire  _T_1418 = bypass_index[4:2] == 3'h1; // @[el2_ifu_mem_ctl.scala 418:114]
  wire  _T_1285 = io_ifu_axi_rid == 3'h1; // @[el2_ifu_mem_ctl.scala 401:91]
  wire  write_fill_data_1 = bus_ifu_wr_en & _T_1285; // @[el2_ifu_mem_ctl.scala 401:73]
  wire  _T_1345 = ic_miss_buff_data_valid[1] & _T_1341; // @[el2_ifu_mem_ctl.scala 407:116]
  wire  ic_miss_buff_data_valid_in_1 = write_fill_data_1 | _T_1345; // @[el2_ifu_mem_ctl.scala 407:88]
  wire  _T_1439 = _T_1418 & ic_miss_buff_data_valid_in_1; // @[Mux.scala 27:72]
  wire  _T_1446 = _T_1438 | _T_1439; // @[Mux.scala 27:72]
  wire  _T_1421 = bypass_index[4:2] == 3'h2; // @[el2_ifu_mem_ctl.scala 418:114]
  wire  _T_1286 = io_ifu_axi_rid == 3'h2; // @[el2_ifu_mem_ctl.scala 401:91]
  wire  write_fill_data_2 = bus_ifu_wr_en & _T_1286; // @[el2_ifu_mem_ctl.scala 401:73]
  wire  _T_1348 = ic_miss_buff_data_valid[2] & _T_1341; // @[el2_ifu_mem_ctl.scala 407:116]
  wire  ic_miss_buff_data_valid_in_2 = write_fill_data_2 | _T_1348; // @[el2_ifu_mem_ctl.scala 407:88]
  wire  _T_1440 = _T_1421 & ic_miss_buff_data_valid_in_2; // @[Mux.scala 27:72]
  wire  _T_1447 = _T_1446 | _T_1440; // @[Mux.scala 27:72]
  wire  _T_1424 = bypass_index[4:2] == 3'h3; // @[el2_ifu_mem_ctl.scala 418:114]
  wire  _T_1287 = io_ifu_axi_rid == 3'h3; // @[el2_ifu_mem_ctl.scala 401:91]
  wire  write_fill_data_3 = bus_ifu_wr_en & _T_1287; // @[el2_ifu_mem_ctl.scala 401:73]
  wire  _T_1351 = ic_miss_buff_data_valid[3] & _T_1341; // @[el2_ifu_mem_ctl.scala 407:116]
  wire  ic_miss_buff_data_valid_in_3 = write_fill_data_3 | _T_1351; // @[el2_ifu_mem_ctl.scala 407:88]
  wire  _T_1441 = _T_1424 & ic_miss_buff_data_valid_in_3; // @[Mux.scala 27:72]
  wire  _T_1448 = _T_1447 | _T_1441; // @[Mux.scala 27:72]
  wire  _T_1427 = bypass_index[4:2] == 3'h4; // @[el2_ifu_mem_ctl.scala 418:114]
  wire  _T_1288 = io_ifu_axi_rid == 3'h4; // @[el2_ifu_mem_ctl.scala 401:91]
  wire  write_fill_data_4 = bus_ifu_wr_en & _T_1288; // @[el2_ifu_mem_ctl.scala 401:73]
  wire  _T_1354 = ic_miss_buff_data_valid[4] & _T_1341; // @[el2_ifu_mem_ctl.scala 407:116]
  wire  ic_miss_buff_data_valid_in_4 = write_fill_data_4 | _T_1354; // @[el2_ifu_mem_ctl.scala 407:88]
  wire  _T_1442 = _T_1427 & ic_miss_buff_data_valid_in_4; // @[Mux.scala 27:72]
  wire  _T_1449 = _T_1448 | _T_1442; // @[Mux.scala 27:72]
  wire  _T_1430 = bypass_index[4:2] == 3'h5; // @[el2_ifu_mem_ctl.scala 418:114]
  wire  _T_1289 = io_ifu_axi_rid == 3'h5; // @[el2_ifu_mem_ctl.scala 401:91]
  wire  write_fill_data_5 = bus_ifu_wr_en & _T_1289; // @[el2_ifu_mem_ctl.scala 401:73]
  wire  _T_1357 = ic_miss_buff_data_valid[5] & _T_1341; // @[el2_ifu_mem_ctl.scala 407:116]
  wire  ic_miss_buff_data_valid_in_5 = write_fill_data_5 | _T_1357; // @[el2_ifu_mem_ctl.scala 407:88]
  wire  _T_1443 = _T_1430 & ic_miss_buff_data_valid_in_5; // @[Mux.scala 27:72]
  wire  _T_1450 = _T_1449 | _T_1443; // @[Mux.scala 27:72]
  wire  _T_1433 = bypass_index[4:2] == 3'h6; // @[el2_ifu_mem_ctl.scala 418:114]
  wire  _T_1290 = io_ifu_axi_rid == 3'h6; // @[el2_ifu_mem_ctl.scala 401:91]
  wire  write_fill_data_6 = bus_ifu_wr_en & _T_1290; // @[el2_ifu_mem_ctl.scala 401:73]
  wire  _T_1360 = ic_miss_buff_data_valid[6] & _T_1341; // @[el2_ifu_mem_ctl.scala 407:116]
  wire  ic_miss_buff_data_valid_in_6 = write_fill_data_6 | _T_1360; // @[el2_ifu_mem_ctl.scala 407:88]
  wire  _T_1444 = _T_1433 & ic_miss_buff_data_valid_in_6; // @[Mux.scala 27:72]
  wire  _T_1451 = _T_1450 | _T_1444; // @[Mux.scala 27:72]
  wire  _T_1436 = bypass_index[4:2] == 3'h7; // @[el2_ifu_mem_ctl.scala 418:114]
  wire  _T_1291 = io_ifu_axi_rid == 3'h7; // @[el2_ifu_mem_ctl.scala 401:91]
  wire  write_fill_data_7 = bus_ifu_wr_en & _T_1291; // @[el2_ifu_mem_ctl.scala 401:73]
  wire  _T_1363 = ic_miss_buff_data_valid[7] & _T_1341; // @[el2_ifu_mem_ctl.scala 407:116]
  wire  ic_miss_buff_data_valid_in_7 = write_fill_data_7 | _T_1363; // @[el2_ifu_mem_ctl.scala 407:88]
  wire  _T_1445 = _T_1436 & ic_miss_buff_data_valid_in_7; // @[Mux.scala 27:72]
  wire  bypass_valid_value_check = _T_1451 | _T_1445; // @[Mux.scala 27:72]
  wire  _T_1454 = ~bypass_index[1]; // @[el2_ifu_mem_ctl.scala 419:58]
  wire  _T_1455 = bypass_valid_value_check & _T_1454; // @[el2_ifu_mem_ctl.scala 419:56]
  wire  _T_1457 = ~bypass_index[0]; // @[el2_ifu_mem_ctl.scala 419:77]
  wire  _T_1458 = _T_1455 & _T_1457; // @[el2_ifu_mem_ctl.scala 419:75]
  wire  _T_1463 = _T_1455 & bypass_index[0]; // @[el2_ifu_mem_ctl.scala 420:75]
  wire  _T_1464 = _T_1458 | _T_1463; // @[el2_ifu_mem_ctl.scala 419:95]
  wire  _T_1466 = bypass_valid_value_check & bypass_index[1]; // @[el2_ifu_mem_ctl.scala 421:56]
  wire  _T_1469 = _T_1466 & _T_1457; // @[el2_ifu_mem_ctl.scala 421:74]
  wire  _T_1470 = _T_1464 | _T_1469; // @[el2_ifu_mem_ctl.scala 420:94]
  wire  _T_1474 = _T_1466 & bypass_index[0]; // @[el2_ifu_mem_ctl.scala 422:51]
  wire [2:0] bypass_index_5_3_inc = bypass_index[4:2] + 3'h1; // @[el2_ifu_mem_ctl.scala 417:70]
  wire  _T_1475 = bypass_index_5_3_inc == 3'h0; // @[el2_ifu_mem_ctl.scala 422:132]
  wire  _T_1491 = _T_1475 & ic_miss_buff_data_valid_in_0; // @[Mux.scala 27:72]
  wire  _T_1477 = bypass_index_5_3_inc == 3'h1; // @[el2_ifu_mem_ctl.scala 422:132]
  wire  _T_1492 = _T_1477 & ic_miss_buff_data_valid_in_1; // @[Mux.scala 27:72]
  wire  _T_1499 = _T_1491 | _T_1492; // @[Mux.scala 27:72]
  wire  _T_1479 = bypass_index_5_3_inc == 3'h2; // @[el2_ifu_mem_ctl.scala 422:132]
  wire  _T_1493 = _T_1479 & ic_miss_buff_data_valid_in_2; // @[Mux.scala 27:72]
  wire  _T_1500 = _T_1499 | _T_1493; // @[Mux.scala 27:72]
  wire  _T_1481 = bypass_index_5_3_inc == 3'h3; // @[el2_ifu_mem_ctl.scala 422:132]
  wire  _T_1494 = _T_1481 & ic_miss_buff_data_valid_in_3; // @[Mux.scala 27:72]
  wire  _T_1501 = _T_1500 | _T_1494; // @[Mux.scala 27:72]
  wire  _T_1483 = bypass_index_5_3_inc == 3'h4; // @[el2_ifu_mem_ctl.scala 422:132]
  wire  _T_1495 = _T_1483 & ic_miss_buff_data_valid_in_4; // @[Mux.scala 27:72]
  wire  _T_1502 = _T_1501 | _T_1495; // @[Mux.scala 27:72]
  wire  _T_1485 = bypass_index_5_3_inc == 3'h5; // @[el2_ifu_mem_ctl.scala 422:132]
  wire  _T_1496 = _T_1485 & ic_miss_buff_data_valid_in_5; // @[Mux.scala 27:72]
  wire  _T_1503 = _T_1502 | _T_1496; // @[Mux.scala 27:72]
  wire  _T_1487 = bypass_index_5_3_inc == 3'h6; // @[el2_ifu_mem_ctl.scala 422:132]
  wire  _T_1497 = _T_1487 & ic_miss_buff_data_valid_in_6; // @[Mux.scala 27:72]
  wire  _T_1504 = _T_1503 | _T_1497; // @[Mux.scala 27:72]
  wire  _T_1489 = bypass_index_5_3_inc == 3'h7; // @[el2_ifu_mem_ctl.scala 422:132]
  wire  _T_1498 = _T_1489 & ic_miss_buff_data_valid_in_7; // @[Mux.scala 27:72]
  wire  _T_1505 = _T_1504 | _T_1498; // @[Mux.scala 27:72]
  wire  _T_1507 = _T_1474 & _T_1505; // @[el2_ifu_mem_ctl.scala 422:69]
  wire  _T_1508 = _T_1470 | _T_1507; // @[el2_ifu_mem_ctl.scala 421:94]
  wire [4:0] _GEN_664 = {{2'd0}, bypass_index[4:2]}; // @[el2_ifu_mem_ctl.scala 423:95]
  wire  _T_1511 = _GEN_664 == 5'h1f; // @[el2_ifu_mem_ctl.scala 423:95]
  wire  _T_1512 = bypass_valid_value_check & _T_1511; // @[el2_ifu_mem_ctl.scala 423:56]
  wire  bypass_data_ready_in = _T_1508 | _T_1512; // @[el2_ifu_mem_ctl.scala 422:181]
  wire  _T_1513 = bypass_data_ready_in & crit_wd_byp_ok_ff; // @[el2_ifu_mem_ctl.scala 427:53]
  wire  _T_1514 = _T_1513 & uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 427:73]
  wire  _T_1516 = _T_1514 & _T_317; // @[el2_ifu_mem_ctl.scala 427:96]
  wire  _T_1518 = _T_1516 & _T_58; // @[el2_ifu_mem_ctl.scala 427:118]
  wire  _T_1520 = crit_wd_byp_ok_ff & _T_17; // @[el2_ifu_mem_ctl.scala 428:73]
  wire  _T_1522 = _T_1520 & _T_317; // @[el2_ifu_mem_ctl.scala 428:96]
  wire  _T_1524 = _T_1522 & _T_58; // @[el2_ifu_mem_ctl.scala 428:118]
  wire  _T_1525 = _T_1518 | _T_1524; // @[el2_ifu_mem_ctl.scala 427:143]
  reg  ic_crit_wd_rdy_new_ff; // @[el2_ifu_mem_ctl.scala 430:58]
  wire  _T_1526 = ic_crit_wd_rdy_new_ff & crit_wd_byp_ok_ff; // @[el2_ifu_mem_ctl.scala 429:54]
  wire  _T_1527 = ~fetch_req_icache_f; // @[el2_ifu_mem_ctl.scala 429:76]
  wire  _T_1528 = _T_1526 & _T_1527; // @[el2_ifu_mem_ctl.scala 429:74]
  wire  _T_1530 = _T_1528 & _T_317; // @[el2_ifu_mem_ctl.scala 429:96]
  wire  ic_crit_wd_rdy_new_in = _T_1525 | _T_1530; // @[el2_ifu_mem_ctl.scala 428:143]
  wire  ic_crit_wd_rdy = ic_crit_wd_rdy_new_in | ic_crit_wd_rdy_new_ff; // @[el2_ifu_mem_ctl.scala 627:43]
  wire  _T_1251 = ic_crit_wd_rdy | _T_2235; // @[el2_ifu_mem_ctl.scala 374:38]
  wire  _T_1253 = _T_1251 | _T_2251; // @[el2_ifu_mem_ctl.scala 374:64]
  wire  _T_1254 = ~_T_1253; // @[el2_ifu_mem_ctl.scala 374:21]
  wire  _T_1255 = ~fetch_req_iccm_f; // @[el2_ifu_mem_ctl.scala 374:98]
  wire  sel_ic_data = _T_1254 & _T_1255; // @[el2_ifu_mem_ctl.scala 374:96]
  wire  _T_2418 = io_ic_tag_perr & sel_ic_data; // @[el2_ifu_mem_ctl.scala 472:44]
  wire  _T_1624 = ifu_fetch_addr_int_f[1] & ifu_fetch_addr_int_f[0]; // @[el2_ifu_mem_ctl.scala 441:31]
  reg [7:0] ic_miss_buff_data_error; // @[el2_ifu_mem_ctl.scala 413:60]
  wire  _T_1568 = _T_1415 & ic_miss_buff_data_error[0]; // @[Mux.scala 27:72]
  wire  _T_1569 = _T_1418 & ic_miss_buff_data_error[1]; // @[Mux.scala 27:72]
  wire  _T_1576 = _T_1568 | _T_1569; // @[Mux.scala 27:72]
  wire  _T_1570 = _T_1421 & ic_miss_buff_data_error[2]; // @[Mux.scala 27:72]
  wire  _T_1577 = _T_1576 | _T_1570; // @[Mux.scala 27:72]
  wire  _T_1571 = _T_1424 & ic_miss_buff_data_error[3]; // @[Mux.scala 27:72]
  wire  _T_1578 = _T_1577 | _T_1571; // @[Mux.scala 27:72]
  wire  _T_1572 = _T_1427 & ic_miss_buff_data_error[4]; // @[Mux.scala 27:72]
  wire  _T_1579 = _T_1578 | _T_1572; // @[Mux.scala 27:72]
  wire  _T_1573 = _T_1430 & ic_miss_buff_data_error[5]; // @[Mux.scala 27:72]
  wire  _T_1580 = _T_1579 | _T_1573; // @[Mux.scala 27:72]
  wire  _T_1574 = _T_1433 & ic_miss_buff_data_error[6]; // @[Mux.scala 27:72]
  wire  _T_1581 = _T_1580 | _T_1574; // @[Mux.scala 27:72]
  wire  _T_1575 = _T_1436 & ic_miss_buff_data_error[7]; // @[Mux.scala 27:72]
  wire  ic_miss_buff_data_error_bypass = _T_1581 | _T_1575; // @[Mux.scala 27:72]
  wire  _T_1607 = _T_2168 & ic_miss_buff_data_error[0]; // @[Mux.scala 27:72]
  wire  _T_1608 = _T_2171 & ic_miss_buff_data_error[1]; // @[Mux.scala 27:72]
  wire  _T_1615 = _T_1607 | _T_1608; // @[Mux.scala 27:72]
  wire  _T_1609 = _T_2174 & ic_miss_buff_data_error[2]; // @[Mux.scala 27:72]
  wire  _T_1616 = _T_1615 | _T_1609; // @[Mux.scala 27:72]
  wire  _T_1610 = _T_2177 & ic_miss_buff_data_error[3]; // @[Mux.scala 27:72]
  wire  _T_1617 = _T_1616 | _T_1610; // @[Mux.scala 27:72]
  wire  _T_1611 = _T_2180 & ic_miss_buff_data_error[4]; // @[Mux.scala 27:72]
  wire  _T_1618 = _T_1617 | _T_1611; // @[Mux.scala 27:72]
  wire  _T_1612 = _T_2183 & ic_miss_buff_data_error[5]; // @[Mux.scala 27:72]
  wire  _T_1619 = _T_1618 | _T_1612; // @[Mux.scala 27:72]
  wire  _T_1613 = _T_2186 & ic_miss_buff_data_error[6]; // @[Mux.scala 27:72]
  wire  _T_1620 = _T_1619 | _T_1613; // @[Mux.scala 27:72]
  wire  _T_1614 = _T_2189 & ic_miss_buff_data_error[7]; // @[Mux.scala 27:72]
  wire  ic_miss_buff_data_error_bypass_inc = _T_1620 | _T_1614; // @[Mux.scala 27:72]
  wire  _T_1625 = ic_miss_buff_data_error_bypass | ic_miss_buff_data_error_bypass_inc; // @[el2_ifu_mem_ctl.scala 443:70]
  wire  ifu_byp_data_err_new = _T_1624 ? ic_miss_buff_data_error_bypass : _T_1625; // @[el2_ifu_mem_ctl.scala 441:56]
  wire  ifc_bus_acc_fault_f = ic_byp_hit_f & ifu_byp_data_err_new; // @[el2_ifu_mem_ctl.scala 385:42]
  wire  _T_2419 = ifc_region_acc_fault_final_f | ifc_bus_acc_fault_f; // @[el2_ifu_mem_ctl.scala 472:91]
  wire  _T_2420 = ~_T_2419; // @[el2_ifu_mem_ctl.scala 472:60]
  wire  ic_rd_parity_final_err = _T_2418 & _T_2420; // @[el2_ifu_mem_ctl.scala 472:58]
  reg  ic_debug_ict_array_sel_ff; // @[Reg.scala 27:20]
  reg  ic_tag_valid_out_1_0; // @[Reg.scala 27:20]
  wire  _T_9691 = _T_4485 ? 1'h0 : ic_tag_valid_out_1_0; // @[el2_ifu_mem_ctl.scala 754:10]
  reg  ic_tag_valid_out_1_1; // @[Reg.scala 27:20]
  wire  _T_9693 = _T_4489 ? 1'h0 : ic_tag_valid_out_1_1; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9946 = _T_9691 | _T_9693; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_2; // @[Reg.scala 27:20]
  wire  _T_9695 = _T_4493 ? 1'h0 : ic_tag_valid_out_1_2; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9947 = _T_9946 | _T_9695; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_3; // @[Reg.scala 27:20]
  wire  _T_9697 = _T_4497 ? 1'h0 : ic_tag_valid_out_1_3; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9948 = _T_9947 | _T_9697; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_4; // @[Reg.scala 27:20]
  wire  _T_9699 = _T_4501 ? 1'h0 : ic_tag_valid_out_1_4; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9949 = _T_9948 | _T_9699; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_5; // @[Reg.scala 27:20]
  wire  _T_9701 = _T_4505 ? 1'h0 : ic_tag_valid_out_1_5; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9950 = _T_9949 | _T_9701; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_6; // @[Reg.scala 27:20]
  wire  _T_9703 = _T_4509 ? 1'h0 : ic_tag_valid_out_1_6; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9951 = _T_9950 | _T_9703; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_7; // @[Reg.scala 27:20]
  wire  _T_9705 = _T_4513 ? 1'h0 : ic_tag_valid_out_1_7; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9952 = _T_9951 | _T_9705; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_8; // @[Reg.scala 27:20]
  wire  _T_9707 = _T_4517 ? 1'h0 : ic_tag_valid_out_1_8; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9953 = _T_9952 | _T_9707; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_9; // @[Reg.scala 27:20]
  wire  _T_9709 = _T_4521 ? 1'h0 : ic_tag_valid_out_1_9; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9954 = _T_9953 | _T_9709; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_10; // @[Reg.scala 27:20]
  wire  _T_9711 = _T_4525 ? 1'h0 : ic_tag_valid_out_1_10; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9955 = _T_9954 | _T_9711; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_11; // @[Reg.scala 27:20]
  wire  _T_9713 = _T_4529 ? 1'h0 : ic_tag_valid_out_1_11; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9956 = _T_9955 | _T_9713; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_12; // @[Reg.scala 27:20]
  wire  _T_9715 = _T_4533 ? 1'h0 : ic_tag_valid_out_1_12; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9957 = _T_9956 | _T_9715; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_13; // @[Reg.scala 27:20]
  wire  _T_9717 = _T_4537 ? 1'h0 : ic_tag_valid_out_1_13; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9958 = _T_9957 | _T_9717; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_14; // @[Reg.scala 27:20]
  wire  _T_9719 = _T_4541 ? 1'h0 : ic_tag_valid_out_1_14; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9959 = _T_9958 | _T_9719; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_15; // @[Reg.scala 27:20]
  wire  _T_9721 = _T_4545 ? 1'h0 : ic_tag_valid_out_1_15; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9960 = _T_9959 | _T_9721; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_16; // @[Reg.scala 27:20]
  wire  _T_9723 = _T_4549 ? 1'h0 : ic_tag_valid_out_1_16; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9961 = _T_9960 | _T_9723; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_17; // @[Reg.scala 27:20]
  wire  _T_9725 = _T_4553 ? 1'h0 : ic_tag_valid_out_1_17; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9962 = _T_9961 | _T_9725; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_18; // @[Reg.scala 27:20]
  wire  _T_9727 = _T_4557 ? 1'h0 : ic_tag_valid_out_1_18; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9963 = _T_9962 | _T_9727; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_19; // @[Reg.scala 27:20]
  wire  _T_9729 = _T_4561 ? 1'h0 : ic_tag_valid_out_1_19; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9964 = _T_9963 | _T_9729; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_20; // @[Reg.scala 27:20]
  wire  _T_9731 = _T_4565 ? 1'h0 : ic_tag_valid_out_1_20; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9965 = _T_9964 | _T_9731; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_21; // @[Reg.scala 27:20]
  wire  _T_9733 = _T_4569 ? 1'h0 : ic_tag_valid_out_1_21; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9966 = _T_9965 | _T_9733; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_22; // @[Reg.scala 27:20]
  wire  _T_9735 = _T_4573 ? 1'h0 : ic_tag_valid_out_1_22; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9967 = _T_9966 | _T_9735; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_23; // @[Reg.scala 27:20]
  wire  _T_9737 = _T_4577 ? 1'h0 : ic_tag_valid_out_1_23; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9968 = _T_9967 | _T_9737; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_24; // @[Reg.scala 27:20]
  wire  _T_9739 = _T_4581 ? 1'h0 : ic_tag_valid_out_1_24; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9969 = _T_9968 | _T_9739; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_25; // @[Reg.scala 27:20]
  wire  _T_9741 = _T_4585 ? 1'h0 : ic_tag_valid_out_1_25; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9970 = _T_9969 | _T_9741; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_26; // @[Reg.scala 27:20]
  wire  _T_9743 = _T_4589 ? 1'h0 : ic_tag_valid_out_1_26; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9971 = _T_9970 | _T_9743; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_27; // @[Reg.scala 27:20]
  wire  _T_9745 = _T_4593 ? 1'h0 : ic_tag_valid_out_1_27; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9972 = _T_9971 | _T_9745; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_28; // @[Reg.scala 27:20]
  wire  _T_9747 = _T_4597 ? 1'h0 : ic_tag_valid_out_1_28; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9973 = _T_9972 | _T_9747; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_29; // @[Reg.scala 27:20]
  wire  _T_9749 = _T_4601 ? 1'h0 : ic_tag_valid_out_1_29; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9974 = _T_9973 | _T_9749; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_30; // @[Reg.scala 27:20]
  wire  _T_9751 = _T_4605 ? 1'h0 : ic_tag_valid_out_1_30; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9975 = _T_9974 | _T_9751; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_31; // @[Reg.scala 27:20]
  wire  _T_9753 = _T_4609 ? 1'h0 : ic_tag_valid_out_1_31; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9976 = _T_9975 | _T_9753; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_32; // @[Reg.scala 27:20]
  wire  _T_9755 = _T_4613 ? 1'h0 : ic_tag_valid_out_1_32; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9977 = _T_9976 | _T_9755; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_33; // @[Reg.scala 27:20]
  wire  _T_9757 = _T_4617 ? 1'h0 : ic_tag_valid_out_1_33; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9978 = _T_9977 | _T_9757; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_34; // @[Reg.scala 27:20]
  wire  _T_9759 = _T_4621 ? 1'h0 : ic_tag_valid_out_1_34; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9979 = _T_9978 | _T_9759; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_35; // @[Reg.scala 27:20]
  wire  _T_9761 = _T_4625 ? 1'h0 : ic_tag_valid_out_1_35; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9980 = _T_9979 | _T_9761; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_36; // @[Reg.scala 27:20]
  wire  _T_9763 = _T_4629 ? 1'h0 : ic_tag_valid_out_1_36; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9981 = _T_9980 | _T_9763; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_37; // @[Reg.scala 27:20]
  wire  _T_9765 = _T_4633 ? 1'h0 : ic_tag_valid_out_1_37; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9982 = _T_9981 | _T_9765; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_38; // @[Reg.scala 27:20]
  wire  _T_9767 = _T_4637 ? 1'h0 : ic_tag_valid_out_1_38; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9983 = _T_9982 | _T_9767; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_39; // @[Reg.scala 27:20]
  wire  _T_9769 = _T_4641 ? 1'h0 : ic_tag_valid_out_1_39; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9984 = _T_9983 | _T_9769; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_40; // @[Reg.scala 27:20]
  wire  _T_9771 = _T_4645 ? 1'h0 : ic_tag_valid_out_1_40; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9985 = _T_9984 | _T_9771; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_41; // @[Reg.scala 27:20]
  wire  _T_9773 = _T_4649 ? 1'h0 : ic_tag_valid_out_1_41; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9986 = _T_9985 | _T_9773; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_42; // @[Reg.scala 27:20]
  wire  _T_9775 = _T_4653 ? 1'h0 : ic_tag_valid_out_1_42; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9987 = _T_9986 | _T_9775; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_43; // @[Reg.scala 27:20]
  wire  _T_9777 = _T_4657 ? 1'h0 : ic_tag_valid_out_1_43; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9988 = _T_9987 | _T_9777; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_44; // @[Reg.scala 27:20]
  wire  _T_9779 = _T_4661 ? 1'h0 : ic_tag_valid_out_1_44; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9989 = _T_9988 | _T_9779; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_45; // @[Reg.scala 27:20]
  wire  _T_9781 = _T_4665 ? 1'h0 : ic_tag_valid_out_1_45; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9990 = _T_9989 | _T_9781; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_46; // @[Reg.scala 27:20]
  wire  _T_9783 = _T_4669 ? 1'h0 : ic_tag_valid_out_1_46; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9991 = _T_9990 | _T_9783; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_47; // @[Reg.scala 27:20]
  wire  _T_9785 = _T_4673 ? 1'h0 : ic_tag_valid_out_1_47; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9992 = _T_9991 | _T_9785; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_48; // @[Reg.scala 27:20]
  wire  _T_9787 = _T_4677 ? 1'h0 : ic_tag_valid_out_1_48; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9993 = _T_9992 | _T_9787; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_49; // @[Reg.scala 27:20]
  wire  _T_9789 = _T_4681 ? 1'h0 : ic_tag_valid_out_1_49; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9994 = _T_9993 | _T_9789; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_50; // @[Reg.scala 27:20]
  wire  _T_9791 = _T_4685 ? 1'h0 : ic_tag_valid_out_1_50; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9995 = _T_9994 | _T_9791; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_51; // @[Reg.scala 27:20]
  wire  _T_9793 = _T_4689 ? 1'h0 : ic_tag_valid_out_1_51; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9996 = _T_9995 | _T_9793; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_52; // @[Reg.scala 27:20]
  wire  _T_9795 = _T_4693 ? 1'h0 : ic_tag_valid_out_1_52; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9997 = _T_9996 | _T_9795; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_53; // @[Reg.scala 27:20]
  wire  _T_9797 = _T_4697 ? 1'h0 : ic_tag_valid_out_1_53; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9998 = _T_9997 | _T_9797; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_54; // @[Reg.scala 27:20]
  wire  _T_9799 = _T_4701 ? 1'h0 : ic_tag_valid_out_1_54; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9999 = _T_9998 | _T_9799; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_55; // @[Reg.scala 27:20]
  wire  _T_9801 = _T_4705 ? 1'h0 : ic_tag_valid_out_1_55; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_10000 = _T_9999 | _T_9801; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_56; // @[Reg.scala 27:20]
  wire  _T_9803 = _T_4709 ? 1'h0 : ic_tag_valid_out_1_56; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_10001 = _T_10000 | _T_9803; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_57; // @[Reg.scala 27:20]
  wire  _T_9805 = _T_4713 ? 1'h0 : ic_tag_valid_out_1_57; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_10002 = _T_10001 | _T_9805; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_58; // @[Reg.scala 27:20]
  wire  _T_9807 = _T_4717 ? 1'h0 : ic_tag_valid_out_1_58; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_10003 = _T_10002 | _T_9807; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_59; // @[Reg.scala 27:20]
  wire  _T_9809 = _T_4721 ? 1'h0 : ic_tag_valid_out_1_59; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_10004 = _T_10003 | _T_9809; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_60; // @[Reg.scala 27:20]
  wire  _T_9811 = _T_4725 ? 1'h0 : ic_tag_valid_out_1_60; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_10005 = _T_10004 | _T_9811; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_61; // @[Reg.scala 27:20]
  wire  _T_9813 = _T_4729 ? 1'h0 : ic_tag_valid_out_1_61; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_10006 = _T_10005 | _T_9813; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_62; // @[Reg.scala 27:20]
  wire  _T_9815 = _T_4733 ? 1'h0 : ic_tag_valid_out_1_62; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_10007 = _T_10006 | _T_9815; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_63; // @[Reg.scala 27:20]
  wire  _T_9817 = _T_4737 ? 1'h0 : ic_tag_valid_out_1_63; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_10008 = _T_10007 | _T_9817; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_64; // @[Reg.scala 27:20]
  wire  _T_9819 = _T_4741 ? 1'h0 : ic_tag_valid_out_1_64; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_10009 = _T_10008 | _T_9819; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_65; // @[Reg.scala 27:20]
  wire  _T_9821 = _T_4745 ? 1'h0 : ic_tag_valid_out_1_65; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_10010 = _T_10009 | _T_9821; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_66; // @[Reg.scala 27:20]
  wire  _T_9823 = _T_4749 ? 1'h0 : ic_tag_valid_out_1_66; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_10011 = _T_10010 | _T_9823; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_67; // @[Reg.scala 27:20]
  wire  _T_9825 = _T_4753 ? 1'h0 : ic_tag_valid_out_1_67; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_10012 = _T_10011 | _T_9825; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_68; // @[Reg.scala 27:20]
  wire  _T_9827 = _T_4757 ? 1'h0 : ic_tag_valid_out_1_68; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_10013 = _T_10012 | _T_9827; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_69; // @[Reg.scala 27:20]
  wire  _T_9829 = _T_4761 ? 1'h0 : ic_tag_valid_out_1_69; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_10014 = _T_10013 | _T_9829; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_70; // @[Reg.scala 27:20]
  wire  _T_9831 = _T_4765 ? 1'h0 : ic_tag_valid_out_1_70; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_10015 = _T_10014 | _T_9831; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_71; // @[Reg.scala 27:20]
  wire  _T_9833 = _T_4769 ? 1'h0 : ic_tag_valid_out_1_71; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_10016 = _T_10015 | _T_9833; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_72; // @[Reg.scala 27:20]
  wire  _T_9835 = _T_4773 ? 1'h0 : ic_tag_valid_out_1_72; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_10017 = _T_10016 | _T_9835; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_73; // @[Reg.scala 27:20]
  wire  _T_9837 = _T_4777 ? 1'h0 : ic_tag_valid_out_1_73; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_10018 = _T_10017 | _T_9837; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_74; // @[Reg.scala 27:20]
  wire  _T_9839 = _T_4781 ? 1'h0 : ic_tag_valid_out_1_74; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_10019 = _T_10018 | _T_9839; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_75; // @[Reg.scala 27:20]
  wire  _T_9841 = _T_4785 ? 1'h0 : ic_tag_valid_out_1_75; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_10020 = _T_10019 | _T_9841; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_76; // @[Reg.scala 27:20]
  wire  _T_9843 = _T_4789 ? 1'h0 : ic_tag_valid_out_1_76; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_10021 = _T_10020 | _T_9843; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_77; // @[Reg.scala 27:20]
  wire  _T_9845 = _T_4793 ? 1'h0 : ic_tag_valid_out_1_77; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_10022 = _T_10021 | _T_9845; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_78; // @[Reg.scala 27:20]
  wire  _T_9847 = _T_4797 ? 1'h0 : ic_tag_valid_out_1_78; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_10023 = _T_10022 | _T_9847; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_79; // @[Reg.scala 27:20]
  wire  _T_9849 = _T_4801 ? 1'h0 : ic_tag_valid_out_1_79; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_10024 = _T_10023 | _T_9849; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_80; // @[Reg.scala 27:20]
  wire  _T_9851 = _T_4805 ? 1'h0 : ic_tag_valid_out_1_80; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_10025 = _T_10024 | _T_9851; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_81; // @[Reg.scala 27:20]
  wire  _T_9853 = _T_4809 ? 1'h0 : ic_tag_valid_out_1_81; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_10026 = _T_10025 | _T_9853; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_82; // @[Reg.scala 27:20]
  wire  _T_9855 = _T_4813 ? 1'h0 : ic_tag_valid_out_1_82; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_10027 = _T_10026 | _T_9855; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_83; // @[Reg.scala 27:20]
  wire  _T_9857 = _T_4817 ? 1'h0 : ic_tag_valid_out_1_83; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_10028 = _T_10027 | _T_9857; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_84; // @[Reg.scala 27:20]
  wire  _T_9859 = _T_4821 ? 1'h0 : ic_tag_valid_out_1_84; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_10029 = _T_10028 | _T_9859; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_85; // @[Reg.scala 27:20]
  wire  _T_9861 = _T_4825 ? 1'h0 : ic_tag_valid_out_1_85; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_10030 = _T_10029 | _T_9861; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_86; // @[Reg.scala 27:20]
  wire  _T_9863 = _T_4829 ? 1'h0 : ic_tag_valid_out_1_86; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_10031 = _T_10030 | _T_9863; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_87; // @[Reg.scala 27:20]
  wire  _T_9865 = _T_4833 ? 1'h0 : ic_tag_valid_out_1_87; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_10032 = _T_10031 | _T_9865; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_88; // @[Reg.scala 27:20]
  wire  _T_9867 = _T_4837 ? 1'h0 : ic_tag_valid_out_1_88; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_10033 = _T_10032 | _T_9867; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_89; // @[Reg.scala 27:20]
  wire  _T_9869 = _T_4841 ? 1'h0 : ic_tag_valid_out_1_89; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_10034 = _T_10033 | _T_9869; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_90; // @[Reg.scala 27:20]
  wire  _T_9871 = _T_4845 ? 1'h0 : ic_tag_valid_out_1_90; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_10035 = _T_10034 | _T_9871; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_91; // @[Reg.scala 27:20]
  wire  _T_9873 = _T_4849 ? 1'h0 : ic_tag_valid_out_1_91; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_10036 = _T_10035 | _T_9873; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_92; // @[Reg.scala 27:20]
  wire  _T_9875 = _T_4853 ? 1'h0 : ic_tag_valid_out_1_92; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_10037 = _T_10036 | _T_9875; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_93; // @[Reg.scala 27:20]
  wire  _T_9877 = _T_4857 ? 1'h0 : ic_tag_valid_out_1_93; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_10038 = _T_10037 | _T_9877; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_94; // @[Reg.scala 27:20]
  wire  _T_9879 = _T_4861 ? 1'h0 : ic_tag_valid_out_1_94; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_10039 = _T_10038 | _T_9879; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_95; // @[Reg.scala 27:20]
  wire  _T_9881 = _T_4865 ? 1'h0 : ic_tag_valid_out_1_95; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_10040 = _T_10039 | _T_9881; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_96; // @[Reg.scala 27:20]
  wire  _T_9883 = _T_4869 ? 1'h0 : ic_tag_valid_out_1_96; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_10041 = _T_10040 | _T_9883; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_97; // @[Reg.scala 27:20]
  wire  _T_9885 = _T_4873 ? 1'h0 : ic_tag_valid_out_1_97; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_10042 = _T_10041 | _T_9885; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_98; // @[Reg.scala 27:20]
  wire  _T_9887 = _T_4877 ? 1'h0 : ic_tag_valid_out_1_98; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_10043 = _T_10042 | _T_9887; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_99; // @[Reg.scala 27:20]
  wire  _T_9889 = _T_4881 ? 1'h0 : ic_tag_valid_out_1_99; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_10044 = _T_10043 | _T_9889; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_100; // @[Reg.scala 27:20]
  wire  _T_9891 = _T_4885 ? 1'h0 : ic_tag_valid_out_1_100; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_10045 = _T_10044 | _T_9891; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_101; // @[Reg.scala 27:20]
  wire  _T_9893 = _T_4889 ? 1'h0 : ic_tag_valid_out_1_101; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_10046 = _T_10045 | _T_9893; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_102; // @[Reg.scala 27:20]
  wire  _T_9895 = _T_4893 ? 1'h0 : ic_tag_valid_out_1_102; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_10047 = _T_10046 | _T_9895; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_103; // @[Reg.scala 27:20]
  wire  _T_9897 = _T_4897 ? 1'h0 : ic_tag_valid_out_1_103; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_10048 = _T_10047 | _T_9897; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_104; // @[Reg.scala 27:20]
  wire  _T_9899 = _T_4901 ? 1'h0 : ic_tag_valid_out_1_104; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_10049 = _T_10048 | _T_9899; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_105; // @[Reg.scala 27:20]
  wire  _T_9901 = _T_4905 ? 1'h0 : ic_tag_valid_out_1_105; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_10050 = _T_10049 | _T_9901; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_106; // @[Reg.scala 27:20]
  wire  _T_9903 = _T_4909 ? 1'h0 : ic_tag_valid_out_1_106; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_10051 = _T_10050 | _T_9903; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_107; // @[Reg.scala 27:20]
  wire  _T_9905 = _T_4913 ? 1'h0 : ic_tag_valid_out_1_107; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_10052 = _T_10051 | _T_9905; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_108; // @[Reg.scala 27:20]
  wire  _T_9907 = _T_4917 ? 1'h0 : ic_tag_valid_out_1_108; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_10053 = _T_10052 | _T_9907; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_109; // @[Reg.scala 27:20]
  wire  _T_9909 = _T_4921 ? 1'h0 : ic_tag_valid_out_1_109; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_10054 = _T_10053 | _T_9909; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_110; // @[Reg.scala 27:20]
  wire  _T_9911 = _T_4925 ? 1'h0 : ic_tag_valid_out_1_110; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_10055 = _T_10054 | _T_9911; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_111; // @[Reg.scala 27:20]
  wire  _T_9913 = _T_4929 ? 1'h0 : ic_tag_valid_out_1_111; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_10056 = _T_10055 | _T_9913; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_112; // @[Reg.scala 27:20]
  wire  _T_9915 = _T_4933 ? 1'h0 : ic_tag_valid_out_1_112; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_10057 = _T_10056 | _T_9915; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_113; // @[Reg.scala 27:20]
  wire  _T_9917 = _T_4937 ? 1'h0 : ic_tag_valid_out_1_113; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_10058 = _T_10057 | _T_9917; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_114; // @[Reg.scala 27:20]
  wire  _T_9919 = _T_4941 ? 1'h0 : ic_tag_valid_out_1_114; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_10059 = _T_10058 | _T_9919; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_115; // @[Reg.scala 27:20]
  wire  _T_9921 = _T_4945 ? 1'h0 : ic_tag_valid_out_1_115; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_10060 = _T_10059 | _T_9921; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_116; // @[Reg.scala 27:20]
  wire  _T_9923 = _T_4949 ? 1'h0 : ic_tag_valid_out_1_116; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_10061 = _T_10060 | _T_9923; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_117; // @[Reg.scala 27:20]
  wire  _T_9925 = _T_4953 ? 1'h0 : ic_tag_valid_out_1_117; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_10062 = _T_10061 | _T_9925; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_118; // @[Reg.scala 27:20]
  wire  _T_9927 = _T_4957 ? 1'h0 : ic_tag_valid_out_1_118; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_10063 = _T_10062 | _T_9927; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_119; // @[Reg.scala 27:20]
  wire  _T_9929 = _T_4961 ? 1'h0 : ic_tag_valid_out_1_119; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_10064 = _T_10063 | _T_9929; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_120; // @[Reg.scala 27:20]
  wire  _T_9931 = _T_4965 ? 1'h0 : ic_tag_valid_out_1_120; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_10065 = _T_10064 | _T_9931; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_121; // @[Reg.scala 27:20]
  wire  _T_9933 = _T_4969 ? 1'h0 : ic_tag_valid_out_1_121; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_10066 = _T_10065 | _T_9933; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_122; // @[Reg.scala 27:20]
  wire  _T_9935 = _T_4973 ? 1'h0 : ic_tag_valid_out_1_122; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_10067 = _T_10066 | _T_9935; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_123; // @[Reg.scala 27:20]
  wire  _T_9937 = _T_4977 ? 1'h0 : ic_tag_valid_out_1_123; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_10068 = _T_10067 | _T_9937; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_124; // @[Reg.scala 27:20]
  wire  _T_9939 = _T_4981 ? 1'h0 : ic_tag_valid_out_1_124; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_10069 = _T_10068 | _T_9939; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_125; // @[Reg.scala 27:20]
  wire  _T_9941 = _T_4985 ? 1'h0 : ic_tag_valid_out_1_125; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_10070 = _T_10069 | _T_9941; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_126; // @[Reg.scala 27:20]
  wire  _T_9943 = _T_4989 ? 1'h0 : ic_tag_valid_out_1_126; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_10071 = _T_10070 | _T_9943; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_1_127; // @[Reg.scala 27:20]
  wire  _T_9945 = _T_4993 ? 1'h0 : ic_tag_valid_out_1_127; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_10072 = _T_10071 | _T_9945; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_0; // @[Reg.scala 27:20]
  wire  _T_9308 = _T_4485 ? 1'h0 : ic_tag_valid_out_0_0; // @[el2_ifu_mem_ctl.scala 754:10]
  reg  ic_tag_valid_out_0_1; // @[Reg.scala 27:20]
  wire  _T_9310 = _T_4489 ? 1'h0 : ic_tag_valid_out_0_1; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9563 = _T_9308 | _T_9310; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_2; // @[Reg.scala 27:20]
  wire  _T_9312 = _T_4493 ? 1'h0 : ic_tag_valid_out_0_2; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9564 = _T_9563 | _T_9312; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_3; // @[Reg.scala 27:20]
  wire  _T_9314 = _T_4497 ? 1'h0 : ic_tag_valid_out_0_3; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9565 = _T_9564 | _T_9314; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_4; // @[Reg.scala 27:20]
  wire  _T_9316 = _T_4501 ? 1'h0 : ic_tag_valid_out_0_4; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9566 = _T_9565 | _T_9316; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_5; // @[Reg.scala 27:20]
  wire  _T_9318 = _T_4505 ? 1'h0 : ic_tag_valid_out_0_5; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9567 = _T_9566 | _T_9318; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_6; // @[Reg.scala 27:20]
  wire  _T_9320 = _T_4509 ? 1'h0 : ic_tag_valid_out_0_6; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9568 = _T_9567 | _T_9320; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_7; // @[Reg.scala 27:20]
  wire  _T_9322 = _T_4513 ? 1'h0 : ic_tag_valid_out_0_7; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9569 = _T_9568 | _T_9322; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_8; // @[Reg.scala 27:20]
  wire  _T_9324 = _T_4517 ? 1'h0 : ic_tag_valid_out_0_8; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9570 = _T_9569 | _T_9324; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_9; // @[Reg.scala 27:20]
  wire  _T_9326 = _T_4521 ? 1'h0 : ic_tag_valid_out_0_9; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9571 = _T_9570 | _T_9326; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_10; // @[Reg.scala 27:20]
  wire  _T_9328 = _T_4525 ? 1'h0 : ic_tag_valid_out_0_10; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9572 = _T_9571 | _T_9328; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_11; // @[Reg.scala 27:20]
  wire  _T_9330 = _T_4529 ? 1'h0 : ic_tag_valid_out_0_11; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9573 = _T_9572 | _T_9330; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_12; // @[Reg.scala 27:20]
  wire  _T_9332 = _T_4533 ? 1'h0 : ic_tag_valid_out_0_12; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9574 = _T_9573 | _T_9332; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_13; // @[Reg.scala 27:20]
  wire  _T_9334 = _T_4537 ? 1'h0 : ic_tag_valid_out_0_13; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9575 = _T_9574 | _T_9334; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_14; // @[Reg.scala 27:20]
  wire  _T_9336 = _T_4541 ? 1'h0 : ic_tag_valid_out_0_14; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9576 = _T_9575 | _T_9336; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_15; // @[Reg.scala 27:20]
  wire  _T_9338 = _T_4545 ? 1'h0 : ic_tag_valid_out_0_15; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9577 = _T_9576 | _T_9338; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_16; // @[Reg.scala 27:20]
  wire  _T_9340 = _T_4549 ? 1'h0 : ic_tag_valid_out_0_16; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9578 = _T_9577 | _T_9340; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_17; // @[Reg.scala 27:20]
  wire  _T_9342 = _T_4553 ? 1'h0 : ic_tag_valid_out_0_17; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9579 = _T_9578 | _T_9342; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_18; // @[Reg.scala 27:20]
  wire  _T_9344 = _T_4557 ? 1'h0 : ic_tag_valid_out_0_18; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9580 = _T_9579 | _T_9344; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_19; // @[Reg.scala 27:20]
  wire  _T_9346 = _T_4561 ? 1'h0 : ic_tag_valid_out_0_19; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9581 = _T_9580 | _T_9346; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_20; // @[Reg.scala 27:20]
  wire  _T_9348 = _T_4565 ? 1'h0 : ic_tag_valid_out_0_20; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9582 = _T_9581 | _T_9348; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_21; // @[Reg.scala 27:20]
  wire  _T_9350 = _T_4569 ? 1'h0 : ic_tag_valid_out_0_21; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9583 = _T_9582 | _T_9350; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_22; // @[Reg.scala 27:20]
  wire  _T_9352 = _T_4573 ? 1'h0 : ic_tag_valid_out_0_22; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9584 = _T_9583 | _T_9352; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_23; // @[Reg.scala 27:20]
  wire  _T_9354 = _T_4577 ? 1'h0 : ic_tag_valid_out_0_23; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9585 = _T_9584 | _T_9354; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_24; // @[Reg.scala 27:20]
  wire  _T_9356 = _T_4581 ? 1'h0 : ic_tag_valid_out_0_24; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9586 = _T_9585 | _T_9356; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_25; // @[Reg.scala 27:20]
  wire  _T_9358 = _T_4585 ? 1'h0 : ic_tag_valid_out_0_25; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9587 = _T_9586 | _T_9358; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_26; // @[Reg.scala 27:20]
  wire  _T_9360 = _T_4589 ? 1'h0 : ic_tag_valid_out_0_26; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9588 = _T_9587 | _T_9360; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_27; // @[Reg.scala 27:20]
  wire  _T_9362 = _T_4593 ? 1'h0 : ic_tag_valid_out_0_27; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9589 = _T_9588 | _T_9362; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_28; // @[Reg.scala 27:20]
  wire  _T_9364 = _T_4597 ? 1'h0 : ic_tag_valid_out_0_28; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9590 = _T_9589 | _T_9364; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_29; // @[Reg.scala 27:20]
  wire  _T_9366 = _T_4601 ? 1'h0 : ic_tag_valid_out_0_29; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9591 = _T_9590 | _T_9366; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_30; // @[Reg.scala 27:20]
  wire  _T_9368 = _T_4605 ? 1'h0 : ic_tag_valid_out_0_30; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9592 = _T_9591 | _T_9368; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_31; // @[Reg.scala 27:20]
  wire  _T_9370 = _T_4609 ? 1'h0 : ic_tag_valid_out_0_31; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9593 = _T_9592 | _T_9370; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_32; // @[Reg.scala 27:20]
  wire  _T_9372 = _T_4613 ? 1'h0 : ic_tag_valid_out_0_32; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9594 = _T_9593 | _T_9372; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_33; // @[Reg.scala 27:20]
  wire  _T_9374 = _T_4617 ? 1'h0 : ic_tag_valid_out_0_33; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9595 = _T_9594 | _T_9374; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_34; // @[Reg.scala 27:20]
  wire  _T_9376 = _T_4621 ? 1'h0 : ic_tag_valid_out_0_34; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9596 = _T_9595 | _T_9376; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_35; // @[Reg.scala 27:20]
  wire  _T_9378 = _T_4625 ? 1'h0 : ic_tag_valid_out_0_35; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9597 = _T_9596 | _T_9378; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_36; // @[Reg.scala 27:20]
  wire  _T_9380 = _T_4629 ? 1'h0 : ic_tag_valid_out_0_36; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9598 = _T_9597 | _T_9380; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_37; // @[Reg.scala 27:20]
  wire  _T_9382 = _T_4633 ? 1'h0 : ic_tag_valid_out_0_37; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9599 = _T_9598 | _T_9382; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_38; // @[Reg.scala 27:20]
  wire  _T_9384 = _T_4637 ? 1'h0 : ic_tag_valid_out_0_38; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9600 = _T_9599 | _T_9384; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_39; // @[Reg.scala 27:20]
  wire  _T_9386 = _T_4641 ? 1'h0 : ic_tag_valid_out_0_39; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9601 = _T_9600 | _T_9386; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_40; // @[Reg.scala 27:20]
  wire  _T_9388 = _T_4645 ? 1'h0 : ic_tag_valid_out_0_40; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9602 = _T_9601 | _T_9388; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_41; // @[Reg.scala 27:20]
  wire  _T_9390 = _T_4649 ? 1'h0 : ic_tag_valid_out_0_41; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9603 = _T_9602 | _T_9390; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_42; // @[Reg.scala 27:20]
  wire  _T_9392 = _T_4653 ? 1'h0 : ic_tag_valid_out_0_42; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9604 = _T_9603 | _T_9392; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_43; // @[Reg.scala 27:20]
  wire  _T_9394 = _T_4657 ? 1'h0 : ic_tag_valid_out_0_43; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9605 = _T_9604 | _T_9394; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_44; // @[Reg.scala 27:20]
  wire  _T_9396 = _T_4661 ? 1'h0 : ic_tag_valid_out_0_44; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9606 = _T_9605 | _T_9396; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_45; // @[Reg.scala 27:20]
  wire  _T_9398 = _T_4665 ? 1'h0 : ic_tag_valid_out_0_45; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9607 = _T_9606 | _T_9398; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_46; // @[Reg.scala 27:20]
  wire  _T_9400 = _T_4669 ? 1'h0 : ic_tag_valid_out_0_46; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9608 = _T_9607 | _T_9400; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_47; // @[Reg.scala 27:20]
  wire  _T_9402 = _T_4673 ? 1'h0 : ic_tag_valid_out_0_47; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9609 = _T_9608 | _T_9402; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_48; // @[Reg.scala 27:20]
  wire  _T_9404 = _T_4677 ? 1'h0 : ic_tag_valid_out_0_48; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9610 = _T_9609 | _T_9404; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_49; // @[Reg.scala 27:20]
  wire  _T_9406 = _T_4681 ? 1'h0 : ic_tag_valid_out_0_49; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9611 = _T_9610 | _T_9406; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_50; // @[Reg.scala 27:20]
  wire  _T_9408 = _T_4685 ? 1'h0 : ic_tag_valid_out_0_50; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9612 = _T_9611 | _T_9408; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_51; // @[Reg.scala 27:20]
  wire  _T_9410 = _T_4689 ? 1'h0 : ic_tag_valid_out_0_51; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9613 = _T_9612 | _T_9410; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_52; // @[Reg.scala 27:20]
  wire  _T_9412 = _T_4693 ? 1'h0 : ic_tag_valid_out_0_52; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9614 = _T_9613 | _T_9412; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_53; // @[Reg.scala 27:20]
  wire  _T_9414 = _T_4697 ? 1'h0 : ic_tag_valid_out_0_53; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9615 = _T_9614 | _T_9414; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_54; // @[Reg.scala 27:20]
  wire  _T_9416 = _T_4701 ? 1'h0 : ic_tag_valid_out_0_54; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9616 = _T_9615 | _T_9416; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_55; // @[Reg.scala 27:20]
  wire  _T_9418 = _T_4705 ? 1'h0 : ic_tag_valid_out_0_55; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9617 = _T_9616 | _T_9418; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_56; // @[Reg.scala 27:20]
  wire  _T_9420 = _T_4709 ? 1'h0 : ic_tag_valid_out_0_56; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9618 = _T_9617 | _T_9420; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_57; // @[Reg.scala 27:20]
  wire  _T_9422 = _T_4713 ? 1'h0 : ic_tag_valid_out_0_57; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9619 = _T_9618 | _T_9422; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_58; // @[Reg.scala 27:20]
  wire  _T_9424 = _T_4717 ? 1'h0 : ic_tag_valid_out_0_58; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9620 = _T_9619 | _T_9424; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_59; // @[Reg.scala 27:20]
  wire  _T_9426 = _T_4721 ? 1'h0 : ic_tag_valid_out_0_59; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9621 = _T_9620 | _T_9426; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_60; // @[Reg.scala 27:20]
  wire  _T_9428 = _T_4725 ? 1'h0 : ic_tag_valid_out_0_60; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9622 = _T_9621 | _T_9428; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_61; // @[Reg.scala 27:20]
  wire  _T_9430 = _T_4729 ? 1'h0 : ic_tag_valid_out_0_61; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9623 = _T_9622 | _T_9430; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_62; // @[Reg.scala 27:20]
  wire  _T_9432 = _T_4733 ? 1'h0 : ic_tag_valid_out_0_62; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9624 = _T_9623 | _T_9432; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_63; // @[Reg.scala 27:20]
  wire  _T_9434 = _T_4737 ? 1'h0 : ic_tag_valid_out_0_63; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9625 = _T_9624 | _T_9434; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_64; // @[Reg.scala 27:20]
  wire  _T_9436 = _T_4741 ? 1'h0 : ic_tag_valid_out_0_64; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9626 = _T_9625 | _T_9436; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_65; // @[Reg.scala 27:20]
  wire  _T_9438 = _T_4745 ? 1'h0 : ic_tag_valid_out_0_65; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9627 = _T_9626 | _T_9438; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_66; // @[Reg.scala 27:20]
  wire  _T_9440 = _T_4749 ? 1'h0 : ic_tag_valid_out_0_66; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9628 = _T_9627 | _T_9440; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_67; // @[Reg.scala 27:20]
  wire  _T_9442 = _T_4753 ? 1'h0 : ic_tag_valid_out_0_67; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9629 = _T_9628 | _T_9442; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_68; // @[Reg.scala 27:20]
  wire  _T_9444 = _T_4757 ? 1'h0 : ic_tag_valid_out_0_68; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9630 = _T_9629 | _T_9444; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_69; // @[Reg.scala 27:20]
  wire  _T_9446 = _T_4761 ? 1'h0 : ic_tag_valid_out_0_69; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9631 = _T_9630 | _T_9446; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_70; // @[Reg.scala 27:20]
  wire  _T_9448 = _T_4765 ? 1'h0 : ic_tag_valid_out_0_70; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9632 = _T_9631 | _T_9448; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_71; // @[Reg.scala 27:20]
  wire  _T_9450 = _T_4769 ? 1'h0 : ic_tag_valid_out_0_71; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9633 = _T_9632 | _T_9450; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_72; // @[Reg.scala 27:20]
  wire  _T_9452 = _T_4773 ? 1'h0 : ic_tag_valid_out_0_72; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9634 = _T_9633 | _T_9452; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_73; // @[Reg.scala 27:20]
  wire  _T_9454 = _T_4777 ? 1'h0 : ic_tag_valid_out_0_73; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9635 = _T_9634 | _T_9454; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_74; // @[Reg.scala 27:20]
  wire  _T_9456 = _T_4781 ? 1'h0 : ic_tag_valid_out_0_74; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9636 = _T_9635 | _T_9456; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_75; // @[Reg.scala 27:20]
  wire  _T_9458 = _T_4785 ? 1'h0 : ic_tag_valid_out_0_75; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9637 = _T_9636 | _T_9458; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_76; // @[Reg.scala 27:20]
  wire  _T_9460 = _T_4789 ? 1'h0 : ic_tag_valid_out_0_76; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9638 = _T_9637 | _T_9460; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_77; // @[Reg.scala 27:20]
  wire  _T_9462 = _T_4793 ? 1'h0 : ic_tag_valid_out_0_77; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9639 = _T_9638 | _T_9462; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_78; // @[Reg.scala 27:20]
  wire  _T_9464 = _T_4797 ? 1'h0 : ic_tag_valid_out_0_78; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9640 = _T_9639 | _T_9464; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_79; // @[Reg.scala 27:20]
  wire  _T_9466 = _T_4801 ? 1'h0 : ic_tag_valid_out_0_79; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9641 = _T_9640 | _T_9466; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_80; // @[Reg.scala 27:20]
  wire  _T_9468 = _T_4805 ? 1'h0 : ic_tag_valid_out_0_80; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9642 = _T_9641 | _T_9468; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_81; // @[Reg.scala 27:20]
  wire  _T_9470 = _T_4809 ? 1'h0 : ic_tag_valid_out_0_81; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9643 = _T_9642 | _T_9470; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_82; // @[Reg.scala 27:20]
  wire  _T_9472 = _T_4813 ? 1'h0 : ic_tag_valid_out_0_82; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9644 = _T_9643 | _T_9472; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_83; // @[Reg.scala 27:20]
  wire  _T_9474 = _T_4817 ? 1'h0 : ic_tag_valid_out_0_83; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9645 = _T_9644 | _T_9474; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_84; // @[Reg.scala 27:20]
  wire  _T_9476 = _T_4821 ? 1'h0 : ic_tag_valid_out_0_84; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9646 = _T_9645 | _T_9476; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_85; // @[Reg.scala 27:20]
  wire  _T_9478 = _T_4825 ? 1'h0 : ic_tag_valid_out_0_85; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9647 = _T_9646 | _T_9478; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_86; // @[Reg.scala 27:20]
  wire  _T_9480 = _T_4829 ? 1'h0 : ic_tag_valid_out_0_86; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9648 = _T_9647 | _T_9480; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_87; // @[Reg.scala 27:20]
  wire  _T_9482 = _T_4833 ? 1'h0 : ic_tag_valid_out_0_87; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9649 = _T_9648 | _T_9482; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_88; // @[Reg.scala 27:20]
  wire  _T_9484 = _T_4837 ? 1'h0 : ic_tag_valid_out_0_88; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9650 = _T_9649 | _T_9484; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_89; // @[Reg.scala 27:20]
  wire  _T_9486 = _T_4841 ? 1'h0 : ic_tag_valid_out_0_89; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9651 = _T_9650 | _T_9486; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_90; // @[Reg.scala 27:20]
  wire  _T_9488 = _T_4845 ? 1'h0 : ic_tag_valid_out_0_90; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9652 = _T_9651 | _T_9488; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_91; // @[Reg.scala 27:20]
  wire  _T_9490 = _T_4849 ? 1'h0 : ic_tag_valid_out_0_91; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9653 = _T_9652 | _T_9490; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_92; // @[Reg.scala 27:20]
  wire  _T_9492 = _T_4853 ? 1'h0 : ic_tag_valid_out_0_92; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9654 = _T_9653 | _T_9492; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_93; // @[Reg.scala 27:20]
  wire  _T_9494 = _T_4857 ? 1'h0 : ic_tag_valid_out_0_93; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9655 = _T_9654 | _T_9494; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_94; // @[Reg.scala 27:20]
  wire  _T_9496 = _T_4861 ? 1'h0 : ic_tag_valid_out_0_94; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9656 = _T_9655 | _T_9496; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_95; // @[Reg.scala 27:20]
  wire  _T_9498 = _T_4865 ? 1'h0 : ic_tag_valid_out_0_95; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9657 = _T_9656 | _T_9498; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_96; // @[Reg.scala 27:20]
  wire  _T_9500 = _T_4869 ? 1'h0 : ic_tag_valid_out_0_96; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9658 = _T_9657 | _T_9500; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_97; // @[Reg.scala 27:20]
  wire  _T_9502 = _T_4873 ? 1'h0 : ic_tag_valid_out_0_97; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9659 = _T_9658 | _T_9502; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_98; // @[Reg.scala 27:20]
  wire  _T_9504 = _T_4877 ? 1'h0 : ic_tag_valid_out_0_98; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9660 = _T_9659 | _T_9504; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_99; // @[Reg.scala 27:20]
  wire  _T_9506 = _T_4881 ? 1'h0 : ic_tag_valid_out_0_99; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9661 = _T_9660 | _T_9506; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_100; // @[Reg.scala 27:20]
  wire  _T_9508 = _T_4885 ? 1'h0 : ic_tag_valid_out_0_100; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9662 = _T_9661 | _T_9508; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_101; // @[Reg.scala 27:20]
  wire  _T_9510 = _T_4889 ? 1'h0 : ic_tag_valid_out_0_101; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9663 = _T_9662 | _T_9510; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_102; // @[Reg.scala 27:20]
  wire  _T_9512 = _T_4893 ? 1'h0 : ic_tag_valid_out_0_102; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9664 = _T_9663 | _T_9512; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_103; // @[Reg.scala 27:20]
  wire  _T_9514 = _T_4897 ? 1'h0 : ic_tag_valid_out_0_103; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9665 = _T_9664 | _T_9514; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_104; // @[Reg.scala 27:20]
  wire  _T_9516 = _T_4901 ? 1'h0 : ic_tag_valid_out_0_104; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9666 = _T_9665 | _T_9516; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_105; // @[Reg.scala 27:20]
  wire  _T_9518 = _T_4905 ? 1'h0 : ic_tag_valid_out_0_105; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9667 = _T_9666 | _T_9518; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_106; // @[Reg.scala 27:20]
  wire  _T_9520 = _T_4909 ? 1'h0 : ic_tag_valid_out_0_106; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9668 = _T_9667 | _T_9520; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_107; // @[Reg.scala 27:20]
  wire  _T_9522 = _T_4913 ? 1'h0 : ic_tag_valid_out_0_107; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9669 = _T_9668 | _T_9522; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_108; // @[Reg.scala 27:20]
  wire  _T_9524 = _T_4917 ? 1'h0 : ic_tag_valid_out_0_108; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9670 = _T_9669 | _T_9524; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_109; // @[Reg.scala 27:20]
  wire  _T_9526 = _T_4921 ? 1'h0 : ic_tag_valid_out_0_109; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9671 = _T_9670 | _T_9526; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_110; // @[Reg.scala 27:20]
  wire  _T_9528 = _T_4925 ? 1'h0 : ic_tag_valid_out_0_110; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9672 = _T_9671 | _T_9528; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_111; // @[Reg.scala 27:20]
  wire  _T_9530 = _T_4929 ? 1'h0 : ic_tag_valid_out_0_111; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9673 = _T_9672 | _T_9530; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_112; // @[Reg.scala 27:20]
  wire  _T_9532 = _T_4933 ? 1'h0 : ic_tag_valid_out_0_112; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9674 = _T_9673 | _T_9532; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_113; // @[Reg.scala 27:20]
  wire  _T_9534 = _T_4937 ? 1'h0 : ic_tag_valid_out_0_113; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9675 = _T_9674 | _T_9534; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_114; // @[Reg.scala 27:20]
  wire  _T_9536 = _T_4941 ? 1'h0 : ic_tag_valid_out_0_114; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9676 = _T_9675 | _T_9536; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_115; // @[Reg.scala 27:20]
  wire  _T_9538 = _T_4945 ? 1'h0 : ic_tag_valid_out_0_115; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9677 = _T_9676 | _T_9538; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_116; // @[Reg.scala 27:20]
  wire  _T_9540 = _T_4949 ? 1'h0 : ic_tag_valid_out_0_116; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9678 = _T_9677 | _T_9540; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_117; // @[Reg.scala 27:20]
  wire  _T_9542 = _T_4953 ? 1'h0 : ic_tag_valid_out_0_117; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9679 = _T_9678 | _T_9542; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_118; // @[Reg.scala 27:20]
  wire  _T_9544 = _T_4957 ? 1'h0 : ic_tag_valid_out_0_118; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9680 = _T_9679 | _T_9544; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_119; // @[Reg.scala 27:20]
  wire  _T_9546 = _T_4961 ? 1'h0 : ic_tag_valid_out_0_119; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9681 = _T_9680 | _T_9546; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_120; // @[Reg.scala 27:20]
  wire  _T_9548 = _T_4965 ? 1'h0 : ic_tag_valid_out_0_120; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9682 = _T_9681 | _T_9548; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_121; // @[Reg.scala 27:20]
  wire  _T_9550 = _T_4969 ? 1'h0 : ic_tag_valid_out_0_121; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9683 = _T_9682 | _T_9550; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_122; // @[Reg.scala 27:20]
  wire  _T_9552 = _T_4973 ? 1'h0 : ic_tag_valid_out_0_122; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9684 = _T_9683 | _T_9552; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_123; // @[Reg.scala 27:20]
  wire  _T_9554 = _T_4977 ? 1'h0 : ic_tag_valid_out_0_123; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9685 = _T_9684 | _T_9554; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_124; // @[Reg.scala 27:20]
  wire  _T_9556 = _T_4981 ? 1'h0 : ic_tag_valid_out_0_124; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9686 = _T_9685 | _T_9556; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_125; // @[Reg.scala 27:20]
  wire  _T_9558 = _T_4985 ? 1'h0 : ic_tag_valid_out_0_125; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9687 = _T_9686 | _T_9558; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_126; // @[Reg.scala 27:20]
  wire  _T_9560 = _T_4989 ? 1'h0 : ic_tag_valid_out_0_126; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9688 = _T_9687 | _T_9560; // @[el2_ifu_mem_ctl.scala 754:91]
  reg  ic_tag_valid_out_0_127; // @[Reg.scala 27:20]
  wire  _T_9562 = _T_4993 ? 1'h0 : ic_tag_valid_out_0_127; // @[el2_ifu_mem_ctl.scala 754:10]
  wire  _T_9689 = _T_9688 | _T_9562; // @[el2_ifu_mem_ctl.scala 754:91]
  wire [1:0] ic_tag_valid_unq = {_T_10072,_T_9689}; // @[Cat.scala 29:58]
  reg [1:0] ic_debug_way_ff; // @[Reg.scala 27:20]
  reg  ic_debug_rd_en_ff; // @[el2_ifu_mem_ctl.scala 827:54]
  wire [1:0] _T_10111 = ic_debug_rd_en_ff ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [1:0] _T_10112 = ic_debug_way_ff & _T_10111; // @[el2_ifu_mem_ctl.scala 808:67]
  wire [1:0] _T_10113 = ic_tag_valid_unq & _T_10112; // @[el2_ifu_mem_ctl.scala 808:48]
  wire  ic_debug_tag_val_rd_out = |_T_10113; // @[el2_ifu_mem_ctl.scala 808:115]
  wire [65:0] _T_1208 = {2'h0,io_ictag_debug_rd_data[25:21],32'h0,io_ictag_debug_rd_data[20:0],1'h0,way_status,3'h0,ic_debug_tag_val_rd_out}; // @[Cat.scala 29:58]
  reg [70:0] _T_1209; // @[el2_ifu_mem_ctl.scala 356:37]
  wire  ifu_wr_cumulative_err = ifu_wr_cumulative_err_data & _T_2553; // @[el2_ifu_mem_ctl.scala 368:80]
  wire  _T_1249 = ~ifu_byp_data_err_new; // @[el2_ifu_mem_ctl.scala 373:98]
  wire  sel_byp_data = _T_1253 & _T_1249; // @[el2_ifu_mem_ctl.scala 373:96]
  wire [63:0] _T_1260 = fetch_req_iccm_f ? 64'hffffffffffffffff : 64'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_1261 = _T_1260 & io_iccm_rd_data; // @[el2_ifu_mem_ctl.scala 380:64]
  wire [63:0] _T_1263 = sel_byp_data ? 64'hffffffffffffffff : 64'h0; // @[Bitwise.scala 72:12]
  wire  _T_2115 = ~ifu_fetch_addr_int_f[0]; // @[el2_ifu_mem_ctl.scala 449:31]
  wire [3:0] byp_fetch_index_inc_0 = {byp_fetch_index_inc,1'h0}; // @[Cat.scala 29:58]
  wire  _T_1629 = byp_fetch_index_inc_0 == 4'h0; // @[el2_ifu_mem_ctl.scala 446:73]
  wire [15:0] _T_1677 = _T_1629 ? ic_miss_buff_data_0[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire  _T_1632 = byp_fetch_index_inc_0 == 4'h1; // @[el2_ifu_mem_ctl.scala 446:73]
  wire [15:0] _T_1678 = _T_1632 ? ic_miss_buff_data_1[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1693 = _T_1677 | _T_1678; // @[Mux.scala 27:72]
  wire  _T_1635 = byp_fetch_index_inc_0 == 4'h2; // @[el2_ifu_mem_ctl.scala 446:73]
  wire [15:0] _T_1679 = _T_1635 ? ic_miss_buff_data_2[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1694 = _T_1693 | _T_1679; // @[Mux.scala 27:72]
  wire  _T_1638 = byp_fetch_index_inc_0 == 4'h3; // @[el2_ifu_mem_ctl.scala 446:73]
  wire [15:0] _T_1680 = _T_1638 ? ic_miss_buff_data_3[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1695 = _T_1694 | _T_1680; // @[Mux.scala 27:72]
  wire  _T_1641 = byp_fetch_index_inc_0 == 4'h4; // @[el2_ifu_mem_ctl.scala 446:73]
  wire [15:0] _T_1681 = _T_1641 ? ic_miss_buff_data_4[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1696 = _T_1695 | _T_1681; // @[Mux.scala 27:72]
  wire  _T_1644 = byp_fetch_index_inc_0 == 4'h5; // @[el2_ifu_mem_ctl.scala 446:73]
  wire [15:0] _T_1682 = _T_1644 ? ic_miss_buff_data_5[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1697 = _T_1696 | _T_1682; // @[Mux.scala 27:72]
  wire  _T_1647 = byp_fetch_index_inc_0 == 4'h6; // @[el2_ifu_mem_ctl.scala 446:73]
  wire [15:0] _T_1683 = _T_1647 ? ic_miss_buff_data_6[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1698 = _T_1697 | _T_1683; // @[Mux.scala 27:72]
  wire  _T_1650 = byp_fetch_index_inc_0 == 4'h7; // @[el2_ifu_mem_ctl.scala 446:73]
  wire [15:0] _T_1684 = _T_1650 ? ic_miss_buff_data_7[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1699 = _T_1698 | _T_1684; // @[Mux.scala 27:72]
  wire  _T_1653 = byp_fetch_index_inc_0 == 4'h8; // @[el2_ifu_mem_ctl.scala 446:73]
  wire [15:0] _T_1685 = _T_1653 ? ic_miss_buff_data_8[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1700 = _T_1699 | _T_1685; // @[Mux.scala 27:72]
  wire  _T_1656 = byp_fetch_index_inc_0 == 4'h9; // @[el2_ifu_mem_ctl.scala 446:73]
  wire [15:0] _T_1686 = _T_1656 ? ic_miss_buff_data_9[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1701 = _T_1700 | _T_1686; // @[Mux.scala 27:72]
  wire  _T_1659 = byp_fetch_index_inc_0 == 4'ha; // @[el2_ifu_mem_ctl.scala 446:73]
  wire [15:0] _T_1687 = _T_1659 ? ic_miss_buff_data_10[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1702 = _T_1701 | _T_1687; // @[Mux.scala 27:72]
  wire  _T_1662 = byp_fetch_index_inc_0 == 4'hb; // @[el2_ifu_mem_ctl.scala 446:73]
  wire [15:0] _T_1688 = _T_1662 ? ic_miss_buff_data_11[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1703 = _T_1702 | _T_1688; // @[Mux.scala 27:72]
  wire  _T_1665 = byp_fetch_index_inc_0 == 4'hc; // @[el2_ifu_mem_ctl.scala 446:73]
  wire [15:0] _T_1689 = _T_1665 ? ic_miss_buff_data_12[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1704 = _T_1703 | _T_1689; // @[Mux.scala 27:72]
  wire  _T_1668 = byp_fetch_index_inc_0 == 4'hd; // @[el2_ifu_mem_ctl.scala 446:73]
  wire [15:0] _T_1690 = _T_1668 ? ic_miss_buff_data_13[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1705 = _T_1704 | _T_1690; // @[Mux.scala 27:72]
  wire  _T_1671 = byp_fetch_index_inc_0 == 4'he; // @[el2_ifu_mem_ctl.scala 446:73]
  wire [15:0] _T_1691 = _T_1671 ? ic_miss_buff_data_14[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1706 = _T_1705 | _T_1691; // @[Mux.scala 27:72]
  wire  _T_1674 = byp_fetch_index_inc_0 == 4'hf; // @[el2_ifu_mem_ctl.scala 446:73]
  wire [15:0] _T_1692 = _T_1674 ? ic_miss_buff_data_15[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1707 = _T_1706 | _T_1692; // @[Mux.scala 27:72]
  wire [3:0] byp_fetch_index_1 = {ifu_fetch_addr_int_f[4:2],1'h1}; // @[Cat.scala 29:58]
  wire  _T_1709 = byp_fetch_index_1 == 4'h0; // @[el2_ifu_mem_ctl.scala 446:179]
  wire [31:0] _T_1757 = _T_1709 ? ic_miss_buff_data_0 : 32'h0; // @[Mux.scala 27:72]
  wire  _T_1712 = byp_fetch_index_1 == 4'h1; // @[el2_ifu_mem_ctl.scala 446:179]
  wire [31:0] _T_1758 = _T_1712 ? ic_miss_buff_data_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1773 = _T_1757 | _T_1758; // @[Mux.scala 27:72]
  wire  _T_1715 = byp_fetch_index_1 == 4'h2; // @[el2_ifu_mem_ctl.scala 446:179]
  wire [31:0] _T_1759 = _T_1715 ? ic_miss_buff_data_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1774 = _T_1773 | _T_1759; // @[Mux.scala 27:72]
  wire  _T_1718 = byp_fetch_index_1 == 4'h3; // @[el2_ifu_mem_ctl.scala 446:179]
  wire [31:0] _T_1760 = _T_1718 ? ic_miss_buff_data_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1775 = _T_1774 | _T_1760; // @[Mux.scala 27:72]
  wire  _T_1721 = byp_fetch_index_1 == 4'h4; // @[el2_ifu_mem_ctl.scala 446:179]
  wire [31:0] _T_1761 = _T_1721 ? ic_miss_buff_data_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1776 = _T_1775 | _T_1761; // @[Mux.scala 27:72]
  wire  _T_1724 = byp_fetch_index_1 == 4'h5; // @[el2_ifu_mem_ctl.scala 446:179]
  wire [31:0] _T_1762 = _T_1724 ? ic_miss_buff_data_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1777 = _T_1776 | _T_1762; // @[Mux.scala 27:72]
  wire  _T_1727 = byp_fetch_index_1 == 4'h6; // @[el2_ifu_mem_ctl.scala 446:179]
  wire [31:0] _T_1763 = _T_1727 ? ic_miss_buff_data_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1778 = _T_1777 | _T_1763; // @[Mux.scala 27:72]
  wire  _T_1730 = byp_fetch_index_1 == 4'h7; // @[el2_ifu_mem_ctl.scala 446:179]
  wire [31:0] _T_1764 = _T_1730 ? ic_miss_buff_data_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1779 = _T_1778 | _T_1764; // @[Mux.scala 27:72]
  wire  _T_1733 = byp_fetch_index_1 == 4'h8; // @[el2_ifu_mem_ctl.scala 446:179]
  wire [31:0] _T_1765 = _T_1733 ? ic_miss_buff_data_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1780 = _T_1779 | _T_1765; // @[Mux.scala 27:72]
  wire  _T_1736 = byp_fetch_index_1 == 4'h9; // @[el2_ifu_mem_ctl.scala 446:179]
  wire [31:0] _T_1766 = _T_1736 ? ic_miss_buff_data_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1781 = _T_1780 | _T_1766; // @[Mux.scala 27:72]
  wire  _T_1739 = byp_fetch_index_1 == 4'ha; // @[el2_ifu_mem_ctl.scala 446:179]
  wire [31:0] _T_1767 = _T_1739 ? ic_miss_buff_data_10 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1782 = _T_1781 | _T_1767; // @[Mux.scala 27:72]
  wire  _T_1742 = byp_fetch_index_1 == 4'hb; // @[el2_ifu_mem_ctl.scala 446:179]
  wire [31:0] _T_1768 = _T_1742 ? ic_miss_buff_data_11 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1783 = _T_1782 | _T_1768; // @[Mux.scala 27:72]
  wire  _T_1745 = byp_fetch_index_1 == 4'hc; // @[el2_ifu_mem_ctl.scala 446:179]
  wire [31:0] _T_1769 = _T_1745 ? ic_miss_buff_data_12 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1784 = _T_1783 | _T_1769; // @[Mux.scala 27:72]
  wire  _T_1748 = byp_fetch_index_1 == 4'hd; // @[el2_ifu_mem_ctl.scala 446:179]
  wire [31:0] _T_1770 = _T_1748 ? ic_miss_buff_data_13 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1785 = _T_1784 | _T_1770; // @[Mux.scala 27:72]
  wire  _T_1751 = byp_fetch_index_1 == 4'he; // @[el2_ifu_mem_ctl.scala 446:179]
  wire [31:0] _T_1771 = _T_1751 ? ic_miss_buff_data_14 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1786 = _T_1785 | _T_1771; // @[Mux.scala 27:72]
  wire  _T_1754 = byp_fetch_index_1 == 4'hf; // @[el2_ifu_mem_ctl.scala 446:179]
  wire [31:0] _T_1772 = _T_1754 ? ic_miss_buff_data_15 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1787 = _T_1786 | _T_1772; // @[Mux.scala 27:72]
  wire [3:0] byp_fetch_index_0 = {ifu_fetch_addr_int_f[4:2],1'h0}; // @[Cat.scala 29:58]
  wire  _T_1789 = byp_fetch_index_0 == 4'h0; // @[el2_ifu_mem_ctl.scala 446:285]
  wire [31:0] _T_1837 = _T_1789 ? ic_miss_buff_data_0 : 32'h0; // @[Mux.scala 27:72]
  wire  _T_1792 = byp_fetch_index_0 == 4'h1; // @[el2_ifu_mem_ctl.scala 446:285]
  wire [31:0] _T_1838 = _T_1792 ? ic_miss_buff_data_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1853 = _T_1837 | _T_1838; // @[Mux.scala 27:72]
  wire  _T_1795 = byp_fetch_index_0 == 4'h2; // @[el2_ifu_mem_ctl.scala 446:285]
  wire [31:0] _T_1839 = _T_1795 ? ic_miss_buff_data_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1854 = _T_1853 | _T_1839; // @[Mux.scala 27:72]
  wire  _T_1798 = byp_fetch_index_0 == 4'h3; // @[el2_ifu_mem_ctl.scala 446:285]
  wire [31:0] _T_1840 = _T_1798 ? ic_miss_buff_data_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1855 = _T_1854 | _T_1840; // @[Mux.scala 27:72]
  wire  _T_1801 = byp_fetch_index_0 == 4'h4; // @[el2_ifu_mem_ctl.scala 446:285]
  wire [31:0] _T_1841 = _T_1801 ? ic_miss_buff_data_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1856 = _T_1855 | _T_1841; // @[Mux.scala 27:72]
  wire  _T_1804 = byp_fetch_index_0 == 4'h5; // @[el2_ifu_mem_ctl.scala 446:285]
  wire [31:0] _T_1842 = _T_1804 ? ic_miss_buff_data_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1857 = _T_1856 | _T_1842; // @[Mux.scala 27:72]
  wire  _T_1807 = byp_fetch_index_0 == 4'h6; // @[el2_ifu_mem_ctl.scala 446:285]
  wire [31:0] _T_1843 = _T_1807 ? ic_miss_buff_data_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1858 = _T_1857 | _T_1843; // @[Mux.scala 27:72]
  wire  _T_1810 = byp_fetch_index_0 == 4'h7; // @[el2_ifu_mem_ctl.scala 446:285]
  wire [31:0] _T_1844 = _T_1810 ? ic_miss_buff_data_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1859 = _T_1858 | _T_1844; // @[Mux.scala 27:72]
  wire  _T_1813 = byp_fetch_index_0 == 4'h8; // @[el2_ifu_mem_ctl.scala 446:285]
  wire [31:0] _T_1845 = _T_1813 ? ic_miss_buff_data_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1860 = _T_1859 | _T_1845; // @[Mux.scala 27:72]
  wire  _T_1816 = byp_fetch_index_0 == 4'h9; // @[el2_ifu_mem_ctl.scala 446:285]
  wire [31:0] _T_1846 = _T_1816 ? ic_miss_buff_data_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1861 = _T_1860 | _T_1846; // @[Mux.scala 27:72]
  wire  _T_1819 = byp_fetch_index_0 == 4'ha; // @[el2_ifu_mem_ctl.scala 446:285]
  wire [31:0] _T_1847 = _T_1819 ? ic_miss_buff_data_10 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1862 = _T_1861 | _T_1847; // @[Mux.scala 27:72]
  wire  _T_1822 = byp_fetch_index_0 == 4'hb; // @[el2_ifu_mem_ctl.scala 446:285]
  wire [31:0] _T_1848 = _T_1822 ? ic_miss_buff_data_11 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1863 = _T_1862 | _T_1848; // @[Mux.scala 27:72]
  wire  _T_1825 = byp_fetch_index_0 == 4'hc; // @[el2_ifu_mem_ctl.scala 446:285]
  wire [31:0] _T_1849 = _T_1825 ? ic_miss_buff_data_12 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1864 = _T_1863 | _T_1849; // @[Mux.scala 27:72]
  wire  _T_1828 = byp_fetch_index_0 == 4'hd; // @[el2_ifu_mem_ctl.scala 446:285]
  wire [31:0] _T_1850 = _T_1828 ? ic_miss_buff_data_13 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1865 = _T_1864 | _T_1850; // @[Mux.scala 27:72]
  wire  _T_1831 = byp_fetch_index_0 == 4'he; // @[el2_ifu_mem_ctl.scala 446:285]
  wire [31:0] _T_1851 = _T_1831 ? ic_miss_buff_data_14 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1866 = _T_1865 | _T_1851; // @[Mux.scala 27:72]
  wire  _T_1834 = byp_fetch_index_0 == 4'hf; // @[el2_ifu_mem_ctl.scala 446:285]
  wire [31:0] _T_1852 = _T_1834 ? ic_miss_buff_data_15 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1867 = _T_1866 | _T_1852; // @[Mux.scala 27:72]
  wire [79:0] _T_1870 = {_T_1707,_T_1787,_T_1867}; // @[Cat.scala 29:58]
  wire [3:0] byp_fetch_index_inc_1 = {byp_fetch_index_inc,1'h1}; // @[Cat.scala 29:58]
  wire  _T_1871 = byp_fetch_index_inc_1 == 4'h0; // @[el2_ifu_mem_ctl.scala 447:73]
  wire [15:0] _T_1919 = _T_1871 ? ic_miss_buff_data_0[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire  _T_1874 = byp_fetch_index_inc_1 == 4'h1; // @[el2_ifu_mem_ctl.scala 447:73]
  wire [15:0] _T_1920 = _T_1874 ? ic_miss_buff_data_1[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1935 = _T_1919 | _T_1920; // @[Mux.scala 27:72]
  wire  _T_1877 = byp_fetch_index_inc_1 == 4'h2; // @[el2_ifu_mem_ctl.scala 447:73]
  wire [15:0] _T_1921 = _T_1877 ? ic_miss_buff_data_2[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1936 = _T_1935 | _T_1921; // @[Mux.scala 27:72]
  wire  _T_1880 = byp_fetch_index_inc_1 == 4'h3; // @[el2_ifu_mem_ctl.scala 447:73]
  wire [15:0] _T_1922 = _T_1880 ? ic_miss_buff_data_3[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1937 = _T_1936 | _T_1922; // @[Mux.scala 27:72]
  wire  _T_1883 = byp_fetch_index_inc_1 == 4'h4; // @[el2_ifu_mem_ctl.scala 447:73]
  wire [15:0] _T_1923 = _T_1883 ? ic_miss_buff_data_4[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1938 = _T_1937 | _T_1923; // @[Mux.scala 27:72]
  wire  _T_1886 = byp_fetch_index_inc_1 == 4'h5; // @[el2_ifu_mem_ctl.scala 447:73]
  wire [15:0] _T_1924 = _T_1886 ? ic_miss_buff_data_5[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1939 = _T_1938 | _T_1924; // @[Mux.scala 27:72]
  wire  _T_1889 = byp_fetch_index_inc_1 == 4'h6; // @[el2_ifu_mem_ctl.scala 447:73]
  wire [15:0] _T_1925 = _T_1889 ? ic_miss_buff_data_6[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1940 = _T_1939 | _T_1925; // @[Mux.scala 27:72]
  wire  _T_1892 = byp_fetch_index_inc_1 == 4'h7; // @[el2_ifu_mem_ctl.scala 447:73]
  wire [15:0] _T_1926 = _T_1892 ? ic_miss_buff_data_7[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1941 = _T_1940 | _T_1926; // @[Mux.scala 27:72]
  wire  _T_1895 = byp_fetch_index_inc_1 == 4'h8; // @[el2_ifu_mem_ctl.scala 447:73]
  wire [15:0] _T_1927 = _T_1895 ? ic_miss_buff_data_8[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1942 = _T_1941 | _T_1927; // @[Mux.scala 27:72]
  wire  _T_1898 = byp_fetch_index_inc_1 == 4'h9; // @[el2_ifu_mem_ctl.scala 447:73]
  wire [15:0] _T_1928 = _T_1898 ? ic_miss_buff_data_9[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1943 = _T_1942 | _T_1928; // @[Mux.scala 27:72]
  wire  _T_1901 = byp_fetch_index_inc_1 == 4'ha; // @[el2_ifu_mem_ctl.scala 447:73]
  wire [15:0] _T_1929 = _T_1901 ? ic_miss_buff_data_10[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1944 = _T_1943 | _T_1929; // @[Mux.scala 27:72]
  wire  _T_1904 = byp_fetch_index_inc_1 == 4'hb; // @[el2_ifu_mem_ctl.scala 447:73]
  wire [15:0] _T_1930 = _T_1904 ? ic_miss_buff_data_11[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1945 = _T_1944 | _T_1930; // @[Mux.scala 27:72]
  wire  _T_1907 = byp_fetch_index_inc_1 == 4'hc; // @[el2_ifu_mem_ctl.scala 447:73]
  wire [15:0] _T_1931 = _T_1907 ? ic_miss_buff_data_12[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1946 = _T_1945 | _T_1931; // @[Mux.scala 27:72]
  wire  _T_1910 = byp_fetch_index_inc_1 == 4'hd; // @[el2_ifu_mem_ctl.scala 447:73]
  wire [15:0] _T_1932 = _T_1910 ? ic_miss_buff_data_13[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1947 = _T_1946 | _T_1932; // @[Mux.scala 27:72]
  wire  _T_1913 = byp_fetch_index_inc_1 == 4'he; // @[el2_ifu_mem_ctl.scala 447:73]
  wire [15:0] _T_1933 = _T_1913 ? ic_miss_buff_data_14[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1948 = _T_1947 | _T_1933; // @[Mux.scala 27:72]
  wire  _T_1916 = byp_fetch_index_inc_1 == 4'hf; // @[el2_ifu_mem_ctl.scala 447:73]
  wire [15:0] _T_1934 = _T_1916 ? ic_miss_buff_data_15[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1949 = _T_1948 | _T_1934; // @[Mux.scala 27:72]
  wire [31:0] _T_1999 = _T_1629 ? ic_miss_buff_data_0 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2000 = _T_1632 ? ic_miss_buff_data_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2015 = _T_1999 | _T_2000; // @[Mux.scala 27:72]
  wire [31:0] _T_2001 = _T_1635 ? ic_miss_buff_data_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2016 = _T_2015 | _T_2001; // @[Mux.scala 27:72]
  wire [31:0] _T_2002 = _T_1638 ? ic_miss_buff_data_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2017 = _T_2016 | _T_2002; // @[Mux.scala 27:72]
  wire [31:0] _T_2003 = _T_1641 ? ic_miss_buff_data_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2018 = _T_2017 | _T_2003; // @[Mux.scala 27:72]
  wire [31:0] _T_2004 = _T_1644 ? ic_miss_buff_data_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2019 = _T_2018 | _T_2004; // @[Mux.scala 27:72]
  wire [31:0] _T_2005 = _T_1647 ? ic_miss_buff_data_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2020 = _T_2019 | _T_2005; // @[Mux.scala 27:72]
  wire [31:0] _T_2006 = _T_1650 ? ic_miss_buff_data_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2021 = _T_2020 | _T_2006; // @[Mux.scala 27:72]
  wire [31:0] _T_2007 = _T_1653 ? ic_miss_buff_data_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2022 = _T_2021 | _T_2007; // @[Mux.scala 27:72]
  wire [31:0] _T_2008 = _T_1656 ? ic_miss_buff_data_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2023 = _T_2022 | _T_2008; // @[Mux.scala 27:72]
  wire [31:0] _T_2009 = _T_1659 ? ic_miss_buff_data_10 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2024 = _T_2023 | _T_2009; // @[Mux.scala 27:72]
  wire [31:0] _T_2010 = _T_1662 ? ic_miss_buff_data_11 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2025 = _T_2024 | _T_2010; // @[Mux.scala 27:72]
  wire [31:0] _T_2011 = _T_1665 ? ic_miss_buff_data_12 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2026 = _T_2025 | _T_2011; // @[Mux.scala 27:72]
  wire [31:0] _T_2012 = _T_1668 ? ic_miss_buff_data_13 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2027 = _T_2026 | _T_2012; // @[Mux.scala 27:72]
  wire [31:0] _T_2013 = _T_1671 ? ic_miss_buff_data_14 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2028 = _T_2027 | _T_2013; // @[Mux.scala 27:72]
  wire [31:0] _T_2014 = _T_1674 ? ic_miss_buff_data_15 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2029 = _T_2028 | _T_2014; // @[Mux.scala 27:72]
  wire [79:0] _T_2112 = {_T_1949,_T_2029,_T_1787}; // @[Cat.scala 29:58]
  wire [79:0] ic_byp_data_only_pre_new = _T_2115 ? _T_1870 : _T_2112; // @[el2_ifu_mem_ctl.scala 445:37]
  wire [79:0] _T_2117 = {16'h0,ic_byp_data_only_pre_new[79:16]}; // @[Cat.scala 29:58]
  wire [79:0] ic_byp_data_only_new = _T_2115 ? ic_byp_data_only_pre_new : _T_2117; // @[el2_ifu_mem_ctl.scala 449:30]
  wire [79:0] _GEN_793 = {{16'd0}, _T_1263}; // @[el2_ifu_mem_ctl.scala 380:109]
  wire [79:0] _T_1264 = _GEN_793 & ic_byp_data_only_new; // @[el2_ifu_mem_ctl.scala 380:109]
  wire [79:0] _GEN_794 = {{16'd0}, _T_1261}; // @[el2_ifu_mem_ctl.scala 380:83]
  wire [79:0] ic_premux_data = _GEN_794 | _T_1264; // @[el2_ifu_mem_ctl.scala 380:83]
  wire  fetch_req_f_qual = io_ic_hit_f & _T_317; // @[el2_ifu_mem_ctl.scala 387:38]
  wire [1:0] _T_1273 = ifc_region_acc_fault_f ? 2'h2 : 2'h0; // @[el2_ifu_mem_ctl.scala 391:8]
  wire [7:0] _T_1370 = {ic_miss_buff_data_valid_in_7,ic_miss_buff_data_valid_in_6,ic_miss_buff_data_valid_in_5,ic_miss_buff_data_valid_in_4,ic_miss_buff_data_valid_in_3,ic_miss_buff_data_valid_in_2,ic_miss_buff_data_valid_in_1,ic_miss_buff_data_valid_in_0}; // @[Cat.scala 29:58]
  wire  _T_1375 = ic_miss_buff_data_error[0] & _T_1341; // @[el2_ifu_mem_ctl.scala 412:32]
  wire  _T_2621 = |io_ifu_axi_rresp; // @[el2_ifu_mem_ctl.scala 623:47]
  wire  _T_2622 = _T_2621 & _T_13; // @[el2_ifu_mem_ctl.scala 623:50]
  wire  bus_ifu_wr_data_error = _T_2622 & miss_pending; // @[el2_ifu_mem_ctl.scala 623:68]
  wire  ic_miss_buff_data_error_in_0 = write_fill_data_0 ? bus_ifu_wr_data_error : _T_1375; // @[el2_ifu_mem_ctl.scala 411:72]
  wire  _T_1379 = ic_miss_buff_data_error[1] & _T_1341; // @[el2_ifu_mem_ctl.scala 412:32]
  wire  ic_miss_buff_data_error_in_1 = write_fill_data_1 ? bus_ifu_wr_data_error : _T_1379; // @[el2_ifu_mem_ctl.scala 411:72]
  wire  _T_1383 = ic_miss_buff_data_error[2] & _T_1341; // @[el2_ifu_mem_ctl.scala 412:32]
  wire  ic_miss_buff_data_error_in_2 = write_fill_data_2 ? bus_ifu_wr_data_error : _T_1383; // @[el2_ifu_mem_ctl.scala 411:72]
  wire  _T_1387 = ic_miss_buff_data_error[3] & _T_1341; // @[el2_ifu_mem_ctl.scala 412:32]
  wire  ic_miss_buff_data_error_in_3 = write_fill_data_3 ? bus_ifu_wr_data_error : _T_1387; // @[el2_ifu_mem_ctl.scala 411:72]
  wire  _T_1391 = ic_miss_buff_data_error[4] & _T_1341; // @[el2_ifu_mem_ctl.scala 412:32]
  wire  ic_miss_buff_data_error_in_4 = write_fill_data_4 ? bus_ifu_wr_data_error : _T_1391; // @[el2_ifu_mem_ctl.scala 411:72]
  wire  _T_1395 = ic_miss_buff_data_error[5] & _T_1341; // @[el2_ifu_mem_ctl.scala 412:32]
  wire  ic_miss_buff_data_error_in_5 = write_fill_data_5 ? bus_ifu_wr_data_error : _T_1395; // @[el2_ifu_mem_ctl.scala 411:72]
  wire  _T_1399 = ic_miss_buff_data_error[6] & _T_1341; // @[el2_ifu_mem_ctl.scala 412:32]
  wire  ic_miss_buff_data_error_in_6 = write_fill_data_6 ? bus_ifu_wr_data_error : _T_1399; // @[el2_ifu_mem_ctl.scala 411:72]
  wire  _T_1403 = ic_miss_buff_data_error[7] & _T_1341; // @[el2_ifu_mem_ctl.scala 412:32]
  wire  ic_miss_buff_data_error_in_7 = write_fill_data_7 ? bus_ifu_wr_data_error : _T_1403; // @[el2_ifu_mem_ctl.scala 411:72]
  wire [7:0] _T_1410 = {ic_miss_buff_data_error_in_7,ic_miss_buff_data_error_in_6,ic_miss_buff_data_error_in_5,ic_miss_buff_data_error_in_4,ic_miss_buff_data_error_in_3,ic_miss_buff_data_error_in_2,ic_miss_buff_data_error_in_1,ic_miss_buff_data_error_in_0}; // @[Cat.scala 29:58]
  reg [5:0] perr_ic_index_ff; // @[Reg.scala 27:20]
  wire  _T_2427 = 3'h0 == perr_state; // @[Conditional.scala 37:30]
  wire  _T_2435 = _T_6 & _T_317; // @[el2_ifu_mem_ctl.scala 492:65]
  wire  _T_2436 = _T_2435 | io_iccm_dma_sb_error; // @[el2_ifu_mem_ctl.scala 492:88]
  wire  _T_2438 = _T_2436 & _T_2549; // @[el2_ifu_mem_ctl.scala 492:112]
  wire  _T_2439 = 3'h1 == perr_state; // @[Conditional.scala 37:30]
  wire  _T_2440 = io_dec_tlu_flush_lower_wb | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 497:50]
  wire  _T_2442 = 3'h2 == perr_state; // @[Conditional.scala 37:30]
  wire  _T_2448 = 3'h4 == perr_state; // @[Conditional.scala 37:30]
  wire  _T_2450 = 3'h3 == perr_state; // @[Conditional.scala 37:30]
  wire  _GEN_38 = _T_2448 | _T_2450; // @[Conditional.scala 39:67]
  wire  _GEN_40 = _T_2442 ? _T_2440 : _GEN_38; // @[Conditional.scala 39:67]
  wire  _GEN_42 = _T_2439 ? _T_2440 : _GEN_40; // @[Conditional.scala 39:67]
  wire  perr_state_en = _T_2427 ? _T_2438 : _GEN_42; // @[Conditional.scala 40:58]
  wire  perr_sb_write_status = _T_2427 & perr_state_en; // @[Conditional.scala 40:58]
  wire  _T_2441 = io_dec_tlu_flush_lower_wb & io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 498:56]
  wire  _GEN_43 = _T_2439 & _T_2441; // @[Conditional.scala 39:67]
  wire  perr_sel_invalidate = _T_2427 ? 1'h0 : _GEN_43; // @[Conditional.scala 40:58]
  wire [1:0] perr_err_inv_way = perr_sel_invalidate ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  reg  dma_sb_err_state_ff; // @[el2_ifu_mem_ctl.scala 483:58]
  wire  _T_2424 = ~dma_sb_err_state_ff; // @[el2_ifu_mem_ctl.scala 482:49]
  wire  _T_2429 = io_ic_error_start & _T_317; // @[el2_ifu_mem_ctl.scala 491:87]
  wire  _T_2443 = io_dec_tlu_flush_err_wb & io_dec_tlu_flush_lower_wb; // @[el2_ifu_mem_ctl.scala 501:54]
  wire  _T_2444 = _T_2443 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 501:84]
  wire  _T_2453 = perr_state == 3'h2; // @[el2_ifu_mem_ctl.scala 522:66]
  wire  _T_2454 = io_dec_tlu_flush_err_wb & _T_2453; // @[el2_ifu_mem_ctl.scala 522:52]
  wire  _T_2456 = _T_2454 & _T_2549; // @[el2_ifu_mem_ctl.scala 522:81]
  wire  _T_2458 = io_dec_tlu_flush_lower_wb | io_dec_tlu_i0_commit_cmt; // @[el2_ifu_mem_ctl.scala 525:59]
  wire  _T_2459 = _T_2458 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 525:86]
  wire  _T_2473 = _T_2458 | io_ifu_fetch_val[0]; // @[el2_ifu_mem_ctl.scala 528:81]
  wire  _T_2474 = _T_2473 | ifu_bp_hit_taken_q_f; // @[el2_ifu_mem_ctl.scala 528:103]
  wire  _T_2475 = _T_2474 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 528:126]
  wire  _T_2495 = _T_2473 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 535:103]
  wire  _T_2502 = ~io_dec_tlu_flush_err_wb; // @[el2_ifu_mem_ctl.scala 540:62]
  wire  _T_2503 = io_dec_tlu_flush_lower_wb & _T_2502; // @[el2_ifu_mem_ctl.scala 540:60]
  wire  _T_2504 = _T_2503 | io_dec_tlu_i0_commit_cmt; // @[el2_ifu_mem_ctl.scala 540:88]
  wire  _T_2505 = _T_2504 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 540:115]
  wire  _GEN_50 = _T_2501 & _T_2459; // @[Conditional.scala 39:67]
  wire  _GEN_53 = _T_2484 ? _T_2495 : _GEN_50; // @[Conditional.scala 39:67]
  wire  _GEN_55 = _T_2484 | _T_2501; // @[Conditional.scala 39:67]
  wire  _GEN_57 = _T_2457 ? _T_2475 : _GEN_53; // @[Conditional.scala 39:67]
  wire  _GEN_59 = _T_2457 | _GEN_55; // @[Conditional.scala 39:67]
  wire  err_stop_state_en = _T_2452 ? _T_2456 : _GEN_57; // @[Conditional.scala 40:58]
  reg  ifu_bus_cmd_valid; // @[Reg.scala 27:20]
  wire  _T_2517 = ic_act_miss_f | ifu_bus_cmd_valid; // @[el2_ifu_mem_ctl.scala 557:64]
  wire  _T_2519 = _T_2517 & _T_2549; // @[el2_ifu_mem_ctl.scala 557:85]
  reg [2:0] bus_cmd_beat_count; // @[Reg.scala 27:20]
  wire  _T_2521 = bus_cmd_beat_count == 3'h7; // @[el2_ifu_mem_ctl.scala 557:133]
  wire  _T_2522 = _T_2521 & ifu_bus_cmd_valid; // @[el2_ifu_mem_ctl.scala 557:164]
  wire  _T_2523 = _T_2522 & io_ifu_axi_arready; // @[el2_ifu_mem_ctl.scala 557:184]
  wire  _T_2524 = _T_2523 & miss_pending; // @[el2_ifu_mem_ctl.scala 557:204]
  wire  _T_2525 = ~_T_2524; // @[el2_ifu_mem_ctl.scala 557:112]
  wire  ifc_bus_ic_req_ff_in = _T_2519 & _T_2525; // @[el2_ifu_mem_ctl.scala 557:110]
  wire  _T_2526 = io_ifu_bus_clk_en | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 558:80]
  wire  ifu_bus_arready = io_ifu_axi_arready & io_ifu_bus_clk_en; // @[el2_ifu_mem_ctl.scala 589:45]
  wire  _T_2543 = io_ifu_axi_arvalid & ifu_bus_arready; // @[el2_ifu_mem_ctl.scala 592:35]
  wire  _T_2544 = _T_2543 & miss_pending; // @[el2_ifu_mem_ctl.scala 592:53]
  wire  bus_cmd_sent = _T_2544 & _T_2549; // @[el2_ifu_mem_ctl.scala 592:68]
  wire [2:0] _T_2534 = ifu_bus_cmd_valid ? 3'h7 : 3'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_2536 = {miss_addr,bus_rd_addr_count,3'h0}; // @[Cat.scala 29:58]
  wire [31:0] _T_2538 = ifu_bus_cmd_valid ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  reg  ifu_bus_arready_unq_ff; // @[Reg.scala 27:20]
  reg  ifu_bus_arvalid_ff; // @[Reg.scala 27:20]
  wire  ifu_bus_arready_ff = ifu_bus_arready_unq_ff & bus_ifu_bus_clk_en_ff; // @[el2_ifu_mem_ctl.scala 590:51]
  wire  _T_2564 = ~scnd_miss_req; // @[el2_ifu_mem_ctl.scala 600:73]
  wire  _T_2565 = _T_2550 & _T_2564; // @[el2_ifu_mem_ctl.scala 600:71]
  wire  _T_2567 = last_data_recieved_ff & _T_1341; // @[el2_ifu_mem_ctl.scala 600:114]
  wire  last_data_recieved_in = _T_2565 | _T_2567; // @[el2_ifu_mem_ctl.scala 600:89]
  wire [2:0] _T_2573 = bus_rd_addr_count + 3'h1; // @[el2_ifu_mem_ctl.scala 605:45]
  wire  _T_2576 = io_ifu_bus_clk_en | ic_act_miss_f; // @[el2_ifu_mem_ctl.scala 606:81]
  wire  _T_2577 = _T_2576 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 606:97]
  wire  _T_2579 = ifu_bus_cmd_valid & io_ifu_axi_arready; // @[el2_ifu_mem_ctl.scala 608:48]
  wire  _T_2580 = _T_2579 & miss_pending; // @[el2_ifu_mem_ctl.scala 608:68]
  wire  bus_inc_cmd_beat_cnt = _T_2580 & _T_2549; // @[el2_ifu_mem_ctl.scala 608:83]
  wire  bus_reset_cmd_beat_cnt_secondlast = ic_act_miss_f & uncacheable_miss_in; // @[el2_ifu_mem_ctl.scala 610:57]
  wire  _T_2584 = ~bus_inc_cmd_beat_cnt; // @[el2_ifu_mem_ctl.scala 611:31]
  wire  _T_2585 = ic_act_miss_f | scnd_miss_req; // @[el2_ifu_mem_ctl.scala 611:71]
  wire  _T_2586 = _T_2585 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 611:87]
  wire  _T_2587 = ~_T_2586; // @[el2_ifu_mem_ctl.scala 611:55]
  wire  bus_hold_cmd_beat_cnt = _T_2584 & _T_2587; // @[el2_ifu_mem_ctl.scala 611:53]
  wire  _T_2588 = bus_inc_cmd_beat_cnt | ic_act_miss_f; // @[el2_ifu_mem_ctl.scala 612:46]
  wire  bus_cmd_beat_en = _T_2588 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 612:62]
  wire [2:0] _T_2591 = bus_cmd_beat_count + 3'h1; // @[el2_ifu_mem_ctl.scala 614:46]
  wire [2:0] _T_2593 = bus_reset_cmd_beat_cnt_secondlast ? 3'h6 : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_2594 = bus_inc_cmd_beat_cnt ? _T_2591 : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_2595 = bus_hold_cmd_beat_cnt ? bus_cmd_beat_count : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_2597 = _T_2593 | _T_2594; // @[Mux.scala 27:72]
  wire [2:0] bus_new_cmd_beat_count = _T_2597 | _T_2595; // @[Mux.scala 27:72]
  wire  _T_2601 = _T_2577 & bus_cmd_beat_en; // @[el2_ifu_mem_ctl.scala 615:125]
  reg  ifc_dma_access_ok_prev; // @[el2_ifu_mem_ctl.scala 626:62]
  wire  _T_2629 = ~iccm_correct_ecc; // @[el2_ifu_mem_ctl.scala 631:50]
  wire  _T_2630 = io_ifc_dma_access_ok & _T_2629; // @[el2_ifu_mem_ctl.scala 631:47]
  wire  _T_2631 = ~io_iccm_dma_sb_error; // @[el2_ifu_mem_ctl.scala 631:70]
  wire  ifc_dma_access_ok_d = _T_2630 & _T_2631; // @[el2_ifu_mem_ctl.scala 631:68]
  wire  _T_2635 = _T_2630 & ifc_dma_access_ok_prev; // @[el2_ifu_mem_ctl.scala 632:72]
  wire  _T_2636 = perr_state == 3'h0; // @[el2_ifu_mem_ctl.scala 632:111]
  wire  _T_2637 = _T_2635 & _T_2636; // @[el2_ifu_mem_ctl.scala 632:97]
  wire  ifc_dma_access_q_ok = _T_2637 & _T_2631; // @[el2_ifu_mem_ctl.scala 632:127]
  wire  _T_2640 = ifc_dma_access_q_ok & io_dma_iccm_req; // @[el2_ifu_mem_ctl.scala 635:40]
  wire  _T_2641 = _T_2640 & io_dma_mem_write; // @[el2_ifu_mem_ctl.scala 635:58]
  wire  _T_2644 = ~io_dma_mem_write; // @[el2_ifu_mem_ctl.scala 636:60]
  wire  _T_2645 = _T_2640 & _T_2644; // @[el2_ifu_mem_ctl.scala 636:58]
  wire  _T_2646 = io_ifc_iccm_access_bf & io_ifc_fetch_req_bf; // @[el2_ifu_mem_ctl.scala 636:104]
  wire [2:0] _T_2651 = io_dma_iccm_req ? 3'h7 : 3'h0; // @[Bitwise.scala 72:12]
  wire [8:0] _T_2757 = {io_dma_mem_wdata[48],io_dma_mem_wdata[46],io_dma_mem_wdata[44],io_dma_mem_wdata[42],io_dma_mem_wdata[40],io_dma_mem_wdata[38],io_dma_mem_wdata[37],io_dma_mem_wdata[35],io_dma_mem_wdata[33]}; // @[el2_lib.scala 268:22]
  wire [17:0] _T_2766 = {io_dma_mem_wdata[63],io_dma_mem_wdata[62],io_dma_mem_wdata[60],io_dma_mem_wdata[59],io_dma_mem_wdata[57],io_dma_mem_wdata[55],io_dma_mem_wdata[53],io_dma_mem_wdata[52],io_dma_mem_wdata[50],_T_2757}; // @[el2_lib.scala 268:22]
  wire  _T_2767 = ^_T_2766; // @[el2_lib.scala 268:29]
  wire [8:0] _T_2775 = {io_dma_mem_wdata[47],io_dma_mem_wdata[46],io_dma_mem_wdata[43],io_dma_mem_wdata[42],io_dma_mem_wdata[39],io_dma_mem_wdata[38],io_dma_mem_wdata[36],io_dma_mem_wdata[35],io_dma_mem_wdata[32]}; // @[el2_lib.scala 268:39]
  wire [17:0] _T_2784 = {io_dma_mem_wdata[63],io_dma_mem_wdata[61],io_dma_mem_wdata[60],io_dma_mem_wdata[58],io_dma_mem_wdata[57],io_dma_mem_wdata[54],io_dma_mem_wdata[53],io_dma_mem_wdata[51],io_dma_mem_wdata[50],_T_2775}; // @[el2_lib.scala 268:39]
  wire  _T_2785 = ^_T_2784; // @[el2_lib.scala 268:46]
  wire [8:0] _T_2793 = {io_dma_mem_wdata[47],io_dma_mem_wdata[46],io_dma_mem_wdata[41],io_dma_mem_wdata[40],io_dma_mem_wdata[39],io_dma_mem_wdata[38],io_dma_mem_wdata[34],io_dma_mem_wdata[33],io_dma_mem_wdata[32]}; // @[el2_lib.scala 268:56]
  wire [17:0] _T_2802 = {io_dma_mem_wdata[62],io_dma_mem_wdata[61],io_dma_mem_wdata[60],io_dma_mem_wdata[56],io_dma_mem_wdata[55],io_dma_mem_wdata[54],io_dma_mem_wdata[53],io_dma_mem_wdata[49],io_dma_mem_wdata[48],_T_2793}; // @[el2_lib.scala 268:56]
  wire  _T_2803 = ^_T_2802; // @[el2_lib.scala 268:63]
  wire [6:0] _T_2809 = {io_dma_mem_wdata[44],io_dma_mem_wdata[43],io_dma_mem_wdata[42],io_dma_mem_wdata[41],io_dma_mem_wdata[40],io_dma_mem_wdata[39],io_dma_mem_wdata[38]}; // @[el2_lib.scala 268:73]
  wire [14:0] _T_2817 = {io_dma_mem_wdata[59],io_dma_mem_wdata[58],io_dma_mem_wdata[57],io_dma_mem_wdata[56],io_dma_mem_wdata[55],io_dma_mem_wdata[54],io_dma_mem_wdata[53],io_dma_mem_wdata[45],_T_2809}; // @[el2_lib.scala 268:73]
  wire  _T_2818 = ^_T_2817; // @[el2_lib.scala 268:80]
  wire [14:0] _T_2832 = {io_dma_mem_wdata[52],io_dma_mem_wdata[51],io_dma_mem_wdata[50],io_dma_mem_wdata[49],io_dma_mem_wdata[48],io_dma_mem_wdata[47],io_dma_mem_wdata[46],io_dma_mem_wdata[45],_T_2809}; // @[el2_lib.scala 268:90]
  wire  _T_2833 = ^_T_2832; // @[el2_lib.scala 268:97]
  wire [5:0] _T_2838 = {io_dma_mem_wdata[37],io_dma_mem_wdata[36],io_dma_mem_wdata[35],io_dma_mem_wdata[34],io_dma_mem_wdata[33],io_dma_mem_wdata[32]}; // @[el2_lib.scala 268:107]
  wire  _T_2839 = ^_T_2838; // @[el2_lib.scala 268:114]
  wire [5:0] _T_2844 = {_T_2767,_T_2785,_T_2803,_T_2818,_T_2833,_T_2839}; // @[Cat.scala 29:58]
  wire  _T_2845 = ^io_dma_mem_wdata[63:32]; // @[el2_lib.scala 269:13]
  wire  _T_2846 = ^_T_2844; // @[el2_lib.scala 269:23]
  wire  _T_2847 = _T_2845 ^ _T_2846; // @[el2_lib.scala 269:18]
  wire [8:0] _T_2953 = {io_dma_mem_wdata[16],io_dma_mem_wdata[14],io_dma_mem_wdata[12],io_dma_mem_wdata[10],io_dma_mem_wdata[8],io_dma_mem_wdata[6],io_dma_mem_wdata[5],io_dma_mem_wdata[3],io_dma_mem_wdata[1]}; // @[el2_lib.scala 268:22]
  wire [17:0] _T_2962 = {io_dma_mem_wdata[31],io_dma_mem_wdata[30],io_dma_mem_wdata[28],io_dma_mem_wdata[27],io_dma_mem_wdata[25],io_dma_mem_wdata[23],io_dma_mem_wdata[21],io_dma_mem_wdata[20],io_dma_mem_wdata[18],_T_2953}; // @[el2_lib.scala 268:22]
  wire  _T_2963 = ^_T_2962; // @[el2_lib.scala 268:29]
  wire [8:0] _T_2971 = {io_dma_mem_wdata[15],io_dma_mem_wdata[14],io_dma_mem_wdata[11],io_dma_mem_wdata[10],io_dma_mem_wdata[7],io_dma_mem_wdata[6],io_dma_mem_wdata[4],io_dma_mem_wdata[3],io_dma_mem_wdata[0]}; // @[el2_lib.scala 268:39]
  wire [17:0] _T_2980 = {io_dma_mem_wdata[31],io_dma_mem_wdata[29],io_dma_mem_wdata[28],io_dma_mem_wdata[26],io_dma_mem_wdata[25],io_dma_mem_wdata[22],io_dma_mem_wdata[21],io_dma_mem_wdata[19],io_dma_mem_wdata[18],_T_2971}; // @[el2_lib.scala 268:39]
  wire  _T_2981 = ^_T_2980; // @[el2_lib.scala 268:46]
  wire [8:0] _T_2989 = {io_dma_mem_wdata[15],io_dma_mem_wdata[14],io_dma_mem_wdata[9],io_dma_mem_wdata[8],io_dma_mem_wdata[7],io_dma_mem_wdata[6],io_dma_mem_wdata[2],io_dma_mem_wdata[1],io_dma_mem_wdata[0]}; // @[el2_lib.scala 268:56]
  wire [17:0] _T_2998 = {io_dma_mem_wdata[30],io_dma_mem_wdata[29],io_dma_mem_wdata[28],io_dma_mem_wdata[24],io_dma_mem_wdata[23],io_dma_mem_wdata[22],io_dma_mem_wdata[21],io_dma_mem_wdata[17],io_dma_mem_wdata[16],_T_2989}; // @[el2_lib.scala 268:56]
  wire  _T_2999 = ^_T_2998; // @[el2_lib.scala 268:63]
  wire [6:0] _T_3005 = {io_dma_mem_wdata[12],io_dma_mem_wdata[11],io_dma_mem_wdata[10],io_dma_mem_wdata[9],io_dma_mem_wdata[8],io_dma_mem_wdata[7],io_dma_mem_wdata[6]}; // @[el2_lib.scala 268:73]
  wire [14:0] _T_3013 = {io_dma_mem_wdata[27],io_dma_mem_wdata[26],io_dma_mem_wdata[25],io_dma_mem_wdata[24],io_dma_mem_wdata[23],io_dma_mem_wdata[22],io_dma_mem_wdata[21],io_dma_mem_wdata[13],_T_3005}; // @[el2_lib.scala 268:73]
  wire  _T_3014 = ^_T_3013; // @[el2_lib.scala 268:80]
  wire [14:0] _T_3028 = {io_dma_mem_wdata[20],io_dma_mem_wdata[19],io_dma_mem_wdata[18],io_dma_mem_wdata[17],io_dma_mem_wdata[16],io_dma_mem_wdata[15],io_dma_mem_wdata[14],io_dma_mem_wdata[13],_T_3005}; // @[el2_lib.scala 268:90]
  wire  _T_3029 = ^_T_3028; // @[el2_lib.scala 268:97]
  wire [5:0] _T_3034 = {io_dma_mem_wdata[5],io_dma_mem_wdata[4],io_dma_mem_wdata[3],io_dma_mem_wdata[2],io_dma_mem_wdata[1],io_dma_mem_wdata[0]}; // @[el2_lib.scala 268:107]
  wire  _T_3035 = ^_T_3034; // @[el2_lib.scala 268:114]
  wire [5:0] _T_3040 = {_T_2963,_T_2981,_T_2999,_T_3014,_T_3029,_T_3035}; // @[Cat.scala 29:58]
  wire  _T_3041 = ^io_dma_mem_wdata[31:0]; // @[el2_lib.scala 269:13]
  wire  _T_3042 = ^_T_3040; // @[el2_lib.scala 269:23]
  wire  _T_3043 = _T_3041 ^ _T_3042; // @[el2_lib.scala 269:18]
  wire [6:0] _T_3044 = {_T_3043,_T_2963,_T_2981,_T_2999,_T_3014,_T_3029,_T_3035}; // @[Cat.scala 29:58]
  wire [13:0] dma_mem_ecc = {_T_2847,_T_2767,_T_2785,_T_2803,_T_2818,_T_2833,_T_2839,_T_3044}; // @[Cat.scala 29:58]
  wire  _T_3046 = ~_T_2640; // @[el2_ifu_mem_ctl.scala 641:45]
  wire  _T_3047 = iccm_correct_ecc & _T_3046; // @[el2_ifu_mem_ctl.scala 641:43]
  reg [38:0] iccm_ecc_corr_data_ff; // @[Reg.scala 27:20]
  wire [77:0] _T_3048 = {iccm_ecc_corr_data_ff,iccm_ecc_corr_data_ff}; // @[Cat.scala 29:58]
  wire [77:0] _T_3055 = {dma_mem_ecc[13:7],io_dma_mem_wdata[63:32],dma_mem_ecc[6:0],io_dma_mem_wdata[31:0]}; // @[Cat.scala 29:58]
  reg [1:0] dma_mem_addr_ff; // @[el2_ifu_mem_ctl.scala 655:53]
  wire  _T_3387 = _T_3299[5:0] == 6'h27; // @[el2_lib.scala 307:41]
  wire  _T_3385 = _T_3299[5:0] == 6'h26; // @[el2_lib.scala 307:41]
  wire  _T_3383 = _T_3299[5:0] == 6'h25; // @[el2_lib.scala 307:41]
  wire  _T_3381 = _T_3299[5:0] == 6'h24; // @[el2_lib.scala 307:41]
  wire  _T_3379 = _T_3299[5:0] == 6'h23; // @[el2_lib.scala 307:41]
  wire  _T_3377 = _T_3299[5:0] == 6'h22; // @[el2_lib.scala 307:41]
  wire  _T_3375 = _T_3299[5:0] == 6'h21; // @[el2_lib.scala 307:41]
  wire  _T_3373 = _T_3299[5:0] == 6'h20; // @[el2_lib.scala 307:41]
  wire  _T_3371 = _T_3299[5:0] == 6'h1f; // @[el2_lib.scala 307:41]
  wire  _T_3369 = _T_3299[5:0] == 6'h1e; // @[el2_lib.scala 307:41]
  wire [9:0] _T_3445 = {_T_3387,_T_3385,_T_3383,_T_3381,_T_3379,_T_3377,_T_3375,_T_3373,_T_3371,_T_3369}; // @[el2_lib.scala 310:69]
  wire  _T_3367 = _T_3299[5:0] == 6'h1d; // @[el2_lib.scala 307:41]
  wire  _T_3365 = _T_3299[5:0] == 6'h1c; // @[el2_lib.scala 307:41]
  wire  _T_3363 = _T_3299[5:0] == 6'h1b; // @[el2_lib.scala 307:41]
  wire  _T_3361 = _T_3299[5:0] == 6'h1a; // @[el2_lib.scala 307:41]
  wire  _T_3359 = _T_3299[5:0] == 6'h19; // @[el2_lib.scala 307:41]
  wire  _T_3357 = _T_3299[5:0] == 6'h18; // @[el2_lib.scala 307:41]
  wire  _T_3355 = _T_3299[5:0] == 6'h17; // @[el2_lib.scala 307:41]
  wire  _T_3353 = _T_3299[5:0] == 6'h16; // @[el2_lib.scala 307:41]
  wire  _T_3351 = _T_3299[5:0] == 6'h15; // @[el2_lib.scala 307:41]
  wire  _T_3349 = _T_3299[5:0] == 6'h14; // @[el2_lib.scala 307:41]
  wire [9:0] _T_3436 = {_T_3367,_T_3365,_T_3363,_T_3361,_T_3359,_T_3357,_T_3355,_T_3353,_T_3351,_T_3349}; // @[el2_lib.scala 310:69]
  wire  _T_3347 = _T_3299[5:0] == 6'h13; // @[el2_lib.scala 307:41]
  wire  _T_3345 = _T_3299[5:0] == 6'h12; // @[el2_lib.scala 307:41]
  wire  _T_3343 = _T_3299[5:0] == 6'h11; // @[el2_lib.scala 307:41]
  wire  _T_3341 = _T_3299[5:0] == 6'h10; // @[el2_lib.scala 307:41]
  wire  _T_3339 = _T_3299[5:0] == 6'hf; // @[el2_lib.scala 307:41]
  wire  _T_3337 = _T_3299[5:0] == 6'he; // @[el2_lib.scala 307:41]
  wire  _T_3335 = _T_3299[5:0] == 6'hd; // @[el2_lib.scala 307:41]
  wire  _T_3333 = _T_3299[5:0] == 6'hc; // @[el2_lib.scala 307:41]
  wire  _T_3331 = _T_3299[5:0] == 6'hb; // @[el2_lib.scala 307:41]
  wire  _T_3329 = _T_3299[5:0] == 6'ha; // @[el2_lib.scala 307:41]
  wire [9:0] _T_3426 = {_T_3347,_T_3345,_T_3343,_T_3341,_T_3339,_T_3337,_T_3335,_T_3333,_T_3331,_T_3329}; // @[el2_lib.scala 310:69]
  wire  _T_3327 = _T_3299[5:0] == 6'h9; // @[el2_lib.scala 307:41]
  wire  _T_3325 = _T_3299[5:0] == 6'h8; // @[el2_lib.scala 307:41]
  wire  _T_3323 = _T_3299[5:0] == 6'h7; // @[el2_lib.scala 307:41]
  wire  _T_3321 = _T_3299[5:0] == 6'h6; // @[el2_lib.scala 307:41]
  wire  _T_3319 = _T_3299[5:0] == 6'h5; // @[el2_lib.scala 307:41]
  wire  _T_3317 = _T_3299[5:0] == 6'h4; // @[el2_lib.scala 307:41]
  wire  _T_3315 = _T_3299[5:0] == 6'h3; // @[el2_lib.scala 307:41]
  wire  _T_3313 = _T_3299[5:0] == 6'h2; // @[el2_lib.scala 307:41]
  wire  _T_3311 = _T_3299[5:0] == 6'h1; // @[el2_lib.scala 307:41]
  wire [18:0] _T_3427 = {_T_3426,_T_3327,_T_3325,_T_3323,_T_3321,_T_3319,_T_3317,_T_3315,_T_3313,_T_3311}; // @[el2_lib.scala 310:69]
  wire [38:0] _T_3447 = {_T_3445,_T_3436,_T_3427}; // @[el2_lib.scala 310:69]
  wire [7:0] _T_3402 = {io_iccm_rd_data_ecc[35],io_iccm_rd_data_ecc[3:1],io_iccm_rd_data_ecc[34],io_iccm_rd_data_ecc[0],io_iccm_rd_data_ecc[33:32]}; // @[Cat.scala 29:58]
  wire [38:0] _T_3408 = {io_iccm_rd_data_ecc[38],io_iccm_rd_data_ecc[31:26],io_iccm_rd_data_ecc[37],io_iccm_rd_data_ecc[25:11],io_iccm_rd_data_ecc[36],io_iccm_rd_data_ecc[10:4],_T_3402}; // @[Cat.scala 29:58]
  wire [38:0] _T_3448 = _T_3447 ^ _T_3408; // @[el2_lib.scala 310:76]
  wire [38:0] _T_3449 = _T_3303 ? _T_3448 : _T_3408; // @[el2_lib.scala 310:31]
  wire [31:0] iccm_corrected_data_0 = {_T_3449[37:32],_T_3449[30:16],_T_3449[14:8],_T_3449[6:4],_T_3449[2]}; // @[Cat.scala 29:58]
  wire  _T_3772 = _T_3684[5:0] == 6'h27; // @[el2_lib.scala 307:41]
  wire  _T_3770 = _T_3684[5:0] == 6'h26; // @[el2_lib.scala 307:41]
  wire  _T_3768 = _T_3684[5:0] == 6'h25; // @[el2_lib.scala 307:41]
  wire  _T_3766 = _T_3684[5:0] == 6'h24; // @[el2_lib.scala 307:41]
  wire  _T_3764 = _T_3684[5:0] == 6'h23; // @[el2_lib.scala 307:41]
  wire  _T_3762 = _T_3684[5:0] == 6'h22; // @[el2_lib.scala 307:41]
  wire  _T_3760 = _T_3684[5:0] == 6'h21; // @[el2_lib.scala 307:41]
  wire  _T_3758 = _T_3684[5:0] == 6'h20; // @[el2_lib.scala 307:41]
  wire  _T_3756 = _T_3684[5:0] == 6'h1f; // @[el2_lib.scala 307:41]
  wire  _T_3754 = _T_3684[5:0] == 6'h1e; // @[el2_lib.scala 307:41]
  wire [9:0] _T_3830 = {_T_3772,_T_3770,_T_3768,_T_3766,_T_3764,_T_3762,_T_3760,_T_3758,_T_3756,_T_3754}; // @[el2_lib.scala 310:69]
  wire  _T_3752 = _T_3684[5:0] == 6'h1d; // @[el2_lib.scala 307:41]
  wire  _T_3750 = _T_3684[5:0] == 6'h1c; // @[el2_lib.scala 307:41]
  wire  _T_3748 = _T_3684[5:0] == 6'h1b; // @[el2_lib.scala 307:41]
  wire  _T_3746 = _T_3684[5:0] == 6'h1a; // @[el2_lib.scala 307:41]
  wire  _T_3744 = _T_3684[5:0] == 6'h19; // @[el2_lib.scala 307:41]
  wire  _T_3742 = _T_3684[5:0] == 6'h18; // @[el2_lib.scala 307:41]
  wire  _T_3740 = _T_3684[5:0] == 6'h17; // @[el2_lib.scala 307:41]
  wire  _T_3738 = _T_3684[5:0] == 6'h16; // @[el2_lib.scala 307:41]
  wire  _T_3736 = _T_3684[5:0] == 6'h15; // @[el2_lib.scala 307:41]
  wire  _T_3734 = _T_3684[5:0] == 6'h14; // @[el2_lib.scala 307:41]
  wire [9:0] _T_3821 = {_T_3752,_T_3750,_T_3748,_T_3746,_T_3744,_T_3742,_T_3740,_T_3738,_T_3736,_T_3734}; // @[el2_lib.scala 310:69]
  wire  _T_3732 = _T_3684[5:0] == 6'h13; // @[el2_lib.scala 307:41]
  wire  _T_3730 = _T_3684[5:0] == 6'h12; // @[el2_lib.scala 307:41]
  wire  _T_3728 = _T_3684[5:0] == 6'h11; // @[el2_lib.scala 307:41]
  wire  _T_3726 = _T_3684[5:0] == 6'h10; // @[el2_lib.scala 307:41]
  wire  _T_3724 = _T_3684[5:0] == 6'hf; // @[el2_lib.scala 307:41]
  wire  _T_3722 = _T_3684[5:0] == 6'he; // @[el2_lib.scala 307:41]
  wire  _T_3720 = _T_3684[5:0] == 6'hd; // @[el2_lib.scala 307:41]
  wire  _T_3718 = _T_3684[5:0] == 6'hc; // @[el2_lib.scala 307:41]
  wire  _T_3716 = _T_3684[5:0] == 6'hb; // @[el2_lib.scala 307:41]
  wire  _T_3714 = _T_3684[5:0] == 6'ha; // @[el2_lib.scala 307:41]
  wire [9:0] _T_3811 = {_T_3732,_T_3730,_T_3728,_T_3726,_T_3724,_T_3722,_T_3720,_T_3718,_T_3716,_T_3714}; // @[el2_lib.scala 310:69]
  wire  _T_3712 = _T_3684[5:0] == 6'h9; // @[el2_lib.scala 307:41]
  wire  _T_3710 = _T_3684[5:0] == 6'h8; // @[el2_lib.scala 307:41]
  wire  _T_3708 = _T_3684[5:0] == 6'h7; // @[el2_lib.scala 307:41]
  wire  _T_3706 = _T_3684[5:0] == 6'h6; // @[el2_lib.scala 307:41]
  wire  _T_3704 = _T_3684[5:0] == 6'h5; // @[el2_lib.scala 307:41]
  wire  _T_3702 = _T_3684[5:0] == 6'h4; // @[el2_lib.scala 307:41]
  wire  _T_3700 = _T_3684[5:0] == 6'h3; // @[el2_lib.scala 307:41]
  wire  _T_3698 = _T_3684[5:0] == 6'h2; // @[el2_lib.scala 307:41]
  wire  _T_3696 = _T_3684[5:0] == 6'h1; // @[el2_lib.scala 307:41]
  wire [18:0] _T_3812 = {_T_3811,_T_3712,_T_3710,_T_3708,_T_3706,_T_3704,_T_3702,_T_3700,_T_3698,_T_3696}; // @[el2_lib.scala 310:69]
  wire [38:0] _T_3832 = {_T_3830,_T_3821,_T_3812}; // @[el2_lib.scala 310:69]
  wire [7:0] _T_3787 = {io_iccm_rd_data_ecc[74],io_iccm_rd_data_ecc[42:40],io_iccm_rd_data_ecc[73],io_iccm_rd_data_ecc[39],io_iccm_rd_data_ecc[72:71]}; // @[Cat.scala 29:58]
  wire [38:0] _T_3793 = {io_iccm_rd_data_ecc[77],io_iccm_rd_data_ecc[70:65],io_iccm_rd_data_ecc[76],io_iccm_rd_data_ecc[64:50],io_iccm_rd_data_ecc[75],io_iccm_rd_data_ecc[49:43],_T_3787}; // @[Cat.scala 29:58]
  wire [38:0] _T_3833 = _T_3832 ^ _T_3793; // @[el2_lib.scala 310:76]
  wire [38:0] _T_3834 = _T_3688 ? _T_3833 : _T_3793; // @[el2_lib.scala 310:31]
  wire [31:0] iccm_corrected_data_1 = {_T_3834[37:32],_T_3834[30:16],_T_3834[14:8],_T_3834[6:4],_T_3834[2]}; // @[Cat.scala 29:58]
  wire [31:0] iccm_dma_rdata_1_muxed = dma_mem_addr_ff[0] ? iccm_corrected_data_0 : iccm_corrected_data_1; // @[el2_ifu_mem_ctl.scala 647:35]
  wire  _T_3307 = ~_T_3299[6]; // @[el2_lib.scala 303:55]
  wire  _T_3308 = _T_3301 & _T_3307; // @[el2_lib.scala 303:53]
  wire  _T_3692 = ~_T_3684[6]; // @[el2_lib.scala 303:55]
  wire  _T_3693 = _T_3686 & _T_3692; // @[el2_lib.scala 303:53]
  wire [1:0] iccm_double_ecc_error = {_T_3308,_T_3693}; // @[Cat.scala 29:58]
  wire  iccm_dma_ecc_error_in = |iccm_double_ecc_error; // @[el2_ifu_mem_ctl.scala 649:53]
  wire [63:0] _T_3059 = {io_dma_mem_addr,io_dma_mem_addr}; // @[Cat.scala 29:58]
  wire [63:0] _T_3060 = {iccm_dma_rdata_1_muxed,_T_3449[37:32],_T_3449[30:16],_T_3449[14:8],_T_3449[6:4],_T_3449[2]}; // @[Cat.scala 29:58]
  reg [2:0] dma_mem_tag_ff; // @[el2_ifu_mem_ctl.scala 651:54]
  reg [2:0] iccm_dma_rtag; // @[el2_ifu_mem_ctl.scala 652:69]
  reg  iccm_dma_rvalid; // @[el2_ifu_mem_ctl.scala 657:71]
  reg [63:0] iccm_dma_rdata; // @[el2_ifu_mem_ctl.scala 661:70]
  wire  _T_3065 = _T_2640 & _T_2629; // @[el2_ifu_mem_ctl.scala 664:65]
  wire  _T_3068 = _T_3046 & iccm_correct_ecc; // @[el2_ifu_mem_ctl.scala 665:50]
  reg [13:0] iccm_ecc_corr_index_ff; // @[Reg.scala 27:20]
  wire [14:0] _T_3069 = {iccm_ecc_corr_index_ff,1'h0}; // @[Cat.scala 29:58]
  wire [15:0] _T_3071 = _T_3068 ? {{1'd0}, _T_3069} : io_ifc_fetch_addr_bf[15:0]; // @[el2_ifu_mem_ctl.scala 665:8]
  wire [31:0] _T_3072 = _T_3065 ? io_dma_mem_addr : {{16'd0}, _T_3071}; // @[el2_ifu_mem_ctl.scala 664:25]
  wire  _T_3461 = _T_3299 == 7'h40; // @[el2_lib.scala 313:62]
  wire  _T_3462 = _T_3449[38] ^ _T_3461; // @[el2_lib.scala 313:44]
  wire [6:0] iccm_corrected_ecc_0 = {_T_3462,_T_3449[31],_T_3449[15],_T_3449[7],_T_3449[3],_T_3449[1:0]}; // @[Cat.scala 29:58]
  wire  _T_3846 = _T_3684 == 7'h40; // @[el2_lib.scala 313:62]
  wire  _T_3847 = _T_3834[38] ^ _T_3846; // @[el2_lib.scala 313:44]
  wire [6:0] iccm_corrected_ecc_1 = {_T_3847,_T_3834[31],_T_3834[15],_T_3834[7],_T_3834[3],_T_3834[1:0]}; // @[Cat.scala 29:58]
  wire  _T_3863 = _T_3 & ifc_iccm_access_f; // @[el2_ifu_mem_ctl.scala 677:58]
  wire [31:0] iccm_corrected_data_f_mux = iccm_single_ecc_error[0] ? iccm_corrected_data_0 : iccm_corrected_data_1; // @[el2_ifu_mem_ctl.scala 679:38]
  wire [6:0] iccm_corrected_ecc_f_mux = iccm_single_ecc_error[0] ? iccm_corrected_ecc_0 : iccm_corrected_ecc_1; // @[el2_ifu_mem_ctl.scala 680:37]
  reg  iccm_rd_ecc_single_err_ff; // @[el2_ifu_mem_ctl.scala 688:62]
  wire  _T_3871 = ~iccm_rd_ecc_single_err_ff; // @[el2_ifu_mem_ctl.scala 682:76]
  wire  _T_3872 = io_iccm_rd_ecc_single_err & _T_3871; // @[el2_ifu_mem_ctl.scala 682:74]
  wire  _T_3874 = _T_3872 & _T_317; // @[el2_ifu_mem_ctl.scala 682:104]
  wire  iccm_ecc_write_status = _T_3874 | io_iccm_dma_sb_error; // @[el2_ifu_mem_ctl.scala 682:127]
  wire  _T_3875 = io_iccm_rd_ecc_single_err | iccm_rd_ecc_single_err_ff; // @[el2_ifu_mem_ctl.scala 683:67]
  wire  iccm_rd_ecc_single_err_hold_in = _T_3875 & _T_317; // @[el2_ifu_mem_ctl.scala 683:96]
  reg [13:0] iccm_rw_addr_f; // @[el2_ifu_mem_ctl.scala 687:51]
  wire [13:0] _T_3880 = iccm_rw_addr_f + 14'h1; // @[el2_ifu_mem_ctl.scala 686:102]
  wire [38:0] _T_3884 = {iccm_corrected_ecc_f_mux,iccm_corrected_data_f_mux}; // @[Cat.scala 29:58]
  wire  _T_3889 = ~io_ifc_fetch_uncacheable_bf; // @[el2_ifu_mem_ctl.scala 691:41]
  wire  _T_3890 = io_ifc_fetch_req_bf & _T_3889; // @[el2_ifu_mem_ctl.scala 691:39]
  wire  _T_3891 = ~io_ifc_iccm_access_bf; // @[el2_ifu_mem_ctl.scala 691:72]
  wire  _T_3892 = _T_3890 & _T_3891; // @[el2_ifu_mem_ctl.scala 691:70]
  wire  _T_3894 = ~miss_state_en; // @[el2_ifu_mem_ctl.scala 692:34]
  wire  _T_3895 = _T_2235 & _T_3894; // @[el2_ifu_mem_ctl.scala 692:32]
  wire  _T_3898 = _T_2251 & _T_3894; // @[el2_ifu_mem_ctl.scala 693:37]
  wire  _T_3899 = _T_3895 | _T_3898; // @[el2_ifu_mem_ctl.scala 692:88]
  wire  _T_3900 = miss_state == 3'h7; // @[el2_ifu_mem_ctl.scala 694:19]
  wire  _T_3902 = _T_3900 & _T_3894; // @[el2_ifu_mem_ctl.scala 694:41]
  wire  _T_3903 = _T_3899 | _T_3902; // @[el2_ifu_mem_ctl.scala 693:88]
  wire  _T_3904 = miss_state == 3'h3; // @[el2_ifu_mem_ctl.scala 695:19]
  wire  _T_3906 = _T_3904 & _T_3894; // @[el2_ifu_mem_ctl.scala 695:35]
  wire  _T_3907 = _T_3903 | _T_3906; // @[el2_ifu_mem_ctl.scala 694:88]
  wire  _T_3910 = _T_2250 & _T_3894; // @[el2_ifu_mem_ctl.scala 696:38]
  wire  _T_3911 = _T_3907 | _T_3910; // @[el2_ifu_mem_ctl.scala 695:88]
  wire  _T_3913 = _T_2251 & miss_state_en; // @[el2_ifu_mem_ctl.scala 697:37]
  wire  _T_3914 = miss_nxtstate == 3'h3; // @[el2_ifu_mem_ctl.scala 697:71]
  wire  _T_3915 = _T_3913 & _T_3914; // @[el2_ifu_mem_ctl.scala 697:54]
  wire  _T_3916 = _T_3911 | _T_3915; // @[el2_ifu_mem_ctl.scala 696:57]
  wire  _T_3917 = ~_T_3916; // @[el2_ifu_mem_ctl.scala 692:5]
  wire  _T_3918 = _T_3892 & _T_3917; // @[el2_ifu_mem_ctl.scala 691:96]
  wire  _T_3919 = io_ifc_fetch_req_bf & io_exu_flush_final; // @[el2_ifu_mem_ctl.scala 698:28]
  wire  _T_3921 = _T_3919 & _T_3889; // @[el2_ifu_mem_ctl.scala 698:50]
  wire  _T_3923 = _T_3921 & _T_3891; // @[el2_ifu_mem_ctl.scala 698:81]
  wire  _T_3932 = ~_T_108; // @[el2_ifu_mem_ctl.scala 701:106]
  wire  _T_3933 = _T_2235 & _T_3932; // @[el2_ifu_mem_ctl.scala 701:104]
  wire  _T_3934 = _T_2251 | _T_3933; // @[el2_ifu_mem_ctl.scala 701:77]
  wire  _T_3938 = ~_T_51; // @[el2_ifu_mem_ctl.scala 701:172]
  wire  _T_3939 = _T_3934 & _T_3938; // @[el2_ifu_mem_ctl.scala 701:170]
  wire  _T_3940 = ~_T_3939; // @[el2_ifu_mem_ctl.scala 701:44]
  wire  _T_3944 = reset_ic_in | reset_ic_ff; // @[el2_ifu_mem_ctl.scala 704:64]
  wire  _T_3945 = ~_T_3944; // @[el2_ifu_mem_ctl.scala 704:50]
  wire  _T_3946 = _T_276 & _T_3945; // @[el2_ifu_mem_ctl.scala 704:48]
  wire  _T_3947 = ~reset_tag_valid_for_miss; // @[el2_ifu_mem_ctl.scala 704:81]
  wire  ic_valid = _T_3946 & _T_3947; // @[el2_ifu_mem_ctl.scala 704:79]
  wire  _T_3949 = debug_c1_clken & io_ic_debug_tag_array; // @[el2_ifu_mem_ctl.scala 705:82]
  reg [6:0] ifu_status_wr_addr_ff; // @[el2_ifu_mem_ctl.scala 708:14]
  wire  _T_3952 = io_ic_debug_wr_en & io_ic_debug_tag_array; // @[el2_ifu_mem_ctl.scala 711:74]
  wire  _T_10094 = bus_ifu_wr_en_ff_q & last_beat; // @[el2_ifu_mem_ctl.scala 785:45]
  wire  way_status_wr_en = _T_10094 | ic_act_hit_f; // @[el2_ifu_mem_ctl.scala 785:58]
  wire  way_status_wr_en_w_debug = way_status_wr_en | _T_3952; // @[el2_ifu_mem_ctl.scala 711:53]
  reg  way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 713:14]
  wire [2:0] _T_3956 = {{2'd0}, io_ic_debug_wr_data[4]}; // @[el2_ifu_mem_ctl.scala 717:10]
  wire  way_status_hit_new = io_ic_rd_hit[0]; // @[el2_ifu_mem_ctl.scala 781:41]
  wire  way_status_new = _T_10094 ? replace_way_mb_any_0 : way_status_hit_new; // @[el2_ifu_mem_ctl.scala 784:26]
  reg [2:0] way_status_new_ff; // @[el2_ifu_mem_ctl.scala 719:14]
  wire  way_status_clken_0 = ifu_status_wr_addr_ff[6:3] == 4'h0; // @[el2_ifu_mem_ctl.scala 721:132]
  wire  way_status_clken_1 = ifu_status_wr_addr_ff[6:3] == 4'h1; // @[el2_ifu_mem_ctl.scala 721:132]
  wire  way_status_clken_2 = ifu_status_wr_addr_ff[6:3] == 4'h2; // @[el2_ifu_mem_ctl.scala 721:132]
  wire  way_status_clken_3 = ifu_status_wr_addr_ff[6:3] == 4'h3; // @[el2_ifu_mem_ctl.scala 721:132]
  wire  way_status_clken_4 = ifu_status_wr_addr_ff[6:3] == 4'h4; // @[el2_ifu_mem_ctl.scala 721:132]
  wire  way_status_clken_5 = ifu_status_wr_addr_ff[6:3] == 4'h5; // @[el2_ifu_mem_ctl.scala 721:132]
  wire  way_status_clken_6 = ifu_status_wr_addr_ff[6:3] == 4'h6; // @[el2_ifu_mem_ctl.scala 721:132]
  wire  way_status_clken_7 = ifu_status_wr_addr_ff[6:3] == 4'h7; // @[el2_ifu_mem_ctl.scala 721:132]
  wire  way_status_clken_8 = ifu_status_wr_addr_ff[6:3] == 4'h8; // @[el2_ifu_mem_ctl.scala 721:132]
  wire  way_status_clken_9 = ifu_status_wr_addr_ff[6:3] == 4'h9; // @[el2_ifu_mem_ctl.scala 721:132]
  wire  way_status_clken_10 = ifu_status_wr_addr_ff[6:3] == 4'ha; // @[el2_ifu_mem_ctl.scala 721:132]
  wire  way_status_clken_11 = ifu_status_wr_addr_ff[6:3] == 4'hb; // @[el2_ifu_mem_ctl.scala 721:132]
  wire  way_status_clken_12 = ifu_status_wr_addr_ff[6:3] == 4'hc; // @[el2_ifu_mem_ctl.scala 721:132]
  wire  way_status_clken_13 = ifu_status_wr_addr_ff[6:3] == 4'hd; // @[el2_ifu_mem_ctl.scala 721:132]
  wire  way_status_clken_14 = ifu_status_wr_addr_ff[6:3] == 4'he; // @[el2_ifu_mem_ctl.scala 721:132]
  wire  way_status_clken_15 = ifu_status_wr_addr_ff[6:3] == 4'hf; // @[el2_ifu_mem_ctl.scala 721:132]
  wire  _T_3973 = ifu_status_wr_addr_ff == 7'h0; // @[el2_ifu_mem_ctl.scala 725:93]
  wire  _T_3974 = _T_3973 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 725:102]
  wire  _T_3975 = _T_3974 & way_status_clken_0; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_3977 = ifu_status_wr_addr_ff == 7'h1; // @[el2_ifu_mem_ctl.scala 725:93]
  wire  _T_3978 = _T_3977 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 725:102]
  wire  _T_3979 = _T_3978 & way_status_clken_0; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_3981 = ifu_status_wr_addr_ff == 7'h2; // @[el2_ifu_mem_ctl.scala 725:93]
  wire  _T_3982 = _T_3981 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 725:102]
  wire  _T_3983 = _T_3982 & way_status_clken_0; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_3985 = ifu_status_wr_addr_ff == 7'h3; // @[el2_ifu_mem_ctl.scala 725:93]
  wire  _T_3986 = _T_3985 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 725:102]
  wire  _T_3987 = _T_3986 & way_status_clken_0; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_3989 = ifu_status_wr_addr_ff == 7'h4; // @[el2_ifu_mem_ctl.scala 725:93]
  wire  _T_3990 = _T_3989 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 725:102]
  wire  _T_3991 = _T_3990 & way_status_clken_0; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_3993 = ifu_status_wr_addr_ff == 7'h5; // @[el2_ifu_mem_ctl.scala 725:93]
  wire  _T_3994 = _T_3993 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 725:102]
  wire  _T_3995 = _T_3994 & way_status_clken_0; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_3997 = ifu_status_wr_addr_ff == 7'h6; // @[el2_ifu_mem_ctl.scala 725:93]
  wire  _T_3998 = _T_3997 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 725:102]
  wire  _T_3999 = _T_3998 & way_status_clken_0; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4001 = ifu_status_wr_addr_ff == 7'h7; // @[el2_ifu_mem_ctl.scala 725:93]
  wire  _T_4002 = _T_4001 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 725:102]
  wire  _T_4003 = _T_4002 & way_status_clken_0; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4007 = _T_3974 & way_status_clken_1; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4011 = _T_3978 & way_status_clken_1; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4015 = _T_3982 & way_status_clken_1; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4019 = _T_3986 & way_status_clken_1; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4023 = _T_3990 & way_status_clken_1; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4027 = _T_3994 & way_status_clken_1; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4031 = _T_3998 & way_status_clken_1; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4035 = _T_4002 & way_status_clken_1; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4039 = _T_3974 & way_status_clken_2; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4043 = _T_3978 & way_status_clken_2; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4047 = _T_3982 & way_status_clken_2; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4051 = _T_3986 & way_status_clken_2; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4055 = _T_3990 & way_status_clken_2; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4059 = _T_3994 & way_status_clken_2; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4063 = _T_3998 & way_status_clken_2; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4067 = _T_4002 & way_status_clken_2; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4071 = _T_3974 & way_status_clken_3; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4075 = _T_3978 & way_status_clken_3; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4079 = _T_3982 & way_status_clken_3; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4083 = _T_3986 & way_status_clken_3; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4087 = _T_3990 & way_status_clken_3; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4091 = _T_3994 & way_status_clken_3; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4095 = _T_3998 & way_status_clken_3; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4099 = _T_4002 & way_status_clken_3; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4103 = _T_3974 & way_status_clken_4; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4107 = _T_3978 & way_status_clken_4; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4111 = _T_3982 & way_status_clken_4; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4115 = _T_3986 & way_status_clken_4; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4119 = _T_3990 & way_status_clken_4; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4123 = _T_3994 & way_status_clken_4; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4127 = _T_3998 & way_status_clken_4; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4131 = _T_4002 & way_status_clken_4; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4135 = _T_3974 & way_status_clken_5; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4139 = _T_3978 & way_status_clken_5; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4143 = _T_3982 & way_status_clken_5; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4147 = _T_3986 & way_status_clken_5; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4151 = _T_3990 & way_status_clken_5; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4155 = _T_3994 & way_status_clken_5; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4159 = _T_3998 & way_status_clken_5; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4163 = _T_4002 & way_status_clken_5; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4167 = _T_3974 & way_status_clken_6; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4171 = _T_3978 & way_status_clken_6; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4175 = _T_3982 & way_status_clken_6; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4179 = _T_3986 & way_status_clken_6; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4183 = _T_3990 & way_status_clken_6; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4187 = _T_3994 & way_status_clken_6; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4191 = _T_3998 & way_status_clken_6; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4195 = _T_4002 & way_status_clken_6; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4199 = _T_3974 & way_status_clken_7; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4203 = _T_3978 & way_status_clken_7; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4207 = _T_3982 & way_status_clken_7; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4211 = _T_3986 & way_status_clken_7; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4215 = _T_3990 & way_status_clken_7; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4219 = _T_3994 & way_status_clken_7; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4223 = _T_3998 & way_status_clken_7; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4227 = _T_4002 & way_status_clken_7; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4231 = _T_3974 & way_status_clken_8; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4235 = _T_3978 & way_status_clken_8; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4239 = _T_3982 & way_status_clken_8; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4243 = _T_3986 & way_status_clken_8; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4247 = _T_3990 & way_status_clken_8; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4251 = _T_3994 & way_status_clken_8; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4255 = _T_3998 & way_status_clken_8; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4259 = _T_4002 & way_status_clken_8; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4263 = _T_3974 & way_status_clken_9; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4267 = _T_3978 & way_status_clken_9; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4271 = _T_3982 & way_status_clken_9; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4275 = _T_3986 & way_status_clken_9; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4279 = _T_3990 & way_status_clken_9; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4283 = _T_3994 & way_status_clken_9; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4287 = _T_3998 & way_status_clken_9; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4291 = _T_4002 & way_status_clken_9; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4295 = _T_3974 & way_status_clken_10; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4299 = _T_3978 & way_status_clken_10; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4303 = _T_3982 & way_status_clken_10; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4307 = _T_3986 & way_status_clken_10; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4311 = _T_3990 & way_status_clken_10; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4315 = _T_3994 & way_status_clken_10; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4319 = _T_3998 & way_status_clken_10; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4323 = _T_4002 & way_status_clken_10; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4327 = _T_3974 & way_status_clken_11; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4331 = _T_3978 & way_status_clken_11; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4335 = _T_3982 & way_status_clken_11; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4339 = _T_3986 & way_status_clken_11; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4343 = _T_3990 & way_status_clken_11; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4347 = _T_3994 & way_status_clken_11; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4351 = _T_3998 & way_status_clken_11; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4355 = _T_4002 & way_status_clken_11; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4359 = _T_3974 & way_status_clken_12; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4363 = _T_3978 & way_status_clken_12; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4367 = _T_3982 & way_status_clken_12; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4371 = _T_3986 & way_status_clken_12; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4375 = _T_3990 & way_status_clken_12; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4379 = _T_3994 & way_status_clken_12; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4383 = _T_3998 & way_status_clken_12; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4387 = _T_4002 & way_status_clken_12; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4391 = _T_3974 & way_status_clken_13; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4395 = _T_3978 & way_status_clken_13; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4399 = _T_3982 & way_status_clken_13; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4403 = _T_3986 & way_status_clken_13; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4407 = _T_3990 & way_status_clken_13; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4411 = _T_3994 & way_status_clken_13; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4415 = _T_3998 & way_status_clken_13; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4419 = _T_4002 & way_status_clken_13; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4423 = _T_3974 & way_status_clken_14; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4427 = _T_3978 & way_status_clken_14; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4431 = _T_3982 & way_status_clken_14; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4435 = _T_3986 & way_status_clken_14; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4439 = _T_3990 & way_status_clken_14; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4443 = _T_3994 & way_status_clken_14; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4447 = _T_3998 & way_status_clken_14; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4451 = _T_4002 & way_status_clken_14; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4455 = _T_3974 & way_status_clken_15; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4459 = _T_3978 & way_status_clken_15; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4463 = _T_3982 & way_status_clken_15; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4467 = _T_3986 & way_status_clken_15; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4471 = _T_3990 & way_status_clken_15; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4475 = _T_3994 & way_status_clken_15; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4479 = _T_3998 & way_status_clken_15; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_4483 = _T_4002 & way_status_clken_15; // @[el2_ifu_mem_ctl.scala 725:124]
  wire  _T_10100 = _T_100 & replace_way_mb_any_1; // @[el2_ifu_mem_ctl.scala 788:84]
  wire  _T_10101 = _T_10100 & miss_pending; // @[el2_ifu_mem_ctl.scala 788:108]
  wire  bus_wren_last_1 = _T_10101 & bus_last_data_beat; // @[el2_ifu_mem_ctl.scala 788:123]
  wire  wren_reset_miss_1 = replace_way_mb_any_1 & reset_tag_valid_for_miss; // @[el2_ifu_mem_ctl.scala 789:84]
  wire  _T_10103 = bus_wren_last_1 | wren_reset_miss_1; // @[el2_ifu_mem_ctl.scala 790:73]
  wire  _T_10098 = _T_100 & replace_way_mb_any_0; // @[el2_ifu_mem_ctl.scala 788:84]
  wire  _T_10099 = _T_10098 & miss_pending; // @[el2_ifu_mem_ctl.scala 788:108]
  wire  bus_wren_last_0 = _T_10099 & bus_last_data_beat; // @[el2_ifu_mem_ctl.scala 788:123]
  wire  wren_reset_miss_0 = replace_way_mb_any_0 & reset_tag_valid_for_miss; // @[el2_ifu_mem_ctl.scala 789:84]
  wire  _T_10102 = bus_wren_last_0 | wren_reset_miss_0; // @[el2_ifu_mem_ctl.scala 790:73]
  wire [1:0] ifu_tag_wren = {_T_10103,_T_10102}; // @[Cat.scala 29:58]
  wire [1:0] _T_10137 = _T_3952 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [1:0] ic_debug_tag_wr_en = _T_10137 & io_ic_debug_way; // @[el2_ifu_mem_ctl.scala 823:90]
  wire [1:0] ifu_tag_wren_w_debug = ifu_tag_wren | ic_debug_tag_wr_en; // @[el2_ifu_mem_ctl.scala 734:45]
  reg [1:0] ifu_tag_wren_ff; // @[el2_ifu_mem_ctl.scala 736:14]
  reg  ic_valid_ff; // @[el2_ifu_mem_ctl.scala 740:14]
  wire  _T_5132 = ifu_ic_rw_int_addr_ff[5:4] == 2'h0; // @[el2_ifu_mem_ctl.scala 744:82]
  wire  _T_5134 = _T_5132 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 744:91]
  wire  _T_5136 = perr_ic_index_ff[5:4] == 2'h0; // @[el2_ifu_mem_ctl.scala 745:74]
  wire  _T_5138 = _T_5136 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 745:83]
  wire  _T_5139 = _T_5134 | _T_5138; // @[el2_ifu_mem_ctl.scala 744:113]
  wire  _T_5140 = _T_5139 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 745:106]
  wire  _T_5144 = _T_5132 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 744:91]
  wire  _T_5148 = _T_5136 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 745:83]
  wire  _T_5149 = _T_5144 | _T_5148; // @[el2_ifu_mem_ctl.scala 744:113]
  wire  _T_5150 = _T_5149 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 745:106]
  wire [1:0] tag_valid_clken_0 = {_T_5140,_T_5150}; // @[Cat.scala 29:58]
  wire  _T_5152 = ifu_ic_rw_int_addr_ff[5:4] == 2'h1; // @[el2_ifu_mem_ctl.scala 744:82]
  wire  _T_5154 = _T_5152 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 744:91]
  wire  _T_5156 = perr_ic_index_ff[5:4] == 2'h1; // @[el2_ifu_mem_ctl.scala 745:74]
  wire  _T_5158 = _T_5156 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 745:83]
  wire  _T_5159 = _T_5154 | _T_5158; // @[el2_ifu_mem_ctl.scala 744:113]
  wire  _T_5160 = _T_5159 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 745:106]
  wire  _T_5164 = _T_5152 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 744:91]
  wire  _T_5168 = _T_5156 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 745:83]
  wire  _T_5169 = _T_5164 | _T_5168; // @[el2_ifu_mem_ctl.scala 744:113]
  wire  _T_5170 = _T_5169 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 745:106]
  wire [1:0] tag_valid_clken_1 = {_T_5160,_T_5170}; // @[Cat.scala 29:58]
  wire  _T_5172 = ifu_ic_rw_int_addr_ff[5:4] == 2'h2; // @[el2_ifu_mem_ctl.scala 744:82]
  wire  _T_5174 = _T_5172 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 744:91]
  wire  _T_5176 = perr_ic_index_ff[5:4] == 2'h2; // @[el2_ifu_mem_ctl.scala 745:74]
  wire  _T_5178 = _T_5176 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 745:83]
  wire  _T_5179 = _T_5174 | _T_5178; // @[el2_ifu_mem_ctl.scala 744:113]
  wire  _T_5180 = _T_5179 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 745:106]
  wire  _T_5184 = _T_5172 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 744:91]
  wire  _T_5188 = _T_5176 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 745:83]
  wire  _T_5189 = _T_5184 | _T_5188; // @[el2_ifu_mem_ctl.scala 744:113]
  wire  _T_5190 = _T_5189 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 745:106]
  wire [1:0] tag_valid_clken_2 = {_T_5180,_T_5190}; // @[Cat.scala 29:58]
  wire  _T_5192 = ifu_ic_rw_int_addr_ff[5:4] == 2'h3; // @[el2_ifu_mem_ctl.scala 744:82]
  wire  _T_5194 = _T_5192 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 744:91]
  wire  _T_5196 = perr_ic_index_ff[5:4] == 2'h3; // @[el2_ifu_mem_ctl.scala 745:74]
  wire  _T_5198 = _T_5196 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 745:83]
  wire  _T_5199 = _T_5194 | _T_5198; // @[el2_ifu_mem_ctl.scala 744:113]
  wire  _T_5200 = _T_5199 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 745:106]
  wire  _T_5204 = _T_5192 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 744:91]
  wire  _T_5208 = _T_5196 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 745:83]
  wire  _T_5209 = _T_5204 | _T_5208; // @[el2_ifu_mem_ctl.scala 744:113]
  wire  _T_5210 = _T_5209 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 745:106]
  wire [1:0] tag_valid_clken_3 = {_T_5200,_T_5210}; // @[Cat.scala 29:58]
  wire  _T_5213 = ic_valid_ff & _T_195; // @[el2_ifu_mem_ctl.scala 750:64]
  wire  _T_5214 = ~perr_sel_invalidate; // @[el2_ifu_mem_ctl.scala 750:91]
  wire  _T_5215 = _T_5213 & _T_5214; // @[el2_ifu_mem_ctl.scala 750:89]
  wire  _T_5218 = _T_4485 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_5219 = perr_ic_index_ff == 6'h0; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_5221 = _T_5219 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_5223 = _T_5221 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_5224 = _T_5218 | _T_5223; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_5234 = _T_4489 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_5235 = perr_ic_index_ff == 6'h1; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_5237 = _T_5235 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_5239 = _T_5237 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_5240 = _T_5234 | _T_5239; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_5250 = _T_4493 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_5251 = perr_ic_index_ff == 6'h2; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_5253 = _T_5251 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_5255 = _T_5253 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_5256 = _T_5250 | _T_5255; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_5266 = _T_4497 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_5267 = perr_ic_index_ff == 6'h3; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_5269 = _T_5267 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_5271 = _T_5269 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_5272 = _T_5266 | _T_5271; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_5282 = _T_4501 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_5283 = perr_ic_index_ff == 6'h4; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_5285 = _T_5283 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_5287 = _T_5285 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_5288 = _T_5282 | _T_5287; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_5298 = _T_4505 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_5299 = perr_ic_index_ff == 6'h5; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_5301 = _T_5299 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_5303 = _T_5301 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_5304 = _T_5298 | _T_5303; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_5314 = _T_4509 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_5315 = perr_ic_index_ff == 6'h6; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_5317 = _T_5315 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_5319 = _T_5317 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_5320 = _T_5314 | _T_5319; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_5330 = _T_4513 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_5331 = perr_ic_index_ff == 6'h7; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_5333 = _T_5331 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_5335 = _T_5333 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_5336 = _T_5330 | _T_5335; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_5346 = _T_4517 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_5347 = perr_ic_index_ff == 6'h8; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_5349 = _T_5347 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_5351 = _T_5349 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_5352 = _T_5346 | _T_5351; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_5362 = _T_4521 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_5363 = perr_ic_index_ff == 6'h9; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_5365 = _T_5363 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_5367 = _T_5365 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_5368 = _T_5362 | _T_5367; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_5378 = _T_4525 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_5379 = perr_ic_index_ff == 6'ha; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_5381 = _T_5379 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_5383 = _T_5381 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_5384 = _T_5378 | _T_5383; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_5394 = _T_4529 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_5395 = perr_ic_index_ff == 6'hb; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_5397 = _T_5395 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_5399 = _T_5397 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_5400 = _T_5394 | _T_5399; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_5410 = _T_4533 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_5411 = perr_ic_index_ff == 6'hc; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_5413 = _T_5411 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_5415 = _T_5413 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_5416 = _T_5410 | _T_5415; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_5426 = _T_4537 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_5427 = perr_ic_index_ff == 6'hd; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_5429 = _T_5427 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_5431 = _T_5429 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_5432 = _T_5426 | _T_5431; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_5442 = _T_4541 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_5443 = perr_ic_index_ff == 6'he; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_5445 = _T_5443 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_5447 = _T_5445 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_5448 = _T_5442 | _T_5447; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_5458 = _T_4545 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_5459 = perr_ic_index_ff == 6'hf; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_5461 = _T_5459 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_5463 = _T_5461 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_5464 = _T_5458 | _T_5463; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_5474 = _T_4549 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_5475 = perr_ic_index_ff == 6'h10; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_5477 = _T_5475 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_5479 = _T_5477 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_5480 = _T_5474 | _T_5479; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_5490 = _T_4553 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_5491 = perr_ic_index_ff == 6'h11; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_5493 = _T_5491 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_5495 = _T_5493 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_5496 = _T_5490 | _T_5495; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_5506 = _T_4557 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_5507 = perr_ic_index_ff == 6'h12; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_5509 = _T_5507 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_5511 = _T_5509 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_5512 = _T_5506 | _T_5511; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_5522 = _T_4561 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_5523 = perr_ic_index_ff == 6'h13; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_5525 = _T_5523 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_5527 = _T_5525 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_5528 = _T_5522 | _T_5527; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_5538 = _T_4565 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_5539 = perr_ic_index_ff == 6'h14; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_5541 = _T_5539 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_5543 = _T_5541 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_5544 = _T_5538 | _T_5543; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_5554 = _T_4569 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_5555 = perr_ic_index_ff == 6'h15; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_5557 = _T_5555 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_5559 = _T_5557 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_5560 = _T_5554 | _T_5559; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_5570 = _T_4573 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_5571 = perr_ic_index_ff == 6'h16; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_5573 = _T_5571 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_5575 = _T_5573 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_5576 = _T_5570 | _T_5575; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_5586 = _T_4577 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_5587 = perr_ic_index_ff == 6'h17; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_5589 = _T_5587 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_5591 = _T_5589 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_5592 = _T_5586 | _T_5591; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_5602 = _T_4581 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_5603 = perr_ic_index_ff == 6'h18; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_5605 = _T_5603 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_5607 = _T_5605 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_5608 = _T_5602 | _T_5607; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_5618 = _T_4585 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_5619 = perr_ic_index_ff == 6'h19; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_5621 = _T_5619 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_5623 = _T_5621 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_5624 = _T_5618 | _T_5623; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_5634 = _T_4589 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_5635 = perr_ic_index_ff == 6'h1a; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_5637 = _T_5635 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_5639 = _T_5637 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_5640 = _T_5634 | _T_5639; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_5650 = _T_4593 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_5651 = perr_ic_index_ff == 6'h1b; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_5653 = _T_5651 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_5655 = _T_5653 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_5656 = _T_5650 | _T_5655; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_5666 = _T_4597 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_5667 = perr_ic_index_ff == 6'h1c; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_5669 = _T_5667 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_5671 = _T_5669 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_5672 = _T_5666 | _T_5671; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_5682 = _T_4601 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_5683 = perr_ic_index_ff == 6'h1d; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_5685 = _T_5683 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_5687 = _T_5685 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_5688 = _T_5682 | _T_5687; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_5698 = _T_4605 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_5699 = perr_ic_index_ff == 6'h1e; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_5701 = _T_5699 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_5703 = _T_5701 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_5704 = _T_5698 | _T_5703; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_5714 = _T_4609 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_5715 = perr_ic_index_ff == 6'h1f; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_5717 = _T_5715 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_5719 = _T_5717 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_5720 = _T_5714 | _T_5719; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_5730 = _T_4485 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_5733 = _T_5219 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_5735 = _T_5733 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_5736 = _T_5730 | _T_5735; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_5746 = _T_4489 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_5749 = _T_5235 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_5751 = _T_5749 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_5752 = _T_5746 | _T_5751; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_5762 = _T_4493 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_5765 = _T_5251 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_5767 = _T_5765 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_5768 = _T_5762 | _T_5767; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_5778 = _T_4497 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_5781 = _T_5267 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_5783 = _T_5781 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_5784 = _T_5778 | _T_5783; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_5794 = _T_4501 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_5797 = _T_5283 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_5799 = _T_5797 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_5800 = _T_5794 | _T_5799; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_5810 = _T_4505 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_5813 = _T_5299 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_5815 = _T_5813 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_5816 = _T_5810 | _T_5815; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_5826 = _T_4509 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_5829 = _T_5315 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_5831 = _T_5829 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_5832 = _T_5826 | _T_5831; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_5842 = _T_4513 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_5845 = _T_5331 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_5847 = _T_5845 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_5848 = _T_5842 | _T_5847; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_5858 = _T_4517 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_5861 = _T_5347 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_5863 = _T_5861 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_5864 = _T_5858 | _T_5863; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_5874 = _T_4521 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_5877 = _T_5363 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_5879 = _T_5877 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_5880 = _T_5874 | _T_5879; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_5890 = _T_4525 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_5893 = _T_5379 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_5895 = _T_5893 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_5896 = _T_5890 | _T_5895; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_5906 = _T_4529 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_5909 = _T_5395 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_5911 = _T_5909 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_5912 = _T_5906 | _T_5911; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_5922 = _T_4533 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_5925 = _T_5411 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_5927 = _T_5925 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_5928 = _T_5922 | _T_5927; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_5938 = _T_4537 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_5941 = _T_5427 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_5943 = _T_5941 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_5944 = _T_5938 | _T_5943; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_5954 = _T_4541 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_5957 = _T_5443 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_5959 = _T_5957 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_5960 = _T_5954 | _T_5959; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_5970 = _T_4545 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_5973 = _T_5459 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_5975 = _T_5973 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_5976 = _T_5970 | _T_5975; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_5986 = _T_4549 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_5989 = _T_5475 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_5991 = _T_5989 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_5992 = _T_5986 | _T_5991; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_6002 = _T_4553 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_6005 = _T_5491 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_6007 = _T_6005 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_6008 = _T_6002 | _T_6007; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_6018 = _T_4557 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_6021 = _T_5507 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_6023 = _T_6021 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_6024 = _T_6018 | _T_6023; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_6034 = _T_4561 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_6037 = _T_5523 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_6039 = _T_6037 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_6040 = _T_6034 | _T_6039; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_6050 = _T_4565 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_6053 = _T_5539 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_6055 = _T_6053 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_6056 = _T_6050 | _T_6055; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_6066 = _T_4569 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_6069 = _T_5555 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_6071 = _T_6069 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_6072 = _T_6066 | _T_6071; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_6082 = _T_4573 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_6085 = _T_5571 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_6087 = _T_6085 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_6088 = _T_6082 | _T_6087; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_6098 = _T_4577 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_6101 = _T_5587 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_6103 = _T_6101 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_6104 = _T_6098 | _T_6103; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_6114 = _T_4581 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_6117 = _T_5603 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_6119 = _T_6117 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_6120 = _T_6114 | _T_6119; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_6130 = _T_4585 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_6133 = _T_5619 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_6135 = _T_6133 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_6136 = _T_6130 | _T_6135; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_6146 = _T_4589 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_6149 = _T_5635 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_6151 = _T_6149 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_6152 = _T_6146 | _T_6151; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_6162 = _T_4593 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_6165 = _T_5651 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_6167 = _T_6165 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_6168 = _T_6162 | _T_6167; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_6178 = _T_4597 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_6181 = _T_5667 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_6183 = _T_6181 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_6184 = _T_6178 | _T_6183; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_6194 = _T_4601 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_6197 = _T_5683 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_6199 = _T_6197 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_6200 = _T_6194 | _T_6199; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_6210 = _T_4605 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_6213 = _T_5699 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_6215 = _T_6213 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_6216 = _T_6210 | _T_6215; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_6226 = _T_4609 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_6229 = _T_5715 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_6231 = _T_6229 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_6232 = _T_6226 | _T_6231; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_6242 = _T_4613 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_6243 = perr_ic_index_ff == 6'h20; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_6245 = _T_6243 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_6247 = _T_6245 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_6248 = _T_6242 | _T_6247; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_6258 = _T_4617 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_6259 = perr_ic_index_ff == 6'h21; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_6261 = _T_6259 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_6263 = _T_6261 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_6264 = _T_6258 | _T_6263; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_6274 = _T_4621 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_6275 = perr_ic_index_ff == 6'h22; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_6277 = _T_6275 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_6279 = _T_6277 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_6280 = _T_6274 | _T_6279; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_6290 = _T_4625 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_6291 = perr_ic_index_ff == 6'h23; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_6293 = _T_6291 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_6295 = _T_6293 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_6296 = _T_6290 | _T_6295; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_6306 = _T_4629 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_6307 = perr_ic_index_ff == 6'h24; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_6309 = _T_6307 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_6311 = _T_6309 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_6312 = _T_6306 | _T_6311; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_6322 = _T_4633 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_6323 = perr_ic_index_ff == 6'h25; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_6325 = _T_6323 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_6327 = _T_6325 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_6328 = _T_6322 | _T_6327; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_6338 = _T_4637 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_6339 = perr_ic_index_ff == 6'h26; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_6341 = _T_6339 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_6343 = _T_6341 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_6344 = _T_6338 | _T_6343; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_6354 = _T_4641 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_6355 = perr_ic_index_ff == 6'h27; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_6357 = _T_6355 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_6359 = _T_6357 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_6360 = _T_6354 | _T_6359; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_6370 = _T_4645 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_6371 = perr_ic_index_ff == 6'h28; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_6373 = _T_6371 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_6375 = _T_6373 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_6376 = _T_6370 | _T_6375; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_6386 = _T_4649 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_6387 = perr_ic_index_ff == 6'h29; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_6389 = _T_6387 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_6391 = _T_6389 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_6392 = _T_6386 | _T_6391; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_6402 = _T_4653 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_6403 = perr_ic_index_ff == 6'h2a; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_6405 = _T_6403 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_6407 = _T_6405 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_6408 = _T_6402 | _T_6407; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_6418 = _T_4657 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_6419 = perr_ic_index_ff == 6'h2b; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_6421 = _T_6419 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_6423 = _T_6421 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_6424 = _T_6418 | _T_6423; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_6434 = _T_4661 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_6435 = perr_ic_index_ff == 6'h2c; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_6437 = _T_6435 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_6439 = _T_6437 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_6440 = _T_6434 | _T_6439; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_6450 = _T_4665 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_6451 = perr_ic_index_ff == 6'h2d; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_6453 = _T_6451 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_6455 = _T_6453 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_6456 = _T_6450 | _T_6455; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_6466 = _T_4669 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_6467 = perr_ic_index_ff == 6'h2e; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_6469 = _T_6467 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_6471 = _T_6469 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_6472 = _T_6466 | _T_6471; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_6482 = _T_4673 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_6483 = perr_ic_index_ff == 6'h2f; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_6485 = _T_6483 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_6487 = _T_6485 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_6488 = _T_6482 | _T_6487; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_6498 = _T_4677 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_6499 = perr_ic_index_ff == 6'h30; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_6501 = _T_6499 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_6503 = _T_6501 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_6504 = _T_6498 | _T_6503; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_6514 = _T_4681 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_6515 = perr_ic_index_ff == 6'h31; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_6517 = _T_6515 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_6519 = _T_6517 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_6520 = _T_6514 | _T_6519; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_6530 = _T_4685 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_6531 = perr_ic_index_ff == 6'h32; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_6533 = _T_6531 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_6535 = _T_6533 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_6536 = _T_6530 | _T_6535; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_6546 = _T_4689 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_6547 = perr_ic_index_ff == 6'h33; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_6549 = _T_6547 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_6551 = _T_6549 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_6552 = _T_6546 | _T_6551; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_6562 = _T_4693 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_6563 = perr_ic_index_ff == 6'h34; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_6565 = _T_6563 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_6567 = _T_6565 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_6568 = _T_6562 | _T_6567; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_6578 = _T_4697 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_6579 = perr_ic_index_ff == 6'h35; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_6581 = _T_6579 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_6583 = _T_6581 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_6584 = _T_6578 | _T_6583; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_6594 = _T_4701 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_6595 = perr_ic_index_ff == 6'h36; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_6597 = _T_6595 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_6599 = _T_6597 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_6600 = _T_6594 | _T_6599; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_6610 = _T_4705 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_6611 = perr_ic_index_ff == 6'h37; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_6613 = _T_6611 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_6615 = _T_6613 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_6616 = _T_6610 | _T_6615; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_6626 = _T_4709 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_6627 = perr_ic_index_ff == 6'h38; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_6629 = _T_6627 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_6631 = _T_6629 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_6632 = _T_6626 | _T_6631; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_6642 = _T_4713 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_6643 = perr_ic_index_ff == 6'h39; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_6645 = _T_6643 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_6647 = _T_6645 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_6648 = _T_6642 | _T_6647; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_6658 = _T_4717 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_6659 = perr_ic_index_ff == 6'h3a; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_6661 = _T_6659 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_6663 = _T_6661 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_6664 = _T_6658 | _T_6663; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_6674 = _T_4721 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_6675 = perr_ic_index_ff == 6'h3b; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_6677 = _T_6675 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_6679 = _T_6677 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_6680 = _T_6674 | _T_6679; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_6690 = _T_4725 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_6691 = perr_ic_index_ff == 6'h3c; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_6693 = _T_6691 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_6695 = _T_6693 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_6696 = _T_6690 | _T_6695; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_6706 = _T_4729 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_6707 = perr_ic_index_ff == 6'h3d; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_6709 = _T_6707 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_6711 = _T_6709 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_6712 = _T_6706 | _T_6711; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_6722 = _T_4733 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_6723 = perr_ic_index_ff == 6'h3e; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_6725 = _T_6723 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_6727 = _T_6725 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_6728 = _T_6722 | _T_6727; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_6738 = _T_4737 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_6739 = perr_ic_index_ff == 6'h3f; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_6741 = _T_6739 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_6743 = _T_6741 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_6744 = _T_6738 | _T_6743; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_6754 = _T_4613 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_6757 = _T_6243 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_6759 = _T_6757 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_6760 = _T_6754 | _T_6759; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_6770 = _T_4617 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_6773 = _T_6259 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_6775 = _T_6773 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_6776 = _T_6770 | _T_6775; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_6786 = _T_4621 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_6789 = _T_6275 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_6791 = _T_6789 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_6792 = _T_6786 | _T_6791; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_6802 = _T_4625 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_6805 = _T_6291 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_6807 = _T_6805 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_6808 = _T_6802 | _T_6807; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_6818 = _T_4629 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_6821 = _T_6307 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_6823 = _T_6821 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_6824 = _T_6818 | _T_6823; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_6834 = _T_4633 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_6837 = _T_6323 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_6839 = _T_6837 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_6840 = _T_6834 | _T_6839; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_6850 = _T_4637 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_6853 = _T_6339 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_6855 = _T_6853 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_6856 = _T_6850 | _T_6855; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_6866 = _T_4641 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_6869 = _T_6355 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_6871 = _T_6869 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_6872 = _T_6866 | _T_6871; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_6882 = _T_4645 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_6885 = _T_6371 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_6887 = _T_6885 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_6888 = _T_6882 | _T_6887; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_6898 = _T_4649 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_6901 = _T_6387 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_6903 = _T_6901 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_6904 = _T_6898 | _T_6903; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_6914 = _T_4653 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_6917 = _T_6403 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_6919 = _T_6917 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_6920 = _T_6914 | _T_6919; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_6930 = _T_4657 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_6933 = _T_6419 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_6935 = _T_6933 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_6936 = _T_6930 | _T_6935; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_6946 = _T_4661 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_6949 = _T_6435 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_6951 = _T_6949 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_6952 = _T_6946 | _T_6951; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_6962 = _T_4665 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_6965 = _T_6451 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_6967 = _T_6965 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_6968 = _T_6962 | _T_6967; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_6978 = _T_4669 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_6981 = _T_6467 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_6983 = _T_6981 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_6984 = _T_6978 | _T_6983; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_6994 = _T_4673 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_6997 = _T_6483 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_6999 = _T_6997 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_7000 = _T_6994 | _T_6999; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_7010 = _T_4677 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_7013 = _T_6499 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_7015 = _T_7013 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_7016 = _T_7010 | _T_7015; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_7026 = _T_4681 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_7029 = _T_6515 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_7031 = _T_7029 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_7032 = _T_7026 | _T_7031; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_7042 = _T_4685 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_7045 = _T_6531 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_7047 = _T_7045 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_7048 = _T_7042 | _T_7047; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_7058 = _T_4689 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_7061 = _T_6547 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_7063 = _T_7061 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_7064 = _T_7058 | _T_7063; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_7074 = _T_4693 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_7077 = _T_6563 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_7079 = _T_7077 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_7080 = _T_7074 | _T_7079; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_7090 = _T_4697 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_7093 = _T_6579 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_7095 = _T_7093 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_7096 = _T_7090 | _T_7095; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_7106 = _T_4701 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_7109 = _T_6595 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_7111 = _T_7109 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_7112 = _T_7106 | _T_7111; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_7122 = _T_4705 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_7125 = _T_6611 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_7127 = _T_7125 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_7128 = _T_7122 | _T_7127; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_7138 = _T_4709 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_7141 = _T_6627 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_7143 = _T_7141 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_7144 = _T_7138 | _T_7143; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_7154 = _T_4713 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_7157 = _T_6643 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_7159 = _T_7157 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_7160 = _T_7154 | _T_7159; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_7170 = _T_4717 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_7173 = _T_6659 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_7175 = _T_7173 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_7176 = _T_7170 | _T_7175; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_7186 = _T_4721 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_7189 = _T_6675 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_7191 = _T_7189 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_7192 = _T_7186 | _T_7191; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_7202 = _T_4725 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_7205 = _T_6691 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_7207 = _T_7205 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_7208 = _T_7202 | _T_7207; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_7218 = _T_4729 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_7221 = _T_6707 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_7223 = _T_7221 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_7224 = _T_7218 | _T_7223; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_7234 = _T_4733 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_7237 = _T_6723 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_7239 = _T_7237 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_7240 = _T_7234 | _T_7239; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_7250 = _T_4737 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_7253 = _T_6739 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_7255 = _T_7253 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_7256 = _T_7250 | _T_7255; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_7266 = _T_4741 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire [6:0] _GEN_796 = {{1'd0}, perr_ic_index_ff}; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_7267 = _GEN_796 == 7'h40; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_7269 = _T_7267 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_7271 = _T_7269 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_7272 = _T_7266 | _T_7271; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_7282 = _T_4745 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_7283 = _GEN_796 == 7'h41; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_7285 = _T_7283 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_7287 = _T_7285 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_7288 = _T_7282 | _T_7287; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_7298 = _T_4749 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_7299 = _GEN_796 == 7'h42; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_7301 = _T_7299 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_7303 = _T_7301 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_7304 = _T_7298 | _T_7303; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_7314 = _T_4753 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_7315 = _GEN_796 == 7'h43; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_7317 = _T_7315 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_7319 = _T_7317 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_7320 = _T_7314 | _T_7319; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_7330 = _T_4757 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_7331 = _GEN_796 == 7'h44; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_7333 = _T_7331 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_7335 = _T_7333 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_7336 = _T_7330 | _T_7335; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_7346 = _T_4761 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_7347 = _GEN_796 == 7'h45; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_7349 = _T_7347 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_7351 = _T_7349 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_7352 = _T_7346 | _T_7351; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_7362 = _T_4765 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_7363 = _GEN_796 == 7'h46; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_7365 = _T_7363 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_7367 = _T_7365 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_7368 = _T_7362 | _T_7367; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_7378 = _T_4769 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_7379 = _GEN_796 == 7'h47; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_7381 = _T_7379 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_7383 = _T_7381 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_7384 = _T_7378 | _T_7383; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_7394 = _T_4773 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_7395 = _GEN_796 == 7'h48; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_7397 = _T_7395 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_7399 = _T_7397 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_7400 = _T_7394 | _T_7399; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_7410 = _T_4777 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_7411 = _GEN_796 == 7'h49; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_7413 = _T_7411 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_7415 = _T_7413 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_7416 = _T_7410 | _T_7415; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_7426 = _T_4781 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_7427 = _GEN_796 == 7'h4a; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_7429 = _T_7427 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_7431 = _T_7429 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_7432 = _T_7426 | _T_7431; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_7442 = _T_4785 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_7443 = _GEN_796 == 7'h4b; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_7445 = _T_7443 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_7447 = _T_7445 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_7448 = _T_7442 | _T_7447; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_7458 = _T_4789 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_7459 = _GEN_796 == 7'h4c; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_7461 = _T_7459 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_7463 = _T_7461 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_7464 = _T_7458 | _T_7463; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_7474 = _T_4793 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_7475 = _GEN_796 == 7'h4d; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_7477 = _T_7475 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_7479 = _T_7477 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_7480 = _T_7474 | _T_7479; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_7490 = _T_4797 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_7491 = _GEN_796 == 7'h4e; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_7493 = _T_7491 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_7495 = _T_7493 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_7496 = _T_7490 | _T_7495; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_7506 = _T_4801 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_7507 = _GEN_796 == 7'h4f; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_7509 = _T_7507 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_7511 = _T_7509 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_7512 = _T_7506 | _T_7511; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_7522 = _T_4805 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_7523 = _GEN_796 == 7'h50; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_7525 = _T_7523 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_7527 = _T_7525 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_7528 = _T_7522 | _T_7527; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_7538 = _T_4809 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_7539 = _GEN_796 == 7'h51; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_7541 = _T_7539 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_7543 = _T_7541 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_7544 = _T_7538 | _T_7543; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_7554 = _T_4813 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_7555 = _GEN_796 == 7'h52; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_7557 = _T_7555 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_7559 = _T_7557 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_7560 = _T_7554 | _T_7559; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_7570 = _T_4817 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_7571 = _GEN_796 == 7'h53; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_7573 = _T_7571 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_7575 = _T_7573 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_7576 = _T_7570 | _T_7575; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_7586 = _T_4821 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_7587 = _GEN_796 == 7'h54; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_7589 = _T_7587 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_7591 = _T_7589 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_7592 = _T_7586 | _T_7591; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_7602 = _T_4825 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_7603 = _GEN_796 == 7'h55; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_7605 = _T_7603 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_7607 = _T_7605 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_7608 = _T_7602 | _T_7607; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_7618 = _T_4829 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_7619 = _GEN_796 == 7'h56; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_7621 = _T_7619 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_7623 = _T_7621 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_7624 = _T_7618 | _T_7623; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_7634 = _T_4833 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_7635 = _GEN_796 == 7'h57; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_7637 = _T_7635 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_7639 = _T_7637 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_7640 = _T_7634 | _T_7639; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_7650 = _T_4837 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_7651 = _GEN_796 == 7'h58; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_7653 = _T_7651 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_7655 = _T_7653 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_7656 = _T_7650 | _T_7655; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_7666 = _T_4841 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_7667 = _GEN_796 == 7'h59; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_7669 = _T_7667 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_7671 = _T_7669 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_7672 = _T_7666 | _T_7671; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_7682 = _T_4845 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_7683 = _GEN_796 == 7'h5a; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_7685 = _T_7683 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_7687 = _T_7685 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_7688 = _T_7682 | _T_7687; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_7698 = _T_4849 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_7699 = _GEN_796 == 7'h5b; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_7701 = _T_7699 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_7703 = _T_7701 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_7704 = _T_7698 | _T_7703; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_7714 = _T_4853 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_7715 = _GEN_796 == 7'h5c; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_7717 = _T_7715 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_7719 = _T_7717 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_7720 = _T_7714 | _T_7719; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_7730 = _T_4857 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_7731 = _GEN_796 == 7'h5d; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_7733 = _T_7731 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_7735 = _T_7733 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_7736 = _T_7730 | _T_7735; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_7746 = _T_4861 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_7747 = _GEN_796 == 7'h5e; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_7749 = _T_7747 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_7751 = _T_7749 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_7752 = _T_7746 | _T_7751; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_7762 = _T_4865 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_7763 = _GEN_796 == 7'h5f; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_7765 = _T_7763 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_7767 = _T_7765 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_7768 = _T_7762 | _T_7767; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_7778 = _T_4741 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_7781 = _T_7267 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_7783 = _T_7781 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_7784 = _T_7778 | _T_7783; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_7794 = _T_4745 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_7797 = _T_7283 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_7799 = _T_7797 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_7800 = _T_7794 | _T_7799; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_7810 = _T_4749 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_7813 = _T_7299 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_7815 = _T_7813 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_7816 = _T_7810 | _T_7815; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_7826 = _T_4753 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_7829 = _T_7315 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_7831 = _T_7829 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_7832 = _T_7826 | _T_7831; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_7842 = _T_4757 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_7845 = _T_7331 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_7847 = _T_7845 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_7848 = _T_7842 | _T_7847; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_7858 = _T_4761 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_7861 = _T_7347 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_7863 = _T_7861 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_7864 = _T_7858 | _T_7863; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_7874 = _T_4765 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_7877 = _T_7363 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_7879 = _T_7877 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_7880 = _T_7874 | _T_7879; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_7890 = _T_4769 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_7893 = _T_7379 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_7895 = _T_7893 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_7896 = _T_7890 | _T_7895; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_7906 = _T_4773 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_7909 = _T_7395 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_7911 = _T_7909 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_7912 = _T_7906 | _T_7911; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_7922 = _T_4777 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_7925 = _T_7411 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_7927 = _T_7925 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_7928 = _T_7922 | _T_7927; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_7938 = _T_4781 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_7941 = _T_7427 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_7943 = _T_7941 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_7944 = _T_7938 | _T_7943; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_7954 = _T_4785 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_7957 = _T_7443 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_7959 = _T_7957 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_7960 = _T_7954 | _T_7959; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_7970 = _T_4789 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_7973 = _T_7459 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_7975 = _T_7973 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_7976 = _T_7970 | _T_7975; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_7986 = _T_4793 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_7989 = _T_7475 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_7991 = _T_7989 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_7992 = _T_7986 | _T_7991; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_8002 = _T_4797 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_8005 = _T_7491 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_8007 = _T_8005 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_8008 = _T_8002 | _T_8007; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_8018 = _T_4801 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_8021 = _T_7507 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_8023 = _T_8021 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_8024 = _T_8018 | _T_8023; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_8034 = _T_4805 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_8037 = _T_7523 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_8039 = _T_8037 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_8040 = _T_8034 | _T_8039; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_8050 = _T_4809 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_8053 = _T_7539 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_8055 = _T_8053 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_8056 = _T_8050 | _T_8055; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_8066 = _T_4813 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_8069 = _T_7555 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_8071 = _T_8069 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_8072 = _T_8066 | _T_8071; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_8082 = _T_4817 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_8085 = _T_7571 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_8087 = _T_8085 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_8088 = _T_8082 | _T_8087; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_8098 = _T_4821 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_8101 = _T_7587 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_8103 = _T_8101 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_8104 = _T_8098 | _T_8103; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_8114 = _T_4825 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_8117 = _T_7603 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_8119 = _T_8117 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_8120 = _T_8114 | _T_8119; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_8130 = _T_4829 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_8133 = _T_7619 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_8135 = _T_8133 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_8136 = _T_8130 | _T_8135; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_8146 = _T_4833 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_8149 = _T_7635 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_8151 = _T_8149 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_8152 = _T_8146 | _T_8151; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_8162 = _T_4837 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_8165 = _T_7651 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_8167 = _T_8165 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_8168 = _T_8162 | _T_8167; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_8178 = _T_4841 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_8181 = _T_7667 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_8183 = _T_8181 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_8184 = _T_8178 | _T_8183; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_8194 = _T_4845 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_8197 = _T_7683 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_8199 = _T_8197 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_8200 = _T_8194 | _T_8199; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_8210 = _T_4849 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_8213 = _T_7699 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_8215 = _T_8213 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_8216 = _T_8210 | _T_8215; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_8226 = _T_4853 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_8229 = _T_7715 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_8231 = _T_8229 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_8232 = _T_8226 | _T_8231; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_8242 = _T_4857 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_8245 = _T_7731 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_8247 = _T_8245 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_8248 = _T_8242 | _T_8247; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_8258 = _T_4861 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_8261 = _T_7747 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_8263 = _T_8261 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_8264 = _T_8258 | _T_8263; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_8274 = _T_4865 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_8277 = _T_7763 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_8279 = _T_8277 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_8280 = _T_8274 | _T_8279; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_8290 = _T_4869 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_8291 = _GEN_796 == 7'h60; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_8293 = _T_8291 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_8295 = _T_8293 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_8296 = _T_8290 | _T_8295; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_8306 = _T_4873 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_8307 = _GEN_796 == 7'h61; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_8309 = _T_8307 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_8311 = _T_8309 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_8312 = _T_8306 | _T_8311; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_8322 = _T_4877 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_8323 = _GEN_796 == 7'h62; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_8325 = _T_8323 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_8327 = _T_8325 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_8328 = _T_8322 | _T_8327; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_8338 = _T_4881 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_8339 = _GEN_796 == 7'h63; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_8341 = _T_8339 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_8343 = _T_8341 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_8344 = _T_8338 | _T_8343; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_8354 = _T_4885 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_8355 = _GEN_796 == 7'h64; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_8357 = _T_8355 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_8359 = _T_8357 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_8360 = _T_8354 | _T_8359; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_8370 = _T_4889 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_8371 = _GEN_796 == 7'h65; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_8373 = _T_8371 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_8375 = _T_8373 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_8376 = _T_8370 | _T_8375; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_8386 = _T_4893 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_8387 = _GEN_796 == 7'h66; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_8389 = _T_8387 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_8391 = _T_8389 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_8392 = _T_8386 | _T_8391; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_8402 = _T_4897 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_8403 = _GEN_796 == 7'h67; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_8405 = _T_8403 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_8407 = _T_8405 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_8408 = _T_8402 | _T_8407; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_8418 = _T_4901 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_8419 = _GEN_796 == 7'h68; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_8421 = _T_8419 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_8423 = _T_8421 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_8424 = _T_8418 | _T_8423; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_8434 = _T_4905 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_8435 = _GEN_796 == 7'h69; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_8437 = _T_8435 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_8439 = _T_8437 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_8440 = _T_8434 | _T_8439; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_8450 = _T_4909 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_8451 = _GEN_796 == 7'h6a; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_8453 = _T_8451 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_8455 = _T_8453 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_8456 = _T_8450 | _T_8455; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_8466 = _T_4913 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_8467 = _GEN_796 == 7'h6b; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_8469 = _T_8467 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_8471 = _T_8469 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_8472 = _T_8466 | _T_8471; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_8482 = _T_4917 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_8483 = _GEN_796 == 7'h6c; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_8485 = _T_8483 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_8487 = _T_8485 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_8488 = _T_8482 | _T_8487; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_8498 = _T_4921 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_8499 = _GEN_796 == 7'h6d; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_8501 = _T_8499 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_8503 = _T_8501 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_8504 = _T_8498 | _T_8503; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_8514 = _T_4925 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_8515 = _GEN_796 == 7'h6e; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_8517 = _T_8515 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_8519 = _T_8517 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_8520 = _T_8514 | _T_8519; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_8530 = _T_4929 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_8531 = _GEN_796 == 7'h6f; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_8533 = _T_8531 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_8535 = _T_8533 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_8536 = _T_8530 | _T_8535; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_8546 = _T_4933 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_8547 = _GEN_796 == 7'h70; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_8549 = _T_8547 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_8551 = _T_8549 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_8552 = _T_8546 | _T_8551; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_8562 = _T_4937 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_8563 = _GEN_796 == 7'h71; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_8565 = _T_8563 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_8567 = _T_8565 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_8568 = _T_8562 | _T_8567; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_8578 = _T_4941 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_8579 = _GEN_796 == 7'h72; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_8581 = _T_8579 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_8583 = _T_8581 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_8584 = _T_8578 | _T_8583; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_8594 = _T_4945 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_8595 = _GEN_796 == 7'h73; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_8597 = _T_8595 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_8599 = _T_8597 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_8600 = _T_8594 | _T_8599; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_8610 = _T_4949 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_8611 = _GEN_796 == 7'h74; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_8613 = _T_8611 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_8615 = _T_8613 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_8616 = _T_8610 | _T_8615; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_8626 = _T_4953 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_8627 = _GEN_796 == 7'h75; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_8629 = _T_8627 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_8631 = _T_8629 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_8632 = _T_8626 | _T_8631; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_8642 = _T_4957 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_8643 = _GEN_796 == 7'h76; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_8645 = _T_8643 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_8647 = _T_8645 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_8648 = _T_8642 | _T_8647; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_8658 = _T_4961 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_8659 = _GEN_796 == 7'h77; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_8661 = _T_8659 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_8663 = _T_8661 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_8664 = _T_8658 | _T_8663; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_8674 = _T_4965 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_8675 = _GEN_796 == 7'h78; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_8677 = _T_8675 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_8679 = _T_8677 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_8680 = _T_8674 | _T_8679; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_8690 = _T_4969 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_8691 = _GEN_796 == 7'h79; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_8693 = _T_8691 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_8695 = _T_8693 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_8696 = _T_8690 | _T_8695; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_8706 = _T_4973 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_8707 = _GEN_796 == 7'h7a; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_8709 = _T_8707 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_8711 = _T_8709 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_8712 = _T_8706 | _T_8711; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_8722 = _T_4977 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_8723 = _GEN_796 == 7'h7b; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_8725 = _T_8723 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_8727 = _T_8725 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_8728 = _T_8722 | _T_8727; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_8738 = _T_4981 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_8739 = _GEN_796 == 7'h7c; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_8741 = _T_8739 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_8743 = _T_8741 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_8744 = _T_8738 | _T_8743; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_8754 = _T_4985 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_8755 = _GEN_796 == 7'h7d; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_8757 = _T_8755 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_8759 = _T_8757 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_8760 = _T_8754 | _T_8759; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_8770 = _T_4989 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_8771 = _GEN_796 == 7'h7e; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_8773 = _T_8771 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_8775 = _T_8773 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_8776 = _T_8770 | _T_8775; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_8786 = _T_4993 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_8787 = _GEN_796 == 7'h7f; // @[el2_ifu_mem_ctl.scala 751:101]
  wire  _T_8789 = _T_8787 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_8791 = _T_8789 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_8792 = _T_8786 | _T_8791; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_8802 = _T_4869 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_8805 = _T_8291 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_8807 = _T_8805 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_8808 = _T_8802 | _T_8807; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_8818 = _T_4873 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_8821 = _T_8307 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_8823 = _T_8821 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_8824 = _T_8818 | _T_8823; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_8834 = _T_4877 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_8837 = _T_8323 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_8839 = _T_8837 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_8840 = _T_8834 | _T_8839; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_8850 = _T_4881 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_8853 = _T_8339 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_8855 = _T_8853 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_8856 = _T_8850 | _T_8855; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_8866 = _T_4885 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_8869 = _T_8355 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_8871 = _T_8869 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_8872 = _T_8866 | _T_8871; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_8882 = _T_4889 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_8885 = _T_8371 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_8887 = _T_8885 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_8888 = _T_8882 | _T_8887; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_8898 = _T_4893 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_8901 = _T_8387 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_8903 = _T_8901 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_8904 = _T_8898 | _T_8903; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_8914 = _T_4897 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_8917 = _T_8403 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_8919 = _T_8917 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_8920 = _T_8914 | _T_8919; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_8930 = _T_4901 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_8933 = _T_8419 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_8935 = _T_8933 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_8936 = _T_8930 | _T_8935; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_8946 = _T_4905 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_8949 = _T_8435 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_8951 = _T_8949 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_8952 = _T_8946 | _T_8951; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_8962 = _T_4909 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_8965 = _T_8451 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_8967 = _T_8965 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_8968 = _T_8962 | _T_8967; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_8978 = _T_4913 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_8981 = _T_8467 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_8983 = _T_8981 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_8984 = _T_8978 | _T_8983; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_8994 = _T_4917 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_8997 = _T_8483 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_8999 = _T_8997 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_9000 = _T_8994 | _T_8999; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_9010 = _T_4921 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_9013 = _T_8499 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_9015 = _T_9013 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_9016 = _T_9010 | _T_9015; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_9026 = _T_4925 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_9029 = _T_8515 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_9031 = _T_9029 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_9032 = _T_9026 | _T_9031; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_9042 = _T_4929 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_9045 = _T_8531 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_9047 = _T_9045 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_9048 = _T_9042 | _T_9047; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_9058 = _T_4933 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_9061 = _T_8547 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_9063 = _T_9061 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_9064 = _T_9058 | _T_9063; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_9074 = _T_4937 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_9077 = _T_8563 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_9079 = _T_9077 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_9080 = _T_9074 | _T_9079; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_9090 = _T_4941 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_9093 = _T_8579 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_9095 = _T_9093 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_9096 = _T_9090 | _T_9095; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_9106 = _T_4945 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_9109 = _T_8595 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_9111 = _T_9109 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_9112 = _T_9106 | _T_9111; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_9122 = _T_4949 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_9125 = _T_8611 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_9127 = _T_9125 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_9128 = _T_9122 | _T_9127; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_9138 = _T_4953 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_9141 = _T_8627 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_9143 = _T_9141 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_9144 = _T_9138 | _T_9143; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_9154 = _T_4957 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_9157 = _T_8643 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_9159 = _T_9157 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_9160 = _T_9154 | _T_9159; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_9170 = _T_4961 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_9173 = _T_8659 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_9175 = _T_9173 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_9176 = _T_9170 | _T_9175; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_9186 = _T_4965 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_9189 = _T_8675 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_9191 = _T_9189 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_9192 = _T_9186 | _T_9191; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_9202 = _T_4969 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_9205 = _T_8691 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_9207 = _T_9205 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_9208 = _T_9202 | _T_9207; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_9218 = _T_4973 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_9221 = _T_8707 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_9223 = _T_9221 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_9224 = _T_9218 | _T_9223; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_9234 = _T_4977 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_9237 = _T_8723 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_9239 = _T_9237 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_9240 = _T_9234 | _T_9239; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_9250 = _T_4981 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_9253 = _T_8739 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_9255 = _T_9253 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_9256 = _T_9250 | _T_9255; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_9266 = _T_4985 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_9269 = _T_8755 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_9271 = _T_9269 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_9272 = _T_9266 | _T_9271; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_9282 = _T_4989 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_9285 = _T_8771 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_9287 = _T_9285 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_9288 = _T_9282 | _T_9287; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_9298 = _T_4993 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:58]
  wire  _T_9301 = _T_8787 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:123]
  wire  _T_9303 = _T_9301 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 751:144]
  wire  _T_9304 = _T_9298 | _T_9303; // @[el2_ifu_mem_ctl.scala 751:80]
  wire  _T_10105 = ~fetch_uncacheable_ff; // @[el2_ifu_mem_ctl.scala 805:63]
  wire  _T_10106 = _T_10105 & ifc_fetch_req_f; // @[el2_ifu_mem_ctl.scala 805:85]
  wire [1:0] _T_10108 = _T_10106 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  reg  _T_10115; // @[el2_ifu_mem_ctl.scala 810:57]
  reg  _T_10116; // @[el2_ifu_mem_ctl.scala 811:56]
  reg  _T_10117; // @[el2_ifu_mem_ctl.scala 812:59]
  wire  _T_10118 = ~ifu_bus_arready_ff; // @[el2_ifu_mem_ctl.scala 813:80]
  wire  _T_10119 = ifu_bus_arvalid_ff & _T_10118; // @[el2_ifu_mem_ctl.scala 813:78]
  wire  _T_10120 = _T_10119 & miss_pending; // @[el2_ifu_mem_ctl.scala 813:100]
  reg  _T_10121; // @[el2_ifu_mem_ctl.scala 813:58]
  reg  _T_10122; // @[el2_ifu_mem_ctl.scala 814:58]
  wire  _T_10125 = io_dec_tlu_ic_diag_pkt_icache_dicawics[15:14] == 2'h3; // @[el2_ifu_mem_ctl.scala 821:71]
  wire  _T_10127 = io_dec_tlu_ic_diag_pkt_icache_dicawics[15:14] == 2'h2; // @[el2_ifu_mem_ctl.scala 821:124]
  wire  _T_10129 = io_dec_tlu_ic_diag_pkt_icache_dicawics[15:14] == 2'h1; // @[el2_ifu_mem_ctl.scala 822:50]
  wire  _T_10131 = io_dec_tlu_ic_diag_pkt_icache_dicawics[15:14] == 2'h0; // @[el2_ifu_mem_ctl.scala 822:103]
  wire [3:0] _T_10134 = {_T_10125,_T_10127,_T_10129,_T_10131}; // @[Cat.scala 29:58]
  wire  ic_debug_ict_array_sel_in = io_ic_debug_rd_en & io_ic_debug_tag_array; // @[el2_ifu_mem_ctl.scala 824:53]
  reg  _T_10145; // @[Reg.scala 27:20]
  assign io_ifu_miss_state_idle = miss_state == 3'h0; // @[el2_ifu_mem_ctl.scala 329:26]
  assign io_ifu_ic_mb_empty = _T_326 | _T_231; // @[el2_ifu_mem_ctl.scala 328:22]
  assign io_ic_dma_active = _T_11 | io_dec_tlu_flush_err_wb; // @[el2_ifu_mem_ctl.scala 192:20]
  assign io_ic_write_stall = write_ic_16_bytes & _T_3940; // @[el2_ifu_mem_ctl.scala 701:21]
  assign io_ifu_pmu_ic_miss = _T_10115; // @[el2_ifu_mem_ctl.scala 810:22]
  assign io_ifu_pmu_ic_hit = _T_10116; // @[el2_ifu_mem_ctl.scala 811:21]
  assign io_ifu_pmu_bus_error = _T_10117; // @[el2_ifu_mem_ctl.scala 812:24]
  assign io_ifu_pmu_bus_busy = _T_10121; // @[el2_ifu_mem_ctl.scala 813:23]
  assign io_ifu_pmu_bus_trxn = _T_10122; // @[el2_ifu_mem_ctl.scala 814:23]
  assign io_ifu_axi_awvalid = 1'h0; // @[el2_ifu_mem_ctl.scala 143:22]
  assign io_ifu_axi_awid = 3'h0; // @[el2_ifu_mem_ctl.scala 142:19]
  assign io_ifu_axi_awaddr = 32'h0; // @[el2_ifu_mem_ctl.scala 137:21]
  assign io_ifu_axi_awregion = 4'h0; // @[el2_ifu_mem_ctl.scala 141:23]
  assign io_ifu_axi_awlen = 8'h0; // @[el2_ifu_mem_ctl.scala 139:20]
  assign io_ifu_axi_awsize = 3'h0; // @[el2_ifu_mem_ctl.scala 150:21]
  assign io_ifu_axi_awburst = 2'h0; // @[el2_ifu_mem_ctl.scala 152:22]
  assign io_ifu_axi_awlock = 1'h0; // @[el2_ifu_mem_ctl.scala 147:21]
  assign io_ifu_axi_awcache = 4'h0; // @[el2_ifu_mem_ctl.scala 145:22]
  assign io_ifu_axi_awprot = 3'h0; // @[el2_ifu_mem_ctl.scala 138:21]
  assign io_ifu_axi_awqos = 4'h0; // @[el2_ifu_mem_ctl.scala 136:20]
  assign io_ifu_axi_wvalid = 1'h0; // @[el2_ifu_mem_ctl.scala 134:21]
  assign io_ifu_axi_wdata = 64'h0; // @[el2_ifu_mem_ctl.scala 135:20]
  assign io_ifu_axi_wstrb = 8'h0; // @[el2_ifu_mem_ctl.scala 144:20]
  assign io_ifu_axi_wlast = 1'h0; // @[el2_ifu_mem_ctl.scala 153:20]
  assign io_ifu_axi_bready = 1'h0; // @[el2_ifu_mem_ctl.scala 148:21]
  assign io_ifu_axi_arvalid = ifu_bus_cmd_valid; // @[el2_ifu_mem_ctl.scala 563:22]
  assign io_ifu_axi_arid = bus_rd_addr_count & _T_2534; // @[el2_ifu_mem_ctl.scala 564:19]
  assign io_ifu_axi_araddr = _T_2536 & _T_2538; // @[el2_ifu_mem_ctl.scala 565:21]
  assign io_ifu_axi_arregion = ifu_ic_req_addr_f[28:25]; // @[el2_ifu_mem_ctl.scala 568:23]
  assign io_ifu_axi_arlen = 8'h0; // @[el2_ifu_mem_ctl.scala 149:20]
  assign io_ifu_axi_arsize = 3'h3; // @[el2_ifu_mem_ctl.scala 566:21]
  assign io_ifu_axi_arburst = 2'h1; // @[el2_ifu_mem_ctl.scala 569:22]
  assign io_ifu_axi_arlock = 1'h0; // @[el2_ifu_mem_ctl.scala 140:21]
  assign io_ifu_axi_arcache = 4'hf; // @[el2_ifu_mem_ctl.scala 567:22]
  assign io_ifu_axi_arprot = 3'h0; // @[el2_ifu_mem_ctl.scala 151:21]
  assign io_ifu_axi_arqos = 4'h0; // @[el2_ifu_mem_ctl.scala 146:20]
  assign io_ifu_axi_rready = 1'h1; // @[el2_ifu_mem_ctl.scala 570:21]
  assign io_iccm_dma_ecc_error = |iccm_double_ecc_error; // @[el2_ifu_mem_ctl.scala 660:25]
  assign io_iccm_dma_rvalid = iccm_dma_rvalid; // @[el2_ifu_mem_ctl.scala 658:22]
  assign io_iccm_dma_rdata = iccm_dma_rdata; // @[el2_ifu_mem_ctl.scala 662:21]
  assign io_iccm_dma_rtag = iccm_dma_rtag; // @[el2_ifu_mem_ctl.scala 653:20]
  assign io_iccm_ready = _T_2637 & _T_2631; // @[el2_ifu_mem_ctl.scala 633:17]
  assign io_ic_rw_addr = _T_338 | _T_339; // @[el2_ifu_mem_ctl.scala 338:17]
  assign io_ic_wr_en = 2'h0; // @[el2_ifu_mem_ctl.scala 700:15]
  assign io_ic_rd_en = _T_3918 | _T_3923; // @[el2_ifu_mem_ctl.scala 691:15]
  assign io_ic_wr_data_0 = ic_wr_16bytes_data[70:0]; // @[el2_ifu_mem_ctl.scala 347:17]
  assign io_ic_wr_data_1 = ic_wr_16bytes_data[141:71]; // @[el2_ifu_mem_ctl.scala 347:17]
  assign io_ic_debug_wr_data = io_dec_tlu_ic_diag_pkt_icache_wrdata; // @[el2_ifu_mem_ctl.scala 348:23]
  assign io_ifu_ic_debug_rd_data = _T_1209; // @[el2_ifu_mem_ctl.scala 356:27]
  assign io_ic_debug_addr = io_dec_tlu_ic_diag_pkt_icache_dicawics[9:0]; // @[el2_ifu_mem_ctl.scala 817:20]
  assign io_ic_debug_rd_en = io_dec_tlu_ic_diag_pkt_icache_rd_valid; // @[el2_ifu_mem_ctl.scala 819:21]
  assign io_ic_debug_wr_en = io_dec_tlu_ic_diag_pkt_icache_wr_valid; // @[el2_ifu_mem_ctl.scala 820:21]
  assign io_ic_debug_tag_array = io_dec_tlu_ic_diag_pkt_icache_dicawics[16]; // @[el2_ifu_mem_ctl.scala 818:25]
  assign io_ic_debug_way = _T_10134[1:0]; // @[el2_ifu_mem_ctl.scala 821:19]
  assign io_ic_tag_valid = ic_tag_valid_unq & _T_10108; // @[el2_ifu_mem_ctl.scala 805:19]
  assign io_iccm_rw_addr = _T_3072[14:0]; // @[el2_ifu_mem_ctl.scala 664:19]
  assign io_iccm_wren = _T_2641 | iccm_correct_ecc; // @[el2_ifu_mem_ctl.scala 635:16]
  assign io_iccm_rden = _T_2645 | _T_2646; // @[el2_ifu_mem_ctl.scala 636:16]
  assign io_iccm_wr_data = _T_3047 ? _T_3048 : _T_3055; // @[el2_ifu_mem_ctl.scala 641:19]
  assign io_iccm_wr_size = _T_2651 & io_dma_mem_sz; // @[el2_ifu_mem_ctl.scala 638:19]
  assign io_ic_hit_f = _T_263 | _T_264; // @[el2_ifu_mem_ctl.scala 290:15]
  assign io_ic_access_fault_f = _T_2419 & _T_317; // @[el2_ifu_mem_ctl.scala 389:24]
  assign io_ic_access_fault_type_f = io_iccm_rd_ecc_double_err ? 2'h1 : _T_1273; // @[el2_ifu_mem_ctl.scala 390:29]
  assign io_iccm_rd_ecc_single_err = _T_3863 & ifc_fetch_req_f; // @[el2_ifu_mem_ctl.scala 677:29]
  assign io_iccm_rd_ecc_double_err = iccm_dma_ecc_error_in & ifc_iccm_access_f; // @[el2_ifu_mem_ctl.scala 678:29]
  assign io_ic_error_start = _T_1197 | ic_rd_parity_final_err; // @[el2_ifu_mem_ctl.scala 350:21]
  assign io_ifu_async_error_start = io_iccm_rd_ecc_single_err | io_ic_error_start; // @[el2_ifu_mem_ctl.scala 191:28]
  assign io_iccm_dma_sb_error = _T_3 & dma_iccm_req_f; // @[el2_ifu_mem_ctl.scala 190:24]
  assign io_ic_fetch_val_f = {1'h0,fetch_req_f_qual}; // @[el2_ifu_mem_ctl.scala 394:21]
  assign io_ic_data_f = io_ic_rd_data[31:0]; // @[el2_ifu_mem_ctl.scala 386:16]
  assign io_ic_premux_data = ic_premux_data[63:0]; // @[el2_ifu_mem_ctl.scala 383:21]
  assign io_ic_sel_premux_data = fetch_req_iccm_f | sel_byp_data; // @[el2_ifu_mem_ctl.scala 384:25]
  assign io_ifu_ic_debug_rd_data_valid = _T_10145; // @[el2_ifu_mem_ctl.scala 828:33]
  assign io_iccm_buf_correct_ecc = iccm_correct_ecc & _T_2424; // @[el2_ifu_mem_ctl.scala 482:27]
  assign io_iccm_correction_state = _T_2452 ? 1'h0 : _GEN_59; // @[el2_ifu_mem_ctl.scala 517:28 el2_ifu_mem_ctl.scala 530:32 el2_ifu_mem_ctl.scala 537:32 el2_ifu_mem_ctl.scala 544:32]
  assign io_ic_miss_buff_ecc = {_T_1193,_T_1190}; // @[el2_ifu_mem_ctl.scala 345:23]
  assign io_ic_wr_ecc = {_T_771,_T_768}; // @[el2_ifu_mem_ctl.scala 343:16]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  flush_final_f = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  ifc_fetch_req_f_raw = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  miss_state = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  scnd_miss_req_q = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  ifu_fetch_addr_int_f = _RAND_4[30:0];
  _RAND_5 = {1{`RANDOM}};
  ifc_iccm_access_f = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  iccm_dma_rvalid_in = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  dma_iccm_req_f = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  perr_state = _RAND_8[2:0];
  _RAND_9 = {1{`RANDOM}};
  err_stop_state = _RAND_9[1:0];
  _RAND_10 = {1{`RANDOM}};
  reset_all_tags = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  ifc_region_acc_fault_final_f = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  ifu_bus_rvalid_unq_ff = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  bus_ifu_bus_clk_en_ff = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  uncacheable_miss_ff = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  bus_data_beat_count = _RAND_15[2:0];
  _RAND_16 = {1{`RANDOM}};
  ic_miss_buff_data_valid = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  imb_ff = _RAND_17[30:0];
  _RAND_18 = {1{`RANDOM}};
  last_data_recieved_ff = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  sel_mb_addr_ff = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  way_status_mb_scnd_ff = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  _T_5128 = _RAND_21[6:0];
  _RAND_22 = {1{`RANDOM}};
  _T_4484 = _RAND_22[2:0];
  _RAND_23 = {1{`RANDOM}};
  _T_4480 = _RAND_23[2:0];
  _RAND_24 = {1{`RANDOM}};
  _T_4476 = _RAND_24[2:0];
  _RAND_25 = {1{`RANDOM}};
  _T_4472 = _RAND_25[2:0];
  _RAND_26 = {1{`RANDOM}};
  _T_4468 = _RAND_26[2:0];
  _RAND_27 = {1{`RANDOM}};
  _T_4464 = _RAND_27[2:0];
  _RAND_28 = {1{`RANDOM}};
  _T_4460 = _RAND_28[2:0];
  _RAND_29 = {1{`RANDOM}};
  _T_4456 = _RAND_29[2:0];
  _RAND_30 = {1{`RANDOM}};
  _T_4452 = _RAND_30[2:0];
  _RAND_31 = {1{`RANDOM}};
  _T_4448 = _RAND_31[2:0];
  _RAND_32 = {1{`RANDOM}};
  _T_4444 = _RAND_32[2:0];
  _RAND_33 = {1{`RANDOM}};
  _T_4440 = _RAND_33[2:0];
  _RAND_34 = {1{`RANDOM}};
  _T_4436 = _RAND_34[2:0];
  _RAND_35 = {1{`RANDOM}};
  _T_4432 = _RAND_35[2:0];
  _RAND_36 = {1{`RANDOM}};
  _T_4428 = _RAND_36[2:0];
  _RAND_37 = {1{`RANDOM}};
  _T_4424 = _RAND_37[2:0];
  _RAND_38 = {1{`RANDOM}};
  _T_4420 = _RAND_38[2:0];
  _RAND_39 = {1{`RANDOM}};
  _T_4416 = _RAND_39[2:0];
  _RAND_40 = {1{`RANDOM}};
  _T_4412 = _RAND_40[2:0];
  _RAND_41 = {1{`RANDOM}};
  _T_4408 = _RAND_41[2:0];
  _RAND_42 = {1{`RANDOM}};
  _T_4404 = _RAND_42[2:0];
  _RAND_43 = {1{`RANDOM}};
  _T_4400 = _RAND_43[2:0];
  _RAND_44 = {1{`RANDOM}};
  _T_4396 = _RAND_44[2:0];
  _RAND_45 = {1{`RANDOM}};
  _T_4392 = _RAND_45[2:0];
  _RAND_46 = {1{`RANDOM}};
  _T_4388 = _RAND_46[2:0];
  _RAND_47 = {1{`RANDOM}};
  _T_4384 = _RAND_47[2:0];
  _RAND_48 = {1{`RANDOM}};
  _T_4380 = _RAND_48[2:0];
  _RAND_49 = {1{`RANDOM}};
  _T_4376 = _RAND_49[2:0];
  _RAND_50 = {1{`RANDOM}};
  _T_4372 = _RAND_50[2:0];
  _RAND_51 = {1{`RANDOM}};
  _T_4368 = _RAND_51[2:0];
  _RAND_52 = {1{`RANDOM}};
  _T_4364 = _RAND_52[2:0];
  _RAND_53 = {1{`RANDOM}};
  _T_4360 = _RAND_53[2:0];
  _RAND_54 = {1{`RANDOM}};
  _T_4356 = _RAND_54[2:0];
  _RAND_55 = {1{`RANDOM}};
  _T_4352 = _RAND_55[2:0];
  _RAND_56 = {1{`RANDOM}};
  _T_4348 = _RAND_56[2:0];
  _RAND_57 = {1{`RANDOM}};
  _T_4344 = _RAND_57[2:0];
  _RAND_58 = {1{`RANDOM}};
  _T_4340 = _RAND_58[2:0];
  _RAND_59 = {1{`RANDOM}};
  _T_4336 = _RAND_59[2:0];
  _RAND_60 = {1{`RANDOM}};
  _T_4332 = _RAND_60[2:0];
  _RAND_61 = {1{`RANDOM}};
  _T_4328 = _RAND_61[2:0];
  _RAND_62 = {1{`RANDOM}};
  _T_4324 = _RAND_62[2:0];
  _RAND_63 = {1{`RANDOM}};
  _T_4320 = _RAND_63[2:0];
  _RAND_64 = {1{`RANDOM}};
  _T_4316 = _RAND_64[2:0];
  _RAND_65 = {1{`RANDOM}};
  _T_4312 = _RAND_65[2:0];
  _RAND_66 = {1{`RANDOM}};
  _T_4308 = _RAND_66[2:0];
  _RAND_67 = {1{`RANDOM}};
  _T_4304 = _RAND_67[2:0];
  _RAND_68 = {1{`RANDOM}};
  _T_4300 = _RAND_68[2:0];
  _RAND_69 = {1{`RANDOM}};
  _T_4296 = _RAND_69[2:0];
  _RAND_70 = {1{`RANDOM}};
  _T_4292 = _RAND_70[2:0];
  _RAND_71 = {1{`RANDOM}};
  _T_4288 = _RAND_71[2:0];
  _RAND_72 = {1{`RANDOM}};
  _T_4284 = _RAND_72[2:0];
  _RAND_73 = {1{`RANDOM}};
  _T_4280 = _RAND_73[2:0];
  _RAND_74 = {1{`RANDOM}};
  _T_4276 = _RAND_74[2:0];
  _RAND_75 = {1{`RANDOM}};
  _T_4272 = _RAND_75[2:0];
  _RAND_76 = {1{`RANDOM}};
  _T_4268 = _RAND_76[2:0];
  _RAND_77 = {1{`RANDOM}};
  _T_4264 = _RAND_77[2:0];
  _RAND_78 = {1{`RANDOM}};
  _T_4260 = _RAND_78[2:0];
  _RAND_79 = {1{`RANDOM}};
  _T_4256 = _RAND_79[2:0];
  _RAND_80 = {1{`RANDOM}};
  _T_4252 = _RAND_80[2:0];
  _RAND_81 = {1{`RANDOM}};
  _T_4248 = _RAND_81[2:0];
  _RAND_82 = {1{`RANDOM}};
  _T_4244 = _RAND_82[2:0];
  _RAND_83 = {1{`RANDOM}};
  _T_4240 = _RAND_83[2:0];
  _RAND_84 = {1{`RANDOM}};
  _T_4236 = _RAND_84[2:0];
  _RAND_85 = {1{`RANDOM}};
  _T_4232 = _RAND_85[2:0];
  _RAND_86 = {1{`RANDOM}};
  _T_4228 = _RAND_86[2:0];
  _RAND_87 = {1{`RANDOM}};
  _T_4224 = _RAND_87[2:0];
  _RAND_88 = {1{`RANDOM}};
  _T_4220 = _RAND_88[2:0];
  _RAND_89 = {1{`RANDOM}};
  _T_4216 = _RAND_89[2:0];
  _RAND_90 = {1{`RANDOM}};
  _T_4212 = _RAND_90[2:0];
  _RAND_91 = {1{`RANDOM}};
  _T_4208 = _RAND_91[2:0];
  _RAND_92 = {1{`RANDOM}};
  _T_4204 = _RAND_92[2:0];
  _RAND_93 = {1{`RANDOM}};
  _T_4200 = _RAND_93[2:0];
  _RAND_94 = {1{`RANDOM}};
  _T_4196 = _RAND_94[2:0];
  _RAND_95 = {1{`RANDOM}};
  _T_4192 = _RAND_95[2:0];
  _RAND_96 = {1{`RANDOM}};
  _T_4188 = _RAND_96[2:0];
  _RAND_97 = {1{`RANDOM}};
  _T_4184 = _RAND_97[2:0];
  _RAND_98 = {1{`RANDOM}};
  _T_4180 = _RAND_98[2:0];
  _RAND_99 = {1{`RANDOM}};
  _T_4176 = _RAND_99[2:0];
  _RAND_100 = {1{`RANDOM}};
  _T_4172 = _RAND_100[2:0];
  _RAND_101 = {1{`RANDOM}};
  _T_4168 = _RAND_101[2:0];
  _RAND_102 = {1{`RANDOM}};
  _T_4164 = _RAND_102[2:0];
  _RAND_103 = {1{`RANDOM}};
  _T_4160 = _RAND_103[2:0];
  _RAND_104 = {1{`RANDOM}};
  _T_4156 = _RAND_104[2:0];
  _RAND_105 = {1{`RANDOM}};
  _T_4152 = _RAND_105[2:0];
  _RAND_106 = {1{`RANDOM}};
  _T_4148 = _RAND_106[2:0];
  _RAND_107 = {1{`RANDOM}};
  _T_4144 = _RAND_107[2:0];
  _RAND_108 = {1{`RANDOM}};
  _T_4140 = _RAND_108[2:0];
  _RAND_109 = {1{`RANDOM}};
  _T_4136 = _RAND_109[2:0];
  _RAND_110 = {1{`RANDOM}};
  _T_4132 = _RAND_110[2:0];
  _RAND_111 = {1{`RANDOM}};
  _T_4128 = _RAND_111[2:0];
  _RAND_112 = {1{`RANDOM}};
  _T_4124 = _RAND_112[2:0];
  _RAND_113 = {1{`RANDOM}};
  _T_4120 = _RAND_113[2:0];
  _RAND_114 = {1{`RANDOM}};
  _T_4116 = _RAND_114[2:0];
  _RAND_115 = {1{`RANDOM}};
  _T_4112 = _RAND_115[2:0];
  _RAND_116 = {1{`RANDOM}};
  _T_4108 = _RAND_116[2:0];
  _RAND_117 = {1{`RANDOM}};
  _T_4104 = _RAND_117[2:0];
  _RAND_118 = {1{`RANDOM}};
  _T_4100 = _RAND_118[2:0];
  _RAND_119 = {1{`RANDOM}};
  _T_4096 = _RAND_119[2:0];
  _RAND_120 = {1{`RANDOM}};
  _T_4092 = _RAND_120[2:0];
  _RAND_121 = {1{`RANDOM}};
  _T_4088 = _RAND_121[2:0];
  _RAND_122 = {1{`RANDOM}};
  _T_4084 = _RAND_122[2:0];
  _RAND_123 = {1{`RANDOM}};
  _T_4080 = _RAND_123[2:0];
  _RAND_124 = {1{`RANDOM}};
  _T_4076 = _RAND_124[2:0];
  _RAND_125 = {1{`RANDOM}};
  _T_4072 = _RAND_125[2:0];
  _RAND_126 = {1{`RANDOM}};
  _T_4068 = _RAND_126[2:0];
  _RAND_127 = {1{`RANDOM}};
  _T_4064 = _RAND_127[2:0];
  _RAND_128 = {1{`RANDOM}};
  _T_4060 = _RAND_128[2:0];
  _RAND_129 = {1{`RANDOM}};
  _T_4056 = _RAND_129[2:0];
  _RAND_130 = {1{`RANDOM}};
  _T_4052 = _RAND_130[2:0];
  _RAND_131 = {1{`RANDOM}};
  _T_4048 = _RAND_131[2:0];
  _RAND_132 = {1{`RANDOM}};
  _T_4044 = _RAND_132[2:0];
  _RAND_133 = {1{`RANDOM}};
  _T_4040 = _RAND_133[2:0];
  _RAND_134 = {1{`RANDOM}};
  _T_4036 = _RAND_134[2:0];
  _RAND_135 = {1{`RANDOM}};
  _T_4032 = _RAND_135[2:0];
  _RAND_136 = {1{`RANDOM}};
  _T_4028 = _RAND_136[2:0];
  _RAND_137 = {1{`RANDOM}};
  _T_4024 = _RAND_137[2:0];
  _RAND_138 = {1{`RANDOM}};
  _T_4020 = _RAND_138[2:0];
  _RAND_139 = {1{`RANDOM}};
  _T_4016 = _RAND_139[2:0];
  _RAND_140 = {1{`RANDOM}};
  _T_4012 = _RAND_140[2:0];
  _RAND_141 = {1{`RANDOM}};
  _T_4008 = _RAND_141[2:0];
  _RAND_142 = {1{`RANDOM}};
  _T_4004 = _RAND_142[2:0];
  _RAND_143 = {1{`RANDOM}};
  _T_4000 = _RAND_143[2:0];
  _RAND_144 = {1{`RANDOM}};
  _T_3996 = _RAND_144[2:0];
  _RAND_145 = {1{`RANDOM}};
  _T_3992 = _RAND_145[2:0];
  _RAND_146 = {1{`RANDOM}};
  _T_3988 = _RAND_146[2:0];
  _RAND_147 = {1{`RANDOM}};
  _T_3984 = _RAND_147[2:0];
  _RAND_148 = {1{`RANDOM}};
  _T_3980 = _RAND_148[2:0];
  _RAND_149 = {1{`RANDOM}};
  _T_3976 = _RAND_149[2:0];
  _RAND_150 = {1{`RANDOM}};
  uncacheable_miss_scnd_ff = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  imb_scnd_ff = _RAND_151[30:0];
  _RAND_152 = {1{`RANDOM}};
  ifu_bus_rid_ff = _RAND_152[2:0];
  _RAND_153 = {1{`RANDOM}};
  ifu_bus_rresp_ff = _RAND_153[1:0];
  _RAND_154 = {1{`RANDOM}};
  ifu_wr_data_comb_err_ff = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  way_status_mb_ff = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  tagv_mb_ff = _RAND_156[1:0];
  _RAND_157 = {1{`RANDOM}};
  reset_ic_ff = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  fetch_uncacheable_ff = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  miss_addr = _RAND_159[25:0];
  _RAND_160 = {1{`RANDOM}};
  ifc_region_acc_fault_f = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  bus_rd_addr_count = _RAND_161[2:0];
  _RAND_162 = {1{`RANDOM}};
  ic_act_miss_f_delayed = _RAND_162[0:0];
  _RAND_163 = {2{`RANDOM}};
  ifu_bus_rdata_ff = _RAND_163[63:0];
  _RAND_164 = {1{`RANDOM}};
  ic_miss_buff_data_0 = _RAND_164[31:0];
  _RAND_165 = {1{`RANDOM}};
  ic_miss_buff_data_1 = _RAND_165[31:0];
  _RAND_166 = {1{`RANDOM}};
  ic_miss_buff_data_2 = _RAND_166[31:0];
  _RAND_167 = {1{`RANDOM}};
  ic_miss_buff_data_3 = _RAND_167[31:0];
  _RAND_168 = {1{`RANDOM}};
  ic_miss_buff_data_4 = _RAND_168[31:0];
  _RAND_169 = {1{`RANDOM}};
  ic_miss_buff_data_5 = _RAND_169[31:0];
  _RAND_170 = {1{`RANDOM}};
  ic_miss_buff_data_6 = _RAND_170[31:0];
  _RAND_171 = {1{`RANDOM}};
  ic_miss_buff_data_7 = _RAND_171[31:0];
  _RAND_172 = {1{`RANDOM}};
  ic_miss_buff_data_8 = _RAND_172[31:0];
  _RAND_173 = {1{`RANDOM}};
  ic_miss_buff_data_9 = _RAND_173[31:0];
  _RAND_174 = {1{`RANDOM}};
  ic_miss_buff_data_10 = _RAND_174[31:0];
  _RAND_175 = {1{`RANDOM}};
  ic_miss_buff_data_11 = _RAND_175[31:0];
  _RAND_176 = {1{`RANDOM}};
  ic_miss_buff_data_12 = _RAND_176[31:0];
  _RAND_177 = {1{`RANDOM}};
  ic_miss_buff_data_13 = _RAND_177[31:0];
  _RAND_178 = {1{`RANDOM}};
  ic_miss_buff_data_14 = _RAND_178[31:0];
  _RAND_179 = {1{`RANDOM}};
  ic_miss_buff_data_15 = _RAND_179[31:0];
  _RAND_180 = {1{`RANDOM}};
  ic_crit_wd_rdy_new_ff = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  ic_miss_buff_data_error = _RAND_181[7:0];
  _RAND_182 = {1{`RANDOM}};
  ic_debug_ict_array_sel_ff = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  ic_tag_valid_out_1_0 = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  ic_tag_valid_out_1_1 = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  ic_tag_valid_out_1_2 = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  ic_tag_valid_out_1_3 = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  ic_tag_valid_out_1_4 = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  ic_tag_valid_out_1_5 = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  ic_tag_valid_out_1_6 = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  ic_tag_valid_out_1_7 = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  ic_tag_valid_out_1_8 = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  ic_tag_valid_out_1_9 = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  ic_tag_valid_out_1_10 = _RAND_193[0:0];
  _RAND_194 = {1{`RANDOM}};
  ic_tag_valid_out_1_11 = _RAND_194[0:0];
  _RAND_195 = {1{`RANDOM}};
  ic_tag_valid_out_1_12 = _RAND_195[0:0];
  _RAND_196 = {1{`RANDOM}};
  ic_tag_valid_out_1_13 = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  ic_tag_valid_out_1_14 = _RAND_197[0:0];
  _RAND_198 = {1{`RANDOM}};
  ic_tag_valid_out_1_15 = _RAND_198[0:0];
  _RAND_199 = {1{`RANDOM}};
  ic_tag_valid_out_1_16 = _RAND_199[0:0];
  _RAND_200 = {1{`RANDOM}};
  ic_tag_valid_out_1_17 = _RAND_200[0:0];
  _RAND_201 = {1{`RANDOM}};
  ic_tag_valid_out_1_18 = _RAND_201[0:0];
  _RAND_202 = {1{`RANDOM}};
  ic_tag_valid_out_1_19 = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  ic_tag_valid_out_1_20 = _RAND_203[0:0];
  _RAND_204 = {1{`RANDOM}};
  ic_tag_valid_out_1_21 = _RAND_204[0:0];
  _RAND_205 = {1{`RANDOM}};
  ic_tag_valid_out_1_22 = _RAND_205[0:0];
  _RAND_206 = {1{`RANDOM}};
  ic_tag_valid_out_1_23 = _RAND_206[0:0];
  _RAND_207 = {1{`RANDOM}};
  ic_tag_valid_out_1_24 = _RAND_207[0:0];
  _RAND_208 = {1{`RANDOM}};
  ic_tag_valid_out_1_25 = _RAND_208[0:0];
  _RAND_209 = {1{`RANDOM}};
  ic_tag_valid_out_1_26 = _RAND_209[0:0];
  _RAND_210 = {1{`RANDOM}};
  ic_tag_valid_out_1_27 = _RAND_210[0:0];
  _RAND_211 = {1{`RANDOM}};
  ic_tag_valid_out_1_28 = _RAND_211[0:0];
  _RAND_212 = {1{`RANDOM}};
  ic_tag_valid_out_1_29 = _RAND_212[0:0];
  _RAND_213 = {1{`RANDOM}};
  ic_tag_valid_out_1_30 = _RAND_213[0:0];
  _RAND_214 = {1{`RANDOM}};
  ic_tag_valid_out_1_31 = _RAND_214[0:0];
  _RAND_215 = {1{`RANDOM}};
  ic_tag_valid_out_1_32 = _RAND_215[0:0];
  _RAND_216 = {1{`RANDOM}};
  ic_tag_valid_out_1_33 = _RAND_216[0:0];
  _RAND_217 = {1{`RANDOM}};
  ic_tag_valid_out_1_34 = _RAND_217[0:0];
  _RAND_218 = {1{`RANDOM}};
  ic_tag_valid_out_1_35 = _RAND_218[0:0];
  _RAND_219 = {1{`RANDOM}};
  ic_tag_valid_out_1_36 = _RAND_219[0:0];
  _RAND_220 = {1{`RANDOM}};
  ic_tag_valid_out_1_37 = _RAND_220[0:0];
  _RAND_221 = {1{`RANDOM}};
  ic_tag_valid_out_1_38 = _RAND_221[0:0];
  _RAND_222 = {1{`RANDOM}};
  ic_tag_valid_out_1_39 = _RAND_222[0:0];
  _RAND_223 = {1{`RANDOM}};
  ic_tag_valid_out_1_40 = _RAND_223[0:0];
  _RAND_224 = {1{`RANDOM}};
  ic_tag_valid_out_1_41 = _RAND_224[0:0];
  _RAND_225 = {1{`RANDOM}};
  ic_tag_valid_out_1_42 = _RAND_225[0:0];
  _RAND_226 = {1{`RANDOM}};
  ic_tag_valid_out_1_43 = _RAND_226[0:0];
  _RAND_227 = {1{`RANDOM}};
  ic_tag_valid_out_1_44 = _RAND_227[0:0];
  _RAND_228 = {1{`RANDOM}};
  ic_tag_valid_out_1_45 = _RAND_228[0:0];
  _RAND_229 = {1{`RANDOM}};
  ic_tag_valid_out_1_46 = _RAND_229[0:0];
  _RAND_230 = {1{`RANDOM}};
  ic_tag_valid_out_1_47 = _RAND_230[0:0];
  _RAND_231 = {1{`RANDOM}};
  ic_tag_valid_out_1_48 = _RAND_231[0:0];
  _RAND_232 = {1{`RANDOM}};
  ic_tag_valid_out_1_49 = _RAND_232[0:0];
  _RAND_233 = {1{`RANDOM}};
  ic_tag_valid_out_1_50 = _RAND_233[0:0];
  _RAND_234 = {1{`RANDOM}};
  ic_tag_valid_out_1_51 = _RAND_234[0:0];
  _RAND_235 = {1{`RANDOM}};
  ic_tag_valid_out_1_52 = _RAND_235[0:0];
  _RAND_236 = {1{`RANDOM}};
  ic_tag_valid_out_1_53 = _RAND_236[0:0];
  _RAND_237 = {1{`RANDOM}};
  ic_tag_valid_out_1_54 = _RAND_237[0:0];
  _RAND_238 = {1{`RANDOM}};
  ic_tag_valid_out_1_55 = _RAND_238[0:0];
  _RAND_239 = {1{`RANDOM}};
  ic_tag_valid_out_1_56 = _RAND_239[0:0];
  _RAND_240 = {1{`RANDOM}};
  ic_tag_valid_out_1_57 = _RAND_240[0:0];
  _RAND_241 = {1{`RANDOM}};
  ic_tag_valid_out_1_58 = _RAND_241[0:0];
  _RAND_242 = {1{`RANDOM}};
  ic_tag_valid_out_1_59 = _RAND_242[0:0];
  _RAND_243 = {1{`RANDOM}};
  ic_tag_valid_out_1_60 = _RAND_243[0:0];
  _RAND_244 = {1{`RANDOM}};
  ic_tag_valid_out_1_61 = _RAND_244[0:0];
  _RAND_245 = {1{`RANDOM}};
  ic_tag_valid_out_1_62 = _RAND_245[0:0];
  _RAND_246 = {1{`RANDOM}};
  ic_tag_valid_out_1_63 = _RAND_246[0:0];
  _RAND_247 = {1{`RANDOM}};
  ic_tag_valid_out_1_64 = _RAND_247[0:0];
  _RAND_248 = {1{`RANDOM}};
  ic_tag_valid_out_1_65 = _RAND_248[0:0];
  _RAND_249 = {1{`RANDOM}};
  ic_tag_valid_out_1_66 = _RAND_249[0:0];
  _RAND_250 = {1{`RANDOM}};
  ic_tag_valid_out_1_67 = _RAND_250[0:0];
  _RAND_251 = {1{`RANDOM}};
  ic_tag_valid_out_1_68 = _RAND_251[0:0];
  _RAND_252 = {1{`RANDOM}};
  ic_tag_valid_out_1_69 = _RAND_252[0:0];
  _RAND_253 = {1{`RANDOM}};
  ic_tag_valid_out_1_70 = _RAND_253[0:0];
  _RAND_254 = {1{`RANDOM}};
  ic_tag_valid_out_1_71 = _RAND_254[0:0];
  _RAND_255 = {1{`RANDOM}};
  ic_tag_valid_out_1_72 = _RAND_255[0:0];
  _RAND_256 = {1{`RANDOM}};
  ic_tag_valid_out_1_73 = _RAND_256[0:0];
  _RAND_257 = {1{`RANDOM}};
  ic_tag_valid_out_1_74 = _RAND_257[0:0];
  _RAND_258 = {1{`RANDOM}};
  ic_tag_valid_out_1_75 = _RAND_258[0:0];
  _RAND_259 = {1{`RANDOM}};
  ic_tag_valid_out_1_76 = _RAND_259[0:0];
  _RAND_260 = {1{`RANDOM}};
  ic_tag_valid_out_1_77 = _RAND_260[0:0];
  _RAND_261 = {1{`RANDOM}};
  ic_tag_valid_out_1_78 = _RAND_261[0:0];
  _RAND_262 = {1{`RANDOM}};
  ic_tag_valid_out_1_79 = _RAND_262[0:0];
  _RAND_263 = {1{`RANDOM}};
  ic_tag_valid_out_1_80 = _RAND_263[0:0];
  _RAND_264 = {1{`RANDOM}};
  ic_tag_valid_out_1_81 = _RAND_264[0:0];
  _RAND_265 = {1{`RANDOM}};
  ic_tag_valid_out_1_82 = _RAND_265[0:0];
  _RAND_266 = {1{`RANDOM}};
  ic_tag_valid_out_1_83 = _RAND_266[0:0];
  _RAND_267 = {1{`RANDOM}};
  ic_tag_valid_out_1_84 = _RAND_267[0:0];
  _RAND_268 = {1{`RANDOM}};
  ic_tag_valid_out_1_85 = _RAND_268[0:0];
  _RAND_269 = {1{`RANDOM}};
  ic_tag_valid_out_1_86 = _RAND_269[0:0];
  _RAND_270 = {1{`RANDOM}};
  ic_tag_valid_out_1_87 = _RAND_270[0:0];
  _RAND_271 = {1{`RANDOM}};
  ic_tag_valid_out_1_88 = _RAND_271[0:0];
  _RAND_272 = {1{`RANDOM}};
  ic_tag_valid_out_1_89 = _RAND_272[0:0];
  _RAND_273 = {1{`RANDOM}};
  ic_tag_valid_out_1_90 = _RAND_273[0:0];
  _RAND_274 = {1{`RANDOM}};
  ic_tag_valid_out_1_91 = _RAND_274[0:0];
  _RAND_275 = {1{`RANDOM}};
  ic_tag_valid_out_1_92 = _RAND_275[0:0];
  _RAND_276 = {1{`RANDOM}};
  ic_tag_valid_out_1_93 = _RAND_276[0:0];
  _RAND_277 = {1{`RANDOM}};
  ic_tag_valid_out_1_94 = _RAND_277[0:0];
  _RAND_278 = {1{`RANDOM}};
  ic_tag_valid_out_1_95 = _RAND_278[0:0];
  _RAND_279 = {1{`RANDOM}};
  ic_tag_valid_out_1_96 = _RAND_279[0:0];
  _RAND_280 = {1{`RANDOM}};
  ic_tag_valid_out_1_97 = _RAND_280[0:0];
  _RAND_281 = {1{`RANDOM}};
  ic_tag_valid_out_1_98 = _RAND_281[0:0];
  _RAND_282 = {1{`RANDOM}};
  ic_tag_valid_out_1_99 = _RAND_282[0:0];
  _RAND_283 = {1{`RANDOM}};
  ic_tag_valid_out_1_100 = _RAND_283[0:0];
  _RAND_284 = {1{`RANDOM}};
  ic_tag_valid_out_1_101 = _RAND_284[0:0];
  _RAND_285 = {1{`RANDOM}};
  ic_tag_valid_out_1_102 = _RAND_285[0:0];
  _RAND_286 = {1{`RANDOM}};
  ic_tag_valid_out_1_103 = _RAND_286[0:0];
  _RAND_287 = {1{`RANDOM}};
  ic_tag_valid_out_1_104 = _RAND_287[0:0];
  _RAND_288 = {1{`RANDOM}};
  ic_tag_valid_out_1_105 = _RAND_288[0:0];
  _RAND_289 = {1{`RANDOM}};
  ic_tag_valid_out_1_106 = _RAND_289[0:0];
  _RAND_290 = {1{`RANDOM}};
  ic_tag_valid_out_1_107 = _RAND_290[0:0];
  _RAND_291 = {1{`RANDOM}};
  ic_tag_valid_out_1_108 = _RAND_291[0:0];
  _RAND_292 = {1{`RANDOM}};
  ic_tag_valid_out_1_109 = _RAND_292[0:0];
  _RAND_293 = {1{`RANDOM}};
  ic_tag_valid_out_1_110 = _RAND_293[0:0];
  _RAND_294 = {1{`RANDOM}};
  ic_tag_valid_out_1_111 = _RAND_294[0:0];
  _RAND_295 = {1{`RANDOM}};
  ic_tag_valid_out_1_112 = _RAND_295[0:0];
  _RAND_296 = {1{`RANDOM}};
  ic_tag_valid_out_1_113 = _RAND_296[0:0];
  _RAND_297 = {1{`RANDOM}};
  ic_tag_valid_out_1_114 = _RAND_297[0:0];
  _RAND_298 = {1{`RANDOM}};
  ic_tag_valid_out_1_115 = _RAND_298[0:0];
  _RAND_299 = {1{`RANDOM}};
  ic_tag_valid_out_1_116 = _RAND_299[0:0];
  _RAND_300 = {1{`RANDOM}};
  ic_tag_valid_out_1_117 = _RAND_300[0:0];
  _RAND_301 = {1{`RANDOM}};
  ic_tag_valid_out_1_118 = _RAND_301[0:0];
  _RAND_302 = {1{`RANDOM}};
  ic_tag_valid_out_1_119 = _RAND_302[0:0];
  _RAND_303 = {1{`RANDOM}};
  ic_tag_valid_out_1_120 = _RAND_303[0:0];
  _RAND_304 = {1{`RANDOM}};
  ic_tag_valid_out_1_121 = _RAND_304[0:0];
  _RAND_305 = {1{`RANDOM}};
  ic_tag_valid_out_1_122 = _RAND_305[0:0];
  _RAND_306 = {1{`RANDOM}};
  ic_tag_valid_out_1_123 = _RAND_306[0:0];
  _RAND_307 = {1{`RANDOM}};
  ic_tag_valid_out_1_124 = _RAND_307[0:0];
  _RAND_308 = {1{`RANDOM}};
  ic_tag_valid_out_1_125 = _RAND_308[0:0];
  _RAND_309 = {1{`RANDOM}};
  ic_tag_valid_out_1_126 = _RAND_309[0:0];
  _RAND_310 = {1{`RANDOM}};
  ic_tag_valid_out_1_127 = _RAND_310[0:0];
  _RAND_311 = {1{`RANDOM}};
  ic_tag_valid_out_0_0 = _RAND_311[0:0];
  _RAND_312 = {1{`RANDOM}};
  ic_tag_valid_out_0_1 = _RAND_312[0:0];
  _RAND_313 = {1{`RANDOM}};
  ic_tag_valid_out_0_2 = _RAND_313[0:0];
  _RAND_314 = {1{`RANDOM}};
  ic_tag_valid_out_0_3 = _RAND_314[0:0];
  _RAND_315 = {1{`RANDOM}};
  ic_tag_valid_out_0_4 = _RAND_315[0:0];
  _RAND_316 = {1{`RANDOM}};
  ic_tag_valid_out_0_5 = _RAND_316[0:0];
  _RAND_317 = {1{`RANDOM}};
  ic_tag_valid_out_0_6 = _RAND_317[0:0];
  _RAND_318 = {1{`RANDOM}};
  ic_tag_valid_out_0_7 = _RAND_318[0:0];
  _RAND_319 = {1{`RANDOM}};
  ic_tag_valid_out_0_8 = _RAND_319[0:0];
  _RAND_320 = {1{`RANDOM}};
  ic_tag_valid_out_0_9 = _RAND_320[0:0];
  _RAND_321 = {1{`RANDOM}};
  ic_tag_valid_out_0_10 = _RAND_321[0:0];
  _RAND_322 = {1{`RANDOM}};
  ic_tag_valid_out_0_11 = _RAND_322[0:0];
  _RAND_323 = {1{`RANDOM}};
  ic_tag_valid_out_0_12 = _RAND_323[0:0];
  _RAND_324 = {1{`RANDOM}};
  ic_tag_valid_out_0_13 = _RAND_324[0:0];
  _RAND_325 = {1{`RANDOM}};
  ic_tag_valid_out_0_14 = _RAND_325[0:0];
  _RAND_326 = {1{`RANDOM}};
  ic_tag_valid_out_0_15 = _RAND_326[0:0];
  _RAND_327 = {1{`RANDOM}};
  ic_tag_valid_out_0_16 = _RAND_327[0:0];
  _RAND_328 = {1{`RANDOM}};
  ic_tag_valid_out_0_17 = _RAND_328[0:0];
  _RAND_329 = {1{`RANDOM}};
  ic_tag_valid_out_0_18 = _RAND_329[0:0];
  _RAND_330 = {1{`RANDOM}};
  ic_tag_valid_out_0_19 = _RAND_330[0:0];
  _RAND_331 = {1{`RANDOM}};
  ic_tag_valid_out_0_20 = _RAND_331[0:0];
  _RAND_332 = {1{`RANDOM}};
  ic_tag_valid_out_0_21 = _RAND_332[0:0];
  _RAND_333 = {1{`RANDOM}};
  ic_tag_valid_out_0_22 = _RAND_333[0:0];
  _RAND_334 = {1{`RANDOM}};
  ic_tag_valid_out_0_23 = _RAND_334[0:0];
  _RAND_335 = {1{`RANDOM}};
  ic_tag_valid_out_0_24 = _RAND_335[0:0];
  _RAND_336 = {1{`RANDOM}};
  ic_tag_valid_out_0_25 = _RAND_336[0:0];
  _RAND_337 = {1{`RANDOM}};
  ic_tag_valid_out_0_26 = _RAND_337[0:0];
  _RAND_338 = {1{`RANDOM}};
  ic_tag_valid_out_0_27 = _RAND_338[0:0];
  _RAND_339 = {1{`RANDOM}};
  ic_tag_valid_out_0_28 = _RAND_339[0:0];
  _RAND_340 = {1{`RANDOM}};
  ic_tag_valid_out_0_29 = _RAND_340[0:0];
  _RAND_341 = {1{`RANDOM}};
  ic_tag_valid_out_0_30 = _RAND_341[0:0];
  _RAND_342 = {1{`RANDOM}};
  ic_tag_valid_out_0_31 = _RAND_342[0:0];
  _RAND_343 = {1{`RANDOM}};
  ic_tag_valid_out_0_32 = _RAND_343[0:0];
  _RAND_344 = {1{`RANDOM}};
  ic_tag_valid_out_0_33 = _RAND_344[0:0];
  _RAND_345 = {1{`RANDOM}};
  ic_tag_valid_out_0_34 = _RAND_345[0:0];
  _RAND_346 = {1{`RANDOM}};
  ic_tag_valid_out_0_35 = _RAND_346[0:0];
  _RAND_347 = {1{`RANDOM}};
  ic_tag_valid_out_0_36 = _RAND_347[0:0];
  _RAND_348 = {1{`RANDOM}};
  ic_tag_valid_out_0_37 = _RAND_348[0:0];
  _RAND_349 = {1{`RANDOM}};
  ic_tag_valid_out_0_38 = _RAND_349[0:0];
  _RAND_350 = {1{`RANDOM}};
  ic_tag_valid_out_0_39 = _RAND_350[0:0];
  _RAND_351 = {1{`RANDOM}};
  ic_tag_valid_out_0_40 = _RAND_351[0:0];
  _RAND_352 = {1{`RANDOM}};
  ic_tag_valid_out_0_41 = _RAND_352[0:0];
  _RAND_353 = {1{`RANDOM}};
  ic_tag_valid_out_0_42 = _RAND_353[0:0];
  _RAND_354 = {1{`RANDOM}};
  ic_tag_valid_out_0_43 = _RAND_354[0:0];
  _RAND_355 = {1{`RANDOM}};
  ic_tag_valid_out_0_44 = _RAND_355[0:0];
  _RAND_356 = {1{`RANDOM}};
  ic_tag_valid_out_0_45 = _RAND_356[0:0];
  _RAND_357 = {1{`RANDOM}};
  ic_tag_valid_out_0_46 = _RAND_357[0:0];
  _RAND_358 = {1{`RANDOM}};
  ic_tag_valid_out_0_47 = _RAND_358[0:0];
  _RAND_359 = {1{`RANDOM}};
  ic_tag_valid_out_0_48 = _RAND_359[0:0];
  _RAND_360 = {1{`RANDOM}};
  ic_tag_valid_out_0_49 = _RAND_360[0:0];
  _RAND_361 = {1{`RANDOM}};
  ic_tag_valid_out_0_50 = _RAND_361[0:0];
  _RAND_362 = {1{`RANDOM}};
  ic_tag_valid_out_0_51 = _RAND_362[0:0];
  _RAND_363 = {1{`RANDOM}};
  ic_tag_valid_out_0_52 = _RAND_363[0:0];
  _RAND_364 = {1{`RANDOM}};
  ic_tag_valid_out_0_53 = _RAND_364[0:0];
  _RAND_365 = {1{`RANDOM}};
  ic_tag_valid_out_0_54 = _RAND_365[0:0];
  _RAND_366 = {1{`RANDOM}};
  ic_tag_valid_out_0_55 = _RAND_366[0:0];
  _RAND_367 = {1{`RANDOM}};
  ic_tag_valid_out_0_56 = _RAND_367[0:0];
  _RAND_368 = {1{`RANDOM}};
  ic_tag_valid_out_0_57 = _RAND_368[0:0];
  _RAND_369 = {1{`RANDOM}};
  ic_tag_valid_out_0_58 = _RAND_369[0:0];
  _RAND_370 = {1{`RANDOM}};
  ic_tag_valid_out_0_59 = _RAND_370[0:0];
  _RAND_371 = {1{`RANDOM}};
  ic_tag_valid_out_0_60 = _RAND_371[0:0];
  _RAND_372 = {1{`RANDOM}};
  ic_tag_valid_out_0_61 = _RAND_372[0:0];
  _RAND_373 = {1{`RANDOM}};
  ic_tag_valid_out_0_62 = _RAND_373[0:0];
  _RAND_374 = {1{`RANDOM}};
  ic_tag_valid_out_0_63 = _RAND_374[0:0];
  _RAND_375 = {1{`RANDOM}};
  ic_tag_valid_out_0_64 = _RAND_375[0:0];
  _RAND_376 = {1{`RANDOM}};
  ic_tag_valid_out_0_65 = _RAND_376[0:0];
  _RAND_377 = {1{`RANDOM}};
  ic_tag_valid_out_0_66 = _RAND_377[0:0];
  _RAND_378 = {1{`RANDOM}};
  ic_tag_valid_out_0_67 = _RAND_378[0:0];
  _RAND_379 = {1{`RANDOM}};
  ic_tag_valid_out_0_68 = _RAND_379[0:0];
  _RAND_380 = {1{`RANDOM}};
  ic_tag_valid_out_0_69 = _RAND_380[0:0];
  _RAND_381 = {1{`RANDOM}};
  ic_tag_valid_out_0_70 = _RAND_381[0:0];
  _RAND_382 = {1{`RANDOM}};
  ic_tag_valid_out_0_71 = _RAND_382[0:0];
  _RAND_383 = {1{`RANDOM}};
  ic_tag_valid_out_0_72 = _RAND_383[0:0];
  _RAND_384 = {1{`RANDOM}};
  ic_tag_valid_out_0_73 = _RAND_384[0:0];
  _RAND_385 = {1{`RANDOM}};
  ic_tag_valid_out_0_74 = _RAND_385[0:0];
  _RAND_386 = {1{`RANDOM}};
  ic_tag_valid_out_0_75 = _RAND_386[0:0];
  _RAND_387 = {1{`RANDOM}};
  ic_tag_valid_out_0_76 = _RAND_387[0:0];
  _RAND_388 = {1{`RANDOM}};
  ic_tag_valid_out_0_77 = _RAND_388[0:0];
  _RAND_389 = {1{`RANDOM}};
  ic_tag_valid_out_0_78 = _RAND_389[0:0];
  _RAND_390 = {1{`RANDOM}};
  ic_tag_valid_out_0_79 = _RAND_390[0:0];
  _RAND_391 = {1{`RANDOM}};
  ic_tag_valid_out_0_80 = _RAND_391[0:0];
  _RAND_392 = {1{`RANDOM}};
  ic_tag_valid_out_0_81 = _RAND_392[0:0];
  _RAND_393 = {1{`RANDOM}};
  ic_tag_valid_out_0_82 = _RAND_393[0:0];
  _RAND_394 = {1{`RANDOM}};
  ic_tag_valid_out_0_83 = _RAND_394[0:0];
  _RAND_395 = {1{`RANDOM}};
  ic_tag_valid_out_0_84 = _RAND_395[0:0];
  _RAND_396 = {1{`RANDOM}};
  ic_tag_valid_out_0_85 = _RAND_396[0:0];
  _RAND_397 = {1{`RANDOM}};
  ic_tag_valid_out_0_86 = _RAND_397[0:0];
  _RAND_398 = {1{`RANDOM}};
  ic_tag_valid_out_0_87 = _RAND_398[0:0];
  _RAND_399 = {1{`RANDOM}};
  ic_tag_valid_out_0_88 = _RAND_399[0:0];
  _RAND_400 = {1{`RANDOM}};
  ic_tag_valid_out_0_89 = _RAND_400[0:0];
  _RAND_401 = {1{`RANDOM}};
  ic_tag_valid_out_0_90 = _RAND_401[0:0];
  _RAND_402 = {1{`RANDOM}};
  ic_tag_valid_out_0_91 = _RAND_402[0:0];
  _RAND_403 = {1{`RANDOM}};
  ic_tag_valid_out_0_92 = _RAND_403[0:0];
  _RAND_404 = {1{`RANDOM}};
  ic_tag_valid_out_0_93 = _RAND_404[0:0];
  _RAND_405 = {1{`RANDOM}};
  ic_tag_valid_out_0_94 = _RAND_405[0:0];
  _RAND_406 = {1{`RANDOM}};
  ic_tag_valid_out_0_95 = _RAND_406[0:0];
  _RAND_407 = {1{`RANDOM}};
  ic_tag_valid_out_0_96 = _RAND_407[0:0];
  _RAND_408 = {1{`RANDOM}};
  ic_tag_valid_out_0_97 = _RAND_408[0:0];
  _RAND_409 = {1{`RANDOM}};
  ic_tag_valid_out_0_98 = _RAND_409[0:0];
  _RAND_410 = {1{`RANDOM}};
  ic_tag_valid_out_0_99 = _RAND_410[0:0];
  _RAND_411 = {1{`RANDOM}};
  ic_tag_valid_out_0_100 = _RAND_411[0:0];
  _RAND_412 = {1{`RANDOM}};
  ic_tag_valid_out_0_101 = _RAND_412[0:0];
  _RAND_413 = {1{`RANDOM}};
  ic_tag_valid_out_0_102 = _RAND_413[0:0];
  _RAND_414 = {1{`RANDOM}};
  ic_tag_valid_out_0_103 = _RAND_414[0:0];
  _RAND_415 = {1{`RANDOM}};
  ic_tag_valid_out_0_104 = _RAND_415[0:0];
  _RAND_416 = {1{`RANDOM}};
  ic_tag_valid_out_0_105 = _RAND_416[0:0];
  _RAND_417 = {1{`RANDOM}};
  ic_tag_valid_out_0_106 = _RAND_417[0:0];
  _RAND_418 = {1{`RANDOM}};
  ic_tag_valid_out_0_107 = _RAND_418[0:0];
  _RAND_419 = {1{`RANDOM}};
  ic_tag_valid_out_0_108 = _RAND_419[0:0];
  _RAND_420 = {1{`RANDOM}};
  ic_tag_valid_out_0_109 = _RAND_420[0:0];
  _RAND_421 = {1{`RANDOM}};
  ic_tag_valid_out_0_110 = _RAND_421[0:0];
  _RAND_422 = {1{`RANDOM}};
  ic_tag_valid_out_0_111 = _RAND_422[0:0];
  _RAND_423 = {1{`RANDOM}};
  ic_tag_valid_out_0_112 = _RAND_423[0:0];
  _RAND_424 = {1{`RANDOM}};
  ic_tag_valid_out_0_113 = _RAND_424[0:0];
  _RAND_425 = {1{`RANDOM}};
  ic_tag_valid_out_0_114 = _RAND_425[0:0];
  _RAND_426 = {1{`RANDOM}};
  ic_tag_valid_out_0_115 = _RAND_426[0:0];
  _RAND_427 = {1{`RANDOM}};
  ic_tag_valid_out_0_116 = _RAND_427[0:0];
  _RAND_428 = {1{`RANDOM}};
  ic_tag_valid_out_0_117 = _RAND_428[0:0];
  _RAND_429 = {1{`RANDOM}};
  ic_tag_valid_out_0_118 = _RAND_429[0:0];
  _RAND_430 = {1{`RANDOM}};
  ic_tag_valid_out_0_119 = _RAND_430[0:0];
  _RAND_431 = {1{`RANDOM}};
  ic_tag_valid_out_0_120 = _RAND_431[0:0];
  _RAND_432 = {1{`RANDOM}};
  ic_tag_valid_out_0_121 = _RAND_432[0:0];
  _RAND_433 = {1{`RANDOM}};
  ic_tag_valid_out_0_122 = _RAND_433[0:0];
  _RAND_434 = {1{`RANDOM}};
  ic_tag_valid_out_0_123 = _RAND_434[0:0];
  _RAND_435 = {1{`RANDOM}};
  ic_tag_valid_out_0_124 = _RAND_435[0:0];
  _RAND_436 = {1{`RANDOM}};
  ic_tag_valid_out_0_125 = _RAND_436[0:0];
  _RAND_437 = {1{`RANDOM}};
  ic_tag_valid_out_0_126 = _RAND_437[0:0];
  _RAND_438 = {1{`RANDOM}};
  ic_tag_valid_out_0_127 = _RAND_438[0:0];
  _RAND_439 = {1{`RANDOM}};
  ic_debug_way_ff = _RAND_439[1:0];
  _RAND_440 = {1{`RANDOM}};
  ic_debug_rd_en_ff = _RAND_440[0:0];
  _RAND_441 = {3{`RANDOM}};
  _T_1209 = _RAND_441[70:0];
  _RAND_442 = {1{`RANDOM}};
  perr_ic_index_ff = _RAND_442[5:0];
  _RAND_443 = {1{`RANDOM}};
  dma_sb_err_state_ff = _RAND_443[0:0];
  _RAND_444 = {1{`RANDOM}};
  ifu_bus_cmd_valid = _RAND_444[0:0];
  _RAND_445 = {1{`RANDOM}};
  bus_cmd_beat_count = _RAND_445[2:0];
  _RAND_446 = {1{`RANDOM}};
  ifu_bus_arready_unq_ff = _RAND_446[0:0];
  _RAND_447 = {1{`RANDOM}};
  ifu_bus_arvalid_ff = _RAND_447[0:0];
  _RAND_448 = {1{`RANDOM}};
  ifc_dma_access_ok_prev = _RAND_448[0:0];
  _RAND_449 = {2{`RANDOM}};
  iccm_ecc_corr_data_ff = _RAND_449[38:0];
  _RAND_450 = {1{`RANDOM}};
  dma_mem_addr_ff = _RAND_450[1:0];
  _RAND_451 = {1{`RANDOM}};
  dma_mem_tag_ff = _RAND_451[2:0];
  _RAND_452 = {1{`RANDOM}};
  iccm_dma_rtag = _RAND_452[2:0];
  _RAND_453 = {1{`RANDOM}};
  iccm_dma_rvalid = _RAND_453[0:0];
  _RAND_454 = {2{`RANDOM}};
  iccm_dma_rdata = _RAND_454[63:0];
  _RAND_455 = {1{`RANDOM}};
  iccm_ecc_corr_index_ff = _RAND_455[13:0];
  _RAND_456 = {1{`RANDOM}};
  iccm_rd_ecc_single_err_ff = _RAND_456[0:0];
  _RAND_457 = {1{`RANDOM}};
  iccm_rw_addr_f = _RAND_457[13:0];
  _RAND_458 = {1{`RANDOM}};
  ifu_status_wr_addr_ff = _RAND_458[6:0];
  _RAND_459 = {1{`RANDOM}};
  way_status_wr_en_ff = _RAND_459[0:0];
  _RAND_460 = {1{`RANDOM}};
  way_status_new_ff = _RAND_460[2:0];
  _RAND_461 = {1{`RANDOM}};
  ifu_tag_wren_ff = _RAND_461[1:0];
  _RAND_462 = {1{`RANDOM}};
  ic_valid_ff = _RAND_462[0:0];
  _RAND_463 = {1{`RANDOM}};
  _T_10115 = _RAND_463[0:0];
  _RAND_464 = {1{`RANDOM}};
  _T_10116 = _RAND_464[0:0];
  _RAND_465 = {1{`RANDOM}};
  _T_10117 = _RAND_465[0:0];
  _RAND_466 = {1{`RANDOM}};
  _T_10121 = _RAND_466[0:0];
  _RAND_467 = {1{`RANDOM}};
  _T_10122 = _RAND_467[0:0];
  _RAND_468 = {1{`RANDOM}};
  _T_10145 = _RAND_468[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      flush_final_f <= 1'h0;
    end else begin
      flush_final_f <= io_exu_flush_final;
    end
    if (reset) begin
      ifc_fetch_req_f_raw <= 1'h0;
    end else begin
      ifc_fetch_req_f_raw <= ifc_fetch_req_qual_bf;
    end
    if (reset) begin
      miss_state <= 3'h0;
    end else if (miss_state_en) begin
      if (_T_24) begin
        if (_T_26) begin
          miss_state <= 3'h1;
        end else begin
          miss_state <= 3'h2;
        end
      end else if (_T_31) begin
        if (_T_36) begin
          miss_state <= 3'h0;
        end else if (_T_40) begin
          miss_state <= 3'h3;
        end else if (_T_47) begin
          miss_state <= 3'h4;
        end else if (_T_51) begin
          miss_state <= 3'h0;
        end else if (_T_61) begin
          miss_state <= 3'h6;
        end else if (_T_71) begin
          miss_state <= 3'h6;
        end else if (_T_79) begin
          miss_state <= 3'h0;
        end else if (_T_84) begin
          miss_state <= 3'h2;
        end else begin
          miss_state <= 3'h0;
        end
      end else if (_T_102) begin
        miss_state <= 3'h0;
      end else if (_T_106) begin
        if (_T_113) begin
          miss_state <= 3'h2;
        end else begin
          miss_state <= 3'h0;
        end
      end else if (_T_121) begin
        if (_T_126) begin
          miss_state <= 3'h2;
        end else begin
          miss_state <= 3'h0;
        end
      end else if (_T_132) begin
        if (_T_137) begin
          miss_state <= 3'h5;
        end else if (_T_143) begin
          miss_state <= 3'h7;
        end else begin
          miss_state <= 3'h0;
        end
      end else if (_T_151) begin
        if (io_dec_tlu_force_halt) begin
          miss_state <= 3'h0;
        end else if (io_exu_flush_final) begin
          if (_T_32) begin
            miss_state <= 3'h0;
          end else begin
            miss_state <= 3'h2;
          end
        end else begin
          miss_state <= 3'h1;
        end
      end else if (_T_160) begin
        if (io_dec_tlu_force_halt) begin
          miss_state <= 3'h0;
        end else if (io_exu_flush_final) begin
          if (_T_32) begin
            miss_state <= 3'h0;
          end else begin
            miss_state <= 3'h2;
          end
        end else begin
          miss_state <= 3'h0;
        end
      end else begin
        miss_state <= 3'h0;
      end
    end
    if (reset) begin
      ifu_fetch_addr_int_f <= 31'h0;
    end else begin
      ifu_fetch_addr_int_f <= io_ifc_fetch_addr_bf;
    end
    if (reset) begin
      ifc_iccm_access_f <= 1'h0;
    end else begin
      ifc_iccm_access_f <= io_ifc_iccm_access_bf;
    end
    if (reset) begin
      ifc_region_acc_fault_final_f <= 1'h0;
    end else begin
      ifc_region_acc_fault_final_f <= io_ifc_region_acc_fault_bf;
    end
    if (reset) begin
      ifu_bus_rvalid_unq_ff <= 1'h0;
    end else if (io_ifu_bus_clk_en) begin
      ifu_bus_rvalid_unq_ff <= io_ifu_axi_rvalid;
    end
    if (reset) begin
      uncacheable_miss_ff <= 1'h0;
    end else if (scnd_miss_req) begin
      uncacheable_miss_ff <= uncacheable_miss_scnd_ff;
    end else if (!(sel_hold_imb)) begin
      uncacheable_miss_ff <= io_ifc_fetch_uncacheable_bf;
    end
    if (scnd_miss_req) begin
      imb_ff <= imb_scnd_ff;
    end else if (!(sel_hold_imb)) begin
      imb_ff <= io_ifc_fetch_addr_bf;
    end
    if (reset) begin
      way_status_mb_scnd_ff <= 1'h0;
    end else if (!(_T_19)) begin
      way_status_mb_scnd_ff <= way_status;
    end
    if (reset) begin
      _T_4484 <= 3'h0;
    end else if (_T_4483) begin
      _T_4484 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4480 <= 3'h0;
    end else if (_T_4479) begin
      _T_4480 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4476 <= 3'h0;
    end else if (_T_4475) begin
      _T_4476 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4472 <= 3'h0;
    end else if (_T_4471) begin
      _T_4472 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4468 <= 3'h0;
    end else if (_T_4467) begin
      _T_4468 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4464 <= 3'h0;
    end else if (_T_4463) begin
      _T_4464 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4460 <= 3'h0;
    end else if (_T_4459) begin
      _T_4460 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4456 <= 3'h0;
    end else if (_T_4455) begin
      _T_4456 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4452 <= 3'h0;
    end else if (_T_4451) begin
      _T_4452 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4448 <= 3'h0;
    end else if (_T_4447) begin
      _T_4448 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4444 <= 3'h0;
    end else if (_T_4443) begin
      _T_4444 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4440 <= 3'h0;
    end else if (_T_4439) begin
      _T_4440 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4436 <= 3'h0;
    end else if (_T_4435) begin
      _T_4436 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4432 <= 3'h0;
    end else if (_T_4431) begin
      _T_4432 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4428 <= 3'h0;
    end else if (_T_4427) begin
      _T_4428 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4424 <= 3'h0;
    end else if (_T_4423) begin
      _T_4424 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4420 <= 3'h0;
    end else if (_T_4419) begin
      _T_4420 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4416 <= 3'h0;
    end else if (_T_4415) begin
      _T_4416 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4412 <= 3'h0;
    end else if (_T_4411) begin
      _T_4412 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4408 <= 3'h0;
    end else if (_T_4407) begin
      _T_4408 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4404 <= 3'h0;
    end else if (_T_4403) begin
      _T_4404 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4400 <= 3'h0;
    end else if (_T_4399) begin
      _T_4400 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4396 <= 3'h0;
    end else if (_T_4395) begin
      _T_4396 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4392 <= 3'h0;
    end else if (_T_4391) begin
      _T_4392 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4388 <= 3'h0;
    end else if (_T_4387) begin
      _T_4388 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4384 <= 3'h0;
    end else if (_T_4383) begin
      _T_4384 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4380 <= 3'h0;
    end else if (_T_4379) begin
      _T_4380 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4376 <= 3'h0;
    end else if (_T_4375) begin
      _T_4376 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4372 <= 3'h0;
    end else if (_T_4371) begin
      _T_4372 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4368 <= 3'h0;
    end else if (_T_4367) begin
      _T_4368 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4364 <= 3'h0;
    end else if (_T_4363) begin
      _T_4364 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4360 <= 3'h0;
    end else if (_T_4359) begin
      _T_4360 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4356 <= 3'h0;
    end else if (_T_4355) begin
      _T_4356 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4352 <= 3'h0;
    end else if (_T_4351) begin
      _T_4352 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4348 <= 3'h0;
    end else if (_T_4347) begin
      _T_4348 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4344 <= 3'h0;
    end else if (_T_4343) begin
      _T_4344 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4340 <= 3'h0;
    end else if (_T_4339) begin
      _T_4340 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4336 <= 3'h0;
    end else if (_T_4335) begin
      _T_4336 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4332 <= 3'h0;
    end else if (_T_4331) begin
      _T_4332 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4328 <= 3'h0;
    end else if (_T_4327) begin
      _T_4328 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4324 <= 3'h0;
    end else if (_T_4323) begin
      _T_4324 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4320 <= 3'h0;
    end else if (_T_4319) begin
      _T_4320 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4316 <= 3'h0;
    end else if (_T_4315) begin
      _T_4316 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4312 <= 3'h0;
    end else if (_T_4311) begin
      _T_4312 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4308 <= 3'h0;
    end else if (_T_4307) begin
      _T_4308 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4304 <= 3'h0;
    end else if (_T_4303) begin
      _T_4304 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4300 <= 3'h0;
    end else if (_T_4299) begin
      _T_4300 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4296 <= 3'h0;
    end else if (_T_4295) begin
      _T_4296 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4292 <= 3'h0;
    end else if (_T_4291) begin
      _T_4292 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4288 <= 3'h0;
    end else if (_T_4287) begin
      _T_4288 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4284 <= 3'h0;
    end else if (_T_4283) begin
      _T_4284 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4280 <= 3'h0;
    end else if (_T_4279) begin
      _T_4280 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4276 <= 3'h0;
    end else if (_T_4275) begin
      _T_4276 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4272 <= 3'h0;
    end else if (_T_4271) begin
      _T_4272 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4268 <= 3'h0;
    end else if (_T_4267) begin
      _T_4268 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4264 <= 3'h0;
    end else if (_T_4263) begin
      _T_4264 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4260 <= 3'h0;
    end else if (_T_4259) begin
      _T_4260 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4256 <= 3'h0;
    end else if (_T_4255) begin
      _T_4256 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4252 <= 3'h0;
    end else if (_T_4251) begin
      _T_4252 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4248 <= 3'h0;
    end else if (_T_4247) begin
      _T_4248 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4244 <= 3'h0;
    end else if (_T_4243) begin
      _T_4244 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4240 <= 3'h0;
    end else if (_T_4239) begin
      _T_4240 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4236 <= 3'h0;
    end else if (_T_4235) begin
      _T_4236 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4232 <= 3'h0;
    end else if (_T_4231) begin
      _T_4232 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4228 <= 3'h0;
    end else if (_T_4227) begin
      _T_4228 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4224 <= 3'h0;
    end else if (_T_4223) begin
      _T_4224 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4220 <= 3'h0;
    end else if (_T_4219) begin
      _T_4220 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4216 <= 3'h0;
    end else if (_T_4215) begin
      _T_4216 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4212 <= 3'h0;
    end else if (_T_4211) begin
      _T_4212 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4208 <= 3'h0;
    end else if (_T_4207) begin
      _T_4208 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4204 <= 3'h0;
    end else if (_T_4203) begin
      _T_4204 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4200 <= 3'h0;
    end else if (_T_4199) begin
      _T_4200 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4196 <= 3'h0;
    end else if (_T_4195) begin
      _T_4196 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4192 <= 3'h0;
    end else if (_T_4191) begin
      _T_4192 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4188 <= 3'h0;
    end else if (_T_4187) begin
      _T_4188 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4184 <= 3'h0;
    end else if (_T_4183) begin
      _T_4184 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4180 <= 3'h0;
    end else if (_T_4179) begin
      _T_4180 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4176 <= 3'h0;
    end else if (_T_4175) begin
      _T_4176 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4172 <= 3'h0;
    end else if (_T_4171) begin
      _T_4172 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4168 <= 3'h0;
    end else if (_T_4167) begin
      _T_4168 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4164 <= 3'h0;
    end else if (_T_4163) begin
      _T_4164 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4160 <= 3'h0;
    end else if (_T_4159) begin
      _T_4160 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4156 <= 3'h0;
    end else if (_T_4155) begin
      _T_4156 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4152 <= 3'h0;
    end else if (_T_4151) begin
      _T_4152 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4148 <= 3'h0;
    end else if (_T_4147) begin
      _T_4148 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4144 <= 3'h0;
    end else if (_T_4143) begin
      _T_4144 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4140 <= 3'h0;
    end else if (_T_4139) begin
      _T_4140 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4136 <= 3'h0;
    end else if (_T_4135) begin
      _T_4136 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4132 <= 3'h0;
    end else if (_T_4131) begin
      _T_4132 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4128 <= 3'h0;
    end else if (_T_4127) begin
      _T_4128 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4124 <= 3'h0;
    end else if (_T_4123) begin
      _T_4124 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4120 <= 3'h0;
    end else if (_T_4119) begin
      _T_4120 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4116 <= 3'h0;
    end else if (_T_4115) begin
      _T_4116 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4112 <= 3'h0;
    end else if (_T_4111) begin
      _T_4112 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4108 <= 3'h0;
    end else if (_T_4107) begin
      _T_4108 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4104 <= 3'h0;
    end else if (_T_4103) begin
      _T_4104 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4100 <= 3'h0;
    end else if (_T_4099) begin
      _T_4100 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4096 <= 3'h0;
    end else if (_T_4095) begin
      _T_4096 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4092 <= 3'h0;
    end else if (_T_4091) begin
      _T_4092 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4088 <= 3'h0;
    end else if (_T_4087) begin
      _T_4088 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4084 <= 3'h0;
    end else if (_T_4083) begin
      _T_4084 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4080 <= 3'h0;
    end else if (_T_4079) begin
      _T_4080 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4076 <= 3'h0;
    end else if (_T_4075) begin
      _T_4076 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4072 <= 3'h0;
    end else if (_T_4071) begin
      _T_4072 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4068 <= 3'h0;
    end else if (_T_4067) begin
      _T_4068 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4064 <= 3'h0;
    end else if (_T_4063) begin
      _T_4064 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4060 <= 3'h0;
    end else if (_T_4059) begin
      _T_4060 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4056 <= 3'h0;
    end else if (_T_4055) begin
      _T_4056 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4052 <= 3'h0;
    end else if (_T_4051) begin
      _T_4052 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4048 <= 3'h0;
    end else if (_T_4047) begin
      _T_4048 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4044 <= 3'h0;
    end else if (_T_4043) begin
      _T_4044 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4040 <= 3'h0;
    end else if (_T_4039) begin
      _T_4040 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4036 <= 3'h0;
    end else if (_T_4035) begin
      _T_4036 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4032 <= 3'h0;
    end else if (_T_4031) begin
      _T_4032 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4028 <= 3'h0;
    end else if (_T_4027) begin
      _T_4028 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4024 <= 3'h0;
    end else if (_T_4023) begin
      _T_4024 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4020 <= 3'h0;
    end else if (_T_4019) begin
      _T_4020 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4016 <= 3'h0;
    end else if (_T_4015) begin
      _T_4016 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4012 <= 3'h0;
    end else if (_T_4011) begin
      _T_4012 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4008 <= 3'h0;
    end else if (_T_4007) begin
      _T_4008 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4004 <= 3'h0;
    end else if (_T_4003) begin
      _T_4004 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4000 <= 3'h0;
    end else if (_T_3999) begin
      _T_4000 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3996 <= 3'h0;
    end else if (_T_3995) begin
      _T_3996 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3992 <= 3'h0;
    end else if (_T_3991) begin
      _T_3992 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3988 <= 3'h0;
    end else if (_T_3987) begin
      _T_3988 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3984 <= 3'h0;
    end else if (_T_3983) begin
      _T_3984 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3980 <= 3'h0;
    end else if (_T_3979) begin
      _T_3980 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3976 <= 3'h0;
    end else if (_T_3975) begin
      _T_3976 <= way_status_new_ff;
    end
    if (reset) begin
      uncacheable_miss_scnd_ff <= 1'h0;
    end else if (!(sel_hold_imb_scnd)) begin
      uncacheable_miss_scnd_ff <= io_ifc_fetch_uncacheable_bf;
    end
    if (reset) begin
      imb_scnd_ff <= 31'h0;
    end else if (!(sel_hold_imb_scnd)) begin
      imb_scnd_ff <= io_ifc_fetch_addr_bf;
    end
    if (reset) begin
      ifu_bus_rid_ff <= 3'h0;
    end else if (io_ifu_bus_clk_en) begin
      ifu_bus_rid_ff <= io_ifu_axi_rid;
    end
    if (reset) begin
      ifu_bus_rresp_ff <= 2'h0;
    end else if (io_ifu_bus_clk_en) begin
      ifu_bus_rresp_ff <= io_ifu_axi_rresp;
    end
    if (reset) begin
      way_status_mb_ff <= 1'h0;
    end else if (_T_278) begin
      way_status_mb_ff <= way_status_mb_scnd_ff;
    end else if (_T_280) begin
      way_status_mb_ff <= replace_way_mb_any_0;
    end else if (!(miss_pending)) begin
      way_status_mb_ff <= way_status;
    end
    if (reset) begin
      tagv_mb_ff <= 2'h0;
    end else if (scnd_miss_req) begin
      tagv_mb_ff <= _T_289;
    end else if (!(miss_pending)) begin
      tagv_mb_ff <= 2'h0;
    end
    reset_ic_ff <= _T_298 & _T_299;
    if (reset) begin
      fetch_uncacheable_ff <= 1'h0;
    end else begin
      fetch_uncacheable_ff <= io_ifc_fetch_uncacheable_bf;
    end
    if (reset) begin
      miss_addr <= 26'h0;
    end else if (_T_231) begin
      miss_addr <= imb_ff[30:5];
    end else if (scnd_miss_req_q) begin
      miss_addr <= imb_scnd_ff[30:5];
    end
    if (reset) begin
      ifc_region_acc_fault_f <= 1'h0;
    end else begin
      ifc_region_acc_fault_f <= io_ifc_region_acc_fault_bf;
    end
    if (reset) begin
      bus_rd_addr_count <= 3'h0;
    end else if (_T_2577) begin
      if (_T_231) begin
        bus_rd_addr_count <= imb_ff[4:2];
      end else if (scnd_miss_req_q) begin
        bus_rd_addr_count <= imb_scnd_ff[4:2];
      end else if (bus_cmd_sent) begin
        bus_rd_addr_count <= _T_2573;
      end
    end
    if (reset) begin
      ifu_bus_rdata_ff <= 64'h0;
    end else if (io_ifu_bus_clk_en) begin
      ifu_bus_rdata_ff <= io_ifu_axi_rdata;
    end
    if (reset) begin
      ic_miss_buff_data_0 <= 32'h0;
    end else if (write_fill_data_0) begin
      ic_miss_buff_data_0 <= io_ifu_axi_rdata[31:0];
    end
    if (reset) begin
      ic_miss_buff_data_1 <= 32'h0;
    end else if (write_fill_data_0) begin
      ic_miss_buff_data_1 <= io_ifu_axi_rdata[63:32];
    end
    if (reset) begin
      ic_miss_buff_data_2 <= 32'h0;
    end else if (write_fill_data_1) begin
      ic_miss_buff_data_2 <= io_ifu_axi_rdata[31:0];
    end
    if (reset) begin
      ic_miss_buff_data_3 <= 32'h0;
    end else if (write_fill_data_1) begin
      ic_miss_buff_data_3 <= io_ifu_axi_rdata[63:32];
    end
    if (reset) begin
      ic_miss_buff_data_4 <= 32'h0;
    end else if (write_fill_data_2) begin
      ic_miss_buff_data_4 <= io_ifu_axi_rdata[31:0];
    end
    if (reset) begin
      ic_miss_buff_data_5 <= 32'h0;
    end else if (write_fill_data_2) begin
      ic_miss_buff_data_5 <= io_ifu_axi_rdata[63:32];
    end
    if (reset) begin
      ic_miss_buff_data_6 <= 32'h0;
    end else if (write_fill_data_3) begin
      ic_miss_buff_data_6 <= io_ifu_axi_rdata[31:0];
    end
    if (reset) begin
      ic_miss_buff_data_7 <= 32'h0;
    end else if (write_fill_data_3) begin
      ic_miss_buff_data_7 <= io_ifu_axi_rdata[63:32];
    end
    if (reset) begin
      ic_miss_buff_data_8 <= 32'h0;
    end else if (write_fill_data_4) begin
      ic_miss_buff_data_8 <= io_ifu_axi_rdata[31:0];
    end
    if (reset) begin
      ic_miss_buff_data_9 <= 32'h0;
    end else if (write_fill_data_4) begin
      ic_miss_buff_data_9 <= io_ifu_axi_rdata[63:32];
    end
    if (reset) begin
      ic_miss_buff_data_10 <= 32'h0;
    end else if (write_fill_data_5) begin
      ic_miss_buff_data_10 <= io_ifu_axi_rdata[31:0];
    end
    if (reset) begin
      ic_miss_buff_data_11 <= 32'h0;
    end else if (write_fill_data_5) begin
      ic_miss_buff_data_11 <= io_ifu_axi_rdata[63:32];
    end
    if (reset) begin
      ic_miss_buff_data_12 <= 32'h0;
    end else if (write_fill_data_6) begin
      ic_miss_buff_data_12 <= io_ifu_axi_rdata[31:0];
    end
    if (reset) begin
      ic_miss_buff_data_13 <= 32'h0;
    end else if (write_fill_data_6) begin
      ic_miss_buff_data_13 <= io_ifu_axi_rdata[63:32];
    end
    if (reset) begin
      ic_miss_buff_data_14 <= 32'h0;
    end else if (write_fill_data_7) begin
      ic_miss_buff_data_14 <= io_ifu_axi_rdata[31:0];
    end
    if (reset) begin
      ic_miss_buff_data_15 <= 32'h0;
    end else if (write_fill_data_7) begin
      ic_miss_buff_data_15 <= io_ifu_axi_rdata[63:32];
    end
    if (reset) begin
      ic_debug_ict_array_sel_ff <= 1'h0;
    end else if (debug_c1_clken) begin
      ic_debug_ict_array_sel_ff <= ic_debug_ict_array_sel_in;
    end
    if (reset) begin
      ic_tag_valid_out_1_0 <= 1'h0;
    end else if (_T_5736) begin
      ic_tag_valid_out_1_0 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_1 <= 1'h0;
    end else if (_T_5752) begin
      ic_tag_valid_out_1_1 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_2 <= 1'h0;
    end else if (_T_5768) begin
      ic_tag_valid_out_1_2 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_3 <= 1'h0;
    end else if (_T_5784) begin
      ic_tag_valid_out_1_3 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_4 <= 1'h0;
    end else if (_T_5800) begin
      ic_tag_valid_out_1_4 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_5 <= 1'h0;
    end else if (_T_5816) begin
      ic_tag_valid_out_1_5 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_6 <= 1'h0;
    end else if (_T_5832) begin
      ic_tag_valid_out_1_6 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_7 <= 1'h0;
    end else if (_T_5848) begin
      ic_tag_valid_out_1_7 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_8 <= 1'h0;
    end else if (_T_5864) begin
      ic_tag_valid_out_1_8 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_9 <= 1'h0;
    end else if (_T_5880) begin
      ic_tag_valid_out_1_9 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_10 <= 1'h0;
    end else if (_T_5896) begin
      ic_tag_valid_out_1_10 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_11 <= 1'h0;
    end else if (_T_5912) begin
      ic_tag_valid_out_1_11 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_12 <= 1'h0;
    end else if (_T_5928) begin
      ic_tag_valid_out_1_12 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_13 <= 1'h0;
    end else if (_T_5944) begin
      ic_tag_valid_out_1_13 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_14 <= 1'h0;
    end else if (_T_5960) begin
      ic_tag_valid_out_1_14 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_15 <= 1'h0;
    end else if (_T_5976) begin
      ic_tag_valid_out_1_15 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_16 <= 1'h0;
    end else if (_T_5992) begin
      ic_tag_valid_out_1_16 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_17 <= 1'h0;
    end else if (_T_6008) begin
      ic_tag_valid_out_1_17 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_18 <= 1'h0;
    end else if (_T_6024) begin
      ic_tag_valid_out_1_18 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_19 <= 1'h0;
    end else if (_T_6040) begin
      ic_tag_valid_out_1_19 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_20 <= 1'h0;
    end else if (_T_6056) begin
      ic_tag_valid_out_1_20 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_21 <= 1'h0;
    end else if (_T_6072) begin
      ic_tag_valid_out_1_21 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_22 <= 1'h0;
    end else if (_T_6088) begin
      ic_tag_valid_out_1_22 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_23 <= 1'h0;
    end else if (_T_6104) begin
      ic_tag_valid_out_1_23 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_24 <= 1'h0;
    end else if (_T_6120) begin
      ic_tag_valid_out_1_24 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_25 <= 1'h0;
    end else if (_T_6136) begin
      ic_tag_valid_out_1_25 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_26 <= 1'h0;
    end else if (_T_6152) begin
      ic_tag_valid_out_1_26 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_27 <= 1'h0;
    end else if (_T_6168) begin
      ic_tag_valid_out_1_27 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_28 <= 1'h0;
    end else if (_T_6184) begin
      ic_tag_valid_out_1_28 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_29 <= 1'h0;
    end else if (_T_6200) begin
      ic_tag_valid_out_1_29 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_30 <= 1'h0;
    end else if (_T_6216) begin
      ic_tag_valid_out_1_30 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_31 <= 1'h0;
    end else if (_T_6232) begin
      ic_tag_valid_out_1_31 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_32 <= 1'h0;
    end else if (_T_6760) begin
      ic_tag_valid_out_1_32 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_33 <= 1'h0;
    end else if (_T_6776) begin
      ic_tag_valid_out_1_33 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_34 <= 1'h0;
    end else if (_T_6792) begin
      ic_tag_valid_out_1_34 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_35 <= 1'h0;
    end else if (_T_6808) begin
      ic_tag_valid_out_1_35 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_36 <= 1'h0;
    end else if (_T_6824) begin
      ic_tag_valid_out_1_36 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_37 <= 1'h0;
    end else if (_T_6840) begin
      ic_tag_valid_out_1_37 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_38 <= 1'h0;
    end else if (_T_6856) begin
      ic_tag_valid_out_1_38 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_39 <= 1'h0;
    end else if (_T_6872) begin
      ic_tag_valid_out_1_39 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_40 <= 1'h0;
    end else if (_T_6888) begin
      ic_tag_valid_out_1_40 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_41 <= 1'h0;
    end else if (_T_6904) begin
      ic_tag_valid_out_1_41 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_42 <= 1'h0;
    end else if (_T_6920) begin
      ic_tag_valid_out_1_42 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_43 <= 1'h0;
    end else if (_T_6936) begin
      ic_tag_valid_out_1_43 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_44 <= 1'h0;
    end else if (_T_6952) begin
      ic_tag_valid_out_1_44 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_45 <= 1'h0;
    end else if (_T_6968) begin
      ic_tag_valid_out_1_45 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_46 <= 1'h0;
    end else if (_T_6984) begin
      ic_tag_valid_out_1_46 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_47 <= 1'h0;
    end else if (_T_7000) begin
      ic_tag_valid_out_1_47 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_48 <= 1'h0;
    end else if (_T_7016) begin
      ic_tag_valid_out_1_48 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_49 <= 1'h0;
    end else if (_T_7032) begin
      ic_tag_valid_out_1_49 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_50 <= 1'h0;
    end else if (_T_7048) begin
      ic_tag_valid_out_1_50 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_51 <= 1'h0;
    end else if (_T_7064) begin
      ic_tag_valid_out_1_51 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_52 <= 1'h0;
    end else if (_T_7080) begin
      ic_tag_valid_out_1_52 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_53 <= 1'h0;
    end else if (_T_7096) begin
      ic_tag_valid_out_1_53 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_54 <= 1'h0;
    end else if (_T_7112) begin
      ic_tag_valid_out_1_54 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_55 <= 1'h0;
    end else if (_T_7128) begin
      ic_tag_valid_out_1_55 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_56 <= 1'h0;
    end else if (_T_7144) begin
      ic_tag_valid_out_1_56 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_57 <= 1'h0;
    end else if (_T_7160) begin
      ic_tag_valid_out_1_57 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_58 <= 1'h0;
    end else if (_T_7176) begin
      ic_tag_valid_out_1_58 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_59 <= 1'h0;
    end else if (_T_7192) begin
      ic_tag_valid_out_1_59 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_60 <= 1'h0;
    end else if (_T_7208) begin
      ic_tag_valid_out_1_60 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_61 <= 1'h0;
    end else if (_T_7224) begin
      ic_tag_valid_out_1_61 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_62 <= 1'h0;
    end else if (_T_7240) begin
      ic_tag_valid_out_1_62 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_63 <= 1'h0;
    end else if (_T_7256) begin
      ic_tag_valid_out_1_63 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_64 <= 1'h0;
    end else if (_T_7784) begin
      ic_tag_valid_out_1_64 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_65 <= 1'h0;
    end else if (_T_7800) begin
      ic_tag_valid_out_1_65 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_66 <= 1'h0;
    end else if (_T_7816) begin
      ic_tag_valid_out_1_66 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_67 <= 1'h0;
    end else if (_T_7832) begin
      ic_tag_valid_out_1_67 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_68 <= 1'h0;
    end else if (_T_7848) begin
      ic_tag_valid_out_1_68 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_69 <= 1'h0;
    end else if (_T_7864) begin
      ic_tag_valid_out_1_69 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_70 <= 1'h0;
    end else if (_T_7880) begin
      ic_tag_valid_out_1_70 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_71 <= 1'h0;
    end else if (_T_7896) begin
      ic_tag_valid_out_1_71 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_72 <= 1'h0;
    end else if (_T_7912) begin
      ic_tag_valid_out_1_72 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_73 <= 1'h0;
    end else if (_T_7928) begin
      ic_tag_valid_out_1_73 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_74 <= 1'h0;
    end else if (_T_7944) begin
      ic_tag_valid_out_1_74 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_75 <= 1'h0;
    end else if (_T_7960) begin
      ic_tag_valid_out_1_75 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_76 <= 1'h0;
    end else if (_T_7976) begin
      ic_tag_valid_out_1_76 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_77 <= 1'h0;
    end else if (_T_7992) begin
      ic_tag_valid_out_1_77 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_78 <= 1'h0;
    end else if (_T_8008) begin
      ic_tag_valid_out_1_78 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_79 <= 1'h0;
    end else if (_T_8024) begin
      ic_tag_valid_out_1_79 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_80 <= 1'h0;
    end else if (_T_8040) begin
      ic_tag_valid_out_1_80 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_81 <= 1'h0;
    end else if (_T_8056) begin
      ic_tag_valid_out_1_81 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_82 <= 1'h0;
    end else if (_T_8072) begin
      ic_tag_valid_out_1_82 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_83 <= 1'h0;
    end else if (_T_8088) begin
      ic_tag_valid_out_1_83 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_84 <= 1'h0;
    end else if (_T_8104) begin
      ic_tag_valid_out_1_84 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_85 <= 1'h0;
    end else if (_T_8120) begin
      ic_tag_valid_out_1_85 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_86 <= 1'h0;
    end else if (_T_8136) begin
      ic_tag_valid_out_1_86 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_87 <= 1'h0;
    end else if (_T_8152) begin
      ic_tag_valid_out_1_87 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_88 <= 1'h0;
    end else if (_T_8168) begin
      ic_tag_valid_out_1_88 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_89 <= 1'h0;
    end else if (_T_8184) begin
      ic_tag_valid_out_1_89 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_90 <= 1'h0;
    end else if (_T_8200) begin
      ic_tag_valid_out_1_90 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_91 <= 1'h0;
    end else if (_T_8216) begin
      ic_tag_valid_out_1_91 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_92 <= 1'h0;
    end else if (_T_8232) begin
      ic_tag_valid_out_1_92 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_93 <= 1'h0;
    end else if (_T_8248) begin
      ic_tag_valid_out_1_93 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_94 <= 1'h0;
    end else if (_T_8264) begin
      ic_tag_valid_out_1_94 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_95 <= 1'h0;
    end else if (_T_8280) begin
      ic_tag_valid_out_1_95 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_96 <= 1'h0;
    end else if (_T_8808) begin
      ic_tag_valid_out_1_96 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_97 <= 1'h0;
    end else if (_T_8824) begin
      ic_tag_valid_out_1_97 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_98 <= 1'h0;
    end else if (_T_8840) begin
      ic_tag_valid_out_1_98 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_99 <= 1'h0;
    end else if (_T_8856) begin
      ic_tag_valid_out_1_99 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_100 <= 1'h0;
    end else if (_T_8872) begin
      ic_tag_valid_out_1_100 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_101 <= 1'h0;
    end else if (_T_8888) begin
      ic_tag_valid_out_1_101 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_102 <= 1'h0;
    end else if (_T_8904) begin
      ic_tag_valid_out_1_102 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_103 <= 1'h0;
    end else if (_T_8920) begin
      ic_tag_valid_out_1_103 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_104 <= 1'h0;
    end else if (_T_8936) begin
      ic_tag_valid_out_1_104 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_105 <= 1'h0;
    end else if (_T_8952) begin
      ic_tag_valid_out_1_105 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_106 <= 1'h0;
    end else if (_T_8968) begin
      ic_tag_valid_out_1_106 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_107 <= 1'h0;
    end else if (_T_8984) begin
      ic_tag_valid_out_1_107 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_108 <= 1'h0;
    end else if (_T_9000) begin
      ic_tag_valid_out_1_108 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_109 <= 1'h0;
    end else if (_T_9016) begin
      ic_tag_valid_out_1_109 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_110 <= 1'h0;
    end else if (_T_9032) begin
      ic_tag_valid_out_1_110 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_111 <= 1'h0;
    end else if (_T_9048) begin
      ic_tag_valid_out_1_111 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_112 <= 1'h0;
    end else if (_T_9064) begin
      ic_tag_valid_out_1_112 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_113 <= 1'h0;
    end else if (_T_9080) begin
      ic_tag_valid_out_1_113 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_114 <= 1'h0;
    end else if (_T_9096) begin
      ic_tag_valid_out_1_114 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_115 <= 1'h0;
    end else if (_T_9112) begin
      ic_tag_valid_out_1_115 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_116 <= 1'h0;
    end else if (_T_9128) begin
      ic_tag_valid_out_1_116 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_117 <= 1'h0;
    end else if (_T_9144) begin
      ic_tag_valid_out_1_117 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_118 <= 1'h0;
    end else if (_T_9160) begin
      ic_tag_valid_out_1_118 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_119 <= 1'h0;
    end else if (_T_9176) begin
      ic_tag_valid_out_1_119 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_120 <= 1'h0;
    end else if (_T_9192) begin
      ic_tag_valid_out_1_120 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_121 <= 1'h0;
    end else if (_T_9208) begin
      ic_tag_valid_out_1_121 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_122 <= 1'h0;
    end else if (_T_9224) begin
      ic_tag_valid_out_1_122 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_123 <= 1'h0;
    end else if (_T_9240) begin
      ic_tag_valid_out_1_123 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_124 <= 1'h0;
    end else if (_T_9256) begin
      ic_tag_valid_out_1_124 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_125 <= 1'h0;
    end else if (_T_9272) begin
      ic_tag_valid_out_1_125 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_126 <= 1'h0;
    end else if (_T_9288) begin
      ic_tag_valid_out_1_126 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_1_127 <= 1'h0;
    end else if (_T_9304) begin
      ic_tag_valid_out_1_127 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_0 <= 1'h0;
    end else if (_T_5224) begin
      ic_tag_valid_out_0_0 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_1 <= 1'h0;
    end else if (_T_5240) begin
      ic_tag_valid_out_0_1 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_2 <= 1'h0;
    end else if (_T_5256) begin
      ic_tag_valid_out_0_2 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_3 <= 1'h0;
    end else if (_T_5272) begin
      ic_tag_valid_out_0_3 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_4 <= 1'h0;
    end else if (_T_5288) begin
      ic_tag_valid_out_0_4 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_5 <= 1'h0;
    end else if (_T_5304) begin
      ic_tag_valid_out_0_5 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_6 <= 1'h0;
    end else if (_T_5320) begin
      ic_tag_valid_out_0_6 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_7 <= 1'h0;
    end else if (_T_5336) begin
      ic_tag_valid_out_0_7 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_8 <= 1'h0;
    end else if (_T_5352) begin
      ic_tag_valid_out_0_8 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_9 <= 1'h0;
    end else if (_T_5368) begin
      ic_tag_valid_out_0_9 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_10 <= 1'h0;
    end else if (_T_5384) begin
      ic_tag_valid_out_0_10 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_11 <= 1'h0;
    end else if (_T_5400) begin
      ic_tag_valid_out_0_11 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_12 <= 1'h0;
    end else if (_T_5416) begin
      ic_tag_valid_out_0_12 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_13 <= 1'h0;
    end else if (_T_5432) begin
      ic_tag_valid_out_0_13 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_14 <= 1'h0;
    end else if (_T_5448) begin
      ic_tag_valid_out_0_14 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_15 <= 1'h0;
    end else if (_T_5464) begin
      ic_tag_valid_out_0_15 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_16 <= 1'h0;
    end else if (_T_5480) begin
      ic_tag_valid_out_0_16 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_17 <= 1'h0;
    end else if (_T_5496) begin
      ic_tag_valid_out_0_17 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_18 <= 1'h0;
    end else if (_T_5512) begin
      ic_tag_valid_out_0_18 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_19 <= 1'h0;
    end else if (_T_5528) begin
      ic_tag_valid_out_0_19 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_20 <= 1'h0;
    end else if (_T_5544) begin
      ic_tag_valid_out_0_20 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_21 <= 1'h0;
    end else if (_T_5560) begin
      ic_tag_valid_out_0_21 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_22 <= 1'h0;
    end else if (_T_5576) begin
      ic_tag_valid_out_0_22 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_23 <= 1'h0;
    end else if (_T_5592) begin
      ic_tag_valid_out_0_23 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_24 <= 1'h0;
    end else if (_T_5608) begin
      ic_tag_valid_out_0_24 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_25 <= 1'h0;
    end else if (_T_5624) begin
      ic_tag_valid_out_0_25 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_26 <= 1'h0;
    end else if (_T_5640) begin
      ic_tag_valid_out_0_26 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_27 <= 1'h0;
    end else if (_T_5656) begin
      ic_tag_valid_out_0_27 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_28 <= 1'h0;
    end else if (_T_5672) begin
      ic_tag_valid_out_0_28 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_29 <= 1'h0;
    end else if (_T_5688) begin
      ic_tag_valid_out_0_29 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_30 <= 1'h0;
    end else if (_T_5704) begin
      ic_tag_valid_out_0_30 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_31 <= 1'h0;
    end else if (_T_5720) begin
      ic_tag_valid_out_0_31 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_32 <= 1'h0;
    end else if (_T_6248) begin
      ic_tag_valid_out_0_32 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_33 <= 1'h0;
    end else if (_T_6264) begin
      ic_tag_valid_out_0_33 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_34 <= 1'h0;
    end else if (_T_6280) begin
      ic_tag_valid_out_0_34 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_35 <= 1'h0;
    end else if (_T_6296) begin
      ic_tag_valid_out_0_35 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_36 <= 1'h0;
    end else if (_T_6312) begin
      ic_tag_valid_out_0_36 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_37 <= 1'h0;
    end else if (_T_6328) begin
      ic_tag_valid_out_0_37 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_38 <= 1'h0;
    end else if (_T_6344) begin
      ic_tag_valid_out_0_38 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_39 <= 1'h0;
    end else if (_T_6360) begin
      ic_tag_valid_out_0_39 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_40 <= 1'h0;
    end else if (_T_6376) begin
      ic_tag_valid_out_0_40 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_41 <= 1'h0;
    end else if (_T_6392) begin
      ic_tag_valid_out_0_41 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_42 <= 1'h0;
    end else if (_T_6408) begin
      ic_tag_valid_out_0_42 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_43 <= 1'h0;
    end else if (_T_6424) begin
      ic_tag_valid_out_0_43 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_44 <= 1'h0;
    end else if (_T_6440) begin
      ic_tag_valid_out_0_44 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_45 <= 1'h0;
    end else if (_T_6456) begin
      ic_tag_valid_out_0_45 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_46 <= 1'h0;
    end else if (_T_6472) begin
      ic_tag_valid_out_0_46 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_47 <= 1'h0;
    end else if (_T_6488) begin
      ic_tag_valid_out_0_47 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_48 <= 1'h0;
    end else if (_T_6504) begin
      ic_tag_valid_out_0_48 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_49 <= 1'h0;
    end else if (_T_6520) begin
      ic_tag_valid_out_0_49 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_50 <= 1'h0;
    end else if (_T_6536) begin
      ic_tag_valid_out_0_50 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_51 <= 1'h0;
    end else if (_T_6552) begin
      ic_tag_valid_out_0_51 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_52 <= 1'h0;
    end else if (_T_6568) begin
      ic_tag_valid_out_0_52 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_53 <= 1'h0;
    end else if (_T_6584) begin
      ic_tag_valid_out_0_53 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_54 <= 1'h0;
    end else if (_T_6600) begin
      ic_tag_valid_out_0_54 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_55 <= 1'h0;
    end else if (_T_6616) begin
      ic_tag_valid_out_0_55 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_56 <= 1'h0;
    end else if (_T_6632) begin
      ic_tag_valid_out_0_56 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_57 <= 1'h0;
    end else if (_T_6648) begin
      ic_tag_valid_out_0_57 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_58 <= 1'h0;
    end else if (_T_6664) begin
      ic_tag_valid_out_0_58 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_59 <= 1'h0;
    end else if (_T_6680) begin
      ic_tag_valid_out_0_59 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_60 <= 1'h0;
    end else if (_T_6696) begin
      ic_tag_valid_out_0_60 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_61 <= 1'h0;
    end else if (_T_6712) begin
      ic_tag_valid_out_0_61 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_62 <= 1'h0;
    end else if (_T_6728) begin
      ic_tag_valid_out_0_62 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_63 <= 1'h0;
    end else if (_T_6744) begin
      ic_tag_valid_out_0_63 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_64 <= 1'h0;
    end else if (_T_7272) begin
      ic_tag_valid_out_0_64 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_65 <= 1'h0;
    end else if (_T_7288) begin
      ic_tag_valid_out_0_65 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_66 <= 1'h0;
    end else if (_T_7304) begin
      ic_tag_valid_out_0_66 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_67 <= 1'h0;
    end else if (_T_7320) begin
      ic_tag_valid_out_0_67 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_68 <= 1'h0;
    end else if (_T_7336) begin
      ic_tag_valid_out_0_68 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_69 <= 1'h0;
    end else if (_T_7352) begin
      ic_tag_valid_out_0_69 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_70 <= 1'h0;
    end else if (_T_7368) begin
      ic_tag_valid_out_0_70 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_71 <= 1'h0;
    end else if (_T_7384) begin
      ic_tag_valid_out_0_71 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_72 <= 1'h0;
    end else if (_T_7400) begin
      ic_tag_valid_out_0_72 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_73 <= 1'h0;
    end else if (_T_7416) begin
      ic_tag_valid_out_0_73 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_74 <= 1'h0;
    end else if (_T_7432) begin
      ic_tag_valid_out_0_74 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_75 <= 1'h0;
    end else if (_T_7448) begin
      ic_tag_valid_out_0_75 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_76 <= 1'h0;
    end else if (_T_7464) begin
      ic_tag_valid_out_0_76 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_77 <= 1'h0;
    end else if (_T_7480) begin
      ic_tag_valid_out_0_77 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_78 <= 1'h0;
    end else if (_T_7496) begin
      ic_tag_valid_out_0_78 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_79 <= 1'h0;
    end else if (_T_7512) begin
      ic_tag_valid_out_0_79 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_80 <= 1'h0;
    end else if (_T_7528) begin
      ic_tag_valid_out_0_80 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_81 <= 1'h0;
    end else if (_T_7544) begin
      ic_tag_valid_out_0_81 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_82 <= 1'h0;
    end else if (_T_7560) begin
      ic_tag_valid_out_0_82 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_83 <= 1'h0;
    end else if (_T_7576) begin
      ic_tag_valid_out_0_83 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_84 <= 1'h0;
    end else if (_T_7592) begin
      ic_tag_valid_out_0_84 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_85 <= 1'h0;
    end else if (_T_7608) begin
      ic_tag_valid_out_0_85 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_86 <= 1'h0;
    end else if (_T_7624) begin
      ic_tag_valid_out_0_86 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_87 <= 1'h0;
    end else if (_T_7640) begin
      ic_tag_valid_out_0_87 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_88 <= 1'h0;
    end else if (_T_7656) begin
      ic_tag_valid_out_0_88 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_89 <= 1'h0;
    end else if (_T_7672) begin
      ic_tag_valid_out_0_89 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_90 <= 1'h0;
    end else if (_T_7688) begin
      ic_tag_valid_out_0_90 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_91 <= 1'h0;
    end else if (_T_7704) begin
      ic_tag_valid_out_0_91 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_92 <= 1'h0;
    end else if (_T_7720) begin
      ic_tag_valid_out_0_92 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_93 <= 1'h0;
    end else if (_T_7736) begin
      ic_tag_valid_out_0_93 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_94 <= 1'h0;
    end else if (_T_7752) begin
      ic_tag_valid_out_0_94 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_95 <= 1'h0;
    end else if (_T_7768) begin
      ic_tag_valid_out_0_95 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_96 <= 1'h0;
    end else if (_T_8296) begin
      ic_tag_valid_out_0_96 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_97 <= 1'h0;
    end else if (_T_8312) begin
      ic_tag_valid_out_0_97 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_98 <= 1'h0;
    end else if (_T_8328) begin
      ic_tag_valid_out_0_98 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_99 <= 1'h0;
    end else if (_T_8344) begin
      ic_tag_valid_out_0_99 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_100 <= 1'h0;
    end else if (_T_8360) begin
      ic_tag_valid_out_0_100 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_101 <= 1'h0;
    end else if (_T_8376) begin
      ic_tag_valid_out_0_101 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_102 <= 1'h0;
    end else if (_T_8392) begin
      ic_tag_valid_out_0_102 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_103 <= 1'h0;
    end else if (_T_8408) begin
      ic_tag_valid_out_0_103 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_104 <= 1'h0;
    end else if (_T_8424) begin
      ic_tag_valid_out_0_104 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_105 <= 1'h0;
    end else if (_T_8440) begin
      ic_tag_valid_out_0_105 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_106 <= 1'h0;
    end else if (_T_8456) begin
      ic_tag_valid_out_0_106 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_107 <= 1'h0;
    end else if (_T_8472) begin
      ic_tag_valid_out_0_107 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_108 <= 1'h0;
    end else if (_T_8488) begin
      ic_tag_valid_out_0_108 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_109 <= 1'h0;
    end else if (_T_8504) begin
      ic_tag_valid_out_0_109 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_110 <= 1'h0;
    end else if (_T_8520) begin
      ic_tag_valid_out_0_110 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_111 <= 1'h0;
    end else if (_T_8536) begin
      ic_tag_valid_out_0_111 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_112 <= 1'h0;
    end else if (_T_8552) begin
      ic_tag_valid_out_0_112 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_113 <= 1'h0;
    end else if (_T_8568) begin
      ic_tag_valid_out_0_113 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_114 <= 1'h0;
    end else if (_T_8584) begin
      ic_tag_valid_out_0_114 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_115 <= 1'h0;
    end else if (_T_8600) begin
      ic_tag_valid_out_0_115 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_116 <= 1'h0;
    end else if (_T_8616) begin
      ic_tag_valid_out_0_116 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_117 <= 1'h0;
    end else if (_T_8632) begin
      ic_tag_valid_out_0_117 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_118 <= 1'h0;
    end else if (_T_8648) begin
      ic_tag_valid_out_0_118 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_119 <= 1'h0;
    end else if (_T_8664) begin
      ic_tag_valid_out_0_119 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_120 <= 1'h0;
    end else if (_T_8680) begin
      ic_tag_valid_out_0_120 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_121 <= 1'h0;
    end else if (_T_8696) begin
      ic_tag_valid_out_0_121 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_122 <= 1'h0;
    end else if (_T_8712) begin
      ic_tag_valid_out_0_122 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_123 <= 1'h0;
    end else if (_T_8728) begin
      ic_tag_valid_out_0_123 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_124 <= 1'h0;
    end else if (_T_8744) begin
      ic_tag_valid_out_0_124 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_125 <= 1'h0;
    end else if (_T_8760) begin
      ic_tag_valid_out_0_125 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_126 <= 1'h0;
    end else if (_T_8776) begin
      ic_tag_valid_out_0_126 <= _T_5215;
    end
    if (reset) begin
      ic_tag_valid_out_0_127 <= 1'h0;
    end else if (_T_8792) begin
      ic_tag_valid_out_0_127 <= _T_5215;
    end
    if (reset) begin
      ic_debug_way_ff <= 2'h0;
    end else if (debug_c1_clken) begin
      ic_debug_way_ff <= io_ic_debug_way;
    end
    if (reset) begin
      _T_1209 <= 71'h0;
    end else if (ic_debug_ict_array_sel_ff) begin
      _T_1209 <= {{5'd0}, _T_1208};
    end else begin
      _T_1209 <= io_ic_debug_rd_data;
    end
    if (reset) begin
      ifu_bus_cmd_valid <= 1'h0;
    end else if (_T_2526) begin
      ifu_bus_cmd_valid <= ifc_bus_ic_req_ff_in;
    end
    if (reset) begin
      bus_cmd_beat_count <= 3'h0;
    end else if (_T_2601) begin
      bus_cmd_beat_count <= bus_new_cmd_beat_count;
    end
    if (reset) begin
      ifu_bus_arready_unq_ff <= 1'h0;
    end else if (io_ifu_bus_clk_en) begin
      ifu_bus_arready_unq_ff <= io_ifu_axi_arready;
    end
    if (reset) begin
      ifu_bus_arvalid_ff <= 1'h0;
    end else if (io_ifu_bus_clk_en) begin
      ifu_bus_arvalid_ff <= io_ifu_axi_arvalid;
    end
  end
  always @(posedge io_free_clk) begin
    if (reset) begin
      scnd_miss_req_q <= 1'h0;
    end else begin
      scnd_miss_req_q <= scnd_miss_req_in;
    end
    if (reset) begin
      iccm_dma_rvalid_in <= 1'h0;
    end else begin
      iccm_dma_rvalid_in <= _T_2645;
    end
    if (reset) begin
      dma_iccm_req_f <= 1'h0;
    end else begin
      dma_iccm_req_f <= io_dma_iccm_req;
    end
    if (reset) begin
      perr_state <= 3'h0;
    end else if (perr_state_en) begin
      if (_T_2427) begin
        if (io_iccm_dma_sb_error) begin
          perr_state <= 3'h4;
        end else if (_T_2429) begin
          perr_state <= 3'h1;
        end else begin
          perr_state <= 3'h2;
        end
      end else if (_T_2439) begin
        perr_state <= 3'h0;
      end else if (_T_2442) begin
        if (_T_2444) begin
          perr_state <= 3'h0;
        end else begin
          perr_state <= 3'h3;
        end
      end else if (_T_2448) begin
        if (io_dec_tlu_force_halt) begin
          perr_state <= 3'h0;
        end else begin
          perr_state <= 3'h3;
        end
      end else begin
        perr_state <= 3'h0;
      end
    end
    if (reset) begin
      err_stop_state <= 2'h0;
    end else if (err_stop_state_en) begin
      if (_T_2452) begin
        err_stop_state <= 2'h1;
      end else if (_T_2457) begin
        if (_T_2459) begin
          err_stop_state <= 2'h0;
        end else if (_T_2480) begin
          err_stop_state <= 2'h3;
        end else if (io_ifu_fetch_val[0]) begin
          err_stop_state <= 2'h2;
        end else begin
          err_stop_state <= 2'h1;
        end
      end else if (_T_2484) begin
        if (_T_2459) begin
          err_stop_state <= 2'h0;
        end else if (io_ifu_fetch_val[0]) begin
          err_stop_state <= 2'h3;
        end else begin
          err_stop_state <= 2'h2;
        end
      end else if (_T_2501) begin
        if (_T_2505) begin
          err_stop_state <= 2'h0;
        end else if (io_dec_tlu_flush_err_wb) begin
          err_stop_state <= 2'h1;
        end else begin
          err_stop_state <= 2'h3;
        end
      end else begin
        err_stop_state <= 2'h0;
      end
    end
    if (reset) begin
      bus_ifu_bus_clk_en_ff <= 1'h0;
    end else begin
      bus_ifu_bus_clk_en_ff <= io_ifu_bus_clk_en;
    end
    if (reset) begin
      bus_data_beat_count <= 3'h0;
    end else begin
      bus_data_beat_count <= bus_new_data_beat_count;
    end
    if (reset) begin
      ic_miss_buff_data_valid <= 8'h0;
    end else begin
      ic_miss_buff_data_valid <= _T_1370;
    end
    if (reset) begin
      last_data_recieved_ff <= 1'h0;
    end else begin
      last_data_recieved_ff <= last_data_recieved_in;
    end
    if (reset) begin
      sel_mb_addr_ff <= 1'h0;
    end else begin
      sel_mb_addr_ff <= sel_mb_addr;
    end
    if (reset) begin
      _T_5128 <= 7'h0;
    end else if (_T_3949) begin
      _T_5128 <= io_ic_debug_addr[9:3];
    end else begin
      _T_5128 <= ifu_ic_rw_int_addr[11:5];
    end
    if (reset) begin
      ifu_wr_data_comb_err_ff <= 1'h0;
    end else begin
      ifu_wr_data_comb_err_ff <= ifu_wr_cumulative_err;
    end
    if (reset) begin
      ic_act_miss_f_delayed <= 1'h0;
    end else begin
      ic_act_miss_f_delayed <= ic_act_miss_f;
    end
    if (reset) begin
      ic_crit_wd_rdy_new_ff <= 1'h0;
    end else begin
      ic_crit_wd_rdy_new_ff <= ic_crit_wd_rdy_new_in;
    end
    if (reset) begin
      ic_miss_buff_data_error <= 8'h0;
    end else begin
      ic_miss_buff_data_error <= _T_1410;
    end
    if (reset) begin
      ic_debug_rd_en_ff <= 1'h0;
    end else begin
      ic_debug_rd_en_ff <= io_ic_debug_rd_en;
    end
    if (reset) begin
      ifc_dma_access_ok_prev <= 1'h0;
    end else begin
      ifc_dma_access_ok_prev <= ifc_dma_access_ok_d;
    end
    if (reset) begin
      iccm_ecc_corr_data_ff <= 39'h0;
    end else if (iccm_ecc_write_status) begin
      iccm_ecc_corr_data_ff <= _T_3884;
    end
    if (reset) begin
      dma_mem_addr_ff <= 2'h0;
    end else begin
      dma_mem_addr_ff <= io_dma_mem_addr[3:2];
    end
    if (reset) begin
      dma_mem_tag_ff <= 3'h0;
    end else begin
      dma_mem_tag_ff <= io_dma_mem_tag;
    end
    if (reset) begin
      iccm_dma_rtag <= 3'h0;
    end else begin
      iccm_dma_rtag <= dma_mem_tag_ff;
    end
    if (reset) begin
      iccm_dma_rvalid <= 1'h0;
    end else begin
      iccm_dma_rvalid <= iccm_dma_rvalid_in;
    end
    if (reset) begin
      iccm_dma_rdata <= 64'h0;
    end else if (iccm_dma_ecc_error_in) begin
      iccm_dma_rdata <= _T_3059;
    end else begin
      iccm_dma_rdata <= _T_3060;
    end
    if (reset) begin
      iccm_ecc_corr_index_ff <= 14'h0;
    end else if (iccm_ecc_write_status) begin
      if (iccm_single_ecc_error[0]) begin
        iccm_ecc_corr_index_ff <= iccm_rw_addr_f;
      end else begin
        iccm_ecc_corr_index_ff <= _T_3880;
      end
    end
    if (reset) begin
      iccm_rd_ecc_single_err_ff <= 1'h0;
    end else begin
      iccm_rd_ecc_single_err_ff <= iccm_rd_ecc_single_err_hold_in;
    end
    if (reset) begin
      iccm_rw_addr_f <= 14'h0;
    end else begin
      iccm_rw_addr_f <= io_iccm_rw_addr[14:1];
    end
    if (reset) begin
      ifu_status_wr_addr_ff <= 7'h0;
    end else if (_T_3949) begin
      ifu_status_wr_addr_ff <= io_ic_debug_addr[9:3];
    end else begin
      ifu_status_wr_addr_ff <= ifu_status_wr_addr[11:5];
    end
    if (reset) begin
      way_status_wr_en_ff <= 1'h0;
    end else begin
      way_status_wr_en_ff <= way_status_wr_en_w_debug;
    end
    if (reset) begin
      way_status_new_ff <= 3'h0;
    end else if (_T_3952) begin
      way_status_new_ff <= _T_3956;
    end else begin
      way_status_new_ff <= {{2'd0}, way_status_new};
    end
    if (reset) begin
      ifu_tag_wren_ff <= 2'h0;
    end else begin
      ifu_tag_wren_ff <= ifu_tag_wren_w_debug;
    end
    if (reset) begin
      ic_valid_ff <= 1'h0;
    end else if (_T_3952) begin
      ic_valid_ff <= io_ic_debug_wr_data[0];
    end else begin
      ic_valid_ff <= ic_valid;
    end
    if (reset) begin
      _T_10145 <= 1'h0;
    end else if (ic_debug_rd_en_ff) begin
      _T_10145 <= ic_debug_rd_en_ff;
    end
  end
  always @(posedge io_active_clk) begin
    if (reset) begin
      reset_all_tags <= 1'h0;
    end else begin
      reset_all_tags <= io_dec_tlu_fence_i_wb;
    end
    if (reset) begin
      perr_ic_index_ff <= 6'h0;
    end else if (perr_sb_write_status) begin
      perr_ic_index_ff <= ifu_ic_rw_int_addr_ff;
    end
    if (reset) begin
      dma_sb_err_state_ff <= 1'h0;
    end else begin
      dma_sb_err_state_ff <= _T_7;
    end
    if (reset) begin
      _T_10115 <= 1'h0;
    end else begin
      _T_10115 <= ic_act_miss_f;
    end
    if (reset) begin
      _T_10116 <= 1'h0;
    end else begin
      _T_10116 <= ic_act_hit_f;
    end
    if (reset) begin
      _T_10117 <= 1'h0;
    end else begin
      _T_10117 <= ifc_bus_acc_fault_f;
    end
    if (reset) begin
      _T_10121 <= 1'h0;
    end else begin
      _T_10121 <= _T_10120;
    end
    if (reset) begin
      _T_10122 <= 1'h0;
    end else begin
      _T_10122 <= bus_cmd_sent;
    end
  end
endmodule
