module el2_ifu_compress_ctl(
  input         clock,
  input         reset,
  input  [15:0] io_din,
  output [31:0] io_dout
);
  wire  _T_1 = io_din[1:0] != 2'h3; // @[el2_ifu_compress_ctl.scala 401:27]
  wire [31:0] _T_3 = {16'h0,io_din}; // @[Cat.scala 29:58]
  wire  _T_5 = |_T_3[12:5]; // @[el2_ifu_compress_ctl.scala 257:29]
  wire [6:0] _T_6 = _T_5 ? 7'h13 : 7'h1f; // @[el2_ifu_compress_ctl.scala 257:20]
  wire [29:0] _T_20 = {_T_3[10:7],_T_3[12:11],_T_3[5],_T_3[6],2'h0,5'h2,3'h0,2'h1,_T_3[4:2],_T_6}; // @[Cat.scala 29:58]
  wire [7:0] _T_30 = {_T_3[6:5],_T_3[12:10],3'h0}; // @[Cat.scala 29:58]
  wire [27:0] _T_38 = {_T_3[6:5],_T_3[12:10],3'h0,2'h1,_T_3[9:7],3'h3,2'h1,_T_3[4:2],7'h7}; // @[Cat.scala 29:58]
  wire [6:0] _T_52 = {_T_3[5],_T_3[12:10],_T_3[6],2'h0}; // @[Cat.scala 29:58]
  wire [26:0] _T_60 = {_T_3[5],_T_3[12:10],_T_3[6],2'h0,2'h1,_T_3[9:7],3'h2,2'h1,_T_3[4:2],7'h3}; // @[Cat.scala 29:58]
  wire [26:0] _T_82 = {_T_3[5],_T_3[12:10],_T_3[6],2'h0,2'h1,_T_3[9:7],3'h2,2'h1,_T_3[4:2],7'h7}; // @[Cat.scala 29:58]
  wire [26:0] _T_113 = {_T_52[6:5],2'h1,_T_3[4:2],2'h1,_T_3[9:7],3'h2,_T_52[4:0],7'h3f}; // @[Cat.scala 29:58]
  wire [27:0] _T_140 = {_T_30[7:5],2'h1,_T_3[4:2],2'h1,_T_3[9:7],3'h3,_T_30[4:0],7'h27}; // @[Cat.scala 29:58]
  wire [26:0] _T_171 = {_T_52[6:5],2'h1,_T_3[4:2],2'h1,_T_3[9:7],3'h2,_T_52[4:0],7'h23}; // @[Cat.scala 29:58]
  wire [26:0] _T_202 = {_T_52[6:5],2'h1,_T_3[4:2],2'h1,_T_3[9:7],3'h2,_T_52[4:0],7'h27}; // @[Cat.scala 29:58]
  wire [6:0] _T_213 = _T_3[12] ? 7'h7f : 7'h0; // @[Bitwise.scala 72:12]
  wire [11:0] _T_215 = {_T_213,_T_3[6:2]}; // @[Cat.scala 29:58]
  wire [31:0] _T_221 = {_T_213,_T_3[6:2],_T_3[11:7],3'h0,_T_3[11:7],7'h13}; // @[Cat.scala 29:58]
  wire [9:0] _T_230 = _T_3[12] ? 10'h3ff : 10'h0; // @[Bitwise.scala 72:12]
  wire [20:0] _T_245 = {_T_230,_T_3[8],_T_3[10:9],_T_3[6],_T_3[7],_T_3[2],_T_3[11],_T_3[5:3],1'h0}; // @[Cat.scala 29:58]
  wire [31:0] _T_308 = {_T_245[20],_T_245[10:1],_T_245[11],_T_245[19:12],5'h1,7'h6f}; // @[Cat.scala 29:58]
  wire [31:0] _T_323 = {_T_213,_T_3[6:2],5'h0,3'h0,_T_3[11:7],7'h13}; // @[Cat.scala 29:58]
  wire  _T_334 = |_T_215; // @[el2_ifu_compress_ctl.scala 294:29]
  wire [6:0] _T_335 = _T_334 ? 7'h37 : 7'h3f; // @[el2_ifu_compress_ctl.scala 294:20]
  wire [14:0] _T_338 = _T_3[12] ? 15'h7fff : 15'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_341 = {_T_338,_T_3[6:2],12'h0}; // @[Cat.scala 29:58]
  wire [31:0] _T_345 = {_T_341[31:12],_T_3[11:7],_T_335}; // @[Cat.scala 29:58]
  wire  _T_353 = _T_3[11:7] == 5'h0; // @[el2_ifu_compress_ctl.scala 296:14]
  wire  _T_355 = _T_3[11:7] == 5'h2; // @[el2_ifu_compress_ctl.scala 296:27]
  wire  _T_356 = _T_353 | _T_355; // @[el2_ifu_compress_ctl.scala 296:21]
  wire [6:0] _T_363 = _T_334 ? 7'h13 : 7'h1f; // @[el2_ifu_compress_ctl.scala 290:20]
  wire [2:0] _T_366 = _T_3[12] ? 3'h7 : 3'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_381 = {_T_366,_T_3[4:3],_T_3[5],_T_3[2],_T_3[6],4'h0,_T_3[11:7],3'h0,_T_3[11:7],_T_363}; // @[Cat.scala 29:58]
  wire [31:0] _T_388_bits = _T_356 ? _T_381 : _T_345; // @[el2_ifu_compress_ctl.scala 296:10]
  wire [25:0] _T_399 = {_T_3[12],_T_3[6:2],2'h1,_T_3[9:7],3'h5,2'h1,_T_3[9:7],7'h13}; // @[Cat.scala 29:58]
  wire [30:0] _GEN_172 = {{5'd0}, _T_399}; // @[el2_ifu_compress_ctl.scala 303:23]
  wire [30:0] _T_411 = _GEN_172 | 31'h40000000; // @[el2_ifu_compress_ctl.scala 303:23]
  wire [31:0] _T_424 = {_T_213,_T_3[6:2],2'h1,_T_3[9:7],3'h7,2'h1,_T_3[9:7],7'h13}; // @[Cat.scala 29:58]
  wire [2:0] _T_428 = {_T_3[12],_T_3[6:5]}; // @[Cat.scala 29:58]
  wire  _T_430 = _T_3[6:5] == 2'h0; // @[el2_ifu_compress_ctl.scala 307:30]
  wire [30:0] _T_431 = _T_430 ? 31'h40000000 : 31'h0; // @[el2_ifu_compress_ctl.scala 307:22]
  wire [6:0] _T_433 = _T_3[12] ? 7'h3b : 7'h33; // @[el2_ifu_compress_ctl.scala 308:22]
  wire [2:0] _GEN_1 = 3'h1 == _T_428 ? 3'h4 : 3'h0; // @[Cat.scala 29:58]
  wire [2:0] _GEN_2 = 3'h2 == _T_428 ? 3'h6 : _GEN_1; // @[Cat.scala 29:58]
  wire [2:0] _GEN_3 = 3'h3 == _T_428 ? 3'h7 : _GEN_2; // @[Cat.scala 29:58]
  wire [2:0] _GEN_4 = 3'h4 == _T_428 ? 3'h0 : _GEN_3; // @[Cat.scala 29:58]
  wire [2:0] _GEN_5 = 3'h5 == _T_428 ? 3'h0 : _GEN_4; // @[Cat.scala 29:58]
  wire [2:0] _GEN_6 = 3'h6 == _T_428 ? 3'h2 : _GEN_5; // @[Cat.scala 29:58]
  wire [2:0] _GEN_7 = 3'h7 == _T_428 ? 3'h3 : _GEN_6; // @[Cat.scala 29:58]
  wire [24:0] _T_443 = {2'h1,_T_3[4:2],2'h1,_T_3[9:7],_GEN_7,2'h1,_T_3[9:7],_T_433}; // @[Cat.scala 29:58]
  wire [30:0] _GEN_173 = {{6'd0}, _T_443}; // @[el2_ifu_compress_ctl.scala 309:43]
  wire [30:0] _T_444 = _GEN_173 | _T_431; // @[el2_ifu_compress_ctl.scala 309:43]
  wire [31:0] _T_445_0 = {{6'd0}, _T_399}; // @[el2_ifu_compress_ctl.scala 311:19 el2_ifu_compress_ctl.scala 311:19]
  wire [31:0] _T_445_1 = {{1'd0}, _T_411}; // @[el2_ifu_compress_ctl.scala 311:19 el2_ifu_compress_ctl.scala 311:19]
  wire [31:0] _GEN_9 = 2'h1 == _T_3[11:10] ? _T_445_1 : _T_445_0; // @[el2_ifu_compress_ctl.scala 226:14]
  wire [31:0] _GEN_10 = 2'h2 == _T_3[11:10] ? _T_424 : _GEN_9; // @[el2_ifu_compress_ctl.scala 226:14]
  wire [31:0] _T_445_3 = {{1'd0}, _T_444}; // @[el2_ifu_compress_ctl.scala 311:19 el2_ifu_compress_ctl.scala 311:19]
  wire [31:0] _GEN_11 = 2'h3 == _T_3[11:10] ? _T_445_3 : _GEN_10; // @[el2_ifu_compress_ctl.scala 226:14]
  wire [31:0] _T_535 = {_T_245[20],_T_245[10:1],_T_245[11],_T_245[19:12],5'h0,7'h6f}; // @[Cat.scala 29:58]
  wire [4:0] _T_544 = _T_3[12] ? 5'h1f : 5'h0; // @[Bitwise.scala 72:12]
  wire [12:0] _T_553 = {_T_544,_T_3[6:5],_T_3[2],_T_3[11:10],_T_3[4:3],1'h0}; // @[Cat.scala 29:58]
  wire [31:0] _T_602 = {_T_553[12],_T_553[10:5],5'h0,2'h1,_T_3[9:7],3'h0,_T_553[4:1],_T_553[11],7'h63}; // @[Cat.scala 29:58]
  wire [31:0] _T_669 = {_T_553[12],_T_553[10:5],5'h0,2'h1,_T_3[9:7],3'h1,_T_553[4:1],_T_553[11],7'h63}; // @[Cat.scala 29:58]
  wire  _T_675 = |_T_3[11:7]; // @[el2_ifu_compress_ctl.scala 317:27]
  wire [6:0] _T_676 = _T_675 ? 7'h3 : 7'h1f; // @[el2_ifu_compress_ctl.scala 317:23]
  wire [25:0] _T_685 = {_T_3[12],_T_3[6:2],_T_3[11:7],3'h1,_T_3[11:7],7'h13}; // @[Cat.scala 29:58]
  wire [28:0] _T_701 = {_T_3[4:2],_T_3[12],_T_3[6:5],3'h0,5'h2,3'h3,_T_3[11:7],7'h7}; // @[Cat.scala 29:58]
  wire [27:0] _T_716 = {_T_3[3:2],_T_3[12],_T_3[6:4],2'h0,5'h2,3'h2,_T_3[11:7],_T_676}; // @[Cat.scala 29:58]
  wire [27:0] _T_731 = {_T_3[3:2],_T_3[12],_T_3[6:4],2'h0,5'h2,3'h2,_T_3[11:7],7'h7}; // @[Cat.scala 29:58]
  wire [24:0] _T_741 = {_T_3[6:2],5'h0,3'h0,_T_3[11:7],7'h33}; // @[Cat.scala 29:58]
  wire [24:0] _T_752 = {_T_3[6:2],_T_3[11:7],3'h0,_T_3[11:7],7'h33}; // @[Cat.scala 29:58]
  wire [24:0] _T_763 = {_T_3[6:2],_T_3[11:7],3'h0,12'h67}; // @[Cat.scala 29:58]
  wire [24:0] _T_765 = {_T_763[24:7],7'h1f}; // @[Cat.scala 29:58]
  wire [24:0] _T_768 = _T_675 ? _T_763 : _T_765; // @[el2_ifu_compress_ctl.scala 338:33]
  wire  _T_774 = |_T_3[6:2]; // @[el2_ifu_compress_ctl.scala 339:27]
  wire [31:0] _T_745_bits = {{7'd0}, _T_741}; // @[el2_ifu_compress_ctl.scala 225:19 el2_ifu_compress_ctl.scala 226:14]
  wire [31:0] _T_772_bits = {{7'd0}, _T_768}; // @[el2_ifu_compress_ctl.scala 225:19 el2_ifu_compress_ctl.scala 226:14]
  wire [31:0] _T_775_bits = _T_774 ? _T_745_bits : _T_772_bits; // @[el2_ifu_compress_ctl.scala 339:22]
  wire [24:0] _T_781 = {_T_3[6:2],_T_3[11:7],3'h0,12'he7}; // @[Cat.scala 29:58]
  wire [24:0] _T_783 = {_T_763[24:7],7'h73}; // @[Cat.scala 29:58]
  wire [24:0] _T_784 = _T_783 | 25'h100000; // @[el2_ifu_compress_ctl.scala 341:46]
  wire [24:0] _T_787 = _T_675 ? _T_781 : _T_784; // @[el2_ifu_compress_ctl.scala 342:33]
  wire [31:0] _T_757_bits = {{7'd0}, _T_752}; // @[el2_ifu_compress_ctl.scala 225:19 el2_ifu_compress_ctl.scala 226:14]
  wire [31:0] _T_791_bits = {{7'd0}, _T_787}; // @[el2_ifu_compress_ctl.scala 225:19 el2_ifu_compress_ctl.scala 226:14]
  wire [31:0] _T_794_bits = _T_774 ? _T_757_bits : _T_791_bits; // @[el2_ifu_compress_ctl.scala 343:25]
  wire [31:0] _T_796_bits = _T_3[12] ? _T_794_bits : _T_775_bits; // @[el2_ifu_compress_ctl.scala 344:10]
  wire [8:0] _T_800 = {_T_3[9:7],_T_3[12:10],3'h0}; // @[Cat.scala 29:58]
  wire [28:0] _T_812 = {_T_800[8:5],_T_3[6:2],5'h2,3'h3,_T_800[4:0],7'h27}; // @[Cat.scala 29:58]
  wire [7:0] _T_820 = {_T_3[8:7],_T_3[12:9],2'h0}; // @[Cat.scala 29:58]
  wire [27:0] _T_832 = {_T_820[7:5],_T_3[6:2],5'h2,3'h2,_T_820[4:0],7'h23}; // @[Cat.scala 29:58]
  wire [27:0] _T_852 = {_T_820[7:5],_T_3[6:2],5'h2,3'h2,_T_820[4:0],7'h27}; // @[Cat.scala 29:58]
  wire [4:0] _T_900 = {_T_3[1:0],_T_3[15:13]}; // @[Cat.scala 29:58]
  wire [31:0] _T_26_bits = {{2'd0}, _T_20}; // @[el2_ifu_compress_ctl.scala 225:19 el2_ifu_compress_ctl.scala 226:14]
  wire [31:0] _T_46_bits = {{4'd0}, _T_38}; // @[el2_ifu_compress_ctl.scala 225:19 el2_ifu_compress_ctl.scala 226:14]
  wire [31:0] _GEN_17 = 5'h1 == _T_900 ? _T_46_bits : _T_26_bits; // @[el2_ifu_compress_ctl.scala 404:19]
  wire [31:0] _T_68_bits = {{5'd0}, _T_60}; // @[el2_ifu_compress_ctl.scala 225:19 el2_ifu_compress_ctl.scala 226:14]
  wire [31:0] _GEN_22 = 5'h2 == _T_900 ? _T_68_bits : _GEN_17; // @[el2_ifu_compress_ctl.scala 404:19]
  wire [31:0] _T_90_bits = {{5'd0}, _T_82}; // @[el2_ifu_compress_ctl.scala 225:19 el2_ifu_compress_ctl.scala 226:14]
  wire [31:0] _GEN_27 = 5'h3 == _T_900 ? _T_90_bits : _GEN_22; // @[el2_ifu_compress_ctl.scala 404:19]
  wire [31:0] _T_121_bits = {{5'd0}, _T_113}; // @[el2_ifu_compress_ctl.scala 225:19 el2_ifu_compress_ctl.scala 226:14]
  wire [31:0] _GEN_32 = 5'h4 == _T_900 ? _T_121_bits : _GEN_27; // @[el2_ifu_compress_ctl.scala 404:19]
  wire [31:0] _T_148_bits = {{4'd0}, _T_140}; // @[el2_ifu_compress_ctl.scala 225:19 el2_ifu_compress_ctl.scala 226:14]
  wire [31:0] _GEN_37 = 5'h5 == _T_900 ? _T_148_bits : _GEN_32; // @[el2_ifu_compress_ctl.scala 404:19]
  wire [31:0] _T_179_bits = {{5'd0}, _T_171}; // @[el2_ifu_compress_ctl.scala 225:19 el2_ifu_compress_ctl.scala 226:14]
  wire [31:0] _GEN_42 = 5'h6 == _T_900 ? _T_179_bits : _GEN_37; // @[el2_ifu_compress_ctl.scala 404:19]
  wire [31:0] _T_210_bits = {{5'd0}, _T_202}; // @[el2_ifu_compress_ctl.scala 225:19 el2_ifu_compress_ctl.scala 226:14]
  wire [31:0] _GEN_47 = 5'h7 == _T_900 ? _T_210_bits : _GEN_42; // @[el2_ifu_compress_ctl.scala 404:19]
  wire [31:0] _GEN_52 = 5'h8 == _T_900 ? _T_221 : _GEN_47; // @[el2_ifu_compress_ctl.scala 404:19]
  wire [31:0] _GEN_57 = 5'h9 == _T_900 ? _T_308 : _GEN_52; // @[el2_ifu_compress_ctl.scala 404:19]
  wire [31:0] _GEN_62 = 5'ha == _T_900 ? _T_323 : _GEN_57; // @[el2_ifu_compress_ctl.scala 404:19]
  wire [31:0] _GEN_67 = 5'hb == _T_900 ? _T_388_bits : _GEN_62; // @[el2_ifu_compress_ctl.scala 404:19]
  wire [31:0] _GEN_72 = 5'hc == _T_900 ? _GEN_11 : _GEN_67; // @[el2_ifu_compress_ctl.scala 404:19]
  wire [31:0] _GEN_77 = 5'hd == _T_900 ? _T_535 : _GEN_72; // @[el2_ifu_compress_ctl.scala 404:19]
  wire [31:0] _GEN_82 = 5'he == _T_900 ? _T_602 : _GEN_77; // @[el2_ifu_compress_ctl.scala 404:19]
  wire [31:0] _GEN_87 = 5'hf == _T_900 ? _T_669 : _GEN_82; // @[el2_ifu_compress_ctl.scala 404:19]
  wire [31:0] _T_690_bits = {{6'd0}, _T_685}; // @[el2_ifu_compress_ctl.scala 225:19 el2_ifu_compress_ctl.scala 226:14]
  wire [31:0] _GEN_92 = 5'h10 == _T_900 ? _T_690_bits : _GEN_87; // @[el2_ifu_compress_ctl.scala 404:19]
  wire [31:0] _T_705_bits = {{3'd0}, _T_701}; // @[el2_ifu_compress_ctl.scala 225:19 el2_ifu_compress_ctl.scala 226:14]
  wire [31:0] _GEN_97 = 5'h11 == _T_900 ? _T_705_bits : _GEN_92; // @[el2_ifu_compress_ctl.scala 404:19]
  wire [31:0] _T_720_bits = {{4'd0}, _T_716}; // @[el2_ifu_compress_ctl.scala 225:19 el2_ifu_compress_ctl.scala 226:14]
  wire [31:0] _GEN_102 = 5'h12 == _T_900 ? _T_720_bits : _GEN_97; // @[el2_ifu_compress_ctl.scala 404:19]
  wire [31:0] _T_735_bits = {{4'd0}, _T_731}; // @[el2_ifu_compress_ctl.scala 225:19 el2_ifu_compress_ctl.scala 226:14]
  wire [31:0] _GEN_107 = 5'h13 == _T_900 ? _T_735_bits : _GEN_102; // @[el2_ifu_compress_ctl.scala 404:19]
  wire [31:0] _GEN_112 = 5'h14 == _T_900 ? _T_796_bits : _GEN_107; // @[el2_ifu_compress_ctl.scala 404:19]
  wire [31:0] _T_816_bits = {{3'd0}, _T_812}; // @[el2_ifu_compress_ctl.scala 225:19 el2_ifu_compress_ctl.scala 226:14]
  wire [31:0] _GEN_117 = 5'h15 == _T_900 ? _T_816_bits : _GEN_112; // @[el2_ifu_compress_ctl.scala 404:19]
  wire [31:0] _T_836_bits = {{4'd0}, _T_832}; // @[el2_ifu_compress_ctl.scala 225:19 el2_ifu_compress_ctl.scala 226:14]
  wire [31:0] _GEN_122 = 5'h16 == _T_900 ? _T_836_bits : _GEN_117; // @[el2_ifu_compress_ctl.scala 404:19]
  wire [31:0] _T_856_bits = {{4'd0}, _T_852}; // @[el2_ifu_compress_ctl.scala 225:19 el2_ifu_compress_ctl.scala 226:14]
  wire [31:0] _GEN_127 = 5'h17 == _T_900 ? _T_856_bits : _GEN_122; // @[el2_ifu_compress_ctl.scala 404:19]
  wire [31:0] _GEN_132 = 5'h18 == _T_900 ? _T_3 : _GEN_127; // @[el2_ifu_compress_ctl.scala 404:19]
  wire [31:0] _GEN_137 = 5'h19 == _T_900 ? _T_3 : _GEN_132; // @[el2_ifu_compress_ctl.scala 404:19]
  wire [31:0] _GEN_142 = 5'h1a == _T_900 ? _T_3 : _GEN_137; // @[el2_ifu_compress_ctl.scala 404:19]
  wire [31:0] _GEN_147 = 5'h1b == _T_900 ? _T_3 : _GEN_142; // @[el2_ifu_compress_ctl.scala 404:19]
  wire [31:0] _GEN_152 = 5'h1c == _T_900 ? _T_3 : _GEN_147; // @[el2_ifu_compress_ctl.scala 404:19]
  wire [31:0] _GEN_157 = 5'h1d == _T_900 ? _T_3 : _GEN_152; // @[el2_ifu_compress_ctl.scala 404:19]
  wire [31:0] _GEN_162 = 5'h1e == _T_900 ? _T_3 : _GEN_157; // @[el2_ifu_compress_ctl.scala 404:19]
  wire [31:0] _GEN_167 = 5'h1f == _T_900 ? _T_3 : _GEN_162; // @[el2_ifu_compress_ctl.scala 404:19]
  assign io_dout = _T_1 ? 32'h0 : _GEN_167; // @[el2_ifu_compress_ctl.scala 404:13]
endmodule
