// NOTE NOTE NOTE NOTE NOTE NOTE NOTE NOTE NOTE NOTE NOTE NOTE NOTE NOTE NOTE NOTE
// This is an automatically generated file by waleedbinehsan on و 17:46:00 PKT ت 29 دسمبر 2020
//
// cmd:    quasar -target=default 
//

`include "common_defines.vh"
`undef ASSERT_ON
`undef TEC_RV_ICG
`define TEC_RV_ICG HDBLVT16_CKGTPLT_V5_12
`define PHYSICAL 1
