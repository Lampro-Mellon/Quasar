module rvclkhdr(
  output  io_l1clk,
  input   io_clk,
  input   io_en,
  input   io_scan_mode
);
  wire  clkhdr_Q; // @[el2_lib.scala 452:26]
  wire  clkhdr_CK; // @[el2_lib.scala 452:26]
  wire  clkhdr_EN; // @[el2_lib.scala 452:26]
  wire  clkhdr_SE; // @[el2_lib.scala 452:26]
  TEC_RV_ICG clkhdr ( // @[el2_lib.scala 452:26]
    .Q(clkhdr_Q),
    .CK(clkhdr_CK),
    .EN(clkhdr_EN),
    .SE(clkhdr_SE)
  );
  assign io_l1clk = clkhdr_Q; // @[el2_lib.scala 453:14]
  assign clkhdr_CK = io_clk; // @[el2_lib.scala 454:18]
  assign clkhdr_EN = io_en; // @[el2_lib.scala 455:18]
  assign clkhdr_SE = io_scan_mode; // @[el2_lib.scala 456:18]
endmodule
module el2_ifu_bp_ctl(
  input          clock,
  input          reset,
  input          io_active_clk,
  input          io_ic_hit_f,
  input  [30:0]  io_ifc_fetch_addr_f,
  input          io_ifc_fetch_req_f,
  input          io_dec_tlu_br0_r_pkt_valid,
  input  [1:0]   io_dec_tlu_br0_r_pkt_hist,
  input          io_dec_tlu_br0_r_pkt_br_error,
  input          io_dec_tlu_br0_r_pkt_br_start_error,
  input          io_dec_tlu_br0_r_pkt_way,
  input          io_dec_tlu_br0_r_pkt_middle,
  input  [7:0]   io_exu_i0_br_fghr_r,
  input  [7:0]   io_exu_i0_br_index_r,
  input          io_dec_tlu_flush_lower_wb,
  input          io_dec_tlu_flush_leak_one_wb,
  input          io_dec_tlu_bpred_disable,
  input          io_exu_mp_pkt_misp,
  input          io_exu_mp_pkt_ataken,
  input          io_exu_mp_pkt_boffset,
  input          io_exu_mp_pkt_pc4,
  input  [1:0]   io_exu_mp_pkt_hist,
  input  [11:0]  io_exu_mp_pkt_toffset,
  input          io_exu_mp_pkt_valid,
  input          io_exu_mp_pkt_br_error,
  input          io_exu_mp_pkt_br_start_error,
  input  [30:0]  io_exu_mp_pkt_prett,
  input          io_exu_mp_pkt_pcall,
  input          io_exu_mp_pkt_pret,
  input          io_exu_mp_pkt_pja,
  input          io_exu_mp_pkt_way,
  input  [7:0]   io_exu_mp_eghr,
  input  [7:0]   io_exu_mp_fghr,
  input  [7:0]   io_exu_mp_index,
  input  [4:0]   io_exu_mp_btag,
  input          io_exu_flush_final,
  output         io_ifu_bp_hit_taken_f,
  output [30:0]  io_ifu_bp_btb_target_f,
  output         io_ifu_bp_inst_mask_f,
  output [7:0]   io_ifu_bp_fghr_f,
  output [1:0]   io_ifu_bp_way_f,
  output [1:0]   io_ifu_bp_ret_f,
  output [1:0]   io_ifu_bp_hist1_f,
  output [1:0]   io_ifu_bp_hist0_f,
  output [1:0]   io_ifu_bp_pc4_f,
  output [1:0]   io_ifu_bp_valid_f,
  output [11:0]  io_ifu_bp_poffset_f,
  input          io_scan_mode,
  output [255:0] io_test
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_576;
  reg [31:0] _RAND_577;
  reg [31:0] _RAND_578;
  reg [31:0] _RAND_579;
  reg [31:0] _RAND_580;
  reg [31:0] _RAND_581;
  reg [31:0] _RAND_582;
  reg [31:0] _RAND_583;
  reg [31:0] _RAND_584;
  reg [31:0] _RAND_585;
  reg [31:0] _RAND_586;
  reg [31:0] _RAND_587;
  reg [31:0] _RAND_588;
  reg [31:0] _RAND_589;
  reg [31:0] _RAND_590;
  reg [31:0] _RAND_591;
  reg [31:0] _RAND_592;
  reg [31:0] _RAND_593;
  reg [31:0] _RAND_594;
  reg [31:0] _RAND_595;
  reg [31:0] _RAND_596;
  reg [31:0] _RAND_597;
  reg [31:0] _RAND_598;
  reg [31:0] _RAND_599;
  reg [31:0] _RAND_600;
  reg [31:0] _RAND_601;
  reg [31:0] _RAND_602;
  reg [31:0] _RAND_603;
  reg [31:0] _RAND_604;
  reg [31:0] _RAND_605;
  reg [31:0] _RAND_606;
  reg [31:0] _RAND_607;
  reg [31:0] _RAND_608;
  reg [31:0] _RAND_609;
  reg [31:0] _RAND_610;
  reg [31:0] _RAND_611;
  reg [31:0] _RAND_612;
  reg [31:0] _RAND_613;
  reg [31:0] _RAND_614;
  reg [31:0] _RAND_615;
  reg [31:0] _RAND_616;
  reg [31:0] _RAND_617;
  reg [31:0] _RAND_618;
  reg [31:0] _RAND_619;
  reg [31:0] _RAND_620;
  reg [31:0] _RAND_621;
  reg [31:0] _RAND_622;
  reg [31:0] _RAND_623;
  reg [31:0] _RAND_624;
  reg [31:0] _RAND_625;
  reg [31:0] _RAND_626;
  reg [31:0] _RAND_627;
  reg [31:0] _RAND_628;
  reg [31:0] _RAND_629;
  reg [31:0] _RAND_630;
  reg [31:0] _RAND_631;
  reg [31:0] _RAND_632;
  reg [31:0] _RAND_633;
  reg [31:0] _RAND_634;
  reg [31:0] _RAND_635;
  reg [31:0] _RAND_636;
  reg [31:0] _RAND_637;
  reg [31:0] _RAND_638;
  reg [31:0] _RAND_639;
  reg [31:0] _RAND_640;
  reg [31:0] _RAND_641;
  reg [31:0] _RAND_642;
  reg [31:0] _RAND_643;
  reg [31:0] _RAND_644;
  reg [31:0] _RAND_645;
  reg [31:0] _RAND_646;
  reg [31:0] _RAND_647;
  reg [31:0] _RAND_648;
  reg [31:0] _RAND_649;
  reg [31:0] _RAND_650;
  reg [31:0] _RAND_651;
  reg [31:0] _RAND_652;
  reg [31:0] _RAND_653;
  reg [31:0] _RAND_654;
  reg [31:0] _RAND_655;
  reg [31:0] _RAND_656;
  reg [31:0] _RAND_657;
  reg [31:0] _RAND_658;
  reg [31:0] _RAND_659;
  reg [31:0] _RAND_660;
  reg [31:0] _RAND_661;
  reg [31:0] _RAND_662;
  reg [31:0] _RAND_663;
  reg [31:0] _RAND_664;
  reg [31:0] _RAND_665;
  reg [31:0] _RAND_666;
  reg [31:0] _RAND_667;
  reg [31:0] _RAND_668;
  reg [31:0] _RAND_669;
  reg [31:0] _RAND_670;
  reg [31:0] _RAND_671;
  reg [31:0] _RAND_672;
  reg [31:0] _RAND_673;
  reg [31:0] _RAND_674;
  reg [31:0] _RAND_675;
  reg [31:0] _RAND_676;
  reg [31:0] _RAND_677;
  reg [31:0] _RAND_678;
  reg [31:0] _RAND_679;
  reg [31:0] _RAND_680;
  reg [31:0] _RAND_681;
  reg [31:0] _RAND_682;
  reg [31:0] _RAND_683;
  reg [31:0] _RAND_684;
  reg [31:0] _RAND_685;
  reg [31:0] _RAND_686;
  reg [31:0] _RAND_687;
  reg [31:0] _RAND_688;
  reg [31:0] _RAND_689;
  reg [31:0] _RAND_690;
  reg [31:0] _RAND_691;
  reg [31:0] _RAND_692;
  reg [31:0] _RAND_693;
  reg [31:0] _RAND_694;
  reg [31:0] _RAND_695;
  reg [31:0] _RAND_696;
  reg [31:0] _RAND_697;
  reg [31:0] _RAND_698;
  reg [31:0] _RAND_699;
  reg [31:0] _RAND_700;
  reg [31:0] _RAND_701;
  reg [31:0] _RAND_702;
  reg [31:0] _RAND_703;
  reg [31:0] _RAND_704;
  reg [31:0] _RAND_705;
  reg [31:0] _RAND_706;
  reg [31:0] _RAND_707;
  reg [31:0] _RAND_708;
  reg [31:0] _RAND_709;
  reg [31:0] _RAND_710;
  reg [31:0] _RAND_711;
  reg [31:0] _RAND_712;
  reg [31:0] _RAND_713;
  reg [31:0] _RAND_714;
  reg [31:0] _RAND_715;
  reg [31:0] _RAND_716;
  reg [31:0] _RAND_717;
  reg [31:0] _RAND_718;
  reg [31:0] _RAND_719;
  reg [31:0] _RAND_720;
  reg [31:0] _RAND_721;
  reg [31:0] _RAND_722;
  reg [31:0] _RAND_723;
  reg [31:0] _RAND_724;
  reg [31:0] _RAND_725;
  reg [31:0] _RAND_726;
  reg [31:0] _RAND_727;
  reg [31:0] _RAND_728;
  reg [31:0] _RAND_729;
  reg [31:0] _RAND_730;
  reg [31:0] _RAND_731;
  reg [31:0] _RAND_732;
  reg [31:0] _RAND_733;
  reg [31:0] _RAND_734;
  reg [31:0] _RAND_735;
  reg [31:0] _RAND_736;
  reg [31:0] _RAND_737;
  reg [31:0] _RAND_738;
  reg [31:0] _RAND_739;
  reg [31:0] _RAND_740;
  reg [31:0] _RAND_741;
  reg [31:0] _RAND_742;
  reg [31:0] _RAND_743;
  reg [31:0] _RAND_744;
  reg [31:0] _RAND_745;
  reg [31:0] _RAND_746;
  reg [31:0] _RAND_747;
  reg [31:0] _RAND_748;
  reg [31:0] _RAND_749;
  reg [31:0] _RAND_750;
  reg [31:0] _RAND_751;
  reg [31:0] _RAND_752;
  reg [31:0] _RAND_753;
  reg [31:0] _RAND_754;
  reg [31:0] _RAND_755;
  reg [31:0] _RAND_756;
  reg [31:0] _RAND_757;
  reg [31:0] _RAND_758;
  reg [31:0] _RAND_759;
  reg [31:0] _RAND_760;
  reg [31:0] _RAND_761;
  reg [31:0] _RAND_762;
  reg [31:0] _RAND_763;
  reg [31:0] _RAND_764;
  reg [31:0] _RAND_765;
  reg [31:0] _RAND_766;
  reg [31:0] _RAND_767;
  reg [31:0] _RAND_768;
  reg [31:0] _RAND_769;
  reg [31:0] _RAND_770;
  reg [31:0] _RAND_771;
  reg [31:0] _RAND_772;
  reg [31:0] _RAND_773;
  reg [31:0] _RAND_774;
  reg [31:0] _RAND_775;
  reg [31:0] _RAND_776;
  reg [31:0] _RAND_777;
  reg [31:0] _RAND_778;
  reg [31:0] _RAND_779;
  reg [31:0] _RAND_780;
  reg [31:0] _RAND_781;
  reg [31:0] _RAND_782;
  reg [31:0] _RAND_783;
  reg [31:0] _RAND_784;
  reg [31:0] _RAND_785;
  reg [31:0] _RAND_786;
  reg [31:0] _RAND_787;
  reg [31:0] _RAND_788;
  reg [31:0] _RAND_789;
  reg [31:0] _RAND_790;
  reg [31:0] _RAND_791;
  reg [31:0] _RAND_792;
  reg [31:0] _RAND_793;
  reg [31:0] _RAND_794;
  reg [31:0] _RAND_795;
  reg [31:0] _RAND_796;
  reg [31:0] _RAND_797;
  reg [31:0] _RAND_798;
  reg [31:0] _RAND_799;
  reg [31:0] _RAND_800;
  reg [31:0] _RAND_801;
  reg [31:0] _RAND_802;
  reg [31:0] _RAND_803;
  reg [31:0] _RAND_804;
  reg [31:0] _RAND_805;
  reg [31:0] _RAND_806;
  reg [31:0] _RAND_807;
  reg [31:0] _RAND_808;
  reg [31:0] _RAND_809;
  reg [31:0] _RAND_810;
  reg [31:0] _RAND_811;
  reg [31:0] _RAND_812;
  reg [31:0] _RAND_813;
  reg [31:0] _RAND_814;
  reg [31:0] _RAND_815;
  reg [31:0] _RAND_816;
  reg [31:0] _RAND_817;
  reg [31:0] _RAND_818;
  reg [31:0] _RAND_819;
  reg [31:0] _RAND_820;
  reg [31:0] _RAND_821;
  reg [31:0] _RAND_822;
  reg [31:0] _RAND_823;
  reg [31:0] _RAND_824;
  reg [31:0] _RAND_825;
  reg [31:0] _RAND_826;
  reg [31:0] _RAND_827;
  reg [31:0] _RAND_828;
  reg [31:0] _RAND_829;
  reg [31:0] _RAND_830;
  reg [31:0] _RAND_831;
  reg [31:0] _RAND_832;
  reg [31:0] _RAND_833;
  reg [31:0] _RAND_834;
  reg [31:0] _RAND_835;
  reg [31:0] _RAND_836;
  reg [31:0] _RAND_837;
  reg [31:0] _RAND_838;
  reg [31:0] _RAND_839;
  reg [31:0] _RAND_840;
  reg [31:0] _RAND_841;
  reg [31:0] _RAND_842;
  reg [31:0] _RAND_843;
  reg [31:0] _RAND_844;
  reg [31:0] _RAND_845;
  reg [31:0] _RAND_846;
  reg [31:0] _RAND_847;
  reg [31:0] _RAND_848;
  reg [31:0] _RAND_849;
  reg [31:0] _RAND_850;
  reg [31:0] _RAND_851;
  reg [31:0] _RAND_852;
  reg [31:0] _RAND_853;
  reg [31:0] _RAND_854;
  reg [31:0] _RAND_855;
  reg [31:0] _RAND_856;
  reg [31:0] _RAND_857;
  reg [31:0] _RAND_858;
  reg [31:0] _RAND_859;
  reg [31:0] _RAND_860;
  reg [31:0] _RAND_861;
  reg [31:0] _RAND_862;
  reg [31:0] _RAND_863;
  reg [31:0] _RAND_864;
  reg [31:0] _RAND_865;
  reg [31:0] _RAND_866;
  reg [31:0] _RAND_867;
  reg [31:0] _RAND_868;
  reg [31:0] _RAND_869;
  reg [31:0] _RAND_870;
  reg [31:0] _RAND_871;
  reg [31:0] _RAND_872;
  reg [31:0] _RAND_873;
  reg [31:0] _RAND_874;
  reg [31:0] _RAND_875;
  reg [31:0] _RAND_876;
  reg [31:0] _RAND_877;
  reg [31:0] _RAND_878;
  reg [31:0] _RAND_879;
  reg [31:0] _RAND_880;
  reg [31:0] _RAND_881;
  reg [31:0] _RAND_882;
  reg [31:0] _RAND_883;
  reg [31:0] _RAND_884;
  reg [31:0] _RAND_885;
  reg [31:0] _RAND_886;
  reg [31:0] _RAND_887;
  reg [31:0] _RAND_888;
  reg [31:0] _RAND_889;
  reg [31:0] _RAND_890;
  reg [31:0] _RAND_891;
  reg [31:0] _RAND_892;
  reg [31:0] _RAND_893;
  reg [31:0] _RAND_894;
  reg [31:0] _RAND_895;
  reg [31:0] _RAND_896;
  reg [31:0] _RAND_897;
  reg [31:0] _RAND_898;
  reg [31:0] _RAND_899;
  reg [31:0] _RAND_900;
  reg [31:0] _RAND_901;
  reg [31:0] _RAND_902;
  reg [31:0] _RAND_903;
  reg [31:0] _RAND_904;
  reg [31:0] _RAND_905;
  reg [31:0] _RAND_906;
  reg [31:0] _RAND_907;
  reg [31:0] _RAND_908;
  reg [31:0] _RAND_909;
  reg [31:0] _RAND_910;
  reg [31:0] _RAND_911;
  reg [31:0] _RAND_912;
  reg [31:0] _RAND_913;
  reg [31:0] _RAND_914;
  reg [31:0] _RAND_915;
  reg [31:0] _RAND_916;
  reg [31:0] _RAND_917;
  reg [31:0] _RAND_918;
  reg [31:0] _RAND_919;
  reg [31:0] _RAND_920;
  reg [31:0] _RAND_921;
  reg [31:0] _RAND_922;
  reg [31:0] _RAND_923;
  reg [31:0] _RAND_924;
  reg [31:0] _RAND_925;
  reg [31:0] _RAND_926;
  reg [31:0] _RAND_927;
  reg [31:0] _RAND_928;
  reg [31:0] _RAND_929;
  reg [31:0] _RAND_930;
  reg [31:0] _RAND_931;
  reg [31:0] _RAND_932;
  reg [31:0] _RAND_933;
  reg [31:0] _RAND_934;
  reg [31:0] _RAND_935;
  reg [31:0] _RAND_936;
  reg [31:0] _RAND_937;
  reg [31:0] _RAND_938;
  reg [31:0] _RAND_939;
  reg [31:0] _RAND_940;
  reg [31:0] _RAND_941;
  reg [31:0] _RAND_942;
  reg [31:0] _RAND_943;
  reg [31:0] _RAND_944;
  reg [31:0] _RAND_945;
  reg [31:0] _RAND_946;
  reg [31:0] _RAND_947;
  reg [31:0] _RAND_948;
  reg [31:0] _RAND_949;
  reg [31:0] _RAND_950;
  reg [31:0] _RAND_951;
  reg [31:0] _RAND_952;
  reg [31:0] _RAND_953;
  reg [31:0] _RAND_954;
  reg [31:0] _RAND_955;
  reg [31:0] _RAND_956;
  reg [31:0] _RAND_957;
  reg [31:0] _RAND_958;
  reg [31:0] _RAND_959;
  reg [31:0] _RAND_960;
  reg [31:0] _RAND_961;
  reg [31:0] _RAND_962;
  reg [31:0] _RAND_963;
  reg [31:0] _RAND_964;
  reg [31:0] _RAND_965;
  reg [31:0] _RAND_966;
  reg [31:0] _RAND_967;
  reg [31:0] _RAND_968;
  reg [31:0] _RAND_969;
  reg [31:0] _RAND_970;
  reg [31:0] _RAND_971;
  reg [31:0] _RAND_972;
  reg [31:0] _RAND_973;
  reg [31:0] _RAND_974;
  reg [31:0] _RAND_975;
  reg [31:0] _RAND_976;
  reg [31:0] _RAND_977;
  reg [31:0] _RAND_978;
  reg [31:0] _RAND_979;
  reg [31:0] _RAND_980;
  reg [31:0] _RAND_981;
  reg [31:0] _RAND_982;
  reg [31:0] _RAND_983;
  reg [31:0] _RAND_984;
  reg [31:0] _RAND_985;
  reg [31:0] _RAND_986;
  reg [31:0] _RAND_987;
  reg [31:0] _RAND_988;
  reg [31:0] _RAND_989;
  reg [31:0] _RAND_990;
  reg [31:0] _RAND_991;
  reg [31:0] _RAND_992;
  reg [31:0] _RAND_993;
  reg [31:0] _RAND_994;
  reg [31:0] _RAND_995;
  reg [31:0] _RAND_996;
  reg [31:0] _RAND_997;
  reg [31:0] _RAND_998;
  reg [31:0] _RAND_999;
  reg [31:0] _RAND_1000;
  reg [31:0] _RAND_1001;
  reg [31:0] _RAND_1002;
  reg [31:0] _RAND_1003;
  reg [31:0] _RAND_1004;
  reg [31:0] _RAND_1005;
  reg [31:0] _RAND_1006;
  reg [31:0] _RAND_1007;
  reg [31:0] _RAND_1008;
  reg [31:0] _RAND_1009;
  reg [31:0] _RAND_1010;
  reg [31:0] _RAND_1011;
  reg [31:0] _RAND_1012;
  reg [31:0] _RAND_1013;
  reg [31:0] _RAND_1014;
  reg [31:0] _RAND_1015;
  reg [31:0] _RAND_1016;
  reg [31:0] _RAND_1017;
  reg [31:0] _RAND_1018;
  reg [31:0] _RAND_1019;
  reg [31:0] _RAND_1020;
  reg [31:0] _RAND_1021;
  reg [31:0] _RAND_1022;
  reg [31:0] _RAND_1023;
  reg [31:0] _RAND_1024;
  reg [31:0] _RAND_1025;
  reg [31:0] _RAND_1026;
  reg [31:0] _RAND_1027;
  reg [31:0] _RAND_1028;
  reg [255:0] _RAND_1029;
  reg [31:0] _RAND_1030;
  reg [31:0] _RAND_1031;
  reg [31:0] _RAND_1032;
  reg [31:0] _RAND_1033;
  reg [31:0] _RAND_1034;
  reg [31:0] _RAND_1035;
  reg [31:0] _RAND_1036;
  reg [31:0] _RAND_1037;
  reg [31:0] _RAND_1038;
`endif // RANDOMIZE_REG_INIT
  wire  rvclkhdr_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_1_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_1_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_1_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_1_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_2_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_2_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_2_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_2_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_3_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_3_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_3_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_3_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_4_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_4_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_4_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_4_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_5_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_5_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_5_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_5_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_6_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_6_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_6_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_6_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_7_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_7_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_7_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_7_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_8_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_8_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_8_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_8_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_9_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_9_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_9_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_9_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_10_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_10_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_10_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_10_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_11_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_11_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_11_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_11_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_12_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_12_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_12_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_12_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_13_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_13_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_13_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_13_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_14_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_14_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_14_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_14_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_15_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_15_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_15_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_15_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_16_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_16_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_16_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_16_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_17_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_17_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_17_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_17_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_18_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_18_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_18_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_18_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_19_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_19_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_19_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_19_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_20_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_20_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_20_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_20_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_21_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_21_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_21_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_21_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_22_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_22_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_22_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_22_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_23_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_23_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_23_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_23_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_24_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_24_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_24_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_24_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_25_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_25_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_25_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_25_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_26_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_26_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_26_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_26_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_27_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_27_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_27_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_27_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_28_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_28_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_28_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_28_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_29_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_29_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_29_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_29_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_30_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_30_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_30_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_30_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_31_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_31_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_31_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_31_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_32_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_32_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_32_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_32_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_33_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_33_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_33_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_33_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_34_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_34_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_34_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_34_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_35_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_35_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_35_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_35_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_36_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_36_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_36_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_36_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_37_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_37_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_37_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_37_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_38_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_38_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_38_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_38_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_39_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_39_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_39_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_39_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_40_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_40_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_40_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_40_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_41_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_41_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_41_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_41_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_42_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_42_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_42_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_42_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_43_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_43_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_43_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_43_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_44_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_44_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_44_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_44_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_45_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_45_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_45_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_45_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_46_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_46_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_46_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_46_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_47_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_47_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_47_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_47_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_48_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_48_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_48_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_48_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_49_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_49_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_49_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_49_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_50_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_50_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_50_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_50_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_51_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_51_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_51_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_51_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_52_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_52_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_52_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_52_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_53_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_53_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_53_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_53_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_54_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_54_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_54_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_54_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_55_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_55_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_55_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_55_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_56_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_56_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_56_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_56_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_57_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_57_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_57_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_57_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_58_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_58_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_58_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_58_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_59_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_59_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_59_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_59_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_60_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_60_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_60_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_60_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_61_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_61_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_61_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_61_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_62_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_62_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_62_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_62_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_63_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_63_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_63_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_63_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_64_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_64_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_64_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_64_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_65_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_65_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_65_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_65_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_66_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_66_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_66_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_66_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_67_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_67_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_67_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_67_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_68_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_68_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_68_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_68_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_69_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_69_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_69_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_69_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_70_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_70_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_70_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_70_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_71_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_71_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_71_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_71_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_72_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_72_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_72_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_72_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_73_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_73_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_73_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_73_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_74_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_74_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_74_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_74_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_75_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_75_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_75_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_75_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_76_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_76_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_76_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_76_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_77_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_77_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_77_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_77_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_78_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_78_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_78_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_78_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_79_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_79_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_79_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_79_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_80_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_80_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_80_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_80_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_81_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_81_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_81_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_81_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_82_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_82_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_82_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_82_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_83_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_83_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_83_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_83_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_84_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_84_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_84_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_84_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_85_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_85_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_85_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_85_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_86_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_86_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_86_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_86_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_87_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_87_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_87_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_87_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_88_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_88_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_88_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_88_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_89_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_89_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_89_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_89_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_90_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_90_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_90_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_90_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_91_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_91_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_91_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_91_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_92_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_92_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_92_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_92_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_93_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_93_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_93_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_93_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_94_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_94_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_94_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_94_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_95_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_95_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_95_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_95_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_96_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_96_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_96_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_96_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_97_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_97_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_97_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_97_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_98_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_98_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_98_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_98_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_99_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_99_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_99_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_99_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_100_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_100_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_100_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_100_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_101_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_101_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_101_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_101_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_102_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_102_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_102_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_102_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_103_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_103_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_103_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_103_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_104_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_104_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_104_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_104_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_105_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_105_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_105_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_105_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_106_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_106_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_106_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_106_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_107_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_107_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_107_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_107_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_108_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_108_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_108_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_108_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_109_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_109_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_109_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_109_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_110_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_110_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_110_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_110_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_111_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_111_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_111_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_111_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_112_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_112_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_112_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_112_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_113_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_113_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_113_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_113_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_114_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_114_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_114_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_114_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_115_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_115_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_115_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_115_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_116_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_116_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_116_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_116_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_117_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_117_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_117_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_117_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_118_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_118_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_118_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_118_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_119_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_119_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_119_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_119_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_120_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_120_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_120_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_120_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_121_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_121_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_121_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_121_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_122_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_122_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_122_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_122_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_123_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_123_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_123_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_123_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_124_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_124_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_124_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_124_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_125_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_125_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_125_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_125_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_126_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_126_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_126_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_126_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_127_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_127_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_127_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_127_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_128_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_128_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_128_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_128_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_129_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_129_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_129_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_129_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_130_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_130_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_130_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_130_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_131_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_131_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_131_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_131_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_132_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_132_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_132_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_132_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_133_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_133_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_133_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_133_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_134_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_134_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_134_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_134_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_135_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_135_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_135_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_135_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_136_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_136_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_136_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_136_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_137_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_137_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_137_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_137_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_138_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_138_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_138_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_138_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_139_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_139_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_139_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_139_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_140_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_140_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_140_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_140_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_141_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_141_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_141_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_141_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_142_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_142_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_142_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_142_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_143_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_143_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_143_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_143_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_144_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_144_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_144_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_144_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_145_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_145_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_145_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_145_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_146_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_146_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_146_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_146_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_147_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_147_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_147_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_147_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_148_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_148_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_148_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_148_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_149_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_149_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_149_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_149_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_150_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_150_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_150_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_150_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_151_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_151_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_151_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_151_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_152_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_152_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_152_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_152_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_153_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_153_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_153_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_153_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_154_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_154_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_154_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_154_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_155_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_155_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_155_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_155_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_156_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_156_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_156_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_156_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_157_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_157_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_157_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_157_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_158_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_158_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_158_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_158_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_159_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_159_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_159_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_159_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_160_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_160_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_160_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_160_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_161_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_161_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_161_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_161_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_162_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_162_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_162_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_162_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_163_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_163_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_163_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_163_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_164_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_164_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_164_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_164_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_165_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_165_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_165_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_165_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_166_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_166_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_166_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_166_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_167_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_167_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_167_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_167_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_168_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_168_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_168_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_168_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_169_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_169_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_169_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_169_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_170_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_170_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_170_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_170_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_171_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_171_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_171_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_171_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_172_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_172_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_172_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_172_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_173_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_173_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_173_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_173_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_174_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_174_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_174_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_174_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_175_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_175_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_175_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_175_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_176_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_176_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_176_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_176_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_177_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_177_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_177_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_177_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_178_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_178_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_178_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_178_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_179_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_179_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_179_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_179_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_180_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_180_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_180_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_180_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_181_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_181_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_181_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_181_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_182_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_182_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_182_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_182_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_183_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_183_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_183_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_183_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_184_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_184_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_184_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_184_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_185_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_185_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_185_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_185_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_186_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_186_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_186_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_186_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_187_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_187_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_187_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_187_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_188_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_188_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_188_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_188_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_189_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_189_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_189_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_189_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_190_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_190_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_190_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_190_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_191_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_191_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_191_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_191_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_192_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_192_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_192_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_192_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_193_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_193_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_193_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_193_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_194_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_194_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_194_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_194_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_195_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_195_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_195_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_195_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_196_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_196_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_196_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_196_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_197_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_197_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_197_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_197_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_198_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_198_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_198_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_198_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_199_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_199_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_199_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_199_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_200_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_200_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_200_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_200_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_201_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_201_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_201_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_201_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_202_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_202_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_202_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_202_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_203_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_203_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_203_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_203_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_204_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_204_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_204_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_204_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_205_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_205_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_205_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_205_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_206_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_206_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_206_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_206_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_207_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_207_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_207_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_207_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_208_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_208_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_208_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_208_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_209_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_209_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_209_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_209_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_210_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_210_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_210_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_210_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_211_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_211_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_211_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_211_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_212_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_212_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_212_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_212_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_213_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_213_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_213_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_213_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_214_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_214_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_214_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_214_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_215_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_215_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_215_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_215_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_216_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_216_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_216_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_216_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_217_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_217_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_217_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_217_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_218_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_218_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_218_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_218_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_219_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_219_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_219_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_219_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_220_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_220_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_220_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_220_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_221_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_221_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_221_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_221_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_222_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_222_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_222_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_222_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_223_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_223_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_223_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_223_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_224_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_224_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_224_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_224_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_225_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_225_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_225_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_225_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_226_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_226_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_226_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_226_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_227_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_227_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_227_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_227_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_228_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_228_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_228_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_228_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_229_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_229_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_229_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_229_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_230_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_230_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_230_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_230_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_231_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_231_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_231_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_231_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_232_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_232_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_232_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_232_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_233_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_233_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_233_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_233_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_234_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_234_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_234_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_234_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_235_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_235_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_235_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_235_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_236_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_236_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_236_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_236_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_237_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_237_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_237_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_237_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_238_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_238_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_238_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_238_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_239_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_239_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_239_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_239_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_240_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_240_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_240_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_240_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_241_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_241_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_241_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_241_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_242_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_242_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_242_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_242_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_243_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_243_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_243_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_243_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_244_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_244_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_244_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_244_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_245_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_245_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_245_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_245_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_246_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_246_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_246_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_246_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_247_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_247_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_247_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_247_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_248_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_248_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_248_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_248_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_249_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_249_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_249_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_249_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_250_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_250_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_250_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_250_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_251_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_251_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_251_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_251_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_252_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_252_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_252_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_252_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_253_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_253_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_253_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_253_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_254_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_254_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_254_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_254_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_255_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_255_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_255_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_255_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_256_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_256_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_256_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_256_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_257_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_257_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_257_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_257_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_258_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_258_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_258_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_258_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_259_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_259_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_259_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_259_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_260_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_260_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_260_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_260_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_261_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_261_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_261_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_261_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_262_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_262_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_262_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_262_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_263_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_263_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_263_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_263_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_264_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_264_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_264_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_264_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_265_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_265_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_265_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_265_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_266_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_266_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_266_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_266_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_267_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_267_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_267_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_267_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_268_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_268_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_268_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_268_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_269_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_269_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_269_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_269_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_270_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_270_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_270_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_270_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_271_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_271_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_271_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_271_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_272_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_272_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_272_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_272_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_273_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_273_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_273_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_273_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_274_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_274_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_274_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_274_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_275_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_275_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_275_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_275_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_276_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_276_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_276_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_276_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_277_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_277_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_277_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_277_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_278_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_278_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_278_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_278_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_279_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_279_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_279_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_279_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_280_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_280_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_280_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_280_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_281_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_281_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_281_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_281_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_282_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_282_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_282_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_282_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_283_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_283_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_283_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_283_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_284_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_284_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_284_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_284_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_285_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_285_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_285_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_285_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_286_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_286_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_286_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_286_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_287_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_287_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_287_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_287_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_288_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_288_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_288_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_288_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_289_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_289_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_289_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_289_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_290_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_290_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_290_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_290_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_291_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_291_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_291_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_291_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_292_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_292_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_292_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_292_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_293_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_293_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_293_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_293_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_294_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_294_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_294_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_294_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_295_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_295_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_295_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_295_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_296_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_296_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_296_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_296_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_297_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_297_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_297_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_297_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_298_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_298_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_298_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_298_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_299_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_299_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_299_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_299_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_300_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_300_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_300_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_300_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_301_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_301_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_301_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_301_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_302_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_302_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_302_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_302_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_303_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_303_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_303_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_303_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_304_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_304_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_304_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_304_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_305_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_305_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_305_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_305_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_306_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_306_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_306_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_306_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_307_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_307_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_307_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_307_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_308_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_308_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_308_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_308_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_309_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_309_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_309_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_309_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_310_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_310_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_310_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_310_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_311_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_311_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_311_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_311_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_312_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_312_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_312_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_312_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_313_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_313_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_313_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_313_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_314_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_314_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_314_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_314_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_315_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_315_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_315_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_315_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_316_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_316_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_316_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_316_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_317_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_317_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_317_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_317_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_318_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_318_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_318_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_318_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_319_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_319_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_319_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_319_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_320_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_320_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_320_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_320_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_321_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_321_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_321_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_321_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_322_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_322_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_322_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_322_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_323_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_323_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_323_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_323_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_324_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_324_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_324_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_324_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_325_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_325_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_325_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_325_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_326_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_326_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_326_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_326_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_327_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_327_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_327_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_327_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_328_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_328_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_328_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_328_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_329_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_329_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_329_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_329_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_330_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_330_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_330_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_330_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_331_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_331_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_331_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_331_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_332_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_332_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_332_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_332_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_333_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_333_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_333_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_333_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_334_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_334_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_334_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_334_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_335_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_335_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_335_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_335_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_336_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_336_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_336_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_336_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_337_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_337_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_337_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_337_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_338_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_338_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_338_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_338_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_339_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_339_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_339_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_339_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_340_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_340_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_340_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_340_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_341_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_341_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_341_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_341_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_342_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_342_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_342_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_342_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_343_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_343_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_343_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_343_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_344_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_344_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_344_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_344_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_345_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_345_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_345_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_345_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_346_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_346_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_346_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_346_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_347_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_347_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_347_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_347_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_348_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_348_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_348_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_348_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_349_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_349_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_349_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_349_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_350_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_350_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_350_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_350_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_351_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_351_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_351_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_351_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_352_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_352_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_352_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_352_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_353_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_353_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_353_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_353_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_354_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_354_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_354_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_354_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_355_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_355_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_355_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_355_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_356_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_356_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_356_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_356_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_357_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_357_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_357_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_357_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_358_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_358_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_358_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_358_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_359_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_359_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_359_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_359_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_360_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_360_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_360_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_360_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_361_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_361_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_361_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_361_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_362_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_362_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_362_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_362_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_363_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_363_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_363_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_363_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_364_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_364_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_364_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_364_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_365_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_365_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_365_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_365_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_366_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_366_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_366_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_366_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_367_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_367_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_367_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_367_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_368_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_368_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_368_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_368_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_369_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_369_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_369_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_369_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_370_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_370_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_370_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_370_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_371_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_371_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_371_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_371_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_372_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_372_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_372_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_372_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_373_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_373_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_373_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_373_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_374_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_374_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_374_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_374_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_375_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_375_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_375_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_375_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_376_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_376_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_376_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_376_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_377_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_377_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_377_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_377_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_378_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_378_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_378_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_378_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_379_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_379_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_379_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_379_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_380_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_380_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_380_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_380_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_381_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_381_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_381_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_381_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_382_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_382_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_382_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_382_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_383_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_383_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_383_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_383_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_384_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_384_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_384_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_384_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_385_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_385_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_385_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_385_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_386_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_386_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_386_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_386_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_387_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_387_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_387_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_387_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_388_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_388_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_388_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_388_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_389_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_389_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_389_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_389_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_390_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_390_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_390_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_390_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_391_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_391_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_391_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_391_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_392_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_392_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_392_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_392_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_393_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_393_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_393_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_393_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_394_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_394_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_394_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_394_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_395_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_395_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_395_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_395_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_396_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_396_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_396_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_396_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_397_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_397_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_397_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_397_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_398_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_398_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_398_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_398_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_399_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_399_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_399_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_399_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_400_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_400_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_400_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_400_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_401_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_401_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_401_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_401_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_402_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_402_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_402_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_402_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_403_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_403_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_403_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_403_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_404_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_404_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_404_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_404_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_405_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_405_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_405_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_405_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_406_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_406_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_406_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_406_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_407_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_407_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_407_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_407_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_408_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_408_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_408_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_408_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_409_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_409_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_409_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_409_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_410_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_410_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_410_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_410_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_411_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_411_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_411_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_411_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_412_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_412_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_412_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_412_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_413_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_413_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_413_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_413_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_414_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_414_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_414_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_414_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_415_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_415_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_415_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_415_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_416_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_416_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_416_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_416_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_417_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_417_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_417_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_417_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_418_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_418_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_418_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_418_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_419_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_419_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_419_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_419_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_420_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_420_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_420_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_420_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_421_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_421_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_421_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_421_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_422_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_422_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_422_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_422_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_423_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_423_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_423_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_423_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_424_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_424_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_424_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_424_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_425_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_425_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_425_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_425_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_426_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_426_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_426_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_426_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_427_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_427_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_427_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_427_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_428_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_428_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_428_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_428_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_429_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_429_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_429_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_429_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_430_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_430_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_430_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_430_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_431_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_431_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_431_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_431_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_432_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_432_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_432_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_432_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_433_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_433_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_433_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_433_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_434_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_434_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_434_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_434_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_435_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_435_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_435_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_435_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_436_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_436_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_436_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_436_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_437_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_437_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_437_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_437_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_438_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_438_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_438_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_438_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_439_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_439_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_439_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_439_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_440_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_440_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_440_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_440_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_441_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_441_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_441_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_441_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_442_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_442_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_442_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_442_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_443_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_443_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_443_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_443_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_444_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_444_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_444_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_444_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_445_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_445_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_445_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_445_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_446_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_446_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_446_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_446_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_447_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_447_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_447_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_447_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_448_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_448_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_448_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_448_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_449_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_449_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_449_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_449_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_450_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_450_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_450_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_450_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_451_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_451_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_451_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_451_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_452_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_452_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_452_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_452_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_453_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_453_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_453_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_453_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_454_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_454_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_454_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_454_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_455_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_455_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_455_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_455_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_456_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_456_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_456_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_456_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_457_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_457_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_457_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_457_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_458_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_458_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_458_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_458_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_459_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_459_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_459_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_459_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_460_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_460_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_460_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_460_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_461_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_461_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_461_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_461_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_462_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_462_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_462_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_462_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_463_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_463_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_463_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_463_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_464_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_464_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_464_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_464_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_465_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_465_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_465_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_465_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_466_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_466_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_466_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_466_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_467_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_467_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_467_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_467_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_468_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_468_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_468_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_468_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_469_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_469_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_469_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_469_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_470_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_470_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_470_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_470_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_471_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_471_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_471_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_471_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_472_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_472_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_472_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_472_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_473_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_473_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_473_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_473_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_474_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_474_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_474_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_474_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_475_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_475_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_475_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_475_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_476_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_476_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_476_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_476_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_477_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_477_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_477_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_477_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_478_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_478_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_478_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_478_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_479_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_479_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_479_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_479_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_480_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_480_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_480_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_480_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_481_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_481_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_481_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_481_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_482_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_482_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_482_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_482_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_483_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_483_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_483_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_483_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_484_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_484_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_484_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_484_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_485_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_485_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_485_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_485_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_486_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_486_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_486_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_486_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_487_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_487_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_487_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_487_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_488_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_488_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_488_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_488_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_489_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_489_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_489_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_489_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_490_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_490_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_490_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_490_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_491_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_491_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_491_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_491_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_492_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_492_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_492_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_492_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_493_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_493_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_493_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_493_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_494_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_494_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_494_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_494_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_495_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_495_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_495_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_495_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_496_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_496_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_496_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_496_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_497_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_497_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_497_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_497_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_498_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_498_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_498_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_498_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_499_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_499_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_499_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_499_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_500_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_500_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_500_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_500_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_501_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_501_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_501_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_501_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_502_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_502_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_502_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_502_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_503_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_503_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_503_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_503_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_504_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_504_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_504_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_504_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_505_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_505_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_505_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_505_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_506_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_506_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_506_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_506_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_507_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_507_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_507_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_507_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_508_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_508_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_508_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_508_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_509_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_509_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_509_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_509_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_510_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_510_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_510_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_510_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_511_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_511_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_511_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_511_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_512_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_512_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_512_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_512_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_513_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_513_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_513_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_513_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_514_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_514_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_514_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_514_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_515_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_515_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_515_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_515_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_516_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_516_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_516_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_516_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_517_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_517_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_517_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_517_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_518_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_518_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_518_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_518_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_519_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_519_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_519_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_519_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_520_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_520_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_520_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_520_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_521_io_l1clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_521_io_clk; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_521_io_en; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_521_io_scan_mode; // @[el2_lib.scala 475:23]
  wire  rvclkhdr_522_io_l1clk; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_522_io_clk; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_522_io_en; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_522_io_scan_mode; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_523_io_l1clk; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_523_io_clk; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_523_io_en; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_523_io_scan_mode; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_524_io_l1clk; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_524_io_clk; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_524_io_en; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_524_io_scan_mode; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_525_io_l1clk; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_525_io_clk; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_525_io_en; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_525_io_scan_mode; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_526_io_l1clk; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_526_io_clk; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_526_io_en; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_526_io_scan_mode; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_527_io_l1clk; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_527_io_clk; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_527_io_en; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_527_io_scan_mode; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_528_io_l1clk; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_528_io_clk; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_528_io_en; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_528_io_scan_mode; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_529_io_l1clk; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_529_io_clk; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_529_io_en; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_529_io_scan_mode; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_530_io_l1clk; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_530_io_clk; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_530_io_en; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_530_io_scan_mode; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_531_io_l1clk; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_531_io_clk; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_531_io_en; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_531_io_scan_mode; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_532_io_l1clk; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_532_io_clk; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_532_io_en; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_532_io_scan_mode; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_533_io_l1clk; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_533_io_clk; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_533_io_en; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_533_io_scan_mode; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_534_io_l1clk; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_534_io_clk; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_534_io_en; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_534_io_scan_mode; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_535_io_l1clk; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_535_io_clk; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_535_io_en; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_535_io_scan_mode; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_536_io_l1clk; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_536_io_clk; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_536_io_en; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_536_io_scan_mode; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_537_io_l1clk; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_537_io_clk; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_537_io_en; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_537_io_scan_mode; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_538_io_l1clk; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_538_io_clk; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_538_io_en; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_538_io_scan_mode; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_539_io_l1clk; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_539_io_clk; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_539_io_en; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_539_io_scan_mode; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_540_io_l1clk; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_540_io_clk; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_540_io_en; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_540_io_scan_mode; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_541_io_l1clk; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_541_io_clk; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_541_io_en; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_541_io_scan_mode; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_542_io_l1clk; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_542_io_clk; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_542_io_en; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_542_io_scan_mode; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_543_io_l1clk; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_543_io_clk; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_543_io_en; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_543_io_scan_mode; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_544_io_l1clk; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_544_io_clk; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_544_io_en; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_544_io_scan_mode; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_545_io_l1clk; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_545_io_clk; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_545_io_en; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_545_io_scan_mode; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_546_io_l1clk; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_546_io_clk; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_546_io_en; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_546_io_scan_mode; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_547_io_l1clk; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_547_io_clk; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_547_io_en; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_547_io_scan_mode; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_548_io_l1clk; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_548_io_clk; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_548_io_en; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_548_io_scan_mode; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_549_io_l1clk; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_549_io_clk; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_549_io_en; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_549_io_scan_mode; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_550_io_l1clk; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_550_io_clk; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_550_io_en; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_550_io_scan_mode; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_551_io_l1clk; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_551_io_clk; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_551_io_en; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_551_io_scan_mode; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_552_io_l1clk; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_552_io_clk; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_552_io_en; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_552_io_scan_mode; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_553_io_l1clk; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_553_io_clk; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_553_io_en; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_553_io_scan_mode; // @[el2_lib.scala 461:22]
  wire  _T_40 = io_dec_tlu_flush_leak_one_wb & io_dec_tlu_flush_lower_wb; // @[el2_ifu_bp_ctl.scala 135:47]
  reg  leak_one_f_d1; // @[el2_ifu_bp_ctl.scala 129:56]
  wire  _T_41 = leak_one_f_d1 & io_dec_tlu_flush_lower_wb; // @[el2_ifu_bp_ctl.scala 135:93]
  wire  leak_one_f = _T_40 | _T_41; // @[el2_ifu_bp_ctl.scala 135:76]
  wire  _T = ~leak_one_f; // @[el2_ifu_bp_ctl.scala 72:46]
  wire  exu_mp_valid = io_exu_mp_pkt_misp & _T; // @[el2_ifu_bp_ctl.scala 72:44]
  wire  dec_tlu_error_wb = io_dec_tlu_br0_r_pkt_br_start_error | io_dec_tlu_br0_r_pkt_br_error; // @[el2_ifu_bp_ctl.scala 94:50]
  wire [7:0] _T_4 = io_ifc_fetch_addr_f[8:1] ^ io_ifc_fetch_addr_f[16:9]; // @[el2_lib.scala 189:47]
  wire [7:0] btb_rd_addr_f = _T_4 ^ io_ifc_fetch_addr_f[24:17]; // @[el2_lib.scala 189:85]
  wire [29:0] fetch_addr_p1_f = io_ifc_fetch_addr_f[30:1] + 30'h1; // @[el2_ifu_bp_ctl.scala 102:51]
  wire [30:0] _T_8 = {fetch_addr_p1_f,1'h0}; // @[Cat.scala 29:58]
  wire [7:0] _T_11 = _T_8[8:1] ^ _T_8[16:9]; // @[el2_lib.scala 189:47]
  wire [7:0] btb_rd_addr_p1_f = _T_11 ^ _T_8[24:17]; // @[el2_lib.scala 189:85]
  wire  _T_143 = ~io_ifc_fetch_addr_f[0]; // @[el2_ifu_bp_ctl.scala 186:40]
  wire  _T_2111 = btb_rd_addr_f == 8'h0; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_0; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2623 = _T_2111 ? btb_bank0_rd_data_way0_out_0 : 22'h0; // @[Mux.scala 27:72]
  wire  _T_2113 = btb_rd_addr_f == 8'h1; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_1; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2624 = _T_2113 ? btb_bank0_rd_data_way0_out_1 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2879 = _T_2623 | _T_2624; // @[Mux.scala 27:72]
  wire  _T_2115 = btb_rd_addr_f == 8'h2; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_2; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2625 = _T_2115 ? btb_bank0_rd_data_way0_out_2 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2880 = _T_2879 | _T_2625; // @[Mux.scala 27:72]
  wire  _T_2117 = btb_rd_addr_f == 8'h3; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_3; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2626 = _T_2117 ? btb_bank0_rd_data_way0_out_3 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2881 = _T_2880 | _T_2626; // @[Mux.scala 27:72]
  wire  _T_2119 = btb_rd_addr_f == 8'h4; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_4; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2627 = _T_2119 ? btb_bank0_rd_data_way0_out_4 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2882 = _T_2881 | _T_2627; // @[Mux.scala 27:72]
  wire  _T_2121 = btb_rd_addr_f == 8'h5; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_5; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2628 = _T_2121 ? btb_bank0_rd_data_way0_out_5 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2883 = _T_2882 | _T_2628; // @[Mux.scala 27:72]
  wire  _T_2123 = btb_rd_addr_f == 8'h6; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_6; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2629 = _T_2123 ? btb_bank0_rd_data_way0_out_6 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2884 = _T_2883 | _T_2629; // @[Mux.scala 27:72]
  wire  _T_2125 = btb_rd_addr_f == 8'h7; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_7; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2630 = _T_2125 ? btb_bank0_rd_data_way0_out_7 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2885 = _T_2884 | _T_2630; // @[Mux.scala 27:72]
  wire  _T_2127 = btb_rd_addr_f == 8'h8; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_8; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2631 = _T_2127 ? btb_bank0_rd_data_way0_out_8 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2886 = _T_2885 | _T_2631; // @[Mux.scala 27:72]
  wire  _T_2129 = btb_rd_addr_f == 8'h9; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_9; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2632 = _T_2129 ? btb_bank0_rd_data_way0_out_9 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2887 = _T_2886 | _T_2632; // @[Mux.scala 27:72]
  wire  _T_2131 = btb_rd_addr_f == 8'ha; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_10; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2633 = _T_2131 ? btb_bank0_rd_data_way0_out_10 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2888 = _T_2887 | _T_2633; // @[Mux.scala 27:72]
  wire  _T_2133 = btb_rd_addr_f == 8'hb; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_11; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2634 = _T_2133 ? btb_bank0_rd_data_way0_out_11 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2889 = _T_2888 | _T_2634; // @[Mux.scala 27:72]
  wire  _T_2135 = btb_rd_addr_f == 8'hc; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_12; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2635 = _T_2135 ? btb_bank0_rd_data_way0_out_12 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2890 = _T_2889 | _T_2635; // @[Mux.scala 27:72]
  wire  _T_2137 = btb_rd_addr_f == 8'hd; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_13; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2636 = _T_2137 ? btb_bank0_rd_data_way0_out_13 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2891 = _T_2890 | _T_2636; // @[Mux.scala 27:72]
  wire  _T_2139 = btb_rd_addr_f == 8'he; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_14; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2637 = _T_2139 ? btb_bank0_rd_data_way0_out_14 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2892 = _T_2891 | _T_2637; // @[Mux.scala 27:72]
  wire  _T_2141 = btb_rd_addr_f == 8'hf; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_15; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2638 = _T_2141 ? btb_bank0_rd_data_way0_out_15 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2893 = _T_2892 | _T_2638; // @[Mux.scala 27:72]
  wire  _T_2143 = btb_rd_addr_f == 8'h10; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_16; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2639 = _T_2143 ? btb_bank0_rd_data_way0_out_16 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2894 = _T_2893 | _T_2639; // @[Mux.scala 27:72]
  wire  _T_2145 = btb_rd_addr_f == 8'h11; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_17; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2640 = _T_2145 ? btb_bank0_rd_data_way0_out_17 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2895 = _T_2894 | _T_2640; // @[Mux.scala 27:72]
  wire  _T_2147 = btb_rd_addr_f == 8'h12; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_18; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2641 = _T_2147 ? btb_bank0_rd_data_way0_out_18 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2896 = _T_2895 | _T_2641; // @[Mux.scala 27:72]
  wire  _T_2149 = btb_rd_addr_f == 8'h13; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_19; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2642 = _T_2149 ? btb_bank0_rd_data_way0_out_19 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2897 = _T_2896 | _T_2642; // @[Mux.scala 27:72]
  wire  _T_2151 = btb_rd_addr_f == 8'h14; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_20; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2643 = _T_2151 ? btb_bank0_rd_data_way0_out_20 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2898 = _T_2897 | _T_2643; // @[Mux.scala 27:72]
  wire  _T_2153 = btb_rd_addr_f == 8'h15; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_21; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2644 = _T_2153 ? btb_bank0_rd_data_way0_out_21 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2899 = _T_2898 | _T_2644; // @[Mux.scala 27:72]
  wire  _T_2155 = btb_rd_addr_f == 8'h16; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_22; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2645 = _T_2155 ? btb_bank0_rd_data_way0_out_22 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2900 = _T_2899 | _T_2645; // @[Mux.scala 27:72]
  wire  _T_2157 = btb_rd_addr_f == 8'h17; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_23; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2646 = _T_2157 ? btb_bank0_rd_data_way0_out_23 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2901 = _T_2900 | _T_2646; // @[Mux.scala 27:72]
  wire  _T_2159 = btb_rd_addr_f == 8'h18; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_24; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2647 = _T_2159 ? btb_bank0_rd_data_way0_out_24 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2902 = _T_2901 | _T_2647; // @[Mux.scala 27:72]
  wire  _T_2161 = btb_rd_addr_f == 8'h19; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_25; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2648 = _T_2161 ? btb_bank0_rd_data_way0_out_25 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2903 = _T_2902 | _T_2648; // @[Mux.scala 27:72]
  wire  _T_2163 = btb_rd_addr_f == 8'h1a; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_26; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2649 = _T_2163 ? btb_bank0_rd_data_way0_out_26 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2904 = _T_2903 | _T_2649; // @[Mux.scala 27:72]
  wire  _T_2165 = btb_rd_addr_f == 8'h1b; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_27; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2650 = _T_2165 ? btb_bank0_rd_data_way0_out_27 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2905 = _T_2904 | _T_2650; // @[Mux.scala 27:72]
  wire  _T_2167 = btb_rd_addr_f == 8'h1c; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_28; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2651 = _T_2167 ? btb_bank0_rd_data_way0_out_28 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2906 = _T_2905 | _T_2651; // @[Mux.scala 27:72]
  wire  _T_2169 = btb_rd_addr_f == 8'h1d; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_29; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2652 = _T_2169 ? btb_bank0_rd_data_way0_out_29 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2907 = _T_2906 | _T_2652; // @[Mux.scala 27:72]
  wire  _T_2171 = btb_rd_addr_f == 8'h1e; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_30; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2653 = _T_2171 ? btb_bank0_rd_data_way0_out_30 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2908 = _T_2907 | _T_2653; // @[Mux.scala 27:72]
  wire  _T_2173 = btb_rd_addr_f == 8'h1f; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_31; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2654 = _T_2173 ? btb_bank0_rd_data_way0_out_31 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2909 = _T_2908 | _T_2654; // @[Mux.scala 27:72]
  wire  _T_2175 = btb_rd_addr_f == 8'h20; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_32; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2655 = _T_2175 ? btb_bank0_rd_data_way0_out_32 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2910 = _T_2909 | _T_2655; // @[Mux.scala 27:72]
  wire  _T_2177 = btb_rd_addr_f == 8'h21; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_33; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2656 = _T_2177 ? btb_bank0_rd_data_way0_out_33 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2911 = _T_2910 | _T_2656; // @[Mux.scala 27:72]
  wire  _T_2179 = btb_rd_addr_f == 8'h22; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_34; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2657 = _T_2179 ? btb_bank0_rd_data_way0_out_34 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2912 = _T_2911 | _T_2657; // @[Mux.scala 27:72]
  wire  _T_2181 = btb_rd_addr_f == 8'h23; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_35; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2658 = _T_2181 ? btb_bank0_rd_data_way0_out_35 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2913 = _T_2912 | _T_2658; // @[Mux.scala 27:72]
  wire  _T_2183 = btb_rd_addr_f == 8'h24; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_36; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2659 = _T_2183 ? btb_bank0_rd_data_way0_out_36 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2914 = _T_2913 | _T_2659; // @[Mux.scala 27:72]
  wire  _T_2185 = btb_rd_addr_f == 8'h25; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_37; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2660 = _T_2185 ? btb_bank0_rd_data_way0_out_37 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2915 = _T_2914 | _T_2660; // @[Mux.scala 27:72]
  wire  _T_2187 = btb_rd_addr_f == 8'h26; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_38; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2661 = _T_2187 ? btb_bank0_rd_data_way0_out_38 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2916 = _T_2915 | _T_2661; // @[Mux.scala 27:72]
  wire  _T_2189 = btb_rd_addr_f == 8'h27; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_39; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2662 = _T_2189 ? btb_bank0_rd_data_way0_out_39 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2917 = _T_2916 | _T_2662; // @[Mux.scala 27:72]
  wire  _T_2191 = btb_rd_addr_f == 8'h28; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_40; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2663 = _T_2191 ? btb_bank0_rd_data_way0_out_40 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2918 = _T_2917 | _T_2663; // @[Mux.scala 27:72]
  wire  _T_2193 = btb_rd_addr_f == 8'h29; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_41; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2664 = _T_2193 ? btb_bank0_rd_data_way0_out_41 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2919 = _T_2918 | _T_2664; // @[Mux.scala 27:72]
  wire  _T_2195 = btb_rd_addr_f == 8'h2a; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_42; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2665 = _T_2195 ? btb_bank0_rd_data_way0_out_42 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2920 = _T_2919 | _T_2665; // @[Mux.scala 27:72]
  wire  _T_2197 = btb_rd_addr_f == 8'h2b; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_43; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2666 = _T_2197 ? btb_bank0_rd_data_way0_out_43 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2921 = _T_2920 | _T_2666; // @[Mux.scala 27:72]
  wire  _T_2199 = btb_rd_addr_f == 8'h2c; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_44; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2667 = _T_2199 ? btb_bank0_rd_data_way0_out_44 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2922 = _T_2921 | _T_2667; // @[Mux.scala 27:72]
  wire  _T_2201 = btb_rd_addr_f == 8'h2d; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_45; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2668 = _T_2201 ? btb_bank0_rd_data_way0_out_45 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2923 = _T_2922 | _T_2668; // @[Mux.scala 27:72]
  wire  _T_2203 = btb_rd_addr_f == 8'h2e; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_46; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2669 = _T_2203 ? btb_bank0_rd_data_way0_out_46 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2924 = _T_2923 | _T_2669; // @[Mux.scala 27:72]
  wire  _T_2205 = btb_rd_addr_f == 8'h2f; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_47; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2670 = _T_2205 ? btb_bank0_rd_data_way0_out_47 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2925 = _T_2924 | _T_2670; // @[Mux.scala 27:72]
  wire  _T_2207 = btb_rd_addr_f == 8'h30; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_48; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2671 = _T_2207 ? btb_bank0_rd_data_way0_out_48 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2926 = _T_2925 | _T_2671; // @[Mux.scala 27:72]
  wire  _T_2209 = btb_rd_addr_f == 8'h31; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_49; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2672 = _T_2209 ? btb_bank0_rd_data_way0_out_49 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2927 = _T_2926 | _T_2672; // @[Mux.scala 27:72]
  wire  _T_2211 = btb_rd_addr_f == 8'h32; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_50; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2673 = _T_2211 ? btb_bank0_rd_data_way0_out_50 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2928 = _T_2927 | _T_2673; // @[Mux.scala 27:72]
  wire  _T_2213 = btb_rd_addr_f == 8'h33; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_51; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2674 = _T_2213 ? btb_bank0_rd_data_way0_out_51 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2929 = _T_2928 | _T_2674; // @[Mux.scala 27:72]
  wire  _T_2215 = btb_rd_addr_f == 8'h34; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_52; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2675 = _T_2215 ? btb_bank0_rd_data_way0_out_52 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2930 = _T_2929 | _T_2675; // @[Mux.scala 27:72]
  wire  _T_2217 = btb_rd_addr_f == 8'h35; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_53; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2676 = _T_2217 ? btb_bank0_rd_data_way0_out_53 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2931 = _T_2930 | _T_2676; // @[Mux.scala 27:72]
  wire  _T_2219 = btb_rd_addr_f == 8'h36; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_54; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2677 = _T_2219 ? btb_bank0_rd_data_way0_out_54 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2932 = _T_2931 | _T_2677; // @[Mux.scala 27:72]
  wire  _T_2221 = btb_rd_addr_f == 8'h37; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_55; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2678 = _T_2221 ? btb_bank0_rd_data_way0_out_55 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2933 = _T_2932 | _T_2678; // @[Mux.scala 27:72]
  wire  _T_2223 = btb_rd_addr_f == 8'h38; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_56; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2679 = _T_2223 ? btb_bank0_rd_data_way0_out_56 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2934 = _T_2933 | _T_2679; // @[Mux.scala 27:72]
  wire  _T_2225 = btb_rd_addr_f == 8'h39; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_57; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2680 = _T_2225 ? btb_bank0_rd_data_way0_out_57 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2935 = _T_2934 | _T_2680; // @[Mux.scala 27:72]
  wire  _T_2227 = btb_rd_addr_f == 8'h3a; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_58; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2681 = _T_2227 ? btb_bank0_rd_data_way0_out_58 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2936 = _T_2935 | _T_2681; // @[Mux.scala 27:72]
  wire  _T_2229 = btb_rd_addr_f == 8'h3b; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_59; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2682 = _T_2229 ? btb_bank0_rd_data_way0_out_59 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2937 = _T_2936 | _T_2682; // @[Mux.scala 27:72]
  wire  _T_2231 = btb_rd_addr_f == 8'h3c; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_60; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2683 = _T_2231 ? btb_bank0_rd_data_way0_out_60 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2938 = _T_2937 | _T_2683; // @[Mux.scala 27:72]
  wire  _T_2233 = btb_rd_addr_f == 8'h3d; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_61; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2684 = _T_2233 ? btb_bank0_rd_data_way0_out_61 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2939 = _T_2938 | _T_2684; // @[Mux.scala 27:72]
  wire  _T_2235 = btb_rd_addr_f == 8'h3e; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_62; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2685 = _T_2235 ? btb_bank0_rd_data_way0_out_62 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2940 = _T_2939 | _T_2685; // @[Mux.scala 27:72]
  wire  _T_2237 = btb_rd_addr_f == 8'h3f; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_63; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2686 = _T_2237 ? btb_bank0_rd_data_way0_out_63 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2941 = _T_2940 | _T_2686; // @[Mux.scala 27:72]
  wire  _T_2239 = btb_rd_addr_f == 8'h40; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_64; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2687 = _T_2239 ? btb_bank0_rd_data_way0_out_64 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2942 = _T_2941 | _T_2687; // @[Mux.scala 27:72]
  wire  _T_2241 = btb_rd_addr_f == 8'h41; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_65; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2688 = _T_2241 ? btb_bank0_rd_data_way0_out_65 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2943 = _T_2942 | _T_2688; // @[Mux.scala 27:72]
  wire  _T_2243 = btb_rd_addr_f == 8'h42; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_66; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2689 = _T_2243 ? btb_bank0_rd_data_way0_out_66 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2944 = _T_2943 | _T_2689; // @[Mux.scala 27:72]
  wire  _T_2245 = btb_rd_addr_f == 8'h43; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_67; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2690 = _T_2245 ? btb_bank0_rd_data_way0_out_67 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2945 = _T_2944 | _T_2690; // @[Mux.scala 27:72]
  wire  _T_2247 = btb_rd_addr_f == 8'h44; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_68; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2691 = _T_2247 ? btb_bank0_rd_data_way0_out_68 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2946 = _T_2945 | _T_2691; // @[Mux.scala 27:72]
  wire  _T_2249 = btb_rd_addr_f == 8'h45; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_69; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2692 = _T_2249 ? btb_bank0_rd_data_way0_out_69 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2947 = _T_2946 | _T_2692; // @[Mux.scala 27:72]
  wire  _T_2251 = btb_rd_addr_f == 8'h46; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_70; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2693 = _T_2251 ? btb_bank0_rd_data_way0_out_70 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2948 = _T_2947 | _T_2693; // @[Mux.scala 27:72]
  wire  _T_2253 = btb_rd_addr_f == 8'h47; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_71; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2694 = _T_2253 ? btb_bank0_rd_data_way0_out_71 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2949 = _T_2948 | _T_2694; // @[Mux.scala 27:72]
  wire  _T_2255 = btb_rd_addr_f == 8'h48; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_72; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2695 = _T_2255 ? btb_bank0_rd_data_way0_out_72 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2950 = _T_2949 | _T_2695; // @[Mux.scala 27:72]
  wire  _T_2257 = btb_rd_addr_f == 8'h49; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_73; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2696 = _T_2257 ? btb_bank0_rd_data_way0_out_73 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2951 = _T_2950 | _T_2696; // @[Mux.scala 27:72]
  wire  _T_2259 = btb_rd_addr_f == 8'h4a; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_74; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2697 = _T_2259 ? btb_bank0_rd_data_way0_out_74 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2952 = _T_2951 | _T_2697; // @[Mux.scala 27:72]
  wire  _T_2261 = btb_rd_addr_f == 8'h4b; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_75; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2698 = _T_2261 ? btb_bank0_rd_data_way0_out_75 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2953 = _T_2952 | _T_2698; // @[Mux.scala 27:72]
  wire  _T_2263 = btb_rd_addr_f == 8'h4c; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_76; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2699 = _T_2263 ? btb_bank0_rd_data_way0_out_76 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2954 = _T_2953 | _T_2699; // @[Mux.scala 27:72]
  wire  _T_2265 = btb_rd_addr_f == 8'h4d; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_77; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2700 = _T_2265 ? btb_bank0_rd_data_way0_out_77 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2955 = _T_2954 | _T_2700; // @[Mux.scala 27:72]
  wire  _T_2267 = btb_rd_addr_f == 8'h4e; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_78; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2701 = _T_2267 ? btb_bank0_rd_data_way0_out_78 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2956 = _T_2955 | _T_2701; // @[Mux.scala 27:72]
  wire  _T_2269 = btb_rd_addr_f == 8'h4f; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_79; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2702 = _T_2269 ? btb_bank0_rd_data_way0_out_79 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2957 = _T_2956 | _T_2702; // @[Mux.scala 27:72]
  wire  _T_2271 = btb_rd_addr_f == 8'h50; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_80; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2703 = _T_2271 ? btb_bank0_rd_data_way0_out_80 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2958 = _T_2957 | _T_2703; // @[Mux.scala 27:72]
  wire  _T_2273 = btb_rd_addr_f == 8'h51; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_81; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2704 = _T_2273 ? btb_bank0_rd_data_way0_out_81 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2959 = _T_2958 | _T_2704; // @[Mux.scala 27:72]
  wire  _T_2275 = btb_rd_addr_f == 8'h52; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_82; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2705 = _T_2275 ? btb_bank0_rd_data_way0_out_82 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2960 = _T_2959 | _T_2705; // @[Mux.scala 27:72]
  wire  _T_2277 = btb_rd_addr_f == 8'h53; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_83; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2706 = _T_2277 ? btb_bank0_rd_data_way0_out_83 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2961 = _T_2960 | _T_2706; // @[Mux.scala 27:72]
  wire  _T_2279 = btb_rd_addr_f == 8'h54; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_84; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2707 = _T_2279 ? btb_bank0_rd_data_way0_out_84 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2962 = _T_2961 | _T_2707; // @[Mux.scala 27:72]
  wire  _T_2281 = btb_rd_addr_f == 8'h55; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_85; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2708 = _T_2281 ? btb_bank0_rd_data_way0_out_85 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2963 = _T_2962 | _T_2708; // @[Mux.scala 27:72]
  wire  _T_2283 = btb_rd_addr_f == 8'h56; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_86; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2709 = _T_2283 ? btb_bank0_rd_data_way0_out_86 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2964 = _T_2963 | _T_2709; // @[Mux.scala 27:72]
  wire  _T_2285 = btb_rd_addr_f == 8'h57; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_87; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2710 = _T_2285 ? btb_bank0_rd_data_way0_out_87 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2965 = _T_2964 | _T_2710; // @[Mux.scala 27:72]
  wire  _T_2287 = btb_rd_addr_f == 8'h58; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_88; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2711 = _T_2287 ? btb_bank0_rd_data_way0_out_88 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2966 = _T_2965 | _T_2711; // @[Mux.scala 27:72]
  wire  _T_2289 = btb_rd_addr_f == 8'h59; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_89; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2712 = _T_2289 ? btb_bank0_rd_data_way0_out_89 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2967 = _T_2966 | _T_2712; // @[Mux.scala 27:72]
  wire  _T_2291 = btb_rd_addr_f == 8'h5a; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_90; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2713 = _T_2291 ? btb_bank0_rd_data_way0_out_90 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2968 = _T_2967 | _T_2713; // @[Mux.scala 27:72]
  wire  _T_2293 = btb_rd_addr_f == 8'h5b; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_91; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2714 = _T_2293 ? btb_bank0_rd_data_way0_out_91 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2969 = _T_2968 | _T_2714; // @[Mux.scala 27:72]
  wire  _T_2295 = btb_rd_addr_f == 8'h5c; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_92; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2715 = _T_2295 ? btb_bank0_rd_data_way0_out_92 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2970 = _T_2969 | _T_2715; // @[Mux.scala 27:72]
  wire  _T_2297 = btb_rd_addr_f == 8'h5d; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_93; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2716 = _T_2297 ? btb_bank0_rd_data_way0_out_93 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2971 = _T_2970 | _T_2716; // @[Mux.scala 27:72]
  wire  _T_2299 = btb_rd_addr_f == 8'h5e; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_94; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2717 = _T_2299 ? btb_bank0_rd_data_way0_out_94 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2972 = _T_2971 | _T_2717; // @[Mux.scala 27:72]
  wire  _T_2301 = btb_rd_addr_f == 8'h5f; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_95; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2718 = _T_2301 ? btb_bank0_rd_data_way0_out_95 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2973 = _T_2972 | _T_2718; // @[Mux.scala 27:72]
  wire  _T_2303 = btb_rd_addr_f == 8'h60; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_96; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2719 = _T_2303 ? btb_bank0_rd_data_way0_out_96 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2974 = _T_2973 | _T_2719; // @[Mux.scala 27:72]
  wire  _T_2305 = btb_rd_addr_f == 8'h61; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_97; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2720 = _T_2305 ? btb_bank0_rd_data_way0_out_97 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2975 = _T_2974 | _T_2720; // @[Mux.scala 27:72]
  wire  _T_2307 = btb_rd_addr_f == 8'h62; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_98; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2721 = _T_2307 ? btb_bank0_rd_data_way0_out_98 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2976 = _T_2975 | _T_2721; // @[Mux.scala 27:72]
  wire  _T_2309 = btb_rd_addr_f == 8'h63; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_99; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2722 = _T_2309 ? btb_bank0_rd_data_way0_out_99 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2977 = _T_2976 | _T_2722; // @[Mux.scala 27:72]
  wire  _T_2311 = btb_rd_addr_f == 8'h64; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_100; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2723 = _T_2311 ? btb_bank0_rd_data_way0_out_100 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2978 = _T_2977 | _T_2723; // @[Mux.scala 27:72]
  wire  _T_2313 = btb_rd_addr_f == 8'h65; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_101; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2724 = _T_2313 ? btb_bank0_rd_data_way0_out_101 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2979 = _T_2978 | _T_2724; // @[Mux.scala 27:72]
  wire  _T_2315 = btb_rd_addr_f == 8'h66; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_102; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2725 = _T_2315 ? btb_bank0_rd_data_way0_out_102 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2980 = _T_2979 | _T_2725; // @[Mux.scala 27:72]
  wire  _T_2317 = btb_rd_addr_f == 8'h67; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_103; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2726 = _T_2317 ? btb_bank0_rd_data_way0_out_103 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2981 = _T_2980 | _T_2726; // @[Mux.scala 27:72]
  wire  _T_2319 = btb_rd_addr_f == 8'h68; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_104; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2727 = _T_2319 ? btb_bank0_rd_data_way0_out_104 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2982 = _T_2981 | _T_2727; // @[Mux.scala 27:72]
  wire  _T_2321 = btb_rd_addr_f == 8'h69; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_105; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2728 = _T_2321 ? btb_bank0_rd_data_way0_out_105 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2983 = _T_2982 | _T_2728; // @[Mux.scala 27:72]
  wire  _T_2323 = btb_rd_addr_f == 8'h6a; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_106; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2729 = _T_2323 ? btb_bank0_rd_data_way0_out_106 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2984 = _T_2983 | _T_2729; // @[Mux.scala 27:72]
  wire  _T_2325 = btb_rd_addr_f == 8'h6b; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_107; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2730 = _T_2325 ? btb_bank0_rd_data_way0_out_107 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2985 = _T_2984 | _T_2730; // @[Mux.scala 27:72]
  wire  _T_2327 = btb_rd_addr_f == 8'h6c; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_108; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2731 = _T_2327 ? btb_bank0_rd_data_way0_out_108 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2986 = _T_2985 | _T_2731; // @[Mux.scala 27:72]
  wire  _T_2329 = btb_rd_addr_f == 8'h6d; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_109; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2732 = _T_2329 ? btb_bank0_rd_data_way0_out_109 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2987 = _T_2986 | _T_2732; // @[Mux.scala 27:72]
  wire  _T_2331 = btb_rd_addr_f == 8'h6e; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_110; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2733 = _T_2331 ? btb_bank0_rd_data_way0_out_110 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2988 = _T_2987 | _T_2733; // @[Mux.scala 27:72]
  wire  _T_2333 = btb_rd_addr_f == 8'h6f; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_111; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2734 = _T_2333 ? btb_bank0_rd_data_way0_out_111 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2989 = _T_2988 | _T_2734; // @[Mux.scala 27:72]
  wire  _T_2335 = btb_rd_addr_f == 8'h70; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_112; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2735 = _T_2335 ? btb_bank0_rd_data_way0_out_112 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2990 = _T_2989 | _T_2735; // @[Mux.scala 27:72]
  wire  _T_2337 = btb_rd_addr_f == 8'h71; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_113; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2736 = _T_2337 ? btb_bank0_rd_data_way0_out_113 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2991 = _T_2990 | _T_2736; // @[Mux.scala 27:72]
  wire  _T_2339 = btb_rd_addr_f == 8'h72; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_114; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2737 = _T_2339 ? btb_bank0_rd_data_way0_out_114 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2992 = _T_2991 | _T_2737; // @[Mux.scala 27:72]
  wire  _T_2341 = btb_rd_addr_f == 8'h73; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_115; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2738 = _T_2341 ? btb_bank0_rd_data_way0_out_115 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2993 = _T_2992 | _T_2738; // @[Mux.scala 27:72]
  wire  _T_2343 = btb_rd_addr_f == 8'h74; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_116; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2739 = _T_2343 ? btb_bank0_rd_data_way0_out_116 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2994 = _T_2993 | _T_2739; // @[Mux.scala 27:72]
  wire  _T_2345 = btb_rd_addr_f == 8'h75; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_117; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2740 = _T_2345 ? btb_bank0_rd_data_way0_out_117 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2995 = _T_2994 | _T_2740; // @[Mux.scala 27:72]
  wire  _T_2347 = btb_rd_addr_f == 8'h76; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_118; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2741 = _T_2347 ? btb_bank0_rd_data_way0_out_118 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2996 = _T_2995 | _T_2741; // @[Mux.scala 27:72]
  wire  _T_2349 = btb_rd_addr_f == 8'h77; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_119; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2742 = _T_2349 ? btb_bank0_rd_data_way0_out_119 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2997 = _T_2996 | _T_2742; // @[Mux.scala 27:72]
  wire  _T_2351 = btb_rd_addr_f == 8'h78; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_120; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2743 = _T_2351 ? btb_bank0_rd_data_way0_out_120 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2998 = _T_2997 | _T_2743; // @[Mux.scala 27:72]
  wire  _T_2353 = btb_rd_addr_f == 8'h79; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_121; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2744 = _T_2353 ? btb_bank0_rd_data_way0_out_121 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2999 = _T_2998 | _T_2744; // @[Mux.scala 27:72]
  wire  _T_2355 = btb_rd_addr_f == 8'h7a; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_122; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2745 = _T_2355 ? btb_bank0_rd_data_way0_out_122 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3000 = _T_2999 | _T_2745; // @[Mux.scala 27:72]
  wire  _T_2357 = btb_rd_addr_f == 8'h7b; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_123; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2746 = _T_2357 ? btb_bank0_rd_data_way0_out_123 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3001 = _T_3000 | _T_2746; // @[Mux.scala 27:72]
  wire  _T_2359 = btb_rd_addr_f == 8'h7c; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_124; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2747 = _T_2359 ? btb_bank0_rd_data_way0_out_124 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3002 = _T_3001 | _T_2747; // @[Mux.scala 27:72]
  wire  _T_2361 = btb_rd_addr_f == 8'h7d; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_125; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2748 = _T_2361 ? btb_bank0_rd_data_way0_out_125 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3003 = _T_3002 | _T_2748; // @[Mux.scala 27:72]
  wire  _T_2363 = btb_rd_addr_f == 8'h7e; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_126; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2749 = _T_2363 ? btb_bank0_rd_data_way0_out_126 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3004 = _T_3003 | _T_2749; // @[Mux.scala 27:72]
  wire  _T_2365 = btb_rd_addr_f == 8'h7f; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_127; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2750 = _T_2365 ? btb_bank0_rd_data_way0_out_127 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3005 = _T_3004 | _T_2750; // @[Mux.scala 27:72]
  wire  _T_2367 = btb_rd_addr_f == 8'h80; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_128; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2751 = _T_2367 ? btb_bank0_rd_data_way0_out_128 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3006 = _T_3005 | _T_2751; // @[Mux.scala 27:72]
  wire  _T_2369 = btb_rd_addr_f == 8'h81; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_129; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2752 = _T_2369 ? btb_bank0_rd_data_way0_out_129 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3007 = _T_3006 | _T_2752; // @[Mux.scala 27:72]
  wire  _T_2371 = btb_rd_addr_f == 8'h82; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_130; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2753 = _T_2371 ? btb_bank0_rd_data_way0_out_130 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3008 = _T_3007 | _T_2753; // @[Mux.scala 27:72]
  wire  _T_2373 = btb_rd_addr_f == 8'h83; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_131; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2754 = _T_2373 ? btb_bank0_rd_data_way0_out_131 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3009 = _T_3008 | _T_2754; // @[Mux.scala 27:72]
  wire  _T_2375 = btb_rd_addr_f == 8'h84; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_132; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2755 = _T_2375 ? btb_bank0_rd_data_way0_out_132 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3010 = _T_3009 | _T_2755; // @[Mux.scala 27:72]
  wire  _T_2377 = btb_rd_addr_f == 8'h85; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_133; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2756 = _T_2377 ? btb_bank0_rd_data_way0_out_133 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3011 = _T_3010 | _T_2756; // @[Mux.scala 27:72]
  wire  _T_2379 = btb_rd_addr_f == 8'h86; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_134; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2757 = _T_2379 ? btb_bank0_rd_data_way0_out_134 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3012 = _T_3011 | _T_2757; // @[Mux.scala 27:72]
  wire  _T_2381 = btb_rd_addr_f == 8'h87; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_135; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2758 = _T_2381 ? btb_bank0_rd_data_way0_out_135 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3013 = _T_3012 | _T_2758; // @[Mux.scala 27:72]
  wire  _T_2383 = btb_rd_addr_f == 8'h88; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_136; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2759 = _T_2383 ? btb_bank0_rd_data_way0_out_136 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3014 = _T_3013 | _T_2759; // @[Mux.scala 27:72]
  wire  _T_2385 = btb_rd_addr_f == 8'h89; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_137; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2760 = _T_2385 ? btb_bank0_rd_data_way0_out_137 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3015 = _T_3014 | _T_2760; // @[Mux.scala 27:72]
  wire  _T_2387 = btb_rd_addr_f == 8'h8a; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_138; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2761 = _T_2387 ? btb_bank0_rd_data_way0_out_138 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3016 = _T_3015 | _T_2761; // @[Mux.scala 27:72]
  wire  _T_2389 = btb_rd_addr_f == 8'h8b; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_139; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2762 = _T_2389 ? btb_bank0_rd_data_way0_out_139 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3017 = _T_3016 | _T_2762; // @[Mux.scala 27:72]
  wire  _T_2391 = btb_rd_addr_f == 8'h8c; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_140; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2763 = _T_2391 ? btb_bank0_rd_data_way0_out_140 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3018 = _T_3017 | _T_2763; // @[Mux.scala 27:72]
  wire  _T_2393 = btb_rd_addr_f == 8'h8d; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_141; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2764 = _T_2393 ? btb_bank0_rd_data_way0_out_141 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3019 = _T_3018 | _T_2764; // @[Mux.scala 27:72]
  wire  _T_2395 = btb_rd_addr_f == 8'h8e; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_142; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2765 = _T_2395 ? btb_bank0_rd_data_way0_out_142 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3020 = _T_3019 | _T_2765; // @[Mux.scala 27:72]
  wire  _T_2397 = btb_rd_addr_f == 8'h8f; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_143; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2766 = _T_2397 ? btb_bank0_rd_data_way0_out_143 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3021 = _T_3020 | _T_2766; // @[Mux.scala 27:72]
  wire  _T_2399 = btb_rd_addr_f == 8'h90; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_144; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2767 = _T_2399 ? btb_bank0_rd_data_way0_out_144 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3022 = _T_3021 | _T_2767; // @[Mux.scala 27:72]
  wire  _T_2401 = btb_rd_addr_f == 8'h91; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_145; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2768 = _T_2401 ? btb_bank0_rd_data_way0_out_145 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3023 = _T_3022 | _T_2768; // @[Mux.scala 27:72]
  wire  _T_2403 = btb_rd_addr_f == 8'h92; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_146; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2769 = _T_2403 ? btb_bank0_rd_data_way0_out_146 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3024 = _T_3023 | _T_2769; // @[Mux.scala 27:72]
  wire  _T_2405 = btb_rd_addr_f == 8'h93; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_147; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2770 = _T_2405 ? btb_bank0_rd_data_way0_out_147 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3025 = _T_3024 | _T_2770; // @[Mux.scala 27:72]
  wire  _T_2407 = btb_rd_addr_f == 8'h94; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_148; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2771 = _T_2407 ? btb_bank0_rd_data_way0_out_148 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3026 = _T_3025 | _T_2771; // @[Mux.scala 27:72]
  wire  _T_2409 = btb_rd_addr_f == 8'h95; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_149; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2772 = _T_2409 ? btb_bank0_rd_data_way0_out_149 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3027 = _T_3026 | _T_2772; // @[Mux.scala 27:72]
  wire  _T_2411 = btb_rd_addr_f == 8'h96; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_150; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2773 = _T_2411 ? btb_bank0_rd_data_way0_out_150 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3028 = _T_3027 | _T_2773; // @[Mux.scala 27:72]
  wire  _T_2413 = btb_rd_addr_f == 8'h97; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_151; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2774 = _T_2413 ? btb_bank0_rd_data_way0_out_151 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3029 = _T_3028 | _T_2774; // @[Mux.scala 27:72]
  wire  _T_2415 = btb_rd_addr_f == 8'h98; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_152; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2775 = _T_2415 ? btb_bank0_rd_data_way0_out_152 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3030 = _T_3029 | _T_2775; // @[Mux.scala 27:72]
  wire  _T_2417 = btb_rd_addr_f == 8'h99; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_153; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2776 = _T_2417 ? btb_bank0_rd_data_way0_out_153 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3031 = _T_3030 | _T_2776; // @[Mux.scala 27:72]
  wire  _T_2419 = btb_rd_addr_f == 8'h9a; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_154; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2777 = _T_2419 ? btb_bank0_rd_data_way0_out_154 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3032 = _T_3031 | _T_2777; // @[Mux.scala 27:72]
  wire  _T_2421 = btb_rd_addr_f == 8'h9b; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_155; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2778 = _T_2421 ? btb_bank0_rd_data_way0_out_155 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3033 = _T_3032 | _T_2778; // @[Mux.scala 27:72]
  wire  _T_2423 = btb_rd_addr_f == 8'h9c; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_156; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2779 = _T_2423 ? btb_bank0_rd_data_way0_out_156 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3034 = _T_3033 | _T_2779; // @[Mux.scala 27:72]
  wire  _T_2425 = btb_rd_addr_f == 8'h9d; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_157; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2780 = _T_2425 ? btb_bank0_rd_data_way0_out_157 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3035 = _T_3034 | _T_2780; // @[Mux.scala 27:72]
  wire  _T_2427 = btb_rd_addr_f == 8'h9e; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_158; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2781 = _T_2427 ? btb_bank0_rd_data_way0_out_158 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3036 = _T_3035 | _T_2781; // @[Mux.scala 27:72]
  wire  _T_2429 = btb_rd_addr_f == 8'h9f; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_159; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2782 = _T_2429 ? btb_bank0_rd_data_way0_out_159 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3037 = _T_3036 | _T_2782; // @[Mux.scala 27:72]
  wire  _T_2431 = btb_rd_addr_f == 8'ha0; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_160; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2783 = _T_2431 ? btb_bank0_rd_data_way0_out_160 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3038 = _T_3037 | _T_2783; // @[Mux.scala 27:72]
  wire  _T_2433 = btb_rd_addr_f == 8'ha1; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_161; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2784 = _T_2433 ? btb_bank0_rd_data_way0_out_161 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3039 = _T_3038 | _T_2784; // @[Mux.scala 27:72]
  wire  _T_2435 = btb_rd_addr_f == 8'ha2; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_162; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2785 = _T_2435 ? btb_bank0_rd_data_way0_out_162 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3040 = _T_3039 | _T_2785; // @[Mux.scala 27:72]
  wire  _T_2437 = btb_rd_addr_f == 8'ha3; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_163; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2786 = _T_2437 ? btb_bank0_rd_data_way0_out_163 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3041 = _T_3040 | _T_2786; // @[Mux.scala 27:72]
  wire  _T_2439 = btb_rd_addr_f == 8'ha4; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_164; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2787 = _T_2439 ? btb_bank0_rd_data_way0_out_164 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3042 = _T_3041 | _T_2787; // @[Mux.scala 27:72]
  wire  _T_2441 = btb_rd_addr_f == 8'ha5; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_165; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2788 = _T_2441 ? btb_bank0_rd_data_way0_out_165 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3043 = _T_3042 | _T_2788; // @[Mux.scala 27:72]
  wire  _T_2443 = btb_rd_addr_f == 8'ha6; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_166; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2789 = _T_2443 ? btb_bank0_rd_data_way0_out_166 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3044 = _T_3043 | _T_2789; // @[Mux.scala 27:72]
  wire  _T_2445 = btb_rd_addr_f == 8'ha7; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_167; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2790 = _T_2445 ? btb_bank0_rd_data_way0_out_167 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3045 = _T_3044 | _T_2790; // @[Mux.scala 27:72]
  wire  _T_2447 = btb_rd_addr_f == 8'ha8; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_168; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2791 = _T_2447 ? btb_bank0_rd_data_way0_out_168 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3046 = _T_3045 | _T_2791; // @[Mux.scala 27:72]
  wire  _T_2449 = btb_rd_addr_f == 8'ha9; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_169; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2792 = _T_2449 ? btb_bank0_rd_data_way0_out_169 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3047 = _T_3046 | _T_2792; // @[Mux.scala 27:72]
  wire  _T_2451 = btb_rd_addr_f == 8'haa; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_170; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2793 = _T_2451 ? btb_bank0_rd_data_way0_out_170 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3048 = _T_3047 | _T_2793; // @[Mux.scala 27:72]
  wire  _T_2453 = btb_rd_addr_f == 8'hab; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_171; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2794 = _T_2453 ? btb_bank0_rd_data_way0_out_171 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3049 = _T_3048 | _T_2794; // @[Mux.scala 27:72]
  wire  _T_2455 = btb_rd_addr_f == 8'hac; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_172; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2795 = _T_2455 ? btb_bank0_rd_data_way0_out_172 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3050 = _T_3049 | _T_2795; // @[Mux.scala 27:72]
  wire  _T_2457 = btb_rd_addr_f == 8'had; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_173; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2796 = _T_2457 ? btb_bank0_rd_data_way0_out_173 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3051 = _T_3050 | _T_2796; // @[Mux.scala 27:72]
  wire  _T_2459 = btb_rd_addr_f == 8'hae; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_174; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2797 = _T_2459 ? btb_bank0_rd_data_way0_out_174 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3052 = _T_3051 | _T_2797; // @[Mux.scala 27:72]
  wire  _T_2461 = btb_rd_addr_f == 8'haf; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_175; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2798 = _T_2461 ? btb_bank0_rd_data_way0_out_175 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3053 = _T_3052 | _T_2798; // @[Mux.scala 27:72]
  wire  _T_2463 = btb_rd_addr_f == 8'hb0; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_176; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2799 = _T_2463 ? btb_bank0_rd_data_way0_out_176 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3054 = _T_3053 | _T_2799; // @[Mux.scala 27:72]
  wire  _T_2465 = btb_rd_addr_f == 8'hb1; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_177; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2800 = _T_2465 ? btb_bank0_rd_data_way0_out_177 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3055 = _T_3054 | _T_2800; // @[Mux.scala 27:72]
  wire  _T_2467 = btb_rd_addr_f == 8'hb2; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_178; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2801 = _T_2467 ? btb_bank0_rd_data_way0_out_178 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3056 = _T_3055 | _T_2801; // @[Mux.scala 27:72]
  wire  _T_2469 = btb_rd_addr_f == 8'hb3; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_179; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2802 = _T_2469 ? btb_bank0_rd_data_way0_out_179 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3057 = _T_3056 | _T_2802; // @[Mux.scala 27:72]
  wire  _T_2471 = btb_rd_addr_f == 8'hb4; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_180; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2803 = _T_2471 ? btb_bank0_rd_data_way0_out_180 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3058 = _T_3057 | _T_2803; // @[Mux.scala 27:72]
  wire  _T_2473 = btb_rd_addr_f == 8'hb5; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_181; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2804 = _T_2473 ? btb_bank0_rd_data_way0_out_181 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3059 = _T_3058 | _T_2804; // @[Mux.scala 27:72]
  wire  _T_2475 = btb_rd_addr_f == 8'hb6; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_182; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2805 = _T_2475 ? btb_bank0_rd_data_way0_out_182 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3060 = _T_3059 | _T_2805; // @[Mux.scala 27:72]
  wire  _T_2477 = btb_rd_addr_f == 8'hb7; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_183; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2806 = _T_2477 ? btb_bank0_rd_data_way0_out_183 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3061 = _T_3060 | _T_2806; // @[Mux.scala 27:72]
  wire  _T_2479 = btb_rd_addr_f == 8'hb8; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_184; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2807 = _T_2479 ? btb_bank0_rd_data_way0_out_184 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3062 = _T_3061 | _T_2807; // @[Mux.scala 27:72]
  wire  _T_2481 = btb_rd_addr_f == 8'hb9; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_185; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2808 = _T_2481 ? btb_bank0_rd_data_way0_out_185 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3063 = _T_3062 | _T_2808; // @[Mux.scala 27:72]
  wire  _T_2483 = btb_rd_addr_f == 8'hba; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_186; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2809 = _T_2483 ? btb_bank0_rd_data_way0_out_186 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3064 = _T_3063 | _T_2809; // @[Mux.scala 27:72]
  wire  _T_2485 = btb_rd_addr_f == 8'hbb; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_187; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2810 = _T_2485 ? btb_bank0_rd_data_way0_out_187 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3065 = _T_3064 | _T_2810; // @[Mux.scala 27:72]
  wire  _T_2487 = btb_rd_addr_f == 8'hbc; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_188; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2811 = _T_2487 ? btb_bank0_rd_data_way0_out_188 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3066 = _T_3065 | _T_2811; // @[Mux.scala 27:72]
  wire  _T_2489 = btb_rd_addr_f == 8'hbd; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_189; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2812 = _T_2489 ? btb_bank0_rd_data_way0_out_189 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3067 = _T_3066 | _T_2812; // @[Mux.scala 27:72]
  wire  _T_2491 = btb_rd_addr_f == 8'hbe; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_190; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2813 = _T_2491 ? btb_bank0_rd_data_way0_out_190 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3068 = _T_3067 | _T_2813; // @[Mux.scala 27:72]
  wire  _T_2493 = btb_rd_addr_f == 8'hbf; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_191; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2814 = _T_2493 ? btb_bank0_rd_data_way0_out_191 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3069 = _T_3068 | _T_2814; // @[Mux.scala 27:72]
  wire  _T_2495 = btb_rd_addr_f == 8'hc0; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_192; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2815 = _T_2495 ? btb_bank0_rd_data_way0_out_192 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3070 = _T_3069 | _T_2815; // @[Mux.scala 27:72]
  wire  _T_2497 = btb_rd_addr_f == 8'hc1; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_193; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2816 = _T_2497 ? btb_bank0_rd_data_way0_out_193 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3071 = _T_3070 | _T_2816; // @[Mux.scala 27:72]
  wire  _T_2499 = btb_rd_addr_f == 8'hc2; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_194; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2817 = _T_2499 ? btb_bank0_rd_data_way0_out_194 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3072 = _T_3071 | _T_2817; // @[Mux.scala 27:72]
  wire  _T_2501 = btb_rd_addr_f == 8'hc3; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_195; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2818 = _T_2501 ? btb_bank0_rd_data_way0_out_195 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3073 = _T_3072 | _T_2818; // @[Mux.scala 27:72]
  wire  _T_2503 = btb_rd_addr_f == 8'hc4; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_196; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2819 = _T_2503 ? btb_bank0_rd_data_way0_out_196 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3074 = _T_3073 | _T_2819; // @[Mux.scala 27:72]
  wire  _T_2505 = btb_rd_addr_f == 8'hc5; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_197; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2820 = _T_2505 ? btb_bank0_rd_data_way0_out_197 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3075 = _T_3074 | _T_2820; // @[Mux.scala 27:72]
  wire  _T_2507 = btb_rd_addr_f == 8'hc6; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_198; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2821 = _T_2507 ? btb_bank0_rd_data_way0_out_198 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3076 = _T_3075 | _T_2821; // @[Mux.scala 27:72]
  wire  _T_2509 = btb_rd_addr_f == 8'hc7; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_199; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2822 = _T_2509 ? btb_bank0_rd_data_way0_out_199 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3077 = _T_3076 | _T_2822; // @[Mux.scala 27:72]
  wire  _T_2511 = btb_rd_addr_f == 8'hc8; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_200; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2823 = _T_2511 ? btb_bank0_rd_data_way0_out_200 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3078 = _T_3077 | _T_2823; // @[Mux.scala 27:72]
  wire  _T_2513 = btb_rd_addr_f == 8'hc9; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_201; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2824 = _T_2513 ? btb_bank0_rd_data_way0_out_201 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3079 = _T_3078 | _T_2824; // @[Mux.scala 27:72]
  wire  _T_2515 = btb_rd_addr_f == 8'hca; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_202; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2825 = _T_2515 ? btb_bank0_rd_data_way0_out_202 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3080 = _T_3079 | _T_2825; // @[Mux.scala 27:72]
  wire  _T_2517 = btb_rd_addr_f == 8'hcb; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_203; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2826 = _T_2517 ? btb_bank0_rd_data_way0_out_203 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3081 = _T_3080 | _T_2826; // @[Mux.scala 27:72]
  wire  _T_2519 = btb_rd_addr_f == 8'hcc; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_204; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2827 = _T_2519 ? btb_bank0_rd_data_way0_out_204 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3082 = _T_3081 | _T_2827; // @[Mux.scala 27:72]
  wire  _T_2521 = btb_rd_addr_f == 8'hcd; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_205; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2828 = _T_2521 ? btb_bank0_rd_data_way0_out_205 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3083 = _T_3082 | _T_2828; // @[Mux.scala 27:72]
  wire  _T_2523 = btb_rd_addr_f == 8'hce; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_206; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2829 = _T_2523 ? btb_bank0_rd_data_way0_out_206 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3084 = _T_3083 | _T_2829; // @[Mux.scala 27:72]
  wire  _T_2525 = btb_rd_addr_f == 8'hcf; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_207; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2830 = _T_2525 ? btb_bank0_rd_data_way0_out_207 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3085 = _T_3084 | _T_2830; // @[Mux.scala 27:72]
  wire  _T_2527 = btb_rd_addr_f == 8'hd0; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_208; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2831 = _T_2527 ? btb_bank0_rd_data_way0_out_208 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3086 = _T_3085 | _T_2831; // @[Mux.scala 27:72]
  wire  _T_2529 = btb_rd_addr_f == 8'hd1; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_209; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2832 = _T_2529 ? btb_bank0_rd_data_way0_out_209 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3087 = _T_3086 | _T_2832; // @[Mux.scala 27:72]
  wire  _T_2531 = btb_rd_addr_f == 8'hd2; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_210; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2833 = _T_2531 ? btb_bank0_rd_data_way0_out_210 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3088 = _T_3087 | _T_2833; // @[Mux.scala 27:72]
  wire  _T_2533 = btb_rd_addr_f == 8'hd3; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_211; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2834 = _T_2533 ? btb_bank0_rd_data_way0_out_211 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3089 = _T_3088 | _T_2834; // @[Mux.scala 27:72]
  wire  _T_2535 = btb_rd_addr_f == 8'hd4; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_212; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2835 = _T_2535 ? btb_bank0_rd_data_way0_out_212 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3090 = _T_3089 | _T_2835; // @[Mux.scala 27:72]
  wire  _T_2537 = btb_rd_addr_f == 8'hd5; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_213; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2836 = _T_2537 ? btb_bank0_rd_data_way0_out_213 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3091 = _T_3090 | _T_2836; // @[Mux.scala 27:72]
  wire  _T_2539 = btb_rd_addr_f == 8'hd6; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_214; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2837 = _T_2539 ? btb_bank0_rd_data_way0_out_214 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3092 = _T_3091 | _T_2837; // @[Mux.scala 27:72]
  wire  _T_2541 = btb_rd_addr_f == 8'hd7; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_215; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2838 = _T_2541 ? btb_bank0_rd_data_way0_out_215 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3093 = _T_3092 | _T_2838; // @[Mux.scala 27:72]
  wire  _T_2543 = btb_rd_addr_f == 8'hd8; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_216; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2839 = _T_2543 ? btb_bank0_rd_data_way0_out_216 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3094 = _T_3093 | _T_2839; // @[Mux.scala 27:72]
  wire  _T_2545 = btb_rd_addr_f == 8'hd9; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_217; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2840 = _T_2545 ? btb_bank0_rd_data_way0_out_217 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3095 = _T_3094 | _T_2840; // @[Mux.scala 27:72]
  wire  _T_2547 = btb_rd_addr_f == 8'hda; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_218; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2841 = _T_2547 ? btb_bank0_rd_data_way0_out_218 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3096 = _T_3095 | _T_2841; // @[Mux.scala 27:72]
  wire  _T_2549 = btb_rd_addr_f == 8'hdb; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_219; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2842 = _T_2549 ? btb_bank0_rd_data_way0_out_219 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3097 = _T_3096 | _T_2842; // @[Mux.scala 27:72]
  wire  _T_2551 = btb_rd_addr_f == 8'hdc; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_220; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2843 = _T_2551 ? btb_bank0_rd_data_way0_out_220 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3098 = _T_3097 | _T_2843; // @[Mux.scala 27:72]
  wire  _T_2553 = btb_rd_addr_f == 8'hdd; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_221; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2844 = _T_2553 ? btb_bank0_rd_data_way0_out_221 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3099 = _T_3098 | _T_2844; // @[Mux.scala 27:72]
  wire  _T_2555 = btb_rd_addr_f == 8'hde; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_222; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2845 = _T_2555 ? btb_bank0_rd_data_way0_out_222 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3100 = _T_3099 | _T_2845; // @[Mux.scala 27:72]
  wire  _T_2557 = btb_rd_addr_f == 8'hdf; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_223; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2846 = _T_2557 ? btb_bank0_rd_data_way0_out_223 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3101 = _T_3100 | _T_2846; // @[Mux.scala 27:72]
  wire  _T_2559 = btb_rd_addr_f == 8'he0; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_224; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2847 = _T_2559 ? btb_bank0_rd_data_way0_out_224 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3102 = _T_3101 | _T_2847; // @[Mux.scala 27:72]
  wire  _T_2561 = btb_rd_addr_f == 8'he1; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_225; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2848 = _T_2561 ? btb_bank0_rd_data_way0_out_225 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3103 = _T_3102 | _T_2848; // @[Mux.scala 27:72]
  wire  _T_2563 = btb_rd_addr_f == 8'he2; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_226; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2849 = _T_2563 ? btb_bank0_rd_data_way0_out_226 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3104 = _T_3103 | _T_2849; // @[Mux.scala 27:72]
  wire  _T_2565 = btb_rd_addr_f == 8'he3; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_227; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2850 = _T_2565 ? btb_bank0_rd_data_way0_out_227 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3105 = _T_3104 | _T_2850; // @[Mux.scala 27:72]
  wire  _T_2567 = btb_rd_addr_f == 8'he4; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_228; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2851 = _T_2567 ? btb_bank0_rd_data_way0_out_228 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3106 = _T_3105 | _T_2851; // @[Mux.scala 27:72]
  wire  _T_2569 = btb_rd_addr_f == 8'he5; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_229; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2852 = _T_2569 ? btb_bank0_rd_data_way0_out_229 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3107 = _T_3106 | _T_2852; // @[Mux.scala 27:72]
  wire  _T_2571 = btb_rd_addr_f == 8'he6; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_230; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2853 = _T_2571 ? btb_bank0_rd_data_way0_out_230 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3108 = _T_3107 | _T_2853; // @[Mux.scala 27:72]
  wire  _T_2573 = btb_rd_addr_f == 8'he7; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_231; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2854 = _T_2573 ? btb_bank0_rd_data_way0_out_231 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3109 = _T_3108 | _T_2854; // @[Mux.scala 27:72]
  wire  _T_2575 = btb_rd_addr_f == 8'he8; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_232; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2855 = _T_2575 ? btb_bank0_rd_data_way0_out_232 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3110 = _T_3109 | _T_2855; // @[Mux.scala 27:72]
  wire  _T_2577 = btb_rd_addr_f == 8'he9; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_233; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2856 = _T_2577 ? btb_bank0_rd_data_way0_out_233 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3111 = _T_3110 | _T_2856; // @[Mux.scala 27:72]
  wire  _T_2579 = btb_rd_addr_f == 8'hea; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_234; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2857 = _T_2579 ? btb_bank0_rd_data_way0_out_234 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3112 = _T_3111 | _T_2857; // @[Mux.scala 27:72]
  wire  _T_2581 = btb_rd_addr_f == 8'heb; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_235; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2858 = _T_2581 ? btb_bank0_rd_data_way0_out_235 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3113 = _T_3112 | _T_2858; // @[Mux.scala 27:72]
  wire  _T_2583 = btb_rd_addr_f == 8'hec; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_236; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2859 = _T_2583 ? btb_bank0_rd_data_way0_out_236 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3114 = _T_3113 | _T_2859; // @[Mux.scala 27:72]
  wire  _T_2585 = btb_rd_addr_f == 8'hed; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_237; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2860 = _T_2585 ? btb_bank0_rd_data_way0_out_237 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3115 = _T_3114 | _T_2860; // @[Mux.scala 27:72]
  wire  _T_2587 = btb_rd_addr_f == 8'hee; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_238; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2861 = _T_2587 ? btb_bank0_rd_data_way0_out_238 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3116 = _T_3115 | _T_2861; // @[Mux.scala 27:72]
  wire  _T_2589 = btb_rd_addr_f == 8'hef; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_239; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2862 = _T_2589 ? btb_bank0_rd_data_way0_out_239 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3117 = _T_3116 | _T_2862; // @[Mux.scala 27:72]
  wire  _T_2591 = btb_rd_addr_f == 8'hf0; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_240; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2863 = _T_2591 ? btb_bank0_rd_data_way0_out_240 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3118 = _T_3117 | _T_2863; // @[Mux.scala 27:72]
  wire  _T_2593 = btb_rd_addr_f == 8'hf1; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_241; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2864 = _T_2593 ? btb_bank0_rd_data_way0_out_241 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3119 = _T_3118 | _T_2864; // @[Mux.scala 27:72]
  wire  _T_2595 = btb_rd_addr_f == 8'hf2; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_242; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2865 = _T_2595 ? btb_bank0_rd_data_way0_out_242 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3120 = _T_3119 | _T_2865; // @[Mux.scala 27:72]
  wire  _T_2597 = btb_rd_addr_f == 8'hf3; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_243; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2866 = _T_2597 ? btb_bank0_rd_data_way0_out_243 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3121 = _T_3120 | _T_2866; // @[Mux.scala 27:72]
  wire  _T_2599 = btb_rd_addr_f == 8'hf4; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_244; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2867 = _T_2599 ? btb_bank0_rd_data_way0_out_244 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3122 = _T_3121 | _T_2867; // @[Mux.scala 27:72]
  wire  _T_2601 = btb_rd_addr_f == 8'hf5; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_245; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2868 = _T_2601 ? btb_bank0_rd_data_way0_out_245 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3123 = _T_3122 | _T_2868; // @[Mux.scala 27:72]
  wire  _T_2603 = btb_rd_addr_f == 8'hf6; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_246; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2869 = _T_2603 ? btb_bank0_rd_data_way0_out_246 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3124 = _T_3123 | _T_2869; // @[Mux.scala 27:72]
  wire  _T_2605 = btb_rd_addr_f == 8'hf7; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_247; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2870 = _T_2605 ? btb_bank0_rd_data_way0_out_247 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3125 = _T_3124 | _T_2870; // @[Mux.scala 27:72]
  wire  _T_2607 = btb_rd_addr_f == 8'hf8; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_248; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2871 = _T_2607 ? btb_bank0_rd_data_way0_out_248 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3126 = _T_3125 | _T_2871; // @[Mux.scala 27:72]
  wire  _T_2609 = btb_rd_addr_f == 8'hf9; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_249; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2872 = _T_2609 ? btb_bank0_rd_data_way0_out_249 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3127 = _T_3126 | _T_2872; // @[Mux.scala 27:72]
  wire  _T_2611 = btb_rd_addr_f == 8'hfa; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_250; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2873 = _T_2611 ? btb_bank0_rd_data_way0_out_250 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3128 = _T_3127 | _T_2873; // @[Mux.scala 27:72]
  wire  _T_2613 = btb_rd_addr_f == 8'hfb; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_251; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2874 = _T_2613 ? btb_bank0_rd_data_way0_out_251 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3129 = _T_3128 | _T_2874; // @[Mux.scala 27:72]
  wire  _T_2615 = btb_rd_addr_f == 8'hfc; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_252; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2875 = _T_2615 ? btb_bank0_rd_data_way0_out_252 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3130 = _T_3129 | _T_2875; // @[Mux.scala 27:72]
  wire  _T_2617 = btb_rd_addr_f == 8'hfd; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_253; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2876 = _T_2617 ? btb_bank0_rd_data_way0_out_253 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3131 = _T_3130 | _T_2876; // @[Mux.scala 27:72]
  wire  _T_2619 = btb_rd_addr_f == 8'hfe; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_254; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2877 = _T_2619 ? btb_bank0_rd_data_way0_out_254 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3132 = _T_3131 | _T_2877; // @[Mux.scala 27:72]
  wire  _T_2621 = btb_rd_addr_f == 8'hff; // @[el2_ifu_bp_ctl.scala 430:77]
  reg [21:0] btb_bank0_rd_data_way0_out_255; // @[el2_lib.scala 481:16]
  wire [21:0] _T_2878 = _T_2621 ? btb_bank0_rd_data_way0_out_255 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] btb_bank0_rd_data_way0_f = _T_3132 | _T_2878; // @[Mux.scala 27:72]
  wire [4:0] _T_25 = io_ifc_fetch_addr_f[13:9] ^ io_ifc_fetch_addr_f[18:14]; // @[el2_lib.scala 180:111]
  wire [4:0] fetch_rd_tag_f = _T_25 ^ io_ifc_fetch_addr_f[23:19]; // @[el2_lib.scala 180:111]
  wire  _T_45 = btb_bank0_rd_data_way0_f[21:17] == fetch_rd_tag_f; // @[el2_ifu_bp_ctl.scala 139:97]
  wire  _T_46 = btb_bank0_rd_data_way0_f[0] & _T_45; // @[el2_ifu_bp_ctl.scala 139:55]
  reg  dec_tlu_way_wb_f; // @[el2_ifu_bp_ctl.scala 130:59]
  wire  _T_19 = io_exu_i0_br_index_r == btb_rd_addr_f; // @[el2_ifu_bp_ctl.scala 114:72]
  wire  branch_error_collision_f = dec_tlu_error_wb & _T_19; // @[el2_ifu_bp_ctl.scala 114:51]
  wire  branch_error_bank_conflict_f = branch_error_collision_f & dec_tlu_error_wb; // @[el2_ifu_bp_ctl.scala 118:63]
  wire  _T_47 = dec_tlu_way_wb_f & branch_error_bank_conflict_f; // @[el2_ifu_bp_ctl.scala 140:44]
  wire  _T_48 = ~_T_47; // @[el2_ifu_bp_ctl.scala 140:25]
  wire  _T_49 = _T_46 & _T_48; // @[el2_ifu_bp_ctl.scala 139:117]
  wire  _T_50 = _T_49 & io_ifc_fetch_req_f; // @[el2_ifu_bp_ctl.scala 140:76]
  wire  tag_match_way0_f = _T_50 & _T; // @[el2_ifu_bp_ctl.scala 140:97]
  wire  _T_81 = btb_bank0_rd_data_way0_f[3] ^ btb_bank0_rd_data_way0_f[4]; // @[el2_ifu_bp_ctl.scala 154:91]
  wire  _T_82 = tag_match_way0_f & _T_81; // @[el2_ifu_bp_ctl.scala 154:56]
  wire  _T_86 = ~_T_81; // @[el2_ifu_bp_ctl.scala 155:58]
  wire  _T_87 = tag_match_way0_f & _T_86; // @[el2_ifu_bp_ctl.scala 155:56]
  wire [1:0] tag_match_way0_expanded_f = {_T_82,_T_87}; // @[Cat.scala 29:58]
  wire [21:0] _T_126 = tag_match_way0_expanded_f[1] ? btb_bank0_rd_data_way0_f : 22'h0; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_0; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3647 = _T_2111 ? btb_bank0_rd_data_way1_out_0 : 22'h0; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_1; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3648 = _T_2113 ? btb_bank0_rd_data_way1_out_1 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3903 = _T_3647 | _T_3648; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_2; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3649 = _T_2115 ? btb_bank0_rd_data_way1_out_2 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3904 = _T_3903 | _T_3649; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_3; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3650 = _T_2117 ? btb_bank0_rd_data_way1_out_3 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3905 = _T_3904 | _T_3650; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_4; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3651 = _T_2119 ? btb_bank0_rd_data_way1_out_4 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3906 = _T_3905 | _T_3651; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_5; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3652 = _T_2121 ? btb_bank0_rd_data_way1_out_5 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3907 = _T_3906 | _T_3652; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_6; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3653 = _T_2123 ? btb_bank0_rd_data_way1_out_6 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3908 = _T_3907 | _T_3653; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_7; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3654 = _T_2125 ? btb_bank0_rd_data_way1_out_7 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3909 = _T_3908 | _T_3654; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_8; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3655 = _T_2127 ? btb_bank0_rd_data_way1_out_8 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3910 = _T_3909 | _T_3655; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_9; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3656 = _T_2129 ? btb_bank0_rd_data_way1_out_9 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3911 = _T_3910 | _T_3656; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_10; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3657 = _T_2131 ? btb_bank0_rd_data_way1_out_10 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3912 = _T_3911 | _T_3657; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_11; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3658 = _T_2133 ? btb_bank0_rd_data_way1_out_11 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3913 = _T_3912 | _T_3658; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_12; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3659 = _T_2135 ? btb_bank0_rd_data_way1_out_12 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3914 = _T_3913 | _T_3659; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_13; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3660 = _T_2137 ? btb_bank0_rd_data_way1_out_13 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3915 = _T_3914 | _T_3660; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_14; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3661 = _T_2139 ? btb_bank0_rd_data_way1_out_14 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3916 = _T_3915 | _T_3661; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_15; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3662 = _T_2141 ? btb_bank0_rd_data_way1_out_15 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3917 = _T_3916 | _T_3662; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_16; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3663 = _T_2143 ? btb_bank0_rd_data_way1_out_16 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3918 = _T_3917 | _T_3663; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_17; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3664 = _T_2145 ? btb_bank0_rd_data_way1_out_17 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3919 = _T_3918 | _T_3664; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_18; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3665 = _T_2147 ? btb_bank0_rd_data_way1_out_18 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3920 = _T_3919 | _T_3665; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_19; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3666 = _T_2149 ? btb_bank0_rd_data_way1_out_19 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3921 = _T_3920 | _T_3666; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_20; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3667 = _T_2151 ? btb_bank0_rd_data_way1_out_20 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3922 = _T_3921 | _T_3667; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_21; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3668 = _T_2153 ? btb_bank0_rd_data_way1_out_21 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3923 = _T_3922 | _T_3668; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_22; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3669 = _T_2155 ? btb_bank0_rd_data_way1_out_22 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3924 = _T_3923 | _T_3669; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_23; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3670 = _T_2157 ? btb_bank0_rd_data_way1_out_23 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3925 = _T_3924 | _T_3670; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_24; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3671 = _T_2159 ? btb_bank0_rd_data_way1_out_24 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3926 = _T_3925 | _T_3671; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_25; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3672 = _T_2161 ? btb_bank0_rd_data_way1_out_25 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3927 = _T_3926 | _T_3672; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_26; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3673 = _T_2163 ? btb_bank0_rd_data_way1_out_26 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3928 = _T_3927 | _T_3673; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_27; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3674 = _T_2165 ? btb_bank0_rd_data_way1_out_27 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3929 = _T_3928 | _T_3674; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_28; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3675 = _T_2167 ? btb_bank0_rd_data_way1_out_28 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3930 = _T_3929 | _T_3675; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_29; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3676 = _T_2169 ? btb_bank0_rd_data_way1_out_29 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3931 = _T_3930 | _T_3676; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_30; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3677 = _T_2171 ? btb_bank0_rd_data_way1_out_30 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3932 = _T_3931 | _T_3677; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_31; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3678 = _T_2173 ? btb_bank0_rd_data_way1_out_31 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3933 = _T_3932 | _T_3678; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_32; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3679 = _T_2175 ? btb_bank0_rd_data_way1_out_32 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3934 = _T_3933 | _T_3679; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_33; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3680 = _T_2177 ? btb_bank0_rd_data_way1_out_33 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3935 = _T_3934 | _T_3680; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_34; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3681 = _T_2179 ? btb_bank0_rd_data_way1_out_34 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3936 = _T_3935 | _T_3681; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_35; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3682 = _T_2181 ? btb_bank0_rd_data_way1_out_35 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3937 = _T_3936 | _T_3682; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_36; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3683 = _T_2183 ? btb_bank0_rd_data_way1_out_36 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3938 = _T_3937 | _T_3683; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_37; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3684 = _T_2185 ? btb_bank0_rd_data_way1_out_37 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3939 = _T_3938 | _T_3684; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_38; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3685 = _T_2187 ? btb_bank0_rd_data_way1_out_38 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3940 = _T_3939 | _T_3685; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_39; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3686 = _T_2189 ? btb_bank0_rd_data_way1_out_39 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3941 = _T_3940 | _T_3686; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_40; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3687 = _T_2191 ? btb_bank0_rd_data_way1_out_40 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3942 = _T_3941 | _T_3687; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_41; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3688 = _T_2193 ? btb_bank0_rd_data_way1_out_41 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3943 = _T_3942 | _T_3688; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_42; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3689 = _T_2195 ? btb_bank0_rd_data_way1_out_42 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3944 = _T_3943 | _T_3689; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_43; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3690 = _T_2197 ? btb_bank0_rd_data_way1_out_43 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3945 = _T_3944 | _T_3690; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_44; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3691 = _T_2199 ? btb_bank0_rd_data_way1_out_44 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3946 = _T_3945 | _T_3691; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_45; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3692 = _T_2201 ? btb_bank0_rd_data_way1_out_45 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3947 = _T_3946 | _T_3692; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_46; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3693 = _T_2203 ? btb_bank0_rd_data_way1_out_46 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3948 = _T_3947 | _T_3693; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_47; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3694 = _T_2205 ? btb_bank0_rd_data_way1_out_47 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3949 = _T_3948 | _T_3694; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_48; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3695 = _T_2207 ? btb_bank0_rd_data_way1_out_48 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3950 = _T_3949 | _T_3695; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_49; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3696 = _T_2209 ? btb_bank0_rd_data_way1_out_49 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3951 = _T_3950 | _T_3696; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_50; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3697 = _T_2211 ? btb_bank0_rd_data_way1_out_50 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3952 = _T_3951 | _T_3697; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_51; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3698 = _T_2213 ? btb_bank0_rd_data_way1_out_51 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3953 = _T_3952 | _T_3698; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_52; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3699 = _T_2215 ? btb_bank0_rd_data_way1_out_52 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3954 = _T_3953 | _T_3699; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_53; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3700 = _T_2217 ? btb_bank0_rd_data_way1_out_53 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3955 = _T_3954 | _T_3700; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_54; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3701 = _T_2219 ? btb_bank0_rd_data_way1_out_54 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3956 = _T_3955 | _T_3701; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_55; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3702 = _T_2221 ? btb_bank0_rd_data_way1_out_55 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3957 = _T_3956 | _T_3702; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_56; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3703 = _T_2223 ? btb_bank0_rd_data_way1_out_56 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3958 = _T_3957 | _T_3703; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_57; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3704 = _T_2225 ? btb_bank0_rd_data_way1_out_57 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3959 = _T_3958 | _T_3704; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_58; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3705 = _T_2227 ? btb_bank0_rd_data_way1_out_58 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3960 = _T_3959 | _T_3705; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_59; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3706 = _T_2229 ? btb_bank0_rd_data_way1_out_59 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3961 = _T_3960 | _T_3706; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_60; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3707 = _T_2231 ? btb_bank0_rd_data_way1_out_60 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3962 = _T_3961 | _T_3707; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_61; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3708 = _T_2233 ? btb_bank0_rd_data_way1_out_61 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3963 = _T_3962 | _T_3708; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_62; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3709 = _T_2235 ? btb_bank0_rd_data_way1_out_62 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3964 = _T_3963 | _T_3709; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_63; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3710 = _T_2237 ? btb_bank0_rd_data_way1_out_63 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3965 = _T_3964 | _T_3710; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_64; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3711 = _T_2239 ? btb_bank0_rd_data_way1_out_64 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3966 = _T_3965 | _T_3711; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_65; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3712 = _T_2241 ? btb_bank0_rd_data_way1_out_65 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3967 = _T_3966 | _T_3712; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_66; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3713 = _T_2243 ? btb_bank0_rd_data_way1_out_66 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3968 = _T_3967 | _T_3713; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_67; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3714 = _T_2245 ? btb_bank0_rd_data_way1_out_67 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3969 = _T_3968 | _T_3714; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_68; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3715 = _T_2247 ? btb_bank0_rd_data_way1_out_68 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3970 = _T_3969 | _T_3715; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_69; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3716 = _T_2249 ? btb_bank0_rd_data_way1_out_69 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3971 = _T_3970 | _T_3716; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_70; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3717 = _T_2251 ? btb_bank0_rd_data_way1_out_70 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3972 = _T_3971 | _T_3717; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_71; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3718 = _T_2253 ? btb_bank0_rd_data_way1_out_71 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3973 = _T_3972 | _T_3718; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_72; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3719 = _T_2255 ? btb_bank0_rd_data_way1_out_72 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3974 = _T_3973 | _T_3719; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_73; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3720 = _T_2257 ? btb_bank0_rd_data_way1_out_73 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3975 = _T_3974 | _T_3720; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_74; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3721 = _T_2259 ? btb_bank0_rd_data_way1_out_74 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3976 = _T_3975 | _T_3721; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_75; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3722 = _T_2261 ? btb_bank0_rd_data_way1_out_75 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3977 = _T_3976 | _T_3722; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_76; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3723 = _T_2263 ? btb_bank0_rd_data_way1_out_76 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3978 = _T_3977 | _T_3723; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_77; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3724 = _T_2265 ? btb_bank0_rd_data_way1_out_77 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3979 = _T_3978 | _T_3724; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_78; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3725 = _T_2267 ? btb_bank0_rd_data_way1_out_78 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3980 = _T_3979 | _T_3725; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_79; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3726 = _T_2269 ? btb_bank0_rd_data_way1_out_79 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3981 = _T_3980 | _T_3726; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_80; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3727 = _T_2271 ? btb_bank0_rd_data_way1_out_80 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3982 = _T_3981 | _T_3727; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_81; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3728 = _T_2273 ? btb_bank0_rd_data_way1_out_81 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3983 = _T_3982 | _T_3728; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_82; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3729 = _T_2275 ? btb_bank0_rd_data_way1_out_82 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3984 = _T_3983 | _T_3729; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_83; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3730 = _T_2277 ? btb_bank0_rd_data_way1_out_83 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3985 = _T_3984 | _T_3730; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_84; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3731 = _T_2279 ? btb_bank0_rd_data_way1_out_84 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3986 = _T_3985 | _T_3731; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_85; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3732 = _T_2281 ? btb_bank0_rd_data_way1_out_85 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3987 = _T_3986 | _T_3732; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_86; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3733 = _T_2283 ? btb_bank0_rd_data_way1_out_86 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3988 = _T_3987 | _T_3733; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_87; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3734 = _T_2285 ? btb_bank0_rd_data_way1_out_87 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3989 = _T_3988 | _T_3734; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_88; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3735 = _T_2287 ? btb_bank0_rd_data_way1_out_88 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3990 = _T_3989 | _T_3735; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_89; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3736 = _T_2289 ? btb_bank0_rd_data_way1_out_89 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3991 = _T_3990 | _T_3736; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_90; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3737 = _T_2291 ? btb_bank0_rd_data_way1_out_90 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3992 = _T_3991 | _T_3737; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_91; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3738 = _T_2293 ? btb_bank0_rd_data_way1_out_91 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3993 = _T_3992 | _T_3738; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_92; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3739 = _T_2295 ? btb_bank0_rd_data_way1_out_92 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3994 = _T_3993 | _T_3739; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_93; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3740 = _T_2297 ? btb_bank0_rd_data_way1_out_93 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3995 = _T_3994 | _T_3740; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_94; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3741 = _T_2299 ? btb_bank0_rd_data_way1_out_94 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3996 = _T_3995 | _T_3741; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_95; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3742 = _T_2301 ? btb_bank0_rd_data_way1_out_95 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3997 = _T_3996 | _T_3742; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_96; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3743 = _T_2303 ? btb_bank0_rd_data_way1_out_96 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3998 = _T_3997 | _T_3743; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_97; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3744 = _T_2305 ? btb_bank0_rd_data_way1_out_97 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3999 = _T_3998 | _T_3744; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_98; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3745 = _T_2307 ? btb_bank0_rd_data_way1_out_98 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4000 = _T_3999 | _T_3745; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_99; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3746 = _T_2309 ? btb_bank0_rd_data_way1_out_99 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4001 = _T_4000 | _T_3746; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_100; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3747 = _T_2311 ? btb_bank0_rd_data_way1_out_100 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4002 = _T_4001 | _T_3747; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_101; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3748 = _T_2313 ? btb_bank0_rd_data_way1_out_101 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4003 = _T_4002 | _T_3748; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_102; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3749 = _T_2315 ? btb_bank0_rd_data_way1_out_102 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4004 = _T_4003 | _T_3749; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_103; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3750 = _T_2317 ? btb_bank0_rd_data_way1_out_103 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4005 = _T_4004 | _T_3750; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_104; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3751 = _T_2319 ? btb_bank0_rd_data_way1_out_104 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4006 = _T_4005 | _T_3751; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_105; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3752 = _T_2321 ? btb_bank0_rd_data_way1_out_105 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4007 = _T_4006 | _T_3752; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_106; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3753 = _T_2323 ? btb_bank0_rd_data_way1_out_106 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4008 = _T_4007 | _T_3753; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_107; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3754 = _T_2325 ? btb_bank0_rd_data_way1_out_107 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4009 = _T_4008 | _T_3754; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_108; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3755 = _T_2327 ? btb_bank0_rd_data_way1_out_108 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4010 = _T_4009 | _T_3755; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_109; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3756 = _T_2329 ? btb_bank0_rd_data_way1_out_109 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4011 = _T_4010 | _T_3756; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_110; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3757 = _T_2331 ? btb_bank0_rd_data_way1_out_110 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4012 = _T_4011 | _T_3757; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_111; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3758 = _T_2333 ? btb_bank0_rd_data_way1_out_111 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4013 = _T_4012 | _T_3758; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_112; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3759 = _T_2335 ? btb_bank0_rd_data_way1_out_112 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4014 = _T_4013 | _T_3759; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_113; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3760 = _T_2337 ? btb_bank0_rd_data_way1_out_113 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4015 = _T_4014 | _T_3760; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_114; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3761 = _T_2339 ? btb_bank0_rd_data_way1_out_114 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4016 = _T_4015 | _T_3761; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_115; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3762 = _T_2341 ? btb_bank0_rd_data_way1_out_115 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4017 = _T_4016 | _T_3762; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_116; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3763 = _T_2343 ? btb_bank0_rd_data_way1_out_116 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4018 = _T_4017 | _T_3763; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_117; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3764 = _T_2345 ? btb_bank0_rd_data_way1_out_117 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4019 = _T_4018 | _T_3764; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_118; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3765 = _T_2347 ? btb_bank0_rd_data_way1_out_118 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4020 = _T_4019 | _T_3765; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_119; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3766 = _T_2349 ? btb_bank0_rd_data_way1_out_119 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4021 = _T_4020 | _T_3766; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_120; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3767 = _T_2351 ? btb_bank0_rd_data_way1_out_120 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4022 = _T_4021 | _T_3767; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_121; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3768 = _T_2353 ? btb_bank0_rd_data_way1_out_121 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4023 = _T_4022 | _T_3768; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_122; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3769 = _T_2355 ? btb_bank0_rd_data_way1_out_122 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4024 = _T_4023 | _T_3769; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_123; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3770 = _T_2357 ? btb_bank0_rd_data_way1_out_123 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4025 = _T_4024 | _T_3770; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_124; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3771 = _T_2359 ? btb_bank0_rd_data_way1_out_124 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4026 = _T_4025 | _T_3771; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_125; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3772 = _T_2361 ? btb_bank0_rd_data_way1_out_125 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4027 = _T_4026 | _T_3772; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_126; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3773 = _T_2363 ? btb_bank0_rd_data_way1_out_126 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4028 = _T_4027 | _T_3773; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_127; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3774 = _T_2365 ? btb_bank0_rd_data_way1_out_127 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4029 = _T_4028 | _T_3774; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_128; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3775 = _T_2367 ? btb_bank0_rd_data_way1_out_128 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4030 = _T_4029 | _T_3775; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_129; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3776 = _T_2369 ? btb_bank0_rd_data_way1_out_129 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4031 = _T_4030 | _T_3776; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_130; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3777 = _T_2371 ? btb_bank0_rd_data_way1_out_130 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4032 = _T_4031 | _T_3777; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_131; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3778 = _T_2373 ? btb_bank0_rd_data_way1_out_131 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4033 = _T_4032 | _T_3778; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_132; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3779 = _T_2375 ? btb_bank0_rd_data_way1_out_132 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4034 = _T_4033 | _T_3779; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_133; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3780 = _T_2377 ? btb_bank0_rd_data_way1_out_133 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4035 = _T_4034 | _T_3780; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_134; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3781 = _T_2379 ? btb_bank0_rd_data_way1_out_134 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4036 = _T_4035 | _T_3781; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_135; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3782 = _T_2381 ? btb_bank0_rd_data_way1_out_135 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4037 = _T_4036 | _T_3782; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_136; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3783 = _T_2383 ? btb_bank0_rd_data_way1_out_136 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4038 = _T_4037 | _T_3783; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_137; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3784 = _T_2385 ? btb_bank0_rd_data_way1_out_137 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4039 = _T_4038 | _T_3784; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_138; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3785 = _T_2387 ? btb_bank0_rd_data_way1_out_138 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4040 = _T_4039 | _T_3785; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_139; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3786 = _T_2389 ? btb_bank0_rd_data_way1_out_139 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4041 = _T_4040 | _T_3786; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_140; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3787 = _T_2391 ? btb_bank0_rd_data_way1_out_140 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4042 = _T_4041 | _T_3787; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_141; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3788 = _T_2393 ? btb_bank0_rd_data_way1_out_141 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4043 = _T_4042 | _T_3788; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_142; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3789 = _T_2395 ? btb_bank0_rd_data_way1_out_142 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4044 = _T_4043 | _T_3789; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_143; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3790 = _T_2397 ? btb_bank0_rd_data_way1_out_143 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4045 = _T_4044 | _T_3790; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_144; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3791 = _T_2399 ? btb_bank0_rd_data_way1_out_144 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4046 = _T_4045 | _T_3791; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_145; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3792 = _T_2401 ? btb_bank0_rd_data_way1_out_145 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4047 = _T_4046 | _T_3792; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_146; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3793 = _T_2403 ? btb_bank0_rd_data_way1_out_146 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4048 = _T_4047 | _T_3793; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_147; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3794 = _T_2405 ? btb_bank0_rd_data_way1_out_147 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4049 = _T_4048 | _T_3794; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_148; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3795 = _T_2407 ? btb_bank0_rd_data_way1_out_148 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4050 = _T_4049 | _T_3795; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_149; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3796 = _T_2409 ? btb_bank0_rd_data_way1_out_149 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4051 = _T_4050 | _T_3796; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_150; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3797 = _T_2411 ? btb_bank0_rd_data_way1_out_150 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4052 = _T_4051 | _T_3797; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_151; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3798 = _T_2413 ? btb_bank0_rd_data_way1_out_151 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4053 = _T_4052 | _T_3798; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_152; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3799 = _T_2415 ? btb_bank0_rd_data_way1_out_152 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4054 = _T_4053 | _T_3799; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_153; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3800 = _T_2417 ? btb_bank0_rd_data_way1_out_153 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4055 = _T_4054 | _T_3800; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_154; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3801 = _T_2419 ? btb_bank0_rd_data_way1_out_154 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4056 = _T_4055 | _T_3801; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_155; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3802 = _T_2421 ? btb_bank0_rd_data_way1_out_155 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4057 = _T_4056 | _T_3802; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_156; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3803 = _T_2423 ? btb_bank0_rd_data_way1_out_156 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4058 = _T_4057 | _T_3803; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_157; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3804 = _T_2425 ? btb_bank0_rd_data_way1_out_157 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4059 = _T_4058 | _T_3804; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_158; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3805 = _T_2427 ? btb_bank0_rd_data_way1_out_158 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4060 = _T_4059 | _T_3805; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_159; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3806 = _T_2429 ? btb_bank0_rd_data_way1_out_159 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4061 = _T_4060 | _T_3806; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_160; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3807 = _T_2431 ? btb_bank0_rd_data_way1_out_160 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4062 = _T_4061 | _T_3807; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_161; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3808 = _T_2433 ? btb_bank0_rd_data_way1_out_161 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4063 = _T_4062 | _T_3808; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_162; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3809 = _T_2435 ? btb_bank0_rd_data_way1_out_162 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4064 = _T_4063 | _T_3809; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_163; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3810 = _T_2437 ? btb_bank0_rd_data_way1_out_163 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4065 = _T_4064 | _T_3810; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_164; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3811 = _T_2439 ? btb_bank0_rd_data_way1_out_164 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4066 = _T_4065 | _T_3811; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_165; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3812 = _T_2441 ? btb_bank0_rd_data_way1_out_165 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4067 = _T_4066 | _T_3812; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_166; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3813 = _T_2443 ? btb_bank0_rd_data_way1_out_166 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4068 = _T_4067 | _T_3813; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_167; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3814 = _T_2445 ? btb_bank0_rd_data_way1_out_167 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4069 = _T_4068 | _T_3814; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_168; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3815 = _T_2447 ? btb_bank0_rd_data_way1_out_168 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4070 = _T_4069 | _T_3815; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_169; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3816 = _T_2449 ? btb_bank0_rd_data_way1_out_169 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4071 = _T_4070 | _T_3816; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_170; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3817 = _T_2451 ? btb_bank0_rd_data_way1_out_170 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4072 = _T_4071 | _T_3817; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_171; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3818 = _T_2453 ? btb_bank0_rd_data_way1_out_171 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4073 = _T_4072 | _T_3818; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_172; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3819 = _T_2455 ? btb_bank0_rd_data_way1_out_172 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4074 = _T_4073 | _T_3819; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_173; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3820 = _T_2457 ? btb_bank0_rd_data_way1_out_173 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4075 = _T_4074 | _T_3820; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_174; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3821 = _T_2459 ? btb_bank0_rd_data_way1_out_174 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4076 = _T_4075 | _T_3821; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_175; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3822 = _T_2461 ? btb_bank0_rd_data_way1_out_175 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4077 = _T_4076 | _T_3822; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_176; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3823 = _T_2463 ? btb_bank0_rd_data_way1_out_176 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4078 = _T_4077 | _T_3823; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_177; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3824 = _T_2465 ? btb_bank0_rd_data_way1_out_177 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4079 = _T_4078 | _T_3824; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_178; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3825 = _T_2467 ? btb_bank0_rd_data_way1_out_178 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4080 = _T_4079 | _T_3825; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_179; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3826 = _T_2469 ? btb_bank0_rd_data_way1_out_179 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4081 = _T_4080 | _T_3826; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_180; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3827 = _T_2471 ? btb_bank0_rd_data_way1_out_180 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4082 = _T_4081 | _T_3827; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_181; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3828 = _T_2473 ? btb_bank0_rd_data_way1_out_181 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4083 = _T_4082 | _T_3828; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_182; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3829 = _T_2475 ? btb_bank0_rd_data_way1_out_182 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4084 = _T_4083 | _T_3829; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_183; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3830 = _T_2477 ? btb_bank0_rd_data_way1_out_183 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4085 = _T_4084 | _T_3830; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_184; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3831 = _T_2479 ? btb_bank0_rd_data_way1_out_184 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4086 = _T_4085 | _T_3831; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_185; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3832 = _T_2481 ? btb_bank0_rd_data_way1_out_185 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4087 = _T_4086 | _T_3832; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_186; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3833 = _T_2483 ? btb_bank0_rd_data_way1_out_186 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4088 = _T_4087 | _T_3833; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_187; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3834 = _T_2485 ? btb_bank0_rd_data_way1_out_187 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4089 = _T_4088 | _T_3834; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_188; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3835 = _T_2487 ? btb_bank0_rd_data_way1_out_188 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4090 = _T_4089 | _T_3835; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_189; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3836 = _T_2489 ? btb_bank0_rd_data_way1_out_189 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4091 = _T_4090 | _T_3836; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_190; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3837 = _T_2491 ? btb_bank0_rd_data_way1_out_190 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4092 = _T_4091 | _T_3837; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_191; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3838 = _T_2493 ? btb_bank0_rd_data_way1_out_191 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4093 = _T_4092 | _T_3838; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_192; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3839 = _T_2495 ? btb_bank0_rd_data_way1_out_192 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4094 = _T_4093 | _T_3839; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_193; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3840 = _T_2497 ? btb_bank0_rd_data_way1_out_193 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4095 = _T_4094 | _T_3840; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_194; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3841 = _T_2499 ? btb_bank0_rd_data_way1_out_194 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4096 = _T_4095 | _T_3841; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_195; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3842 = _T_2501 ? btb_bank0_rd_data_way1_out_195 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4097 = _T_4096 | _T_3842; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_196; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3843 = _T_2503 ? btb_bank0_rd_data_way1_out_196 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4098 = _T_4097 | _T_3843; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_197; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3844 = _T_2505 ? btb_bank0_rd_data_way1_out_197 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4099 = _T_4098 | _T_3844; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_198; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3845 = _T_2507 ? btb_bank0_rd_data_way1_out_198 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4100 = _T_4099 | _T_3845; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_199; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3846 = _T_2509 ? btb_bank0_rd_data_way1_out_199 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4101 = _T_4100 | _T_3846; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_200; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3847 = _T_2511 ? btb_bank0_rd_data_way1_out_200 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4102 = _T_4101 | _T_3847; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_201; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3848 = _T_2513 ? btb_bank0_rd_data_way1_out_201 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4103 = _T_4102 | _T_3848; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_202; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3849 = _T_2515 ? btb_bank0_rd_data_way1_out_202 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4104 = _T_4103 | _T_3849; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_203; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3850 = _T_2517 ? btb_bank0_rd_data_way1_out_203 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4105 = _T_4104 | _T_3850; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_204; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3851 = _T_2519 ? btb_bank0_rd_data_way1_out_204 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4106 = _T_4105 | _T_3851; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_205; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3852 = _T_2521 ? btb_bank0_rd_data_way1_out_205 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4107 = _T_4106 | _T_3852; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_206; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3853 = _T_2523 ? btb_bank0_rd_data_way1_out_206 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4108 = _T_4107 | _T_3853; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_207; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3854 = _T_2525 ? btb_bank0_rd_data_way1_out_207 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4109 = _T_4108 | _T_3854; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_208; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3855 = _T_2527 ? btb_bank0_rd_data_way1_out_208 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4110 = _T_4109 | _T_3855; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_209; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3856 = _T_2529 ? btb_bank0_rd_data_way1_out_209 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4111 = _T_4110 | _T_3856; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_210; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3857 = _T_2531 ? btb_bank0_rd_data_way1_out_210 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4112 = _T_4111 | _T_3857; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_211; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3858 = _T_2533 ? btb_bank0_rd_data_way1_out_211 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4113 = _T_4112 | _T_3858; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_212; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3859 = _T_2535 ? btb_bank0_rd_data_way1_out_212 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4114 = _T_4113 | _T_3859; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_213; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3860 = _T_2537 ? btb_bank0_rd_data_way1_out_213 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4115 = _T_4114 | _T_3860; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_214; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3861 = _T_2539 ? btb_bank0_rd_data_way1_out_214 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4116 = _T_4115 | _T_3861; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_215; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3862 = _T_2541 ? btb_bank0_rd_data_way1_out_215 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4117 = _T_4116 | _T_3862; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_216; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3863 = _T_2543 ? btb_bank0_rd_data_way1_out_216 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4118 = _T_4117 | _T_3863; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_217; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3864 = _T_2545 ? btb_bank0_rd_data_way1_out_217 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4119 = _T_4118 | _T_3864; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_218; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3865 = _T_2547 ? btb_bank0_rd_data_way1_out_218 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4120 = _T_4119 | _T_3865; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_219; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3866 = _T_2549 ? btb_bank0_rd_data_way1_out_219 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4121 = _T_4120 | _T_3866; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_220; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3867 = _T_2551 ? btb_bank0_rd_data_way1_out_220 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4122 = _T_4121 | _T_3867; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_221; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3868 = _T_2553 ? btb_bank0_rd_data_way1_out_221 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4123 = _T_4122 | _T_3868; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_222; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3869 = _T_2555 ? btb_bank0_rd_data_way1_out_222 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4124 = _T_4123 | _T_3869; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_223; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3870 = _T_2557 ? btb_bank0_rd_data_way1_out_223 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4125 = _T_4124 | _T_3870; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_224; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3871 = _T_2559 ? btb_bank0_rd_data_way1_out_224 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4126 = _T_4125 | _T_3871; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_225; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3872 = _T_2561 ? btb_bank0_rd_data_way1_out_225 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4127 = _T_4126 | _T_3872; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_226; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3873 = _T_2563 ? btb_bank0_rd_data_way1_out_226 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4128 = _T_4127 | _T_3873; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_227; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3874 = _T_2565 ? btb_bank0_rd_data_way1_out_227 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4129 = _T_4128 | _T_3874; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_228; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3875 = _T_2567 ? btb_bank0_rd_data_way1_out_228 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4130 = _T_4129 | _T_3875; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_229; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3876 = _T_2569 ? btb_bank0_rd_data_way1_out_229 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4131 = _T_4130 | _T_3876; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_230; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3877 = _T_2571 ? btb_bank0_rd_data_way1_out_230 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4132 = _T_4131 | _T_3877; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_231; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3878 = _T_2573 ? btb_bank0_rd_data_way1_out_231 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4133 = _T_4132 | _T_3878; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_232; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3879 = _T_2575 ? btb_bank0_rd_data_way1_out_232 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4134 = _T_4133 | _T_3879; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_233; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3880 = _T_2577 ? btb_bank0_rd_data_way1_out_233 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4135 = _T_4134 | _T_3880; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_234; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3881 = _T_2579 ? btb_bank0_rd_data_way1_out_234 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4136 = _T_4135 | _T_3881; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_235; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3882 = _T_2581 ? btb_bank0_rd_data_way1_out_235 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4137 = _T_4136 | _T_3882; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_236; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3883 = _T_2583 ? btb_bank0_rd_data_way1_out_236 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4138 = _T_4137 | _T_3883; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_237; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3884 = _T_2585 ? btb_bank0_rd_data_way1_out_237 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4139 = _T_4138 | _T_3884; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_238; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3885 = _T_2587 ? btb_bank0_rd_data_way1_out_238 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4140 = _T_4139 | _T_3885; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_239; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3886 = _T_2589 ? btb_bank0_rd_data_way1_out_239 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4141 = _T_4140 | _T_3886; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_240; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3887 = _T_2591 ? btb_bank0_rd_data_way1_out_240 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4142 = _T_4141 | _T_3887; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_241; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3888 = _T_2593 ? btb_bank0_rd_data_way1_out_241 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4143 = _T_4142 | _T_3888; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_242; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3889 = _T_2595 ? btb_bank0_rd_data_way1_out_242 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4144 = _T_4143 | _T_3889; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_243; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3890 = _T_2597 ? btb_bank0_rd_data_way1_out_243 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4145 = _T_4144 | _T_3890; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_244; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3891 = _T_2599 ? btb_bank0_rd_data_way1_out_244 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4146 = _T_4145 | _T_3891; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_245; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3892 = _T_2601 ? btb_bank0_rd_data_way1_out_245 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4147 = _T_4146 | _T_3892; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_246; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3893 = _T_2603 ? btb_bank0_rd_data_way1_out_246 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4148 = _T_4147 | _T_3893; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_247; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3894 = _T_2605 ? btb_bank0_rd_data_way1_out_247 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4149 = _T_4148 | _T_3894; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_248; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3895 = _T_2607 ? btb_bank0_rd_data_way1_out_248 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4150 = _T_4149 | _T_3895; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_249; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3896 = _T_2609 ? btb_bank0_rd_data_way1_out_249 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4151 = _T_4150 | _T_3896; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_250; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3897 = _T_2611 ? btb_bank0_rd_data_way1_out_250 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4152 = _T_4151 | _T_3897; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_251; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3898 = _T_2613 ? btb_bank0_rd_data_way1_out_251 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4153 = _T_4152 | _T_3898; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_252; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3899 = _T_2615 ? btb_bank0_rd_data_way1_out_252 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4154 = _T_4153 | _T_3899; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_253; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3900 = _T_2617 ? btb_bank0_rd_data_way1_out_253 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4155 = _T_4154 | _T_3900; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_254; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3901 = _T_2619 ? btb_bank0_rd_data_way1_out_254 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4156 = _T_4155 | _T_3901; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_255; // @[el2_lib.scala 481:16]
  wire [21:0] _T_3902 = _T_2621 ? btb_bank0_rd_data_way1_out_255 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] btb_bank0_rd_data_way1_f = _T_4156 | _T_3902; // @[Mux.scala 27:72]
  wire  _T_54 = btb_bank0_rd_data_way1_f[21:17] == fetch_rd_tag_f; // @[el2_ifu_bp_ctl.scala 143:97]
  wire  _T_55 = btb_bank0_rd_data_way1_f[0] & _T_54; // @[el2_ifu_bp_ctl.scala 143:55]
  wire  _T_58 = _T_55 & _T_48; // @[el2_ifu_bp_ctl.scala 143:117]
  wire  _T_59 = _T_58 & io_ifc_fetch_req_f; // @[el2_ifu_bp_ctl.scala 144:76]
  wire  tag_match_way1_f = _T_59 & _T; // @[el2_ifu_bp_ctl.scala 144:97]
  wire  _T_90 = btb_bank0_rd_data_way1_f[3] ^ btb_bank0_rd_data_way1_f[4]; // @[el2_ifu_bp_ctl.scala 157:91]
  wire  _T_91 = tag_match_way1_f & _T_90; // @[el2_ifu_bp_ctl.scala 157:56]
  wire  _T_95 = ~_T_90; // @[el2_ifu_bp_ctl.scala 158:58]
  wire  _T_96 = tag_match_way1_f & _T_95; // @[el2_ifu_bp_ctl.scala 158:56]
  wire [1:0] tag_match_way1_expanded_f = {_T_91,_T_96}; // @[Cat.scala 29:58]
  wire [21:0] _T_127 = tag_match_way1_expanded_f[1] ? btb_bank0_rd_data_way1_f : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] btb_bank0o_rd_data_f = _T_126 | _T_127; // @[Mux.scala 27:72]
  wire [21:0] _T_145 = _T_143 ? btb_bank0o_rd_data_f : 22'h0; // @[Mux.scala 27:72]
  wire  _T_4159 = btb_rd_addr_p1_f == 8'h0; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4671 = _T_4159 ? btb_bank0_rd_data_way0_out_0 : 22'h0; // @[Mux.scala 27:72]
  wire  _T_4161 = btb_rd_addr_p1_f == 8'h1; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4672 = _T_4161 ? btb_bank0_rd_data_way0_out_1 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4927 = _T_4671 | _T_4672; // @[Mux.scala 27:72]
  wire  _T_4163 = btb_rd_addr_p1_f == 8'h2; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4673 = _T_4163 ? btb_bank0_rd_data_way0_out_2 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4928 = _T_4927 | _T_4673; // @[Mux.scala 27:72]
  wire  _T_4165 = btb_rd_addr_p1_f == 8'h3; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4674 = _T_4165 ? btb_bank0_rd_data_way0_out_3 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4929 = _T_4928 | _T_4674; // @[Mux.scala 27:72]
  wire  _T_4167 = btb_rd_addr_p1_f == 8'h4; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4675 = _T_4167 ? btb_bank0_rd_data_way0_out_4 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4930 = _T_4929 | _T_4675; // @[Mux.scala 27:72]
  wire  _T_4169 = btb_rd_addr_p1_f == 8'h5; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4676 = _T_4169 ? btb_bank0_rd_data_way0_out_5 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4931 = _T_4930 | _T_4676; // @[Mux.scala 27:72]
  wire  _T_4171 = btb_rd_addr_p1_f == 8'h6; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4677 = _T_4171 ? btb_bank0_rd_data_way0_out_6 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4932 = _T_4931 | _T_4677; // @[Mux.scala 27:72]
  wire  _T_4173 = btb_rd_addr_p1_f == 8'h7; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4678 = _T_4173 ? btb_bank0_rd_data_way0_out_7 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4933 = _T_4932 | _T_4678; // @[Mux.scala 27:72]
  wire  _T_4175 = btb_rd_addr_p1_f == 8'h8; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4679 = _T_4175 ? btb_bank0_rd_data_way0_out_8 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4934 = _T_4933 | _T_4679; // @[Mux.scala 27:72]
  wire  _T_4177 = btb_rd_addr_p1_f == 8'h9; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4680 = _T_4177 ? btb_bank0_rd_data_way0_out_9 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4935 = _T_4934 | _T_4680; // @[Mux.scala 27:72]
  wire  _T_4179 = btb_rd_addr_p1_f == 8'ha; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4681 = _T_4179 ? btb_bank0_rd_data_way0_out_10 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4936 = _T_4935 | _T_4681; // @[Mux.scala 27:72]
  wire  _T_4181 = btb_rd_addr_p1_f == 8'hb; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4682 = _T_4181 ? btb_bank0_rd_data_way0_out_11 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4937 = _T_4936 | _T_4682; // @[Mux.scala 27:72]
  wire  _T_4183 = btb_rd_addr_p1_f == 8'hc; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4683 = _T_4183 ? btb_bank0_rd_data_way0_out_12 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4938 = _T_4937 | _T_4683; // @[Mux.scala 27:72]
  wire  _T_4185 = btb_rd_addr_p1_f == 8'hd; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4684 = _T_4185 ? btb_bank0_rd_data_way0_out_13 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4939 = _T_4938 | _T_4684; // @[Mux.scala 27:72]
  wire  _T_4187 = btb_rd_addr_p1_f == 8'he; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4685 = _T_4187 ? btb_bank0_rd_data_way0_out_14 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4940 = _T_4939 | _T_4685; // @[Mux.scala 27:72]
  wire  _T_4189 = btb_rd_addr_p1_f == 8'hf; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4686 = _T_4189 ? btb_bank0_rd_data_way0_out_15 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4941 = _T_4940 | _T_4686; // @[Mux.scala 27:72]
  wire  _T_4191 = btb_rd_addr_p1_f == 8'h10; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4687 = _T_4191 ? btb_bank0_rd_data_way0_out_16 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4942 = _T_4941 | _T_4687; // @[Mux.scala 27:72]
  wire  _T_4193 = btb_rd_addr_p1_f == 8'h11; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4688 = _T_4193 ? btb_bank0_rd_data_way0_out_17 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4943 = _T_4942 | _T_4688; // @[Mux.scala 27:72]
  wire  _T_4195 = btb_rd_addr_p1_f == 8'h12; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4689 = _T_4195 ? btb_bank0_rd_data_way0_out_18 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4944 = _T_4943 | _T_4689; // @[Mux.scala 27:72]
  wire  _T_4197 = btb_rd_addr_p1_f == 8'h13; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4690 = _T_4197 ? btb_bank0_rd_data_way0_out_19 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4945 = _T_4944 | _T_4690; // @[Mux.scala 27:72]
  wire  _T_4199 = btb_rd_addr_p1_f == 8'h14; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4691 = _T_4199 ? btb_bank0_rd_data_way0_out_20 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4946 = _T_4945 | _T_4691; // @[Mux.scala 27:72]
  wire  _T_4201 = btb_rd_addr_p1_f == 8'h15; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4692 = _T_4201 ? btb_bank0_rd_data_way0_out_21 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4947 = _T_4946 | _T_4692; // @[Mux.scala 27:72]
  wire  _T_4203 = btb_rd_addr_p1_f == 8'h16; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4693 = _T_4203 ? btb_bank0_rd_data_way0_out_22 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4948 = _T_4947 | _T_4693; // @[Mux.scala 27:72]
  wire  _T_4205 = btb_rd_addr_p1_f == 8'h17; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4694 = _T_4205 ? btb_bank0_rd_data_way0_out_23 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4949 = _T_4948 | _T_4694; // @[Mux.scala 27:72]
  wire  _T_4207 = btb_rd_addr_p1_f == 8'h18; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4695 = _T_4207 ? btb_bank0_rd_data_way0_out_24 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4950 = _T_4949 | _T_4695; // @[Mux.scala 27:72]
  wire  _T_4209 = btb_rd_addr_p1_f == 8'h19; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4696 = _T_4209 ? btb_bank0_rd_data_way0_out_25 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4951 = _T_4950 | _T_4696; // @[Mux.scala 27:72]
  wire  _T_4211 = btb_rd_addr_p1_f == 8'h1a; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4697 = _T_4211 ? btb_bank0_rd_data_way0_out_26 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4952 = _T_4951 | _T_4697; // @[Mux.scala 27:72]
  wire  _T_4213 = btb_rd_addr_p1_f == 8'h1b; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4698 = _T_4213 ? btb_bank0_rd_data_way0_out_27 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4953 = _T_4952 | _T_4698; // @[Mux.scala 27:72]
  wire  _T_4215 = btb_rd_addr_p1_f == 8'h1c; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4699 = _T_4215 ? btb_bank0_rd_data_way0_out_28 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4954 = _T_4953 | _T_4699; // @[Mux.scala 27:72]
  wire  _T_4217 = btb_rd_addr_p1_f == 8'h1d; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4700 = _T_4217 ? btb_bank0_rd_data_way0_out_29 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4955 = _T_4954 | _T_4700; // @[Mux.scala 27:72]
  wire  _T_4219 = btb_rd_addr_p1_f == 8'h1e; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4701 = _T_4219 ? btb_bank0_rd_data_way0_out_30 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4956 = _T_4955 | _T_4701; // @[Mux.scala 27:72]
  wire  _T_4221 = btb_rd_addr_p1_f == 8'h1f; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4702 = _T_4221 ? btb_bank0_rd_data_way0_out_31 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4957 = _T_4956 | _T_4702; // @[Mux.scala 27:72]
  wire  _T_4223 = btb_rd_addr_p1_f == 8'h20; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4703 = _T_4223 ? btb_bank0_rd_data_way0_out_32 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4958 = _T_4957 | _T_4703; // @[Mux.scala 27:72]
  wire  _T_4225 = btb_rd_addr_p1_f == 8'h21; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4704 = _T_4225 ? btb_bank0_rd_data_way0_out_33 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4959 = _T_4958 | _T_4704; // @[Mux.scala 27:72]
  wire  _T_4227 = btb_rd_addr_p1_f == 8'h22; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4705 = _T_4227 ? btb_bank0_rd_data_way0_out_34 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4960 = _T_4959 | _T_4705; // @[Mux.scala 27:72]
  wire  _T_4229 = btb_rd_addr_p1_f == 8'h23; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4706 = _T_4229 ? btb_bank0_rd_data_way0_out_35 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4961 = _T_4960 | _T_4706; // @[Mux.scala 27:72]
  wire  _T_4231 = btb_rd_addr_p1_f == 8'h24; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4707 = _T_4231 ? btb_bank0_rd_data_way0_out_36 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4962 = _T_4961 | _T_4707; // @[Mux.scala 27:72]
  wire  _T_4233 = btb_rd_addr_p1_f == 8'h25; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4708 = _T_4233 ? btb_bank0_rd_data_way0_out_37 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4963 = _T_4962 | _T_4708; // @[Mux.scala 27:72]
  wire  _T_4235 = btb_rd_addr_p1_f == 8'h26; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4709 = _T_4235 ? btb_bank0_rd_data_way0_out_38 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4964 = _T_4963 | _T_4709; // @[Mux.scala 27:72]
  wire  _T_4237 = btb_rd_addr_p1_f == 8'h27; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4710 = _T_4237 ? btb_bank0_rd_data_way0_out_39 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4965 = _T_4964 | _T_4710; // @[Mux.scala 27:72]
  wire  _T_4239 = btb_rd_addr_p1_f == 8'h28; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4711 = _T_4239 ? btb_bank0_rd_data_way0_out_40 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4966 = _T_4965 | _T_4711; // @[Mux.scala 27:72]
  wire  _T_4241 = btb_rd_addr_p1_f == 8'h29; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4712 = _T_4241 ? btb_bank0_rd_data_way0_out_41 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4967 = _T_4966 | _T_4712; // @[Mux.scala 27:72]
  wire  _T_4243 = btb_rd_addr_p1_f == 8'h2a; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4713 = _T_4243 ? btb_bank0_rd_data_way0_out_42 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4968 = _T_4967 | _T_4713; // @[Mux.scala 27:72]
  wire  _T_4245 = btb_rd_addr_p1_f == 8'h2b; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4714 = _T_4245 ? btb_bank0_rd_data_way0_out_43 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4969 = _T_4968 | _T_4714; // @[Mux.scala 27:72]
  wire  _T_4247 = btb_rd_addr_p1_f == 8'h2c; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4715 = _T_4247 ? btb_bank0_rd_data_way0_out_44 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4970 = _T_4969 | _T_4715; // @[Mux.scala 27:72]
  wire  _T_4249 = btb_rd_addr_p1_f == 8'h2d; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4716 = _T_4249 ? btb_bank0_rd_data_way0_out_45 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4971 = _T_4970 | _T_4716; // @[Mux.scala 27:72]
  wire  _T_4251 = btb_rd_addr_p1_f == 8'h2e; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4717 = _T_4251 ? btb_bank0_rd_data_way0_out_46 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4972 = _T_4971 | _T_4717; // @[Mux.scala 27:72]
  wire  _T_4253 = btb_rd_addr_p1_f == 8'h2f; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4718 = _T_4253 ? btb_bank0_rd_data_way0_out_47 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4973 = _T_4972 | _T_4718; // @[Mux.scala 27:72]
  wire  _T_4255 = btb_rd_addr_p1_f == 8'h30; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4719 = _T_4255 ? btb_bank0_rd_data_way0_out_48 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4974 = _T_4973 | _T_4719; // @[Mux.scala 27:72]
  wire  _T_4257 = btb_rd_addr_p1_f == 8'h31; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4720 = _T_4257 ? btb_bank0_rd_data_way0_out_49 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4975 = _T_4974 | _T_4720; // @[Mux.scala 27:72]
  wire  _T_4259 = btb_rd_addr_p1_f == 8'h32; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4721 = _T_4259 ? btb_bank0_rd_data_way0_out_50 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4976 = _T_4975 | _T_4721; // @[Mux.scala 27:72]
  wire  _T_4261 = btb_rd_addr_p1_f == 8'h33; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4722 = _T_4261 ? btb_bank0_rd_data_way0_out_51 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4977 = _T_4976 | _T_4722; // @[Mux.scala 27:72]
  wire  _T_4263 = btb_rd_addr_p1_f == 8'h34; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4723 = _T_4263 ? btb_bank0_rd_data_way0_out_52 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4978 = _T_4977 | _T_4723; // @[Mux.scala 27:72]
  wire  _T_4265 = btb_rd_addr_p1_f == 8'h35; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4724 = _T_4265 ? btb_bank0_rd_data_way0_out_53 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4979 = _T_4978 | _T_4724; // @[Mux.scala 27:72]
  wire  _T_4267 = btb_rd_addr_p1_f == 8'h36; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4725 = _T_4267 ? btb_bank0_rd_data_way0_out_54 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4980 = _T_4979 | _T_4725; // @[Mux.scala 27:72]
  wire  _T_4269 = btb_rd_addr_p1_f == 8'h37; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4726 = _T_4269 ? btb_bank0_rd_data_way0_out_55 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4981 = _T_4980 | _T_4726; // @[Mux.scala 27:72]
  wire  _T_4271 = btb_rd_addr_p1_f == 8'h38; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4727 = _T_4271 ? btb_bank0_rd_data_way0_out_56 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4982 = _T_4981 | _T_4727; // @[Mux.scala 27:72]
  wire  _T_4273 = btb_rd_addr_p1_f == 8'h39; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4728 = _T_4273 ? btb_bank0_rd_data_way0_out_57 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4983 = _T_4982 | _T_4728; // @[Mux.scala 27:72]
  wire  _T_4275 = btb_rd_addr_p1_f == 8'h3a; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4729 = _T_4275 ? btb_bank0_rd_data_way0_out_58 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4984 = _T_4983 | _T_4729; // @[Mux.scala 27:72]
  wire  _T_4277 = btb_rd_addr_p1_f == 8'h3b; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4730 = _T_4277 ? btb_bank0_rd_data_way0_out_59 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4985 = _T_4984 | _T_4730; // @[Mux.scala 27:72]
  wire  _T_4279 = btb_rd_addr_p1_f == 8'h3c; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4731 = _T_4279 ? btb_bank0_rd_data_way0_out_60 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4986 = _T_4985 | _T_4731; // @[Mux.scala 27:72]
  wire  _T_4281 = btb_rd_addr_p1_f == 8'h3d; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4732 = _T_4281 ? btb_bank0_rd_data_way0_out_61 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4987 = _T_4986 | _T_4732; // @[Mux.scala 27:72]
  wire  _T_4283 = btb_rd_addr_p1_f == 8'h3e; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4733 = _T_4283 ? btb_bank0_rd_data_way0_out_62 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4988 = _T_4987 | _T_4733; // @[Mux.scala 27:72]
  wire  _T_4285 = btb_rd_addr_p1_f == 8'h3f; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4734 = _T_4285 ? btb_bank0_rd_data_way0_out_63 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4989 = _T_4988 | _T_4734; // @[Mux.scala 27:72]
  wire  _T_4287 = btb_rd_addr_p1_f == 8'h40; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4735 = _T_4287 ? btb_bank0_rd_data_way0_out_64 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4990 = _T_4989 | _T_4735; // @[Mux.scala 27:72]
  wire  _T_4289 = btb_rd_addr_p1_f == 8'h41; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4736 = _T_4289 ? btb_bank0_rd_data_way0_out_65 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4991 = _T_4990 | _T_4736; // @[Mux.scala 27:72]
  wire  _T_4291 = btb_rd_addr_p1_f == 8'h42; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4737 = _T_4291 ? btb_bank0_rd_data_way0_out_66 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4992 = _T_4991 | _T_4737; // @[Mux.scala 27:72]
  wire  _T_4293 = btb_rd_addr_p1_f == 8'h43; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4738 = _T_4293 ? btb_bank0_rd_data_way0_out_67 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4993 = _T_4992 | _T_4738; // @[Mux.scala 27:72]
  wire  _T_4295 = btb_rd_addr_p1_f == 8'h44; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4739 = _T_4295 ? btb_bank0_rd_data_way0_out_68 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4994 = _T_4993 | _T_4739; // @[Mux.scala 27:72]
  wire  _T_4297 = btb_rd_addr_p1_f == 8'h45; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4740 = _T_4297 ? btb_bank0_rd_data_way0_out_69 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4995 = _T_4994 | _T_4740; // @[Mux.scala 27:72]
  wire  _T_4299 = btb_rd_addr_p1_f == 8'h46; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4741 = _T_4299 ? btb_bank0_rd_data_way0_out_70 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4996 = _T_4995 | _T_4741; // @[Mux.scala 27:72]
  wire  _T_4301 = btb_rd_addr_p1_f == 8'h47; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4742 = _T_4301 ? btb_bank0_rd_data_way0_out_71 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4997 = _T_4996 | _T_4742; // @[Mux.scala 27:72]
  wire  _T_4303 = btb_rd_addr_p1_f == 8'h48; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4743 = _T_4303 ? btb_bank0_rd_data_way0_out_72 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4998 = _T_4997 | _T_4743; // @[Mux.scala 27:72]
  wire  _T_4305 = btb_rd_addr_p1_f == 8'h49; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4744 = _T_4305 ? btb_bank0_rd_data_way0_out_73 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4999 = _T_4998 | _T_4744; // @[Mux.scala 27:72]
  wire  _T_4307 = btb_rd_addr_p1_f == 8'h4a; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4745 = _T_4307 ? btb_bank0_rd_data_way0_out_74 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5000 = _T_4999 | _T_4745; // @[Mux.scala 27:72]
  wire  _T_4309 = btb_rd_addr_p1_f == 8'h4b; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4746 = _T_4309 ? btb_bank0_rd_data_way0_out_75 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5001 = _T_5000 | _T_4746; // @[Mux.scala 27:72]
  wire  _T_4311 = btb_rd_addr_p1_f == 8'h4c; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4747 = _T_4311 ? btb_bank0_rd_data_way0_out_76 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5002 = _T_5001 | _T_4747; // @[Mux.scala 27:72]
  wire  _T_4313 = btb_rd_addr_p1_f == 8'h4d; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4748 = _T_4313 ? btb_bank0_rd_data_way0_out_77 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5003 = _T_5002 | _T_4748; // @[Mux.scala 27:72]
  wire  _T_4315 = btb_rd_addr_p1_f == 8'h4e; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4749 = _T_4315 ? btb_bank0_rd_data_way0_out_78 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5004 = _T_5003 | _T_4749; // @[Mux.scala 27:72]
  wire  _T_4317 = btb_rd_addr_p1_f == 8'h4f; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4750 = _T_4317 ? btb_bank0_rd_data_way0_out_79 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5005 = _T_5004 | _T_4750; // @[Mux.scala 27:72]
  wire  _T_4319 = btb_rd_addr_p1_f == 8'h50; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4751 = _T_4319 ? btb_bank0_rd_data_way0_out_80 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5006 = _T_5005 | _T_4751; // @[Mux.scala 27:72]
  wire  _T_4321 = btb_rd_addr_p1_f == 8'h51; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4752 = _T_4321 ? btb_bank0_rd_data_way0_out_81 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5007 = _T_5006 | _T_4752; // @[Mux.scala 27:72]
  wire  _T_4323 = btb_rd_addr_p1_f == 8'h52; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4753 = _T_4323 ? btb_bank0_rd_data_way0_out_82 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5008 = _T_5007 | _T_4753; // @[Mux.scala 27:72]
  wire  _T_4325 = btb_rd_addr_p1_f == 8'h53; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4754 = _T_4325 ? btb_bank0_rd_data_way0_out_83 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5009 = _T_5008 | _T_4754; // @[Mux.scala 27:72]
  wire  _T_4327 = btb_rd_addr_p1_f == 8'h54; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4755 = _T_4327 ? btb_bank0_rd_data_way0_out_84 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5010 = _T_5009 | _T_4755; // @[Mux.scala 27:72]
  wire  _T_4329 = btb_rd_addr_p1_f == 8'h55; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4756 = _T_4329 ? btb_bank0_rd_data_way0_out_85 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5011 = _T_5010 | _T_4756; // @[Mux.scala 27:72]
  wire  _T_4331 = btb_rd_addr_p1_f == 8'h56; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4757 = _T_4331 ? btb_bank0_rd_data_way0_out_86 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5012 = _T_5011 | _T_4757; // @[Mux.scala 27:72]
  wire  _T_4333 = btb_rd_addr_p1_f == 8'h57; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4758 = _T_4333 ? btb_bank0_rd_data_way0_out_87 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5013 = _T_5012 | _T_4758; // @[Mux.scala 27:72]
  wire  _T_4335 = btb_rd_addr_p1_f == 8'h58; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4759 = _T_4335 ? btb_bank0_rd_data_way0_out_88 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5014 = _T_5013 | _T_4759; // @[Mux.scala 27:72]
  wire  _T_4337 = btb_rd_addr_p1_f == 8'h59; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4760 = _T_4337 ? btb_bank0_rd_data_way0_out_89 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5015 = _T_5014 | _T_4760; // @[Mux.scala 27:72]
  wire  _T_4339 = btb_rd_addr_p1_f == 8'h5a; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4761 = _T_4339 ? btb_bank0_rd_data_way0_out_90 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5016 = _T_5015 | _T_4761; // @[Mux.scala 27:72]
  wire  _T_4341 = btb_rd_addr_p1_f == 8'h5b; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4762 = _T_4341 ? btb_bank0_rd_data_way0_out_91 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5017 = _T_5016 | _T_4762; // @[Mux.scala 27:72]
  wire  _T_4343 = btb_rd_addr_p1_f == 8'h5c; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4763 = _T_4343 ? btb_bank0_rd_data_way0_out_92 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5018 = _T_5017 | _T_4763; // @[Mux.scala 27:72]
  wire  _T_4345 = btb_rd_addr_p1_f == 8'h5d; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4764 = _T_4345 ? btb_bank0_rd_data_way0_out_93 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5019 = _T_5018 | _T_4764; // @[Mux.scala 27:72]
  wire  _T_4347 = btb_rd_addr_p1_f == 8'h5e; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4765 = _T_4347 ? btb_bank0_rd_data_way0_out_94 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5020 = _T_5019 | _T_4765; // @[Mux.scala 27:72]
  wire  _T_4349 = btb_rd_addr_p1_f == 8'h5f; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4766 = _T_4349 ? btb_bank0_rd_data_way0_out_95 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5021 = _T_5020 | _T_4766; // @[Mux.scala 27:72]
  wire  _T_4351 = btb_rd_addr_p1_f == 8'h60; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4767 = _T_4351 ? btb_bank0_rd_data_way0_out_96 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5022 = _T_5021 | _T_4767; // @[Mux.scala 27:72]
  wire  _T_4353 = btb_rd_addr_p1_f == 8'h61; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4768 = _T_4353 ? btb_bank0_rd_data_way0_out_97 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5023 = _T_5022 | _T_4768; // @[Mux.scala 27:72]
  wire  _T_4355 = btb_rd_addr_p1_f == 8'h62; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4769 = _T_4355 ? btb_bank0_rd_data_way0_out_98 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5024 = _T_5023 | _T_4769; // @[Mux.scala 27:72]
  wire  _T_4357 = btb_rd_addr_p1_f == 8'h63; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4770 = _T_4357 ? btb_bank0_rd_data_way0_out_99 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5025 = _T_5024 | _T_4770; // @[Mux.scala 27:72]
  wire  _T_4359 = btb_rd_addr_p1_f == 8'h64; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4771 = _T_4359 ? btb_bank0_rd_data_way0_out_100 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5026 = _T_5025 | _T_4771; // @[Mux.scala 27:72]
  wire  _T_4361 = btb_rd_addr_p1_f == 8'h65; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4772 = _T_4361 ? btb_bank0_rd_data_way0_out_101 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5027 = _T_5026 | _T_4772; // @[Mux.scala 27:72]
  wire  _T_4363 = btb_rd_addr_p1_f == 8'h66; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4773 = _T_4363 ? btb_bank0_rd_data_way0_out_102 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5028 = _T_5027 | _T_4773; // @[Mux.scala 27:72]
  wire  _T_4365 = btb_rd_addr_p1_f == 8'h67; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4774 = _T_4365 ? btb_bank0_rd_data_way0_out_103 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5029 = _T_5028 | _T_4774; // @[Mux.scala 27:72]
  wire  _T_4367 = btb_rd_addr_p1_f == 8'h68; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4775 = _T_4367 ? btb_bank0_rd_data_way0_out_104 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5030 = _T_5029 | _T_4775; // @[Mux.scala 27:72]
  wire  _T_4369 = btb_rd_addr_p1_f == 8'h69; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4776 = _T_4369 ? btb_bank0_rd_data_way0_out_105 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5031 = _T_5030 | _T_4776; // @[Mux.scala 27:72]
  wire  _T_4371 = btb_rd_addr_p1_f == 8'h6a; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4777 = _T_4371 ? btb_bank0_rd_data_way0_out_106 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5032 = _T_5031 | _T_4777; // @[Mux.scala 27:72]
  wire  _T_4373 = btb_rd_addr_p1_f == 8'h6b; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4778 = _T_4373 ? btb_bank0_rd_data_way0_out_107 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5033 = _T_5032 | _T_4778; // @[Mux.scala 27:72]
  wire  _T_4375 = btb_rd_addr_p1_f == 8'h6c; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4779 = _T_4375 ? btb_bank0_rd_data_way0_out_108 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5034 = _T_5033 | _T_4779; // @[Mux.scala 27:72]
  wire  _T_4377 = btb_rd_addr_p1_f == 8'h6d; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4780 = _T_4377 ? btb_bank0_rd_data_way0_out_109 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5035 = _T_5034 | _T_4780; // @[Mux.scala 27:72]
  wire  _T_4379 = btb_rd_addr_p1_f == 8'h6e; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4781 = _T_4379 ? btb_bank0_rd_data_way0_out_110 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5036 = _T_5035 | _T_4781; // @[Mux.scala 27:72]
  wire  _T_4381 = btb_rd_addr_p1_f == 8'h6f; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4782 = _T_4381 ? btb_bank0_rd_data_way0_out_111 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5037 = _T_5036 | _T_4782; // @[Mux.scala 27:72]
  wire  _T_4383 = btb_rd_addr_p1_f == 8'h70; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4783 = _T_4383 ? btb_bank0_rd_data_way0_out_112 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5038 = _T_5037 | _T_4783; // @[Mux.scala 27:72]
  wire  _T_4385 = btb_rd_addr_p1_f == 8'h71; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4784 = _T_4385 ? btb_bank0_rd_data_way0_out_113 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5039 = _T_5038 | _T_4784; // @[Mux.scala 27:72]
  wire  _T_4387 = btb_rd_addr_p1_f == 8'h72; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4785 = _T_4387 ? btb_bank0_rd_data_way0_out_114 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5040 = _T_5039 | _T_4785; // @[Mux.scala 27:72]
  wire  _T_4389 = btb_rd_addr_p1_f == 8'h73; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4786 = _T_4389 ? btb_bank0_rd_data_way0_out_115 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5041 = _T_5040 | _T_4786; // @[Mux.scala 27:72]
  wire  _T_4391 = btb_rd_addr_p1_f == 8'h74; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4787 = _T_4391 ? btb_bank0_rd_data_way0_out_116 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5042 = _T_5041 | _T_4787; // @[Mux.scala 27:72]
  wire  _T_4393 = btb_rd_addr_p1_f == 8'h75; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4788 = _T_4393 ? btb_bank0_rd_data_way0_out_117 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5043 = _T_5042 | _T_4788; // @[Mux.scala 27:72]
  wire  _T_4395 = btb_rd_addr_p1_f == 8'h76; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4789 = _T_4395 ? btb_bank0_rd_data_way0_out_118 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5044 = _T_5043 | _T_4789; // @[Mux.scala 27:72]
  wire  _T_4397 = btb_rd_addr_p1_f == 8'h77; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4790 = _T_4397 ? btb_bank0_rd_data_way0_out_119 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5045 = _T_5044 | _T_4790; // @[Mux.scala 27:72]
  wire  _T_4399 = btb_rd_addr_p1_f == 8'h78; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4791 = _T_4399 ? btb_bank0_rd_data_way0_out_120 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5046 = _T_5045 | _T_4791; // @[Mux.scala 27:72]
  wire  _T_4401 = btb_rd_addr_p1_f == 8'h79; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4792 = _T_4401 ? btb_bank0_rd_data_way0_out_121 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5047 = _T_5046 | _T_4792; // @[Mux.scala 27:72]
  wire  _T_4403 = btb_rd_addr_p1_f == 8'h7a; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4793 = _T_4403 ? btb_bank0_rd_data_way0_out_122 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5048 = _T_5047 | _T_4793; // @[Mux.scala 27:72]
  wire  _T_4405 = btb_rd_addr_p1_f == 8'h7b; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4794 = _T_4405 ? btb_bank0_rd_data_way0_out_123 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5049 = _T_5048 | _T_4794; // @[Mux.scala 27:72]
  wire  _T_4407 = btb_rd_addr_p1_f == 8'h7c; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4795 = _T_4407 ? btb_bank0_rd_data_way0_out_124 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5050 = _T_5049 | _T_4795; // @[Mux.scala 27:72]
  wire  _T_4409 = btb_rd_addr_p1_f == 8'h7d; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4796 = _T_4409 ? btb_bank0_rd_data_way0_out_125 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5051 = _T_5050 | _T_4796; // @[Mux.scala 27:72]
  wire  _T_4411 = btb_rd_addr_p1_f == 8'h7e; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4797 = _T_4411 ? btb_bank0_rd_data_way0_out_126 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5052 = _T_5051 | _T_4797; // @[Mux.scala 27:72]
  wire  _T_4413 = btb_rd_addr_p1_f == 8'h7f; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4798 = _T_4413 ? btb_bank0_rd_data_way0_out_127 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5053 = _T_5052 | _T_4798; // @[Mux.scala 27:72]
  wire  _T_4415 = btb_rd_addr_p1_f == 8'h80; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4799 = _T_4415 ? btb_bank0_rd_data_way0_out_128 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5054 = _T_5053 | _T_4799; // @[Mux.scala 27:72]
  wire  _T_4417 = btb_rd_addr_p1_f == 8'h81; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4800 = _T_4417 ? btb_bank0_rd_data_way0_out_129 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5055 = _T_5054 | _T_4800; // @[Mux.scala 27:72]
  wire  _T_4419 = btb_rd_addr_p1_f == 8'h82; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4801 = _T_4419 ? btb_bank0_rd_data_way0_out_130 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5056 = _T_5055 | _T_4801; // @[Mux.scala 27:72]
  wire  _T_4421 = btb_rd_addr_p1_f == 8'h83; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4802 = _T_4421 ? btb_bank0_rd_data_way0_out_131 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5057 = _T_5056 | _T_4802; // @[Mux.scala 27:72]
  wire  _T_4423 = btb_rd_addr_p1_f == 8'h84; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4803 = _T_4423 ? btb_bank0_rd_data_way0_out_132 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5058 = _T_5057 | _T_4803; // @[Mux.scala 27:72]
  wire  _T_4425 = btb_rd_addr_p1_f == 8'h85; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4804 = _T_4425 ? btb_bank0_rd_data_way0_out_133 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5059 = _T_5058 | _T_4804; // @[Mux.scala 27:72]
  wire  _T_4427 = btb_rd_addr_p1_f == 8'h86; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4805 = _T_4427 ? btb_bank0_rd_data_way0_out_134 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5060 = _T_5059 | _T_4805; // @[Mux.scala 27:72]
  wire  _T_4429 = btb_rd_addr_p1_f == 8'h87; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4806 = _T_4429 ? btb_bank0_rd_data_way0_out_135 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5061 = _T_5060 | _T_4806; // @[Mux.scala 27:72]
  wire  _T_4431 = btb_rd_addr_p1_f == 8'h88; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4807 = _T_4431 ? btb_bank0_rd_data_way0_out_136 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5062 = _T_5061 | _T_4807; // @[Mux.scala 27:72]
  wire  _T_4433 = btb_rd_addr_p1_f == 8'h89; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4808 = _T_4433 ? btb_bank0_rd_data_way0_out_137 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5063 = _T_5062 | _T_4808; // @[Mux.scala 27:72]
  wire  _T_4435 = btb_rd_addr_p1_f == 8'h8a; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4809 = _T_4435 ? btb_bank0_rd_data_way0_out_138 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5064 = _T_5063 | _T_4809; // @[Mux.scala 27:72]
  wire  _T_4437 = btb_rd_addr_p1_f == 8'h8b; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4810 = _T_4437 ? btb_bank0_rd_data_way0_out_139 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5065 = _T_5064 | _T_4810; // @[Mux.scala 27:72]
  wire  _T_4439 = btb_rd_addr_p1_f == 8'h8c; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4811 = _T_4439 ? btb_bank0_rd_data_way0_out_140 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5066 = _T_5065 | _T_4811; // @[Mux.scala 27:72]
  wire  _T_4441 = btb_rd_addr_p1_f == 8'h8d; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4812 = _T_4441 ? btb_bank0_rd_data_way0_out_141 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5067 = _T_5066 | _T_4812; // @[Mux.scala 27:72]
  wire  _T_4443 = btb_rd_addr_p1_f == 8'h8e; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4813 = _T_4443 ? btb_bank0_rd_data_way0_out_142 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5068 = _T_5067 | _T_4813; // @[Mux.scala 27:72]
  wire  _T_4445 = btb_rd_addr_p1_f == 8'h8f; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4814 = _T_4445 ? btb_bank0_rd_data_way0_out_143 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5069 = _T_5068 | _T_4814; // @[Mux.scala 27:72]
  wire  _T_4447 = btb_rd_addr_p1_f == 8'h90; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4815 = _T_4447 ? btb_bank0_rd_data_way0_out_144 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5070 = _T_5069 | _T_4815; // @[Mux.scala 27:72]
  wire  _T_4449 = btb_rd_addr_p1_f == 8'h91; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4816 = _T_4449 ? btb_bank0_rd_data_way0_out_145 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5071 = _T_5070 | _T_4816; // @[Mux.scala 27:72]
  wire  _T_4451 = btb_rd_addr_p1_f == 8'h92; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4817 = _T_4451 ? btb_bank0_rd_data_way0_out_146 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5072 = _T_5071 | _T_4817; // @[Mux.scala 27:72]
  wire  _T_4453 = btb_rd_addr_p1_f == 8'h93; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4818 = _T_4453 ? btb_bank0_rd_data_way0_out_147 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5073 = _T_5072 | _T_4818; // @[Mux.scala 27:72]
  wire  _T_4455 = btb_rd_addr_p1_f == 8'h94; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4819 = _T_4455 ? btb_bank0_rd_data_way0_out_148 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5074 = _T_5073 | _T_4819; // @[Mux.scala 27:72]
  wire  _T_4457 = btb_rd_addr_p1_f == 8'h95; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4820 = _T_4457 ? btb_bank0_rd_data_way0_out_149 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5075 = _T_5074 | _T_4820; // @[Mux.scala 27:72]
  wire  _T_4459 = btb_rd_addr_p1_f == 8'h96; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4821 = _T_4459 ? btb_bank0_rd_data_way0_out_150 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5076 = _T_5075 | _T_4821; // @[Mux.scala 27:72]
  wire  _T_4461 = btb_rd_addr_p1_f == 8'h97; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4822 = _T_4461 ? btb_bank0_rd_data_way0_out_151 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5077 = _T_5076 | _T_4822; // @[Mux.scala 27:72]
  wire  _T_4463 = btb_rd_addr_p1_f == 8'h98; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4823 = _T_4463 ? btb_bank0_rd_data_way0_out_152 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5078 = _T_5077 | _T_4823; // @[Mux.scala 27:72]
  wire  _T_4465 = btb_rd_addr_p1_f == 8'h99; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4824 = _T_4465 ? btb_bank0_rd_data_way0_out_153 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5079 = _T_5078 | _T_4824; // @[Mux.scala 27:72]
  wire  _T_4467 = btb_rd_addr_p1_f == 8'h9a; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4825 = _T_4467 ? btb_bank0_rd_data_way0_out_154 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5080 = _T_5079 | _T_4825; // @[Mux.scala 27:72]
  wire  _T_4469 = btb_rd_addr_p1_f == 8'h9b; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4826 = _T_4469 ? btb_bank0_rd_data_way0_out_155 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5081 = _T_5080 | _T_4826; // @[Mux.scala 27:72]
  wire  _T_4471 = btb_rd_addr_p1_f == 8'h9c; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4827 = _T_4471 ? btb_bank0_rd_data_way0_out_156 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5082 = _T_5081 | _T_4827; // @[Mux.scala 27:72]
  wire  _T_4473 = btb_rd_addr_p1_f == 8'h9d; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4828 = _T_4473 ? btb_bank0_rd_data_way0_out_157 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5083 = _T_5082 | _T_4828; // @[Mux.scala 27:72]
  wire  _T_4475 = btb_rd_addr_p1_f == 8'h9e; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4829 = _T_4475 ? btb_bank0_rd_data_way0_out_158 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5084 = _T_5083 | _T_4829; // @[Mux.scala 27:72]
  wire  _T_4477 = btb_rd_addr_p1_f == 8'h9f; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4830 = _T_4477 ? btb_bank0_rd_data_way0_out_159 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5085 = _T_5084 | _T_4830; // @[Mux.scala 27:72]
  wire  _T_4479 = btb_rd_addr_p1_f == 8'ha0; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4831 = _T_4479 ? btb_bank0_rd_data_way0_out_160 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5086 = _T_5085 | _T_4831; // @[Mux.scala 27:72]
  wire  _T_4481 = btb_rd_addr_p1_f == 8'ha1; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4832 = _T_4481 ? btb_bank0_rd_data_way0_out_161 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5087 = _T_5086 | _T_4832; // @[Mux.scala 27:72]
  wire  _T_4483 = btb_rd_addr_p1_f == 8'ha2; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4833 = _T_4483 ? btb_bank0_rd_data_way0_out_162 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5088 = _T_5087 | _T_4833; // @[Mux.scala 27:72]
  wire  _T_4485 = btb_rd_addr_p1_f == 8'ha3; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4834 = _T_4485 ? btb_bank0_rd_data_way0_out_163 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5089 = _T_5088 | _T_4834; // @[Mux.scala 27:72]
  wire  _T_4487 = btb_rd_addr_p1_f == 8'ha4; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4835 = _T_4487 ? btb_bank0_rd_data_way0_out_164 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5090 = _T_5089 | _T_4835; // @[Mux.scala 27:72]
  wire  _T_4489 = btb_rd_addr_p1_f == 8'ha5; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4836 = _T_4489 ? btb_bank0_rd_data_way0_out_165 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5091 = _T_5090 | _T_4836; // @[Mux.scala 27:72]
  wire  _T_4491 = btb_rd_addr_p1_f == 8'ha6; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4837 = _T_4491 ? btb_bank0_rd_data_way0_out_166 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5092 = _T_5091 | _T_4837; // @[Mux.scala 27:72]
  wire  _T_4493 = btb_rd_addr_p1_f == 8'ha7; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4838 = _T_4493 ? btb_bank0_rd_data_way0_out_167 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5093 = _T_5092 | _T_4838; // @[Mux.scala 27:72]
  wire  _T_4495 = btb_rd_addr_p1_f == 8'ha8; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4839 = _T_4495 ? btb_bank0_rd_data_way0_out_168 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5094 = _T_5093 | _T_4839; // @[Mux.scala 27:72]
  wire  _T_4497 = btb_rd_addr_p1_f == 8'ha9; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4840 = _T_4497 ? btb_bank0_rd_data_way0_out_169 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5095 = _T_5094 | _T_4840; // @[Mux.scala 27:72]
  wire  _T_4499 = btb_rd_addr_p1_f == 8'haa; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4841 = _T_4499 ? btb_bank0_rd_data_way0_out_170 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5096 = _T_5095 | _T_4841; // @[Mux.scala 27:72]
  wire  _T_4501 = btb_rd_addr_p1_f == 8'hab; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4842 = _T_4501 ? btb_bank0_rd_data_way0_out_171 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5097 = _T_5096 | _T_4842; // @[Mux.scala 27:72]
  wire  _T_4503 = btb_rd_addr_p1_f == 8'hac; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4843 = _T_4503 ? btb_bank0_rd_data_way0_out_172 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5098 = _T_5097 | _T_4843; // @[Mux.scala 27:72]
  wire  _T_4505 = btb_rd_addr_p1_f == 8'had; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4844 = _T_4505 ? btb_bank0_rd_data_way0_out_173 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5099 = _T_5098 | _T_4844; // @[Mux.scala 27:72]
  wire  _T_4507 = btb_rd_addr_p1_f == 8'hae; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4845 = _T_4507 ? btb_bank0_rd_data_way0_out_174 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5100 = _T_5099 | _T_4845; // @[Mux.scala 27:72]
  wire  _T_4509 = btb_rd_addr_p1_f == 8'haf; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4846 = _T_4509 ? btb_bank0_rd_data_way0_out_175 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5101 = _T_5100 | _T_4846; // @[Mux.scala 27:72]
  wire  _T_4511 = btb_rd_addr_p1_f == 8'hb0; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4847 = _T_4511 ? btb_bank0_rd_data_way0_out_176 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5102 = _T_5101 | _T_4847; // @[Mux.scala 27:72]
  wire  _T_4513 = btb_rd_addr_p1_f == 8'hb1; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4848 = _T_4513 ? btb_bank0_rd_data_way0_out_177 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5103 = _T_5102 | _T_4848; // @[Mux.scala 27:72]
  wire  _T_4515 = btb_rd_addr_p1_f == 8'hb2; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4849 = _T_4515 ? btb_bank0_rd_data_way0_out_178 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5104 = _T_5103 | _T_4849; // @[Mux.scala 27:72]
  wire  _T_4517 = btb_rd_addr_p1_f == 8'hb3; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4850 = _T_4517 ? btb_bank0_rd_data_way0_out_179 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5105 = _T_5104 | _T_4850; // @[Mux.scala 27:72]
  wire  _T_4519 = btb_rd_addr_p1_f == 8'hb4; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4851 = _T_4519 ? btb_bank0_rd_data_way0_out_180 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5106 = _T_5105 | _T_4851; // @[Mux.scala 27:72]
  wire  _T_4521 = btb_rd_addr_p1_f == 8'hb5; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4852 = _T_4521 ? btb_bank0_rd_data_way0_out_181 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5107 = _T_5106 | _T_4852; // @[Mux.scala 27:72]
  wire  _T_4523 = btb_rd_addr_p1_f == 8'hb6; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4853 = _T_4523 ? btb_bank0_rd_data_way0_out_182 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5108 = _T_5107 | _T_4853; // @[Mux.scala 27:72]
  wire  _T_4525 = btb_rd_addr_p1_f == 8'hb7; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4854 = _T_4525 ? btb_bank0_rd_data_way0_out_183 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5109 = _T_5108 | _T_4854; // @[Mux.scala 27:72]
  wire  _T_4527 = btb_rd_addr_p1_f == 8'hb8; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4855 = _T_4527 ? btb_bank0_rd_data_way0_out_184 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5110 = _T_5109 | _T_4855; // @[Mux.scala 27:72]
  wire  _T_4529 = btb_rd_addr_p1_f == 8'hb9; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4856 = _T_4529 ? btb_bank0_rd_data_way0_out_185 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5111 = _T_5110 | _T_4856; // @[Mux.scala 27:72]
  wire  _T_4531 = btb_rd_addr_p1_f == 8'hba; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4857 = _T_4531 ? btb_bank0_rd_data_way0_out_186 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5112 = _T_5111 | _T_4857; // @[Mux.scala 27:72]
  wire  _T_4533 = btb_rd_addr_p1_f == 8'hbb; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4858 = _T_4533 ? btb_bank0_rd_data_way0_out_187 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5113 = _T_5112 | _T_4858; // @[Mux.scala 27:72]
  wire  _T_4535 = btb_rd_addr_p1_f == 8'hbc; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4859 = _T_4535 ? btb_bank0_rd_data_way0_out_188 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5114 = _T_5113 | _T_4859; // @[Mux.scala 27:72]
  wire  _T_4537 = btb_rd_addr_p1_f == 8'hbd; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4860 = _T_4537 ? btb_bank0_rd_data_way0_out_189 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5115 = _T_5114 | _T_4860; // @[Mux.scala 27:72]
  wire  _T_4539 = btb_rd_addr_p1_f == 8'hbe; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4861 = _T_4539 ? btb_bank0_rd_data_way0_out_190 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5116 = _T_5115 | _T_4861; // @[Mux.scala 27:72]
  wire  _T_4541 = btb_rd_addr_p1_f == 8'hbf; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4862 = _T_4541 ? btb_bank0_rd_data_way0_out_191 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5117 = _T_5116 | _T_4862; // @[Mux.scala 27:72]
  wire  _T_4543 = btb_rd_addr_p1_f == 8'hc0; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4863 = _T_4543 ? btb_bank0_rd_data_way0_out_192 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5118 = _T_5117 | _T_4863; // @[Mux.scala 27:72]
  wire  _T_4545 = btb_rd_addr_p1_f == 8'hc1; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4864 = _T_4545 ? btb_bank0_rd_data_way0_out_193 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5119 = _T_5118 | _T_4864; // @[Mux.scala 27:72]
  wire  _T_4547 = btb_rd_addr_p1_f == 8'hc2; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4865 = _T_4547 ? btb_bank0_rd_data_way0_out_194 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5120 = _T_5119 | _T_4865; // @[Mux.scala 27:72]
  wire  _T_4549 = btb_rd_addr_p1_f == 8'hc3; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4866 = _T_4549 ? btb_bank0_rd_data_way0_out_195 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5121 = _T_5120 | _T_4866; // @[Mux.scala 27:72]
  wire  _T_4551 = btb_rd_addr_p1_f == 8'hc4; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4867 = _T_4551 ? btb_bank0_rd_data_way0_out_196 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5122 = _T_5121 | _T_4867; // @[Mux.scala 27:72]
  wire  _T_4553 = btb_rd_addr_p1_f == 8'hc5; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4868 = _T_4553 ? btb_bank0_rd_data_way0_out_197 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5123 = _T_5122 | _T_4868; // @[Mux.scala 27:72]
  wire  _T_4555 = btb_rd_addr_p1_f == 8'hc6; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4869 = _T_4555 ? btb_bank0_rd_data_way0_out_198 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5124 = _T_5123 | _T_4869; // @[Mux.scala 27:72]
  wire  _T_4557 = btb_rd_addr_p1_f == 8'hc7; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4870 = _T_4557 ? btb_bank0_rd_data_way0_out_199 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5125 = _T_5124 | _T_4870; // @[Mux.scala 27:72]
  wire  _T_4559 = btb_rd_addr_p1_f == 8'hc8; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4871 = _T_4559 ? btb_bank0_rd_data_way0_out_200 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5126 = _T_5125 | _T_4871; // @[Mux.scala 27:72]
  wire  _T_4561 = btb_rd_addr_p1_f == 8'hc9; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4872 = _T_4561 ? btb_bank0_rd_data_way0_out_201 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5127 = _T_5126 | _T_4872; // @[Mux.scala 27:72]
  wire  _T_4563 = btb_rd_addr_p1_f == 8'hca; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4873 = _T_4563 ? btb_bank0_rd_data_way0_out_202 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5128 = _T_5127 | _T_4873; // @[Mux.scala 27:72]
  wire  _T_4565 = btb_rd_addr_p1_f == 8'hcb; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4874 = _T_4565 ? btb_bank0_rd_data_way0_out_203 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5129 = _T_5128 | _T_4874; // @[Mux.scala 27:72]
  wire  _T_4567 = btb_rd_addr_p1_f == 8'hcc; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4875 = _T_4567 ? btb_bank0_rd_data_way0_out_204 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5130 = _T_5129 | _T_4875; // @[Mux.scala 27:72]
  wire  _T_4569 = btb_rd_addr_p1_f == 8'hcd; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4876 = _T_4569 ? btb_bank0_rd_data_way0_out_205 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5131 = _T_5130 | _T_4876; // @[Mux.scala 27:72]
  wire  _T_4571 = btb_rd_addr_p1_f == 8'hce; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4877 = _T_4571 ? btb_bank0_rd_data_way0_out_206 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5132 = _T_5131 | _T_4877; // @[Mux.scala 27:72]
  wire  _T_4573 = btb_rd_addr_p1_f == 8'hcf; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4878 = _T_4573 ? btb_bank0_rd_data_way0_out_207 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5133 = _T_5132 | _T_4878; // @[Mux.scala 27:72]
  wire  _T_4575 = btb_rd_addr_p1_f == 8'hd0; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4879 = _T_4575 ? btb_bank0_rd_data_way0_out_208 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5134 = _T_5133 | _T_4879; // @[Mux.scala 27:72]
  wire  _T_4577 = btb_rd_addr_p1_f == 8'hd1; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4880 = _T_4577 ? btb_bank0_rd_data_way0_out_209 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5135 = _T_5134 | _T_4880; // @[Mux.scala 27:72]
  wire  _T_4579 = btb_rd_addr_p1_f == 8'hd2; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4881 = _T_4579 ? btb_bank0_rd_data_way0_out_210 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5136 = _T_5135 | _T_4881; // @[Mux.scala 27:72]
  wire  _T_4581 = btb_rd_addr_p1_f == 8'hd3; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4882 = _T_4581 ? btb_bank0_rd_data_way0_out_211 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5137 = _T_5136 | _T_4882; // @[Mux.scala 27:72]
  wire  _T_4583 = btb_rd_addr_p1_f == 8'hd4; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4883 = _T_4583 ? btb_bank0_rd_data_way0_out_212 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5138 = _T_5137 | _T_4883; // @[Mux.scala 27:72]
  wire  _T_4585 = btb_rd_addr_p1_f == 8'hd5; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4884 = _T_4585 ? btb_bank0_rd_data_way0_out_213 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5139 = _T_5138 | _T_4884; // @[Mux.scala 27:72]
  wire  _T_4587 = btb_rd_addr_p1_f == 8'hd6; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4885 = _T_4587 ? btb_bank0_rd_data_way0_out_214 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5140 = _T_5139 | _T_4885; // @[Mux.scala 27:72]
  wire  _T_4589 = btb_rd_addr_p1_f == 8'hd7; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4886 = _T_4589 ? btb_bank0_rd_data_way0_out_215 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5141 = _T_5140 | _T_4886; // @[Mux.scala 27:72]
  wire  _T_4591 = btb_rd_addr_p1_f == 8'hd8; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4887 = _T_4591 ? btb_bank0_rd_data_way0_out_216 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5142 = _T_5141 | _T_4887; // @[Mux.scala 27:72]
  wire  _T_4593 = btb_rd_addr_p1_f == 8'hd9; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4888 = _T_4593 ? btb_bank0_rd_data_way0_out_217 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5143 = _T_5142 | _T_4888; // @[Mux.scala 27:72]
  wire  _T_4595 = btb_rd_addr_p1_f == 8'hda; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4889 = _T_4595 ? btb_bank0_rd_data_way0_out_218 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5144 = _T_5143 | _T_4889; // @[Mux.scala 27:72]
  wire  _T_4597 = btb_rd_addr_p1_f == 8'hdb; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4890 = _T_4597 ? btb_bank0_rd_data_way0_out_219 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5145 = _T_5144 | _T_4890; // @[Mux.scala 27:72]
  wire  _T_4599 = btb_rd_addr_p1_f == 8'hdc; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4891 = _T_4599 ? btb_bank0_rd_data_way0_out_220 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5146 = _T_5145 | _T_4891; // @[Mux.scala 27:72]
  wire  _T_4601 = btb_rd_addr_p1_f == 8'hdd; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4892 = _T_4601 ? btb_bank0_rd_data_way0_out_221 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5147 = _T_5146 | _T_4892; // @[Mux.scala 27:72]
  wire  _T_4603 = btb_rd_addr_p1_f == 8'hde; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4893 = _T_4603 ? btb_bank0_rd_data_way0_out_222 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5148 = _T_5147 | _T_4893; // @[Mux.scala 27:72]
  wire  _T_4605 = btb_rd_addr_p1_f == 8'hdf; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4894 = _T_4605 ? btb_bank0_rd_data_way0_out_223 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5149 = _T_5148 | _T_4894; // @[Mux.scala 27:72]
  wire  _T_4607 = btb_rd_addr_p1_f == 8'he0; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4895 = _T_4607 ? btb_bank0_rd_data_way0_out_224 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5150 = _T_5149 | _T_4895; // @[Mux.scala 27:72]
  wire  _T_4609 = btb_rd_addr_p1_f == 8'he1; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4896 = _T_4609 ? btb_bank0_rd_data_way0_out_225 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5151 = _T_5150 | _T_4896; // @[Mux.scala 27:72]
  wire  _T_4611 = btb_rd_addr_p1_f == 8'he2; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4897 = _T_4611 ? btb_bank0_rd_data_way0_out_226 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5152 = _T_5151 | _T_4897; // @[Mux.scala 27:72]
  wire  _T_4613 = btb_rd_addr_p1_f == 8'he3; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4898 = _T_4613 ? btb_bank0_rd_data_way0_out_227 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5153 = _T_5152 | _T_4898; // @[Mux.scala 27:72]
  wire  _T_4615 = btb_rd_addr_p1_f == 8'he4; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4899 = _T_4615 ? btb_bank0_rd_data_way0_out_228 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5154 = _T_5153 | _T_4899; // @[Mux.scala 27:72]
  wire  _T_4617 = btb_rd_addr_p1_f == 8'he5; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4900 = _T_4617 ? btb_bank0_rd_data_way0_out_229 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5155 = _T_5154 | _T_4900; // @[Mux.scala 27:72]
  wire  _T_4619 = btb_rd_addr_p1_f == 8'he6; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4901 = _T_4619 ? btb_bank0_rd_data_way0_out_230 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5156 = _T_5155 | _T_4901; // @[Mux.scala 27:72]
  wire  _T_4621 = btb_rd_addr_p1_f == 8'he7; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4902 = _T_4621 ? btb_bank0_rd_data_way0_out_231 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5157 = _T_5156 | _T_4902; // @[Mux.scala 27:72]
  wire  _T_4623 = btb_rd_addr_p1_f == 8'he8; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4903 = _T_4623 ? btb_bank0_rd_data_way0_out_232 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5158 = _T_5157 | _T_4903; // @[Mux.scala 27:72]
  wire  _T_4625 = btb_rd_addr_p1_f == 8'he9; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4904 = _T_4625 ? btb_bank0_rd_data_way0_out_233 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5159 = _T_5158 | _T_4904; // @[Mux.scala 27:72]
  wire  _T_4627 = btb_rd_addr_p1_f == 8'hea; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4905 = _T_4627 ? btb_bank0_rd_data_way0_out_234 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5160 = _T_5159 | _T_4905; // @[Mux.scala 27:72]
  wire  _T_4629 = btb_rd_addr_p1_f == 8'heb; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4906 = _T_4629 ? btb_bank0_rd_data_way0_out_235 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5161 = _T_5160 | _T_4906; // @[Mux.scala 27:72]
  wire  _T_4631 = btb_rd_addr_p1_f == 8'hec; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4907 = _T_4631 ? btb_bank0_rd_data_way0_out_236 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5162 = _T_5161 | _T_4907; // @[Mux.scala 27:72]
  wire  _T_4633 = btb_rd_addr_p1_f == 8'hed; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4908 = _T_4633 ? btb_bank0_rd_data_way0_out_237 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5163 = _T_5162 | _T_4908; // @[Mux.scala 27:72]
  wire  _T_4635 = btb_rd_addr_p1_f == 8'hee; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4909 = _T_4635 ? btb_bank0_rd_data_way0_out_238 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5164 = _T_5163 | _T_4909; // @[Mux.scala 27:72]
  wire  _T_4637 = btb_rd_addr_p1_f == 8'hef; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4910 = _T_4637 ? btb_bank0_rd_data_way0_out_239 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5165 = _T_5164 | _T_4910; // @[Mux.scala 27:72]
  wire  _T_4639 = btb_rd_addr_p1_f == 8'hf0; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4911 = _T_4639 ? btb_bank0_rd_data_way0_out_240 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5166 = _T_5165 | _T_4911; // @[Mux.scala 27:72]
  wire  _T_4641 = btb_rd_addr_p1_f == 8'hf1; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4912 = _T_4641 ? btb_bank0_rd_data_way0_out_241 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5167 = _T_5166 | _T_4912; // @[Mux.scala 27:72]
  wire  _T_4643 = btb_rd_addr_p1_f == 8'hf2; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4913 = _T_4643 ? btb_bank0_rd_data_way0_out_242 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5168 = _T_5167 | _T_4913; // @[Mux.scala 27:72]
  wire  _T_4645 = btb_rd_addr_p1_f == 8'hf3; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4914 = _T_4645 ? btb_bank0_rd_data_way0_out_243 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5169 = _T_5168 | _T_4914; // @[Mux.scala 27:72]
  wire  _T_4647 = btb_rd_addr_p1_f == 8'hf4; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4915 = _T_4647 ? btb_bank0_rd_data_way0_out_244 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5170 = _T_5169 | _T_4915; // @[Mux.scala 27:72]
  wire  _T_4649 = btb_rd_addr_p1_f == 8'hf5; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4916 = _T_4649 ? btb_bank0_rd_data_way0_out_245 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5171 = _T_5170 | _T_4916; // @[Mux.scala 27:72]
  wire  _T_4651 = btb_rd_addr_p1_f == 8'hf6; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4917 = _T_4651 ? btb_bank0_rd_data_way0_out_246 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5172 = _T_5171 | _T_4917; // @[Mux.scala 27:72]
  wire  _T_4653 = btb_rd_addr_p1_f == 8'hf7; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4918 = _T_4653 ? btb_bank0_rd_data_way0_out_247 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5173 = _T_5172 | _T_4918; // @[Mux.scala 27:72]
  wire  _T_4655 = btb_rd_addr_p1_f == 8'hf8; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4919 = _T_4655 ? btb_bank0_rd_data_way0_out_248 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5174 = _T_5173 | _T_4919; // @[Mux.scala 27:72]
  wire  _T_4657 = btb_rd_addr_p1_f == 8'hf9; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4920 = _T_4657 ? btb_bank0_rd_data_way0_out_249 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5175 = _T_5174 | _T_4920; // @[Mux.scala 27:72]
  wire  _T_4659 = btb_rd_addr_p1_f == 8'hfa; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4921 = _T_4659 ? btb_bank0_rd_data_way0_out_250 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5176 = _T_5175 | _T_4921; // @[Mux.scala 27:72]
  wire  _T_4661 = btb_rd_addr_p1_f == 8'hfb; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4922 = _T_4661 ? btb_bank0_rd_data_way0_out_251 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5177 = _T_5176 | _T_4922; // @[Mux.scala 27:72]
  wire  _T_4663 = btb_rd_addr_p1_f == 8'hfc; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4923 = _T_4663 ? btb_bank0_rd_data_way0_out_252 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5178 = _T_5177 | _T_4923; // @[Mux.scala 27:72]
  wire  _T_4665 = btb_rd_addr_p1_f == 8'hfd; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4924 = _T_4665 ? btb_bank0_rd_data_way0_out_253 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5179 = _T_5178 | _T_4924; // @[Mux.scala 27:72]
  wire  _T_4667 = btb_rd_addr_p1_f == 8'hfe; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4925 = _T_4667 ? btb_bank0_rd_data_way0_out_254 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5180 = _T_5179 | _T_4925; // @[Mux.scala 27:72]
  wire  _T_4669 = btb_rd_addr_p1_f == 8'hff; // @[el2_ifu_bp_ctl.scala 434:83]
  wire [21:0] _T_4926 = _T_4669 ? btb_bank0_rd_data_way0_out_255 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] btb_bank0_rd_data_way0_p1_f = _T_5180 | _T_4926; // @[Mux.scala 27:72]
  wire [4:0] _T_31 = _T_8[13:9] ^ _T_8[18:14]; // @[el2_lib.scala 180:111]
  wire [4:0] fetch_rd_tag_p1_f = _T_31 ^ _T_8[23:19]; // @[el2_lib.scala 180:111]
  wire  _T_63 = btb_bank0_rd_data_way0_p1_f[21:17] == fetch_rd_tag_p1_f; // @[el2_ifu_bp_ctl.scala 147:106]
  wire  _T_64 = btb_bank0_rd_data_way0_p1_f[0] & _T_63; // @[el2_ifu_bp_ctl.scala 147:61]
  wire  _T_67 = _T_64 & _T_48; // @[el2_ifu_bp_ctl.scala 147:129]
  wire  _T_68 = _T_67 & io_ifc_fetch_req_f; // @[el2_ifu_bp_ctl.scala 148:56]
  wire  tag_match_way0_p1_f = _T_68 & _T; // @[el2_ifu_bp_ctl.scala 148:77]
  wire  _T_99 = btb_bank0_rd_data_way0_p1_f[3] ^ btb_bank0_rd_data_way0_p1_f[4]; // @[el2_ifu_bp_ctl.scala 160:100]
  wire  _T_100 = tag_match_way0_p1_f & _T_99; // @[el2_ifu_bp_ctl.scala 160:62]
  wire  _T_104 = ~_T_99; // @[el2_ifu_bp_ctl.scala 161:64]
  wire  _T_105 = tag_match_way0_p1_f & _T_104; // @[el2_ifu_bp_ctl.scala 161:62]
  wire [1:0] tag_match_way0_expanded_p1_f = {_T_100,_T_105}; // @[Cat.scala 29:58]
  wire [21:0] _T_133 = tag_match_way0_expanded_p1_f[0] ? btb_bank0_rd_data_way0_p1_f : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5695 = _T_4159 ? btb_bank0_rd_data_way1_out_0 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5696 = _T_4161 ? btb_bank0_rd_data_way1_out_1 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5951 = _T_5695 | _T_5696; // @[Mux.scala 27:72]
  wire [21:0] _T_5697 = _T_4163 ? btb_bank0_rd_data_way1_out_2 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5952 = _T_5951 | _T_5697; // @[Mux.scala 27:72]
  wire [21:0] _T_5698 = _T_4165 ? btb_bank0_rd_data_way1_out_3 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5953 = _T_5952 | _T_5698; // @[Mux.scala 27:72]
  wire [21:0] _T_5699 = _T_4167 ? btb_bank0_rd_data_way1_out_4 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5954 = _T_5953 | _T_5699; // @[Mux.scala 27:72]
  wire [21:0] _T_5700 = _T_4169 ? btb_bank0_rd_data_way1_out_5 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5955 = _T_5954 | _T_5700; // @[Mux.scala 27:72]
  wire [21:0] _T_5701 = _T_4171 ? btb_bank0_rd_data_way1_out_6 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5956 = _T_5955 | _T_5701; // @[Mux.scala 27:72]
  wire [21:0] _T_5702 = _T_4173 ? btb_bank0_rd_data_way1_out_7 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5957 = _T_5956 | _T_5702; // @[Mux.scala 27:72]
  wire [21:0] _T_5703 = _T_4175 ? btb_bank0_rd_data_way1_out_8 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5958 = _T_5957 | _T_5703; // @[Mux.scala 27:72]
  wire [21:0] _T_5704 = _T_4177 ? btb_bank0_rd_data_way1_out_9 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5959 = _T_5958 | _T_5704; // @[Mux.scala 27:72]
  wire [21:0] _T_5705 = _T_4179 ? btb_bank0_rd_data_way1_out_10 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5960 = _T_5959 | _T_5705; // @[Mux.scala 27:72]
  wire [21:0] _T_5706 = _T_4181 ? btb_bank0_rd_data_way1_out_11 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5961 = _T_5960 | _T_5706; // @[Mux.scala 27:72]
  wire [21:0] _T_5707 = _T_4183 ? btb_bank0_rd_data_way1_out_12 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5962 = _T_5961 | _T_5707; // @[Mux.scala 27:72]
  wire [21:0] _T_5708 = _T_4185 ? btb_bank0_rd_data_way1_out_13 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5963 = _T_5962 | _T_5708; // @[Mux.scala 27:72]
  wire [21:0] _T_5709 = _T_4187 ? btb_bank0_rd_data_way1_out_14 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5964 = _T_5963 | _T_5709; // @[Mux.scala 27:72]
  wire [21:0] _T_5710 = _T_4189 ? btb_bank0_rd_data_way1_out_15 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5965 = _T_5964 | _T_5710; // @[Mux.scala 27:72]
  wire [21:0] _T_5711 = _T_4191 ? btb_bank0_rd_data_way1_out_16 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5966 = _T_5965 | _T_5711; // @[Mux.scala 27:72]
  wire [21:0] _T_5712 = _T_4193 ? btb_bank0_rd_data_way1_out_17 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5967 = _T_5966 | _T_5712; // @[Mux.scala 27:72]
  wire [21:0] _T_5713 = _T_4195 ? btb_bank0_rd_data_way1_out_18 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5968 = _T_5967 | _T_5713; // @[Mux.scala 27:72]
  wire [21:0] _T_5714 = _T_4197 ? btb_bank0_rd_data_way1_out_19 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5969 = _T_5968 | _T_5714; // @[Mux.scala 27:72]
  wire [21:0] _T_5715 = _T_4199 ? btb_bank0_rd_data_way1_out_20 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5970 = _T_5969 | _T_5715; // @[Mux.scala 27:72]
  wire [21:0] _T_5716 = _T_4201 ? btb_bank0_rd_data_way1_out_21 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5971 = _T_5970 | _T_5716; // @[Mux.scala 27:72]
  wire [21:0] _T_5717 = _T_4203 ? btb_bank0_rd_data_way1_out_22 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5972 = _T_5971 | _T_5717; // @[Mux.scala 27:72]
  wire [21:0] _T_5718 = _T_4205 ? btb_bank0_rd_data_way1_out_23 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5973 = _T_5972 | _T_5718; // @[Mux.scala 27:72]
  wire [21:0] _T_5719 = _T_4207 ? btb_bank0_rd_data_way1_out_24 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5974 = _T_5973 | _T_5719; // @[Mux.scala 27:72]
  wire [21:0] _T_5720 = _T_4209 ? btb_bank0_rd_data_way1_out_25 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5975 = _T_5974 | _T_5720; // @[Mux.scala 27:72]
  wire [21:0] _T_5721 = _T_4211 ? btb_bank0_rd_data_way1_out_26 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5976 = _T_5975 | _T_5721; // @[Mux.scala 27:72]
  wire [21:0] _T_5722 = _T_4213 ? btb_bank0_rd_data_way1_out_27 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5977 = _T_5976 | _T_5722; // @[Mux.scala 27:72]
  wire [21:0] _T_5723 = _T_4215 ? btb_bank0_rd_data_way1_out_28 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5978 = _T_5977 | _T_5723; // @[Mux.scala 27:72]
  wire [21:0] _T_5724 = _T_4217 ? btb_bank0_rd_data_way1_out_29 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5979 = _T_5978 | _T_5724; // @[Mux.scala 27:72]
  wire [21:0] _T_5725 = _T_4219 ? btb_bank0_rd_data_way1_out_30 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5980 = _T_5979 | _T_5725; // @[Mux.scala 27:72]
  wire [21:0] _T_5726 = _T_4221 ? btb_bank0_rd_data_way1_out_31 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5981 = _T_5980 | _T_5726; // @[Mux.scala 27:72]
  wire [21:0] _T_5727 = _T_4223 ? btb_bank0_rd_data_way1_out_32 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5982 = _T_5981 | _T_5727; // @[Mux.scala 27:72]
  wire [21:0] _T_5728 = _T_4225 ? btb_bank0_rd_data_way1_out_33 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5983 = _T_5982 | _T_5728; // @[Mux.scala 27:72]
  wire [21:0] _T_5729 = _T_4227 ? btb_bank0_rd_data_way1_out_34 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5984 = _T_5983 | _T_5729; // @[Mux.scala 27:72]
  wire [21:0] _T_5730 = _T_4229 ? btb_bank0_rd_data_way1_out_35 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5985 = _T_5984 | _T_5730; // @[Mux.scala 27:72]
  wire [21:0] _T_5731 = _T_4231 ? btb_bank0_rd_data_way1_out_36 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5986 = _T_5985 | _T_5731; // @[Mux.scala 27:72]
  wire [21:0] _T_5732 = _T_4233 ? btb_bank0_rd_data_way1_out_37 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5987 = _T_5986 | _T_5732; // @[Mux.scala 27:72]
  wire [21:0] _T_5733 = _T_4235 ? btb_bank0_rd_data_way1_out_38 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5988 = _T_5987 | _T_5733; // @[Mux.scala 27:72]
  wire [21:0] _T_5734 = _T_4237 ? btb_bank0_rd_data_way1_out_39 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5989 = _T_5988 | _T_5734; // @[Mux.scala 27:72]
  wire [21:0] _T_5735 = _T_4239 ? btb_bank0_rd_data_way1_out_40 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5990 = _T_5989 | _T_5735; // @[Mux.scala 27:72]
  wire [21:0] _T_5736 = _T_4241 ? btb_bank0_rd_data_way1_out_41 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5991 = _T_5990 | _T_5736; // @[Mux.scala 27:72]
  wire [21:0] _T_5737 = _T_4243 ? btb_bank0_rd_data_way1_out_42 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5992 = _T_5991 | _T_5737; // @[Mux.scala 27:72]
  wire [21:0] _T_5738 = _T_4245 ? btb_bank0_rd_data_way1_out_43 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5993 = _T_5992 | _T_5738; // @[Mux.scala 27:72]
  wire [21:0] _T_5739 = _T_4247 ? btb_bank0_rd_data_way1_out_44 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5994 = _T_5993 | _T_5739; // @[Mux.scala 27:72]
  wire [21:0] _T_5740 = _T_4249 ? btb_bank0_rd_data_way1_out_45 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5995 = _T_5994 | _T_5740; // @[Mux.scala 27:72]
  wire [21:0] _T_5741 = _T_4251 ? btb_bank0_rd_data_way1_out_46 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5996 = _T_5995 | _T_5741; // @[Mux.scala 27:72]
  wire [21:0] _T_5742 = _T_4253 ? btb_bank0_rd_data_way1_out_47 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5997 = _T_5996 | _T_5742; // @[Mux.scala 27:72]
  wire [21:0] _T_5743 = _T_4255 ? btb_bank0_rd_data_way1_out_48 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5998 = _T_5997 | _T_5743; // @[Mux.scala 27:72]
  wire [21:0] _T_5744 = _T_4257 ? btb_bank0_rd_data_way1_out_49 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5999 = _T_5998 | _T_5744; // @[Mux.scala 27:72]
  wire [21:0] _T_5745 = _T_4259 ? btb_bank0_rd_data_way1_out_50 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6000 = _T_5999 | _T_5745; // @[Mux.scala 27:72]
  wire [21:0] _T_5746 = _T_4261 ? btb_bank0_rd_data_way1_out_51 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6001 = _T_6000 | _T_5746; // @[Mux.scala 27:72]
  wire [21:0] _T_5747 = _T_4263 ? btb_bank0_rd_data_way1_out_52 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6002 = _T_6001 | _T_5747; // @[Mux.scala 27:72]
  wire [21:0] _T_5748 = _T_4265 ? btb_bank0_rd_data_way1_out_53 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6003 = _T_6002 | _T_5748; // @[Mux.scala 27:72]
  wire [21:0] _T_5749 = _T_4267 ? btb_bank0_rd_data_way1_out_54 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6004 = _T_6003 | _T_5749; // @[Mux.scala 27:72]
  wire [21:0] _T_5750 = _T_4269 ? btb_bank0_rd_data_way1_out_55 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6005 = _T_6004 | _T_5750; // @[Mux.scala 27:72]
  wire [21:0] _T_5751 = _T_4271 ? btb_bank0_rd_data_way1_out_56 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6006 = _T_6005 | _T_5751; // @[Mux.scala 27:72]
  wire [21:0] _T_5752 = _T_4273 ? btb_bank0_rd_data_way1_out_57 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6007 = _T_6006 | _T_5752; // @[Mux.scala 27:72]
  wire [21:0] _T_5753 = _T_4275 ? btb_bank0_rd_data_way1_out_58 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6008 = _T_6007 | _T_5753; // @[Mux.scala 27:72]
  wire [21:0] _T_5754 = _T_4277 ? btb_bank0_rd_data_way1_out_59 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6009 = _T_6008 | _T_5754; // @[Mux.scala 27:72]
  wire [21:0] _T_5755 = _T_4279 ? btb_bank0_rd_data_way1_out_60 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6010 = _T_6009 | _T_5755; // @[Mux.scala 27:72]
  wire [21:0] _T_5756 = _T_4281 ? btb_bank0_rd_data_way1_out_61 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6011 = _T_6010 | _T_5756; // @[Mux.scala 27:72]
  wire [21:0] _T_5757 = _T_4283 ? btb_bank0_rd_data_way1_out_62 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6012 = _T_6011 | _T_5757; // @[Mux.scala 27:72]
  wire [21:0] _T_5758 = _T_4285 ? btb_bank0_rd_data_way1_out_63 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6013 = _T_6012 | _T_5758; // @[Mux.scala 27:72]
  wire [21:0] _T_5759 = _T_4287 ? btb_bank0_rd_data_way1_out_64 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6014 = _T_6013 | _T_5759; // @[Mux.scala 27:72]
  wire [21:0] _T_5760 = _T_4289 ? btb_bank0_rd_data_way1_out_65 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6015 = _T_6014 | _T_5760; // @[Mux.scala 27:72]
  wire [21:0] _T_5761 = _T_4291 ? btb_bank0_rd_data_way1_out_66 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6016 = _T_6015 | _T_5761; // @[Mux.scala 27:72]
  wire [21:0] _T_5762 = _T_4293 ? btb_bank0_rd_data_way1_out_67 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6017 = _T_6016 | _T_5762; // @[Mux.scala 27:72]
  wire [21:0] _T_5763 = _T_4295 ? btb_bank0_rd_data_way1_out_68 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6018 = _T_6017 | _T_5763; // @[Mux.scala 27:72]
  wire [21:0] _T_5764 = _T_4297 ? btb_bank0_rd_data_way1_out_69 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6019 = _T_6018 | _T_5764; // @[Mux.scala 27:72]
  wire [21:0] _T_5765 = _T_4299 ? btb_bank0_rd_data_way1_out_70 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6020 = _T_6019 | _T_5765; // @[Mux.scala 27:72]
  wire [21:0] _T_5766 = _T_4301 ? btb_bank0_rd_data_way1_out_71 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6021 = _T_6020 | _T_5766; // @[Mux.scala 27:72]
  wire [21:0] _T_5767 = _T_4303 ? btb_bank0_rd_data_way1_out_72 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6022 = _T_6021 | _T_5767; // @[Mux.scala 27:72]
  wire [21:0] _T_5768 = _T_4305 ? btb_bank0_rd_data_way1_out_73 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6023 = _T_6022 | _T_5768; // @[Mux.scala 27:72]
  wire [21:0] _T_5769 = _T_4307 ? btb_bank0_rd_data_way1_out_74 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6024 = _T_6023 | _T_5769; // @[Mux.scala 27:72]
  wire [21:0] _T_5770 = _T_4309 ? btb_bank0_rd_data_way1_out_75 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6025 = _T_6024 | _T_5770; // @[Mux.scala 27:72]
  wire [21:0] _T_5771 = _T_4311 ? btb_bank0_rd_data_way1_out_76 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6026 = _T_6025 | _T_5771; // @[Mux.scala 27:72]
  wire [21:0] _T_5772 = _T_4313 ? btb_bank0_rd_data_way1_out_77 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6027 = _T_6026 | _T_5772; // @[Mux.scala 27:72]
  wire [21:0] _T_5773 = _T_4315 ? btb_bank0_rd_data_way1_out_78 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6028 = _T_6027 | _T_5773; // @[Mux.scala 27:72]
  wire [21:0] _T_5774 = _T_4317 ? btb_bank0_rd_data_way1_out_79 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6029 = _T_6028 | _T_5774; // @[Mux.scala 27:72]
  wire [21:0] _T_5775 = _T_4319 ? btb_bank0_rd_data_way1_out_80 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6030 = _T_6029 | _T_5775; // @[Mux.scala 27:72]
  wire [21:0] _T_5776 = _T_4321 ? btb_bank0_rd_data_way1_out_81 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6031 = _T_6030 | _T_5776; // @[Mux.scala 27:72]
  wire [21:0] _T_5777 = _T_4323 ? btb_bank0_rd_data_way1_out_82 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6032 = _T_6031 | _T_5777; // @[Mux.scala 27:72]
  wire [21:0] _T_5778 = _T_4325 ? btb_bank0_rd_data_way1_out_83 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6033 = _T_6032 | _T_5778; // @[Mux.scala 27:72]
  wire [21:0] _T_5779 = _T_4327 ? btb_bank0_rd_data_way1_out_84 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6034 = _T_6033 | _T_5779; // @[Mux.scala 27:72]
  wire [21:0] _T_5780 = _T_4329 ? btb_bank0_rd_data_way1_out_85 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6035 = _T_6034 | _T_5780; // @[Mux.scala 27:72]
  wire [21:0] _T_5781 = _T_4331 ? btb_bank0_rd_data_way1_out_86 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6036 = _T_6035 | _T_5781; // @[Mux.scala 27:72]
  wire [21:0] _T_5782 = _T_4333 ? btb_bank0_rd_data_way1_out_87 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6037 = _T_6036 | _T_5782; // @[Mux.scala 27:72]
  wire [21:0] _T_5783 = _T_4335 ? btb_bank0_rd_data_way1_out_88 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6038 = _T_6037 | _T_5783; // @[Mux.scala 27:72]
  wire [21:0] _T_5784 = _T_4337 ? btb_bank0_rd_data_way1_out_89 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6039 = _T_6038 | _T_5784; // @[Mux.scala 27:72]
  wire [21:0] _T_5785 = _T_4339 ? btb_bank0_rd_data_way1_out_90 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6040 = _T_6039 | _T_5785; // @[Mux.scala 27:72]
  wire [21:0] _T_5786 = _T_4341 ? btb_bank0_rd_data_way1_out_91 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6041 = _T_6040 | _T_5786; // @[Mux.scala 27:72]
  wire [21:0] _T_5787 = _T_4343 ? btb_bank0_rd_data_way1_out_92 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6042 = _T_6041 | _T_5787; // @[Mux.scala 27:72]
  wire [21:0] _T_5788 = _T_4345 ? btb_bank0_rd_data_way1_out_93 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6043 = _T_6042 | _T_5788; // @[Mux.scala 27:72]
  wire [21:0] _T_5789 = _T_4347 ? btb_bank0_rd_data_way1_out_94 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6044 = _T_6043 | _T_5789; // @[Mux.scala 27:72]
  wire [21:0] _T_5790 = _T_4349 ? btb_bank0_rd_data_way1_out_95 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6045 = _T_6044 | _T_5790; // @[Mux.scala 27:72]
  wire [21:0] _T_5791 = _T_4351 ? btb_bank0_rd_data_way1_out_96 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6046 = _T_6045 | _T_5791; // @[Mux.scala 27:72]
  wire [21:0] _T_5792 = _T_4353 ? btb_bank0_rd_data_way1_out_97 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6047 = _T_6046 | _T_5792; // @[Mux.scala 27:72]
  wire [21:0] _T_5793 = _T_4355 ? btb_bank0_rd_data_way1_out_98 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6048 = _T_6047 | _T_5793; // @[Mux.scala 27:72]
  wire [21:0] _T_5794 = _T_4357 ? btb_bank0_rd_data_way1_out_99 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6049 = _T_6048 | _T_5794; // @[Mux.scala 27:72]
  wire [21:0] _T_5795 = _T_4359 ? btb_bank0_rd_data_way1_out_100 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6050 = _T_6049 | _T_5795; // @[Mux.scala 27:72]
  wire [21:0] _T_5796 = _T_4361 ? btb_bank0_rd_data_way1_out_101 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6051 = _T_6050 | _T_5796; // @[Mux.scala 27:72]
  wire [21:0] _T_5797 = _T_4363 ? btb_bank0_rd_data_way1_out_102 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6052 = _T_6051 | _T_5797; // @[Mux.scala 27:72]
  wire [21:0] _T_5798 = _T_4365 ? btb_bank0_rd_data_way1_out_103 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6053 = _T_6052 | _T_5798; // @[Mux.scala 27:72]
  wire [21:0] _T_5799 = _T_4367 ? btb_bank0_rd_data_way1_out_104 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6054 = _T_6053 | _T_5799; // @[Mux.scala 27:72]
  wire [21:0] _T_5800 = _T_4369 ? btb_bank0_rd_data_way1_out_105 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6055 = _T_6054 | _T_5800; // @[Mux.scala 27:72]
  wire [21:0] _T_5801 = _T_4371 ? btb_bank0_rd_data_way1_out_106 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6056 = _T_6055 | _T_5801; // @[Mux.scala 27:72]
  wire [21:0] _T_5802 = _T_4373 ? btb_bank0_rd_data_way1_out_107 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6057 = _T_6056 | _T_5802; // @[Mux.scala 27:72]
  wire [21:0] _T_5803 = _T_4375 ? btb_bank0_rd_data_way1_out_108 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6058 = _T_6057 | _T_5803; // @[Mux.scala 27:72]
  wire [21:0] _T_5804 = _T_4377 ? btb_bank0_rd_data_way1_out_109 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6059 = _T_6058 | _T_5804; // @[Mux.scala 27:72]
  wire [21:0] _T_5805 = _T_4379 ? btb_bank0_rd_data_way1_out_110 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6060 = _T_6059 | _T_5805; // @[Mux.scala 27:72]
  wire [21:0] _T_5806 = _T_4381 ? btb_bank0_rd_data_way1_out_111 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6061 = _T_6060 | _T_5806; // @[Mux.scala 27:72]
  wire [21:0] _T_5807 = _T_4383 ? btb_bank0_rd_data_way1_out_112 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6062 = _T_6061 | _T_5807; // @[Mux.scala 27:72]
  wire [21:0] _T_5808 = _T_4385 ? btb_bank0_rd_data_way1_out_113 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6063 = _T_6062 | _T_5808; // @[Mux.scala 27:72]
  wire [21:0] _T_5809 = _T_4387 ? btb_bank0_rd_data_way1_out_114 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6064 = _T_6063 | _T_5809; // @[Mux.scala 27:72]
  wire [21:0] _T_5810 = _T_4389 ? btb_bank0_rd_data_way1_out_115 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6065 = _T_6064 | _T_5810; // @[Mux.scala 27:72]
  wire [21:0] _T_5811 = _T_4391 ? btb_bank0_rd_data_way1_out_116 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6066 = _T_6065 | _T_5811; // @[Mux.scala 27:72]
  wire [21:0] _T_5812 = _T_4393 ? btb_bank0_rd_data_way1_out_117 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6067 = _T_6066 | _T_5812; // @[Mux.scala 27:72]
  wire [21:0] _T_5813 = _T_4395 ? btb_bank0_rd_data_way1_out_118 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6068 = _T_6067 | _T_5813; // @[Mux.scala 27:72]
  wire [21:0] _T_5814 = _T_4397 ? btb_bank0_rd_data_way1_out_119 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6069 = _T_6068 | _T_5814; // @[Mux.scala 27:72]
  wire [21:0] _T_5815 = _T_4399 ? btb_bank0_rd_data_way1_out_120 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6070 = _T_6069 | _T_5815; // @[Mux.scala 27:72]
  wire [21:0] _T_5816 = _T_4401 ? btb_bank0_rd_data_way1_out_121 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6071 = _T_6070 | _T_5816; // @[Mux.scala 27:72]
  wire [21:0] _T_5817 = _T_4403 ? btb_bank0_rd_data_way1_out_122 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6072 = _T_6071 | _T_5817; // @[Mux.scala 27:72]
  wire [21:0] _T_5818 = _T_4405 ? btb_bank0_rd_data_way1_out_123 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6073 = _T_6072 | _T_5818; // @[Mux.scala 27:72]
  wire [21:0] _T_5819 = _T_4407 ? btb_bank0_rd_data_way1_out_124 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6074 = _T_6073 | _T_5819; // @[Mux.scala 27:72]
  wire [21:0] _T_5820 = _T_4409 ? btb_bank0_rd_data_way1_out_125 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6075 = _T_6074 | _T_5820; // @[Mux.scala 27:72]
  wire [21:0] _T_5821 = _T_4411 ? btb_bank0_rd_data_way1_out_126 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6076 = _T_6075 | _T_5821; // @[Mux.scala 27:72]
  wire [21:0] _T_5822 = _T_4413 ? btb_bank0_rd_data_way1_out_127 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6077 = _T_6076 | _T_5822; // @[Mux.scala 27:72]
  wire [21:0] _T_5823 = _T_4415 ? btb_bank0_rd_data_way1_out_128 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6078 = _T_6077 | _T_5823; // @[Mux.scala 27:72]
  wire [21:0] _T_5824 = _T_4417 ? btb_bank0_rd_data_way1_out_129 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6079 = _T_6078 | _T_5824; // @[Mux.scala 27:72]
  wire [21:0] _T_5825 = _T_4419 ? btb_bank0_rd_data_way1_out_130 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6080 = _T_6079 | _T_5825; // @[Mux.scala 27:72]
  wire [21:0] _T_5826 = _T_4421 ? btb_bank0_rd_data_way1_out_131 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6081 = _T_6080 | _T_5826; // @[Mux.scala 27:72]
  wire [21:0] _T_5827 = _T_4423 ? btb_bank0_rd_data_way1_out_132 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6082 = _T_6081 | _T_5827; // @[Mux.scala 27:72]
  wire [21:0] _T_5828 = _T_4425 ? btb_bank0_rd_data_way1_out_133 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6083 = _T_6082 | _T_5828; // @[Mux.scala 27:72]
  wire [21:0] _T_5829 = _T_4427 ? btb_bank0_rd_data_way1_out_134 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6084 = _T_6083 | _T_5829; // @[Mux.scala 27:72]
  wire [21:0] _T_5830 = _T_4429 ? btb_bank0_rd_data_way1_out_135 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6085 = _T_6084 | _T_5830; // @[Mux.scala 27:72]
  wire [21:0] _T_5831 = _T_4431 ? btb_bank0_rd_data_way1_out_136 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6086 = _T_6085 | _T_5831; // @[Mux.scala 27:72]
  wire [21:0] _T_5832 = _T_4433 ? btb_bank0_rd_data_way1_out_137 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6087 = _T_6086 | _T_5832; // @[Mux.scala 27:72]
  wire [21:0] _T_5833 = _T_4435 ? btb_bank0_rd_data_way1_out_138 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6088 = _T_6087 | _T_5833; // @[Mux.scala 27:72]
  wire [21:0] _T_5834 = _T_4437 ? btb_bank0_rd_data_way1_out_139 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6089 = _T_6088 | _T_5834; // @[Mux.scala 27:72]
  wire [21:0] _T_5835 = _T_4439 ? btb_bank0_rd_data_way1_out_140 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6090 = _T_6089 | _T_5835; // @[Mux.scala 27:72]
  wire [21:0] _T_5836 = _T_4441 ? btb_bank0_rd_data_way1_out_141 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6091 = _T_6090 | _T_5836; // @[Mux.scala 27:72]
  wire [21:0] _T_5837 = _T_4443 ? btb_bank0_rd_data_way1_out_142 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6092 = _T_6091 | _T_5837; // @[Mux.scala 27:72]
  wire [21:0] _T_5838 = _T_4445 ? btb_bank0_rd_data_way1_out_143 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6093 = _T_6092 | _T_5838; // @[Mux.scala 27:72]
  wire [21:0] _T_5839 = _T_4447 ? btb_bank0_rd_data_way1_out_144 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6094 = _T_6093 | _T_5839; // @[Mux.scala 27:72]
  wire [21:0] _T_5840 = _T_4449 ? btb_bank0_rd_data_way1_out_145 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6095 = _T_6094 | _T_5840; // @[Mux.scala 27:72]
  wire [21:0] _T_5841 = _T_4451 ? btb_bank0_rd_data_way1_out_146 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6096 = _T_6095 | _T_5841; // @[Mux.scala 27:72]
  wire [21:0] _T_5842 = _T_4453 ? btb_bank0_rd_data_way1_out_147 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6097 = _T_6096 | _T_5842; // @[Mux.scala 27:72]
  wire [21:0] _T_5843 = _T_4455 ? btb_bank0_rd_data_way1_out_148 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6098 = _T_6097 | _T_5843; // @[Mux.scala 27:72]
  wire [21:0] _T_5844 = _T_4457 ? btb_bank0_rd_data_way1_out_149 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6099 = _T_6098 | _T_5844; // @[Mux.scala 27:72]
  wire [21:0] _T_5845 = _T_4459 ? btb_bank0_rd_data_way1_out_150 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6100 = _T_6099 | _T_5845; // @[Mux.scala 27:72]
  wire [21:0] _T_5846 = _T_4461 ? btb_bank0_rd_data_way1_out_151 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6101 = _T_6100 | _T_5846; // @[Mux.scala 27:72]
  wire [21:0] _T_5847 = _T_4463 ? btb_bank0_rd_data_way1_out_152 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6102 = _T_6101 | _T_5847; // @[Mux.scala 27:72]
  wire [21:0] _T_5848 = _T_4465 ? btb_bank0_rd_data_way1_out_153 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6103 = _T_6102 | _T_5848; // @[Mux.scala 27:72]
  wire [21:0] _T_5849 = _T_4467 ? btb_bank0_rd_data_way1_out_154 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6104 = _T_6103 | _T_5849; // @[Mux.scala 27:72]
  wire [21:0] _T_5850 = _T_4469 ? btb_bank0_rd_data_way1_out_155 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6105 = _T_6104 | _T_5850; // @[Mux.scala 27:72]
  wire [21:0] _T_5851 = _T_4471 ? btb_bank0_rd_data_way1_out_156 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6106 = _T_6105 | _T_5851; // @[Mux.scala 27:72]
  wire [21:0] _T_5852 = _T_4473 ? btb_bank0_rd_data_way1_out_157 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6107 = _T_6106 | _T_5852; // @[Mux.scala 27:72]
  wire [21:0] _T_5853 = _T_4475 ? btb_bank0_rd_data_way1_out_158 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6108 = _T_6107 | _T_5853; // @[Mux.scala 27:72]
  wire [21:0] _T_5854 = _T_4477 ? btb_bank0_rd_data_way1_out_159 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6109 = _T_6108 | _T_5854; // @[Mux.scala 27:72]
  wire [21:0] _T_5855 = _T_4479 ? btb_bank0_rd_data_way1_out_160 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6110 = _T_6109 | _T_5855; // @[Mux.scala 27:72]
  wire [21:0] _T_5856 = _T_4481 ? btb_bank0_rd_data_way1_out_161 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6111 = _T_6110 | _T_5856; // @[Mux.scala 27:72]
  wire [21:0] _T_5857 = _T_4483 ? btb_bank0_rd_data_way1_out_162 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6112 = _T_6111 | _T_5857; // @[Mux.scala 27:72]
  wire [21:0] _T_5858 = _T_4485 ? btb_bank0_rd_data_way1_out_163 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6113 = _T_6112 | _T_5858; // @[Mux.scala 27:72]
  wire [21:0] _T_5859 = _T_4487 ? btb_bank0_rd_data_way1_out_164 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6114 = _T_6113 | _T_5859; // @[Mux.scala 27:72]
  wire [21:0] _T_5860 = _T_4489 ? btb_bank0_rd_data_way1_out_165 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6115 = _T_6114 | _T_5860; // @[Mux.scala 27:72]
  wire [21:0] _T_5861 = _T_4491 ? btb_bank0_rd_data_way1_out_166 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6116 = _T_6115 | _T_5861; // @[Mux.scala 27:72]
  wire [21:0] _T_5862 = _T_4493 ? btb_bank0_rd_data_way1_out_167 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6117 = _T_6116 | _T_5862; // @[Mux.scala 27:72]
  wire [21:0] _T_5863 = _T_4495 ? btb_bank0_rd_data_way1_out_168 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6118 = _T_6117 | _T_5863; // @[Mux.scala 27:72]
  wire [21:0] _T_5864 = _T_4497 ? btb_bank0_rd_data_way1_out_169 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6119 = _T_6118 | _T_5864; // @[Mux.scala 27:72]
  wire [21:0] _T_5865 = _T_4499 ? btb_bank0_rd_data_way1_out_170 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6120 = _T_6119 | _T_5865; // @[Mux.scala 27:72]
  wire [21:0] _T_5866 = _T_4501 ? btb_bank0_rd_data_way1_out_171 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6121 = _T_6120 | _T_5866; // @[Mux.scala 27:72]
  wire [21:0] _T_5867 = _T_4503 ? btb_bank0_rd_data_way1_out_172 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6122 = _T_6121 | _T_5867; // @[Mux.scala 27:72]
  wire [21:0] _T_5868 = _T_4505 ? btb_bank0_rd_data_way1_out_173 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6123 = _T_6122 | _T_5868; // @[Mux.scala 27:72]
  wire [21:0] _T_5869 = _T_4507 ? btb_bank0_rd_data_way1_out_174 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6124 = _T_6123 | _T_5869; // @[Mux.scala 27:72]
  wire [21:0] _T_5870 = _T_4509 ? btb_bank0_rd_data_way1_out_175 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6125 = _T_6124 | _T_5870; // @[Mux.scala 27:72]
  wire [21:0] _T_5871 = _T_4511 ? btb_bank0_rd_data_way1_out_176 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6126 = _T_6125 | _T_5871; // @[Mux.scala 27:72]
  wire [21:0] _T_5872 = _T_4513 ? btb_bank0_rd_data_way1_out_177 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6127 = _T_6126 | _T_5872; // @[Mux.scala 27:72]
  wire [21:0] _T_5873 = _T_4515 ? btb_bank0_rd_data_way1_out_178 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6128 = _T_6127 | _T_5873; // @[Mux.scala 27:72]
  wire [21:0] _T_5874 = _T_4517 ? btb_bank0_rd_data_way1_out_179 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6129 = _T_6128 | _T_5874; // @[Mux.scala 27:72]
  wire [21:0] _T_5875 = _T_4519 ? btb_bank0_rd_data_way1_out_180 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6130 = _T_6129 | _T_5875; // @[Mux.scala 27:72]
  wire [21:0] _T_5876 = _T_4521 ? btb_bank0_rd_data_way1_out_181 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6131 = _T_6130 | _T_5876; // @[Mux.scala 27:72]
  wire [21:0] _T_5877 = _T_4523 ? btb_bank0_rd_data_way1_out_182 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6132 = _T_6131 | _T_5877; // @[Mux.scala 27:72]
  wire [21:0] _T_5878 = _T_4525 ? btb_bank0_rd_data_way1_out_183 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6133 = _T_6132 | _T_5878; // @[Mux.scala 27:72]
  wire [21:0] _T_5879 = _T_4527 ? btb_bank0_rd_data_way1_out_184 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6134 = _T_6133 | _T_5879; // @[Mux.scala 27:72]
  wire [21:0] _T_5880 = _T_4529 ? btb_bank0_rd_data_way1_out_185 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6135 = _T_6134 | _T_5880; // @[Mux.scala 27:72]
  wire [21:0] _T_5881 = _T_4531 ? btb_bank0_rd_data_way1_out_186 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6136 = _T_6135 | _T_5881; // @[Mux.scala 27:72]
  wire [21:0] _T_5882 = _T_4533 ? btb_bank0_rd_data_way1_out_187 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6137 = _T_6136 | _T_5882; // @[Mux.scala 27:72]
  wire [21:0] _T_5883 = _T_4535 ? btb_bank0_rd_data_way1_out_188 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6138 = _T_6137 | _T_5883; // @[Mux.scala 27:72]
  wire [21:0] _T_5884 = _T_4537 ? btb_bank0_rd_data_way1_out_189 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6139 = _T_6138 | _T_5884; // @[Mux.scala 27:72]
  wire [21:0] _T_5885 = _T_4539 ? btb_bank0_rd_data_way1_out_190 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6140 = _T_6139 | _T_5885; // @[Mux.scala 27:72]
  wire [21:0] _T_5886 = _T_4541 ? btb_bank0_rd_data_way1_out_191 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6141 = _T_6140 | _T_5886; // @[Mux.scala 27:72]
  wire [21:0] _T_5887 = _T_4543 ? btb_bank0_rd_data_way1_out_192 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6142 = _T_6141 | _T_5887; // @[Mux.scala 27:72]
  wire [21:0] _T_5888 = _T_4545 ? btb_bank0_rd_data_way1_out_193 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6143 = _T_6142 | _T_5888; // @[Mux.scala 27:72]
  wire [21:0] _T_5889 = _T_4547 ? btb_bank0_rd_data_way1_out_194 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6144 = _T_6143 | _T_5889; // @[Mux.scala 27:72]
  wire [21:0] _T_5890 = _T_4549 ? btb_bank0_rd_data_way1_out_195 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6145 = _T_6144 | _T_5890; // @[Mux.scala 27:72]
  wire [21:0] _T_5891 = _T_4551 ? btb_bank0_rd_data_way1_out_196 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6146 = _T_6145 | _T_5891; // @[Mux.scala 27:72]
  wire [21:0] _T_5892 = _T_4553 ? btb_bank0_rd_data_way1_out_197 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6147 = _T_6146 | _T_5892; // @[Mux.scala 27:72]
  wire [21:0] _T_5893 = _T_4555 ? btb_bank0_rd_data_way1_out_198 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6148 = _T_6147 | _T_5893; // @[Mux.scala 27:72]
  wire [21:0] _T_5894 = _T_4557 ? btb_bank0_rd_data_way1_out_199 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6149 = _T_6148 | _T_5894; // @[Mux.scala 27:72]
  wire [21:0] _T_5895 = _T_4559 ? btb_bank0_rd_data_way1_out_200 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6150 = _T_6149 | _T_5895; // @[Mux.scala 27:72]
  wire [21:0] _T_5896 = _T_4561 ? btb_bank0_rd_data_way1_out_201 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6151 = _T_6150 | _T_5896; // @[Mux.scala 27:72]
  wire [21:0] _T_5897 = _T_4563 ? btb_bank0_rd_data_way1_out_202 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6152 = _T_6151 | _T_5897; // @[Mux.scala 27:72]
  wire [21:0] _T_5898 = _T_4565 ? btb_bank0_rd_data_way1_out_203 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6153 = _T_6152 | _T_5898; // @[Mux.scala 27:72]
  wire [21:0] _T_5899 = _T_4567 ? btb_bank0_rd_data_way1_out_204 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6154 = _T_6153 | _T_5899; // @[Mux.scala 27:72]
  wire [21:0] _T_5900 = _T_4569 ? btb_bank0_rd_data_way1_out_205 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6155 = _T_6154 | _T_5900; // @[Mux.scala 27:72]
  wire [21:0] _T_5901 = _T_4571 ? btb_bank0_rd_data_way1_out_206 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6156 = _T_6155 | _T_5901; // @[Mux.scala 27:72]
  wire [21:0] _T_5902 = _T_4573 ? btb_bank0_rd_data_way1_out_207 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6157 = _T_6156 | _T_5902; // @[Mux.scala 27:72]
  wire [21:0] _T_5903 = _T_4575 ? btb_bank0_rd_data_way1_out_208 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6158 = _T_6157 | _T_5903; // @[Mux.scala 27:72]
  wire [21:0] _T_5904 = _T_4577 ? btb_bank0_rd_data_way1_out_209 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6159 = _T_6158 | _T_5904; // @[Mux.scala 27:72]
  wire [21:0] _T_5905 = _T_4579 ? btb_bank0_rd_data_way1_out_210 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6160 = _T_6159 | _T_5905; // @[Mux.scala 27:72]
  wire [21:0] _T_5906 = _T_4581 ? btb_bank0_rd_data_way1_out_211 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6161 = _T_6160 | _T_5906; // @[Mux.scala 27:72]
  wire [21:0] _T_5907 = _T_4583 ? btb_bank0_rd_data_way1_out_212 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6162 = _T_6161 | _T_5907; // @[Mux.scala 27:72]
  wire [21:0] _T_5908 = _T_4585 ? btb_bank0_rd_data_way1_out_213 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6163 = _T_6162 | _T_5908; // @[Mux.scala 27:72]
  wire [21:0] _T_5909 = _T_4587 ? btb_bank0_rd_data_way1_out_214 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6164 = _T_6163 | _T_5909; // @[Mux.scala 27:72]
  wire [21:0] _T_5910 = _T_4589 ? btb_bank0_rd_data_way1_out_215 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6165 = _T_6164 | _T_5910; // @[Mux.scala 27:72]
  wire [21:0] _T_5911 = _T_4591 ? btb_bank0_rd_data_way1_out_216 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6166 = _T_6165 | _T_5911; // @[Mux.scala 27:72]
  wire [21:0] _T_5912 = _T_4593 ? btb_bank0_rd_data_way1_out_217 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6167 = _T_6166 | _T_5912; // @[Mux.scala 27:72]
  wire [21:0] _T_5913 = _T_4595 ? btb_bank0_rd_data_way1_out_218 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6168 = _T_6167 | _T_5913; // @[Mux.scala 27:72]
  wire [21:0] _T_5914 = _T_4597 ? btb_bank0_rd_data_way1_out_219 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6169 = _T_6168 | _T_5914; // @[Mux.scala 27:72]
  wire [21:0] _T_5915 = _T_4599 ? btb_bank0_rd_data_way1_out_220 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6170 = _T_6169 | _T_5915; // @[Mux.scala 27:72]
  wire [21:0] _T_5916 = _T_4601 ? btb_bank0_rd_data_way1_out_221 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6171 = _T_6170 | _T_5916; // @[Mux.scala 27:72]
  wire [21:0] _T_5917 = _T_4603 ? btb_bank0_rd_data_way1_out_222 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6172 = _T_6171 | _T_5917; // @[Mux.scala 27:72]
  wire [21:0] _T_5918 = _T_4605 ? btb_bank0_rd_data_way1_out_223 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6173 = _T_6172 | _T_5918; // @[Mux.scala 27:72]
  wire [21:0] _T_5919 = _T_4607 ? btb_bank0_rd_data_way1_out_224 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6174 = _T_6173 | _T_5919; // @[Mux.scala 27:72]
  wire [21:0] _T_5920 = _T_4609 ? btb_bank0_rd_data_way1_out_225 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6175 = _T_6174 | _T_5920; // @[Mux.scala 27:72]
  wire [21:0] _T_5921 = _T_4611 ? btb_bank0_rd_data_way1_out_226 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6176 = _T_6175 | _T_5921; // @[Mux.scala 27:72]
  wire [21:0] _T_5922 = _T_4613 ? btb_bank0_rd_data_way1_out_227 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6177 = _T_6176 | _T_5922; // @[Mux.scala 27:72]
  wire [21:0] _T_5923 = _T_4615 ? btb_bank0_rd_data_way1_out_228 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6178 = _T_6177 | _T_5923; // @[Mux.scala 27:72]
  wire [21:0] _T_5924 = _T_4617 ? btb_bank0_rd_data_way1_out_229 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6179 = _T_6178 | _T_5924; // @[Mux.scala 27:72]
  wire [21:0] _T_5925 = _T_4619 ? btb_bank0_rd_data_way1_out_230 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6180 = _T_6179 | _T_5925; // @[Mux.scala 27:72]
  wire [21:0] _T_5926 = _T_4621 ? btb_bank0_rd_data_way1_out_231 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6181 = _T_6180 | _T_5926; // @[Mux.scala 27:72]
  wire [21:0] _T_5927 = _T_4623 ? btb_bank0_rd_data_way1_out_232 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6182 = _T_6181 | _T_5927; // @[Mux.scala 27:72]
  wire [21:0] _T_5928 = _T_4625 ? btb_bank0_rd_data_way1_out_233 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6183 = _T_6182 | _T_5928; // @[Mux.scala 27:72]
  wire [21:0] _T_5929 = _T_4627 ? btb_bank0_rd_data_way1_out_234 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6184 = _T_6183 | _T_5929; // @[Mux.scala 27:72]
  wire [21:0] _T_5930 = _T_4629 ? btb_bank0_rd_data_way1_out_235 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6185 = _T_6184 | _T_5930; // @[Mux.scala 27:72]
  wire [21:0] _T_5931 = _T_4631 ? btb_bank0_rd_data_way1_out_236 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6186 = _T_6185 | _T_5931; // @[Mux.scala 27:72]
  wire [21:0] _T_5932 = _T_4633 ? btb_bank0_rd_data_way1_out_237 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6187 = _T_6186 | _T_5932; // @[Mux.scala 27:72]
  wire [21:0] _T_5933 = _T_4635 ? btb_bank0_rd_data_way1_out_238 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6188 = _T_6187 | _T_5933; // @[Mux.scala 27:72]
  wire [21:0] _T_5934 = _T_4637 ? btb_bank0_rd_data_way1_out_239 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6189 = _T_6188 | _T_5934; // @[Mux.scala 27:72]
  wire [21:0] _T_5935 = _T_4639 ? btb_bank0_rd_data_way1_out_240 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6190 = _T_6189 | _T_5935; // @[Mux.scala 27:72]
  wire [21:0] _T_5936 = _T_4641 ? btb_bank0_rd_data_way1_out_241 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6191 = _T_6190 | _T_5936; // @[Mux.scala 27:72]
  wire [21:0] _T_5937 = _T_4643 ? btb_bank0_rd_data_way1_out_242 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6192 = _T_6191 | _T_5937; // @[Mux.scala 27:72]
  wire [21:0] _T_5938 = _T_4645 ? btb_bank0_rd_data_way1_out_243 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6193 = _T_6192 | _T_5938; // @[Mux.scala 27:72]
  wire [21:0] _T_5939 = _T_4647 ? btb_bank0_rd_data_way1_out_244 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6194 = _T_6193 | _T_5939; // @[Mux.scala 27:72]
  wire [21:0] _T_5940 = _T_4649 ? btb_bank0_rd_data_way1_out_245 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6195 = _T_6194 | _T_5940; // @[Mux.scala 27:72]
  wire [21:0] _T_5941 = _T_4651 ? btb_bank0_rd_data_way1_out_246 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6196 = _T_6195 | _T_5941; // @[Mux.scala 27:72]
  wire [21:0] _T_5942 = _T_4653 ? btb_bank0_rd_data_way1_out_247 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6197 = _T_6196 | _T_5942; // @[Mux.scala 27:72]
  wire [21:0] _T_5943 = _T_4655 ? btb_bank0_rd_data_way1_out_248 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6198 = _T_6197 | _T_5943; // @[Mux.scala 27:72]
  wire [21:0] _T_5944 = _T_4657 ? btb_bank0_rd_data_way1_out_249 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6199 = _T_6198 | _T_5944; // @[Mux.scala 27:72]
  wire [21:0] _T_5945 = _T_4659 ? btb_bank0_rd_data_way1_out_250 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6200 = _T_6199 | _T_5945; // @[Mux.scala 27:72]
  wire [21:0] _T_5946 = _T_4661 ? btb_bank0_rd_data_way1_out_251 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6201 = _T_6200 | _T_5946; // @[Mux.scala 27:72]
  wire [21:0] _T_5947 = _T_4663 ? btb_bank0_rd_data_way1_out_252 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6202 = _T_6201 | _T_5947; // @[Mux.scala 27:72]
  wire [21:0] _T_5948 = _T_4665 ? btb_bank0_rd_data_way1_out_253 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6203 = _T_6202 | _T_5948; // @[Mux.scala 27:72]
  wire [21:0] _T_5949 = _T_4667 ? btb_bank0_rd_data_way1_out_254 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6204 = _T_6203 | _T_5949; // @[Mux.scala 27:72]
  wire [21:0] _T_5950 = _T_4669 ? btb_bank0_rd_data_way1_out_255 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] btb_bank0_rd_data_way1_p1_f = _T_6204 | _T_5950; // @[Mux.scala 27:72]
  wire  _T_72 = btb_bank0_rd_data_way1_p1_f[21:17] == fetch_rd_tag_p1_f; // @[el2_ifu_bp_ctl.scala 150:106]
  wire  _T_73 = btb_bank0_rd_data_way1_p1_f[0] & _T_72; // @[el2_ifu_bp_ctl.scala 150:61]
  wire  _T_76 = _T_73 & _T_48; // @[el2_ifu_bp_ctl.scala 150:129]
  wire  _T_77 = _T_76 & io_ifc_fetch_req_f; // @[el2_ifu_bp_ctl.scala 151:56]
  wire  tag_match_way1_p1_f = _T_77 & _T; // @[el2_ifu_bp_ctl.scala 151:77]
  wire  _T_108 = btb_bank0_rd_data_way1_p1_f[3] ^ btb_bank0_rd_data_way1_p1_f[4]; // @[el2_ifu_bp_ctl.scala 163:100]
  wire  _T_109 = tag_match_way1_p1_f & _T_108; // @[el2_ifu_bp_ctl.scala 163:62]
  wire  _T_113 = ~_T_108; // @[el2_ifu_bp_ctl.scala 164:64]
  wire  _T_114 = tag_match_way1_p1_f & _T_113; // @[el2_ifu_bp_ctl.scala 164:62]
  wire [1:0] tag_match_way1_expanded_p1_f = {_T_109,_T_114}; // @[Cat.scala 29:58]
  wire [21:0] _T_134 = tag_match_way1_expanded_p1_f[0] ? btb_bank0_rd_data_way1_p1_f : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] btb_bank0e_rd_data_p1_f = _T_133 | _T_134; // @[Mux.scala 27:72]
  wire [21:0] _T_146 = io_ifc_fetch_addr_f[0] ? btb_bank0e_rd_data_p1_f : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] btb_vbank1_rd_data_f = _T_145 | _T_146; // @[Mux.scala 27:72]
  wire  _T_242 = btb_vbank1_rd_data_f[2] | btb_vbank1_rd_data_f[1]; // @[el2_ifu_bp_ctl.scala 276:59]
  wire [21:0] _T_119 = tag_match_way0_expanded_f[0] ? btb_bank0_rd_data_way0_f : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_120 = tag_match_way1_expanded_f[0] ? btb_bank0_rd_data_way1_f : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] btb_bank0e_rd_data_f = _T_119 | _T_120; // @[Mux.scala 27:72]
  wire [21:0] _T_139 = _T_143 ? btb_bank0e_rd_data_f : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_140 = io_ifc_fetch_addr_f[0] ? btb_bank0o_rd_data_f : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] btb_vbank0_rd_data_f = _T_139 | _T_140; // @[Mux.scala 27:72]
  wire  _T_245 = btb_vbank0_rd_data_f[2] | btb_vbank0_rd_data_f[1]; // @[el2_ifu_bp_ctl.scala 277:59]
  wire [1:0] bht_force_taken_f = {_T_242,_T_245}; // @[Cat.scala 29:58]
  wire [9:0] _T_569 = {btb_rd_addr_f,2'h0}; // @[Cat.scala 29:58]
  reg [7:0] fghr; // @[el2_ifu_bp_ctl.scala 335:44]
  wire [7:0] bht_rd_addr_hashed_f = _T_569[9:2] ^ fghr; // @[el2_lib.scala 194:35]
  wire  _T_21407 = bht_rd_addr_hashed_f == 8'h0; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_0; // @[Reg.scala 27:20]
  wire [1:0] _T_21919 = _T_21407 ? bht_bank_rd_data_out_1_0 : 2'h0; // @[Mux.scala 27:72]
  wire  _T_21409 = bht_rd_addr_hashed_f == 8'h1; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_1; // @[Reg.scala 27:20]
  wire [1:0] _T_21920 = _T_21409 ? bht_bank_rd_data_out_1_1 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22175 = _T_21919 | _T_21920; // @[Mux.scala 27:72]
  wire  _T_21411 = bht_rd_addr_hashed_f == 8'h2; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_2; // @[Reg.scala 27:20]
  wire [1:0] _T_21921 = _T_21411 ? bht_bank_rd_data_out_1_2 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22176 = _T_22175 | _T_21921; // @[Mux.scala 27:72]
  wire  _T_21413 = bht_rd_addr_hashed_f == 8'h3; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_3; // @[Reg.scala 27:20]
  wire [1:0] _T_21922 = _T_21413 ? bht_bank_rd_data_out_1_3 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22177 = _T_22176 | _T_21922; // @[Mux.scala 27:72]
  wire  _T_21415 = bht_rd_addr_hashed_f == 8'h4; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_4; // @[Reg.scala 27:20]
  wire [1:0] _T_21923 = _T_21415 ? bht_bank_rd_data_out_1_4 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22178 = _T_22177 | _T_21923; // @[Mux.scala 27:72]
  wire  _T_21417 = bht_rd_addr_hashed_f == 8'h5; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_5; // @[Reg.scala 27:20]
  wire [1:0] _T_21924 = _T_21417 ? bht_bank_rd_data_out_1_5 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22179 = _T_22178 | _T_21924; // @[Mux.scala 27:72]
  wire  _T_21419 = bht_rd_addr_hashed_f == 8'h6; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_6; // @[Reg.scala 27:20]
  wire [1:0] _T_21925 = _T_21419 ? bht_bank_rd_data_out_1_6 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22180 = _T_22179 | _T_21925; // @[Mux.scala 27:72]
  wire  _T_21421 = bht_rd_addr_hashed_f == 8'h7; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_7; // @[Reg.scala 27:20]
  wire [1:0] _T_21926 = _T_21421 ? bht_bank_rd_data_out_1_7 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22181 = _T_22180 | _T_21926; // @[Mux.scala 27:72]
  wire  _T_21423 = bht_rd_addr_hashed_f == 8'h8; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_8; // @[Reg.scala 27:20]
  wire [1:0] _T_21927 = _T_21423 ? bht_bank_rd_data_out_1_8 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22182 = _T_22181 | _T_21927; // @[Mux.scala 27:72]
  wire  _T_21425 = bht_rd_addr_hashed_f == 8'h9; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_9; // @[Reg.scala 27:20]
  wire [1:0] _T_21928 = _T_21425 ? bht_bank_rd_data_out_1_9 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22183 = _T_22182 | _T_21928; // @[Mux.scala 27:72]
  wire  _T_21427 = bht_rd_addr_hashed_f == 8'ha; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_10; // @[Reg.scala 27:20]
  wire [1:0] _T_21929 = _T_21427 ? bht_bank_rd_data_out_1_10 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22184 = _T_22183 | _T_21929; // @[Mux.scala 27:72]
  wire  _T_21429 = bht_rd_addr_hashed_f == 8'hb; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_11; // @[Reg.scala 27:20]
  wire [1:0] _T_21930 = _T_21429 ? bht_bank_rd_data_out_1_11 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22185 = _T_22184 | _T_21930; // @[Mux.scala 27:72]
  wire  _T_21431 = bht_rd_addr_hashed_f == 8'hc; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_12; // @[Reg.scala 27:20]
  wire [1:0] _T_21931 = _T_21431 ? bht_bank_rd_data_out_1_12 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22186 = _T_22185 | _T_21931; // @[Mux.scala 27:72]
  wire  _T_21433 = bht_rd_addr_hashed_f == 8'hd; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_13; // @[Reg.scala 27:20]
  wire [1:0] _T_21932 = _T_21433 ? bht_bank_rd_data_out_1_13 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22187 = _T_22186 | _T_21932; // @[Mux.scala 27:72]
  wire  _T_21435 = bht_rd_addr_hashed_f == 8'he; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_14; // @[Reg.scala 27:20]
  wire [1:0] _T_21933 = _T_21435 ? bht_bank_rd_data_out_1_14 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22188 = _T_22187 | _T_21933; // @[Mux.scala 27:72]
  wire  _T_21437 = bht_rd_addr_hashed_f == 8'hf; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_15; // @[Reg.scala 27:20]
  wire [1:0] _T_21934 = _T_21437 ? bht_bank_rd_data_out_1_15 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22189 = _T_22188 | _T_21934; // @[Mux.scala 27:72]
  wire  _T_21439 = bht_rd_addr_hashed_f == 8'h10; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_16; // @[Reg.scala 27:20]
  wire [1:0] _T_21935 = _T_21439 ? bht_bank_rd_data_out_1_16 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22190 = _T_22189 | _T_21935; // @[Mux.scala 27:72]
  wire  _T_21441 = bht_rd_addr_hashed_f == 8'h11; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_17; // @[Reg.scala 27:20]
  wire [1:0] _T_21936 = _T_21441 ? bht_bank_rd_data_out_1_17 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22191 = _T_22190 | _T_21936; // @[Mux.scala 27:72]
  wire  _T_21443 = bht_rd_addr_hashed_f == 8'h12; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_18; // @[Reg.scala 27:20]
  wire [1:0] _T_21937 = _T_21443 ? bht_bank_rd_data_out_1_18 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22192 = _T_22191 | _T_21937; // @[Mux.scala 27:72]
  wire  _T_21445 = bht_rd_addr_hashed_f == 8'h13; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_19; // @[Reg.scala 27:20]
  wire [1:0] _T_21938 = _T_21445 ? bht_bank_rd_data_out_1_19 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22193 = _T_22192 | _T_21938; // @[Mux.scala 27:72]
  wire  _T_21447 = bht_rd_addr_hashed_f == 8'h14; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_20; // @[Reg.scala 27:20]
  wire [1:0] _T_21939 = _T_21447 ? bht_bank_rd_data_out_1_20 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22194 = _T_22193 | _T_21939; // @[Mux.scala 27:72]
  wire  _T_21449 = bht_rd_addr_hashed_f == 8'h15; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_21; // @[Reg.scala 27:20]
  wire [1:0] _T_21940 = _T_21449 ? bht_bank_rd_data_out_1_21 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22195 = _T_22194 | _T_21940; // @[Mux.scala 27:72]
  wire  _T_21451 = bht_rd_addr_hashed_f == 8'h16; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_22; // @[Reg.scala 27:20]
  wire [1:0] _T_21941 = _T_21451 ? bht_bank_rd_data_out_1_22 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22196 = _T_22195 | _T_21941; // @[Mux.scala 27:72]
  wire  _T_21453 = bht_rd_addr_hashed_f == 8'h17; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_23; // @[Reg.scala 27:20]
  wire [1:0] _T_21942 = _T_21453 ? bht_bank_rd_data_out_1_23 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22197 = _T_22196 | _T_21942; // @[Mux.scala 27:72]
  wire  _T_21455 = bht_rd_addr_hashed_f == 8'h18; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_24; // @[Reg.scala 27:20]
  wire [1:0] _T_21943 = _T_21455 ? bht_bank_rd_data_out_1_24 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22198 = _T_22197 | _T_21943; // @[Mux.scala 27:72]
  wire  _T_21457 = bht_rd_addr_hashed_f == 8'h19; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_25; // @[Reg.scala 27:20]
  wire [1:0] _T_21944 = _T_21457 ? bht_bank_rd_data_out_1_25 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22199 = _T_22198 | _T_21944; // @[Mux.scala 27:72]
  wire  _T_21459 = bht_rd_addr_hashed_f == 8'h1a; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_26; // @[Reg.scala 27:20]
  wire [1:0] _T_21945 = _T_21459 ? bht_bank_rd_data_out_1_26 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22200 = _T_22199 | _T_21945; // @[Mux.scala 27:72]
  wire  _T_21461 = bht_rd_addr_hashed_f == 8'h1b; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_27; // @[Reg.scala 27:20]
  wire [1:0] _T_21946 = _T_21461 ? bht_bank_rd_data_out_1_27 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22201 = _T_22200 | _T_21946; // @[Mux.scala 27:72]
  wire  _T_21463 = bht_rd_addr_hashed_f == 8'h1c; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_28; // @[Reg.scala 27:20]
  wire [1:0] _T_21947 = _T_21463 ? bht_bank_rd_data_out_1_28 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22202 = _T_22201 | _T_21947; // @[Mux.scala 27:72]
  wire  _T_21465 = bht_rd_addr_hashed_f == 8'h1d; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_29; // @[Reg.scala 27:20]
  wire [1:0] _T_21948 = _T_21465 ? bht_bank_rd_data_out_1_29 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22203 = _T_22202 | _T_21948; // @[Mux.scala 27:72]
  wire  _T_21467 = bht_rd_addr_hashed_f == 8'h1e; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_30; // @[Reg.scala 27:20]
  wire [1:0] _T_21949 = _T_21467 ? bht_bank_rd_data_out_1_30 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22204 = _T_22203 | _T_21949; // @[Mux.scala 27:72]
  wire  _T_21469 = bht_rd_addr_hashed_f == 8'h1f; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_31; // @[Reg.scala 27:20]
  wire [1:0] _T_21950 = _T_21469 ? bht_bank_rd_data_out_1_31 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22205 = _T_22204 | _T_21950; // @[Mux.scala 27:72]
  wire  _T_21471 = bht_rd_addr_hashed_f == 8'h20; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_32; // @[Reg.scala 27:20]
  wire [1:0] _T_21951 = _T_21471 ? bht_bank_rd_data_out_1_32 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22206 = _T_22205 | _T_21951; // @[Mux.scala 27:72]
  wire  _T_21473 = bht_rd_addr_hashed_f == 8'h21; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_33; // @[Reg.scala 27:20]
  wire [1:0] _T_21952 = _T_21473 ? bht_bank_rd_data_out_1_33 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22207 = _T_22206 | _T_21952; // @[Mux.scala 27:72]
  wire  _T_21475 = bht_rd_addr_hashed_f == 8'h22; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_34; // @[Reg.scala 27:20]
  wire [1:0] _T_21953 = _T_21475 ? bht_bank_rd_data_out_1_34 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22208 = _T_22207 | _T_21953; // @[Mux.scala 27:72]
  wire  _T_21477 = bht_rd_addr_hashed_f == 8'h23; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_35; // @[Reg.scala 27:20]
  wire [1:0] _T_21954 = _T_21477 ? bht_bank_rd_data_out_1_35 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22209 = _T_22208 | _T_21954; // @[Mux.scala 27:72]
  wire  _T_21479 = bht_rd_addr_hashed_f == 8'h24; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_36; // @[Reg.scala 27:20]
  wire [1:0] _T_21955 = _T_21479 ? bht_bank_rd_data_out_1_36 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22210 = _T_22209 | _T_21955; // @[Mux.scala 27:72]
  wire  _T_21481 = bht_rd_addr_hashed_f == 8'h25; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_37; // @[Reg.scala 27:20]
  wire [1:0] _T_21956 = _T_21481 ? bht_bank_rd_data_out_1_37 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22211 = _T_22210 | _T_21956; // @[Mux.scala 27:72]
  wire  _T_21483 = bht_rd_addr_hashed_f == 8'h26; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_38; // @[Reg.scala 27:20]
  wire [1:0] _T_21957 = _T_21483 ? bht_bank_rd_data_out_1_38 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22212 = _T_22211 | _T_21957; // @[Mux.scala 27:72]
  wire  _T_21485 = bht_rd_addr_hashed_f == 8'h27; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_39; // @[Reg.scala 27:20]
  wire [1:0] _T_21958 = _T_21485 ? bht_bank_rd_data_out_1_39 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22213 = _T_22212 | _T_21958; // @[Mux.scala 27:72]
  wire  _T_21487 = bht_rd_addr_hashed_f == 8'h28; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_40; // @[Reg.scala 27:20]
  wire [1:0] _T_21959 = _T_21487 ? bht_bank_rd_data_out_1_40 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22214 = _T_22213 | _T_21959; // @[Mux.scala 27:72]
  wire  _T_21489 = bht_rd_addr_hashed_f == 8'h29; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_41; // @[Reg.scala 27:20]
  wire [1:0] _T_21960 = _T_21489 ? bht_bank_rd_data_out_1_41 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22215 = _T_22214 | _T_21960; // @[Mux.scala 27:72]
  wire  _T_21491 = bht_rd_addr_hashed_f == 8'h2a; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_42; // @[Reg.scala 27:20]
  wire [1:0] _T_21961 = _T_21491 ? bht_bank_rd_data_out_1_42 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22216 = _T_22215 | _T_21961; // @[Mux.scala 27:72]
  wire  _T_21493 = bht_rd_addr_hashed_f == 8'h2b; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_43; // @[Reg.scala 27:20]
  wire [1:0] _T_21962 = _T_21493 ? bht_bank_rd_data_out_1_43 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22217 = _T_22216 | _T_21962; // @[Mux.scala 27:72]
  wire  _T_21495 = bht_rd_addr_hashed_f == 8'h2c; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_44; // @[Reg.scala 27:20]
  wire [1:0] _T_21963 = _T_21495 ? bht_bank_rd_data_out_1_44 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22218 = _T_22217 | _T_21963; // @[Mux.scala 27:72]
  wire  _T_21497 = bht_rd_addr_hashed_f == 8'h2d; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_45; // @[Reg.scala 27:20]
  wire [1:0] _T_21964 = _T_21497 ? bht_bank_rd_data_out_1_45 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22219 = _T_22218 | _T_21964; // @[Mux.scala 27:72]
  wire  _T_21499 = bht_rd_addr_hashed_f == 8'h2e; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_46; // @[Reg.scala 27:20]
  wire [1:0] _T_21965 = _T_21499 ? bht_bank_rd_data_out_1_46 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22220 = _T_22219 | _T_21965; // @[Mux.scala 27:72]
  wire  _T_21501 = bht_rd_addr_hashed_f == 8'h2f; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_47; // @[Reg.scala 27:20]
  wire [1:0] _T_21966 = _T_21501 ? bht_bank_rd_data_out_1_47 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22221 = _T_22220 | _T_21966; // @[Mux.scala 27:72]
  wire  _T_21503 = bht_rd_addr_hashed_f == 8'h30; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_48; // @[Reg.scala 27:20]
  wire [1:0] _T_21967 = _T_21503 ? bht_bank_rd_data_out_1_48 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22222 = _T_22221 | _T_21967; // @[Mux.scala 27:72]
  wire  _T_21505 = bht_rd_addr_hashed_f == 8'h31; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_49; // @[Reg.scala 27:20]
  wire [1:0] _T_21968 = _T_21505 ? bht_bank_rd_data_out_1_49 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22223 = _T_22222 | _T_21968; // @[Mux.scala 27:72]
  wire  _T_21507 = bht_rd_addr_hashed_f == 8'h32; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_50; // @[Reg.scala 27:20]
  wire [1:0] _T_21969 = _T_21507 ? bht_bank_rd_data_out_1_50 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22224 = _T_22223 | _T_21969; // @[Mux.scala 27:72]
  wire  _T_21509 = bht_rd_addr_hashed_f == 8'h33; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_51; // @[Reg.scala 27:20]
  wire [1:0] _T_21970 = _T_21509 ? bht_bank_rd_data_out_1_51 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22225 = _T_22224 | _T_21970; // @[Mux.scala 27:72]
  wire  _T_21511 = bht_rd_addr_hashed_f == 8'h34; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_52; // @[Reg.scala 27:20]
  wire [1:0] _T_21971 = _T_21511 ? bht_bank_rd_data_out_1_52 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22226 = _T_22225 | _T_21971; // @[Mux.scala 27:72]
  wire  _T_21513 = bht_rd_addr_hashed_f == 8'h35; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_53; // @[Reg.scala 27:20]
  wire [1:0] _T_21972 = _T_21513 ? bht_bank_rd_data_out_1_53 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22227 = _T_22226 | _T_21972; // @[Mux.scala 27:72]
  wire  _T_21515 = bht_rd_addr_hashed_f == 8'h36; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_54; // @[Reg.scala 27:20]
  wire [1:0] _T_21973 = _T_21515 ? bht_bank_rd_data_out_1_54 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22228 = _T_22227 | _T_21973; // @[Mux.scala 27:72]
  wire  _T_21517 = bht_rd_addr_hashed_f == 8'h37; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_55; // @[Reg.scala 27:20]
  wire [1:0] _T_21974 = _T_21517 ? bht_bank_rd_data_out_1_55 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22229 = _T_22228 | _T_21974; // @[Mux.scala 27:72]
  wire  _T_21519 = bht_rd_addr_hashed_f == 8'h38; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_56; // @[Reg.scala 27:20]
  wire [1:0] _T_21975 = _T_21519 ? bht_bank_rd_data_out_1_56 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22230 = _T_22229 | _T_21975; // @[Mux.scala 27:72]
  wire  _T_21521 = bht_rd_addr_hashed_f == 8'h39; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_57; // @[Reg.scala 27:20]
  wire [1:0] _T_21976 = _T_21521 ? bht_bank_rd_data_out_1_57 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22231 = _T_22230 | _T_21976; // @[Mux.scala 27:72]
  wire  _T_21523 = bht_rd_addr_hashed_f == 8'h3a; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_58; // @[Reg.scala 27:20]
  wire [1:0] _T_21977 = _T_21523 ? bht_bank_rd_data_out_1_58 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22232 = _T_22231 | _T_21977; // @[Mux.scala 27:72]
  wire  _T_21525 = bht_rd_addr_hashed_f == 8'h3b; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_59; // @[Reg.scala 27:20]
  wire [1:0] _T_21978 = _T_21525 ? bht_bank_rd_data_out_1_59 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22233 = _T_22232 | _T_21978; // @[Mux.scala 27:72]
  wire  _T_21527 = bht_rd_addr_hashed_f == 8'h3c; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_60; // @[Reg.scala 27:20]
  wire [1:0] _T_21979 = _T_21527 ? bht_bank_rd_data_out_1_60 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22234 = _T_22233 | _T_21979; // @[Mux.scala 27:72]
  wire  _T_21529 = bht_rd_addr_hashed_f == 8'h3d; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_61; // @[Reg.scala 27:20]
  wire [1:0] _T_21980 = _T_21529 ? bht_bank_rd_data_out_1_61 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22235 = _T_22234 | _T_21980; // @[Mux.scala 27:72]
  wire  _T_21531 = bht_rd_addr_hashed_f == 8'h3e; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_62; // @[Reg.scala 27:20]
  wire [1:0] _T_21981 = _T_21531 ? bht_bank_rd_data_out_1_62 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22236 = _T_22235 | _T_21981; // @[Mux.scala 27:72]
  wire  _T_21533 = bht_rd_addr_hashed_f == 8'h3f; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_63; // @[Reg.scala 27:20]
  wire [1:0] _T_21982 = _T_21533 ? bht_bank_rd_data_out_1_63 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22237 = _T_22236 | _T_21982; // @[Mux.scala 27:72]
  wire  _T_21535 = bht_rd_addr_hashed_f == 8'h40; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_64; // @[Reg.scala 27:20]
  wire [1:0] _T_21983 = _T_21535 ? bht_bank_rd_data_out_1_64 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22238 = _T_22237 | _T_21983; // @[Mux.scala 27:72]
  wire  _T_21537 = bht_rd_addr_hashed_f == 8'h41; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_65; // @[Reg.scala 27:20]
  wire [1:0] _T_21984 = _T_21537 ? bht_bank_rd_data_out_1_65 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22239 = _T_22238 | _T_21984; // @[Mux.scala 27:72]
  wire  _T_21539 = bht_rd_addr_hashed_f == 8'h42; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_66; // @[Reg.scala 27:20]
  wire [1:0] _T_21985 = _T_21539 ? bht_bank_rd_data_out_1_66 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22240 = _T_22239 | _T_21985; // @[Mux.scala 27:72]
  wire  _T_21541 = bht_rd_addr_hashed_f == 8'h43; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_67; // @[Reg.scala 27:20]
  wire [1:0] _T_21986 = _T_21541 ? bht_bank_rd_data_out_1_67 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22241 = _T_22240 | _T_21986; // @[Mux.scala 27:72]
  wire  _T_21543 = bht_rd_addr_hashed_f == 8'h44; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_68; // @[Reg.scala 27:20]
  wire [1:0] _T_21987 = _T_21543 ? bht_bank_rd_data_out_1_68 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22242 = _T_22241 | _T_21987; // @[Mux.scala 27:72]
  wire  _T_21545 = bht_rd_addr_hashed_f == 8'h45; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_69; // @[Reg.scala 27:20]
  wire [1:0] _T_21988 = _T_21545 ? bht_bank_rd_data_out_1_69 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22243 = _T_22242 | _T_21988; // @[Mux.scala 27:72]
  wire  _T_21547 = bht_rd_addr_hashed_f == 8'h46; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_70; // @[Reg.scala 27:20]
  wire [1:0] _T_21989 = _T_21547 ? bht_bank_rd_data_out_1_70 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22244 = _T_22243 | _T_21989; // @[Mux.scala 27:72]
  wire  _T_21549 = bht_rd_addr_hashed_f == 8'h47; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_71; // @[Reg.scala 27:20]
  wire [1:0] _T_21990 = _T_21549 ? bht_bank_rd_data_out_1_71 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22245 = _T_22244 | _T_21990; // @[Mux.scala 27:72]
  wire  _T_21551 = bht_rd_addr_hashed_f == 8'h48; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_72; // @[Reg.scala 27:20]
  wire [1:0] _T_21991 = _T_21551 ? bht_bank_rd_data_out_1_72 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22246 = _T_22245 | _T_21991; // @[Mux.scala 27:72]
  wire  _T_21553 = bht_rd_addr_hashed_f == 8'h49; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_73; // @[Reg.scala 27:20]
  wire [1:0] _T_21992 = _T_21553 ? bht_bank_rd_data_out_1_73 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22247 = _T_22246 | _T_21992; // @[Mux.scala 27:72]
  wire  _T_21555 = bht_rd_addr_hashed_f == 8'h4a; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_74; // @[Reg.scala 27:20]
  wire [1:0] _T_21993 = _T_21555 ? bht_bank_rd_data_out_1_74 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22248 = _T_22247 | _T_21993; // @[Mux.scala 27:72]
  wire  _T_21557 = bht_rd_addr_hashed_f == 8'h4b; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_75; // @[Reg.scala 27:20]
  wire [1:0] _T_21994 = _T_21557 ? bht_bank_rd_data_out_1_75 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22249 = _T_22248 | _T_21994; // @[Mux.scala 27:72]
  wire  _T_21559 = bht_rd_addr_hashed_f == 8'h4c; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_76; // @[Reg.scala 27:20]
  wire [1:0] _T_21995 = _T_21559 ? bht_bank_rd_data_out_1_76 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22250 = _T_22249 | _T_21995; // @[Mux.scala 27:72]
  wire  _T_21561 = bht_rd_addr_hashed_f == 8'h4d; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_77; // @[Reg.scala 27:20]
  wire [1:0] _T_21996 = _T_21561 ? bht_bank_rd_data_out_1_77 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22251 = _T_22250 | _T_21996; // @[Mux.scala 27:72]
  wire  _T_21563 = bht_rd_addr_hashed_f == 8'h4e; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_78; // @[Reg.scala 27:20]
  wire [1:0] _T_21997 = _T_21563 ? bht_bank_rd_data_out_1_78 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22252 = _T_22251 | _T_21997; // @[Mux.scala 27:72]
  wire  _T_21565 = bht_rd_addr_hashed_f == 8'h4f; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_79; // @[Reg.scala 27:20]
  wire [1:0] _T_21998 = _T_21565 ? bht_bank_rd_data_out_1_79 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22253 = _T_22252 | _T_21998; // @[Mux.scala 27:72]
  wire  _T_21567 = bht_rd_addr_hashed_f == 8'h50; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_80; // @[Reg.scala 27:20]
  wire [1:0] _T_21999 = _T_21567 ? bht_bank_rd_data_out_1_80 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22254 = _T_22253 | _T_21999; // @[Mux.scala 27:72]
  wire  _T_21569 = bht_rd_addr_hashed_f == 8'h51; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_81; // @[Reg.scala 27:20]
  wire [1:0] _T_22000 = _T_21569 ? bht_bank_rd_data_out_1_81 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22255 = _T_22254 | _T_22000; // @[Mux.scala 27:72]
  wire  _T_21571 = bht_rd_addr_hashed_f == 8'h52; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_82; // @[Reg.scala 27:20]
  wire [1:0] _T_22001 = _T_21571 ? bht_bank_rd_data_out_1_82 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22256 = _T_22255 | _T_22001; // @[Mux.scala 27:72]
  wire  _T_21573 = bht_rd_addr_hashed_f == 8'h53; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_83; // @[Reg.scala 27:20]
  wire [1:0] _T_22002 = _T_21573 ? bht_bank_rd_data_out_1_83 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22257 = _T_22256 | _T_22002; // @[Mux.scala 27:72]
  wire  _T_21575 = bht_rd_addr_hashed_f == 8'h54; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_84; // @[Reg.scala 27:20]
  wire [1:0] _T_22003 = _T_21575 ? bht_bank_rd_data_out_1_84 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22258 = _T_22257 | _T_22003; // @[Mux.scala 27:72]
  wire  _T_21577 = bht_rd_addr_hashed_f == 8'h55; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_85; // @[Reg.scala 27:20]
  wire [1:0] _T_22004 = _T_21577 ? bht_bank_rd_data_out_1_85 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22259 = _T_22258 | _T_22004; // @[Mux.scala 27:72]
  wire  _T_21579 = bht_rd_addr_hashed_f == 8'h56; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_86; // @[Reg.scala 27:20]
  wire [1:0] _T_22005 = _T_21579 ? bht_bank_rd_data_out_1_86 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22260 = _T_22259 | _T_22005; // @[Mux.scala 27:72]
  wire  _T_21581 = bht_rd_addr_hashed_f == 8'h57; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_87; // @[Reg.scala 27:20]
  wire [1:0] _T_22006 = _T_21581 ? bht_bank_rd_data_out_1_87 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22261 = _T_22260 | _T_22006; // @[Mux.scala 27:72]
  wire  _T_21583 = bht_rd_addr_hashed_f == 8'h58; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_88; // @[Reg.scala 27:20]
  wire [1:0] _T_22007 = _T_21583 ? bht_bank_rd_data_out_1_88 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22262 = _T_22261 | _T_22007; // @[Mux.scala 27:72]
  wire  _T_21585 = bht_rd_addr_hashed_f == 8'h59; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_89; // @[Reg.scala 27:20]
  wire [1:0] _T_22008 = _T_21585 ? bht_bank_rd_data_out_1_89 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22263 = _T_22262 | _T_22008; // @[Mux.scala 27:72]
  wire  _T_21587 = bht_rd_addr_hashed_f == 8'h5a; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_90; // @[Reg.scala 27:20]
  wire [1:0] _T_22009 = _T_21587 ? bht_bank_rd_data_out_1_90 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22264 = _T_22263 | _T_22009; // @[Mux.scala 27:72]
  wire  _T_21589 = bht_rd_addr_hashed_f == 8'h5b; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_91; // @[Reg.scala 27:20]
  wire [1:0] _T_22010 = _T_21589 ? bht_bank_rd_data_out_1_91 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22265 = _T_22264 | _T_22010; // @[Mux.scala 27:72]
  wire  _T_21591 = bht_rd_addr_hashed_f == 8'h5c; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_92; // @[Reg.scala 27:20]
  wire [1:0] _T_22011 = _T_21591 ? bht_bank_rd_data_out_1_92 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22266 = _T_22265 | _T_22011; // @[Mux.scala 27:72]
  wire  _T_21593 = bht_rd_addr_hashed_f == 8'h5d; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_93; // @[Reg.scala 27:20]
  wire [1:0] _T_22012 = _T_21593 ? bht_bank_rd_data_out_1_93 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22267 = _T_22266 | _T_22012; // @[Mux.scala 27:72]
  wire  _T_21595 = bht_rd_addr_hashed_f == 8'h5e; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_94; // @[Reg.scala 27:20]
  wire [1:0] _T_22013 = _T_21595 ? bht_bank_rd_data_out_1_94 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22268 = _T_22267 | _T_22013; // @[Mux.scala 27:72]
  wire  _T_21597 = bht_rd_addr_hashed_f == 8'h5f; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_95; // @[Reg.scala 27:20]
  wire [1:0] _T_22014 = _T_21597 ? bht_bank_rd_data_out_1_95 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22269 = _T_22268 | _T_22014; // @[Mux.scala 27:72]
  wire  _T_21599 = bht_rd_addr_hashed_f == 8'h60; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_96; // @[Reg.scala 27:20]
  wire [1:0] _T_22015 = _T_21599 ? bht_bank_rd_data_out_1_96 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22270 = _T_22269 | _T_22015; // @[Mux.scala 27:72]
  wire  _T_21601 = bht_rd_addr_hashed_f == 8'h61; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_97; // @[Reg.scala 27:20]
  wire [1:0] _T_22016 = _T_21601 ? bht_bank_rd_data_out_1_97 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22271 = _T_22270 | _T_22016; // @[Mux.scala 27:72]
  wire  _T_21603 = bht_rd_addr_hashed_f == 8'h62; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_98; // @[Reg.scala 27:20]
  wire [1:0] _T_22017 = _T_21603 ? bht_bank_rd_data_out_1_98 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22272 = _T_22271 | _T_22017; // @[Mux.scala 27:72]
  wire  _T_21605 = bht_rd_addr_hashed_f == 8'h63; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_99; // @[Reg.scala 27:20]
  wire [1:0] _T_22018 = _T_21605 ? bht_bank_rd_data_out_1_99 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22273 = _T_22272 | _T_22018; // @[Mux.scala 27:72]
  wire  _T_21607 = bht_rd_addr_hashed_f == 8'h64; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_100; // @[Reg.scala 27:20]
  wire [1:0] _T_22019 = _T_21607 ? bht_bank_rd_data_out_1_100 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22274 = _T_22273 | _T_22019; // @[Mux.scala 27:72]
  wire  _T_21609 = bht_rd_addr_hashed_f == 8'h65; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_101; // @[Reg.scala 27:20]
  wire [1:0] _T_22020 = _T_21609 ? bht_bank_rd_data_out_1_101 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22275 = _T_22274 | _T_22020; // @[Mux.scala 27:72]
  wire  _T_21611 = bht_rd_addr_hashed_f == 8'h66; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_102; // @[Reg.scala 27:20]
  wire [1:0] _T_22021 = _T_21611 ? bht_bank_rd_data_out_1_102 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22276 = _T_22275 | _T_22021; // @[Mux.scala 27:72]
  wire  _T_21613 = bht_rd_addr_hashed_f == 8'h67; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_103; // @[Reg.scala 27:20]
  wire [1:0] _T_22022 = _T_21613 ? bht_bank_rd_data_out_1_103 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22277 = _T_22276 | _T_22022; // @[Mux.scala 27:72]
  wire  _T_21615 = bht_rd_addr_hashed_f == 8'h68; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_104; // @[Reg.scala 27:20]
  wire [1:0] _T_22023 = _T_21615 ? bht_bank_rd_data_out_1_104 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22278 = _T_22277 | _T_22023; // @[Mux.scala 27:72]
  wire  _T_21617 = bht_rd_addr_hashed_f == 8'h69; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_105; // @[Reg.scala 27:20]
  wire [1:0] _T_22024 = _T_21617 ? bht_bank_rd_data_out_1_105 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22279 = _T_22278 | _T_22024; // @[Mux.scala 27:72]
  wire  _T_21619 = bht_rd_addr_hashed_f == 8'h6a; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_106; // @[Reg.scala 27:20]
  wire [1:0] _T_22025 = _T_21619 ? bht_bank_rd_data_out_1_106 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22280 = _T_22279 | _T_22025; // @[Mux.scala 27:72]
  wire  _T_21621 = bht_rd_addr_hashed_f == 8'h6b; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_107; // @[Reg.scala 27:20]
  wire [1:0] _T_22026 = _T_21621 ? bht_bank_rd_data_out_1_107 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22281 = _T_22280 | _T_22026; // @[Mux.scala 27:72]
  wire  _T_21623 = bht_rd_addr_hashed_f == 8'h6c; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_108; // @[Reg.scala 27:20]
  wire [1:0] _T_22027 = _T_21623 ? bht_bank_rd_data_out_1_108 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22282 = _T_22281 | _T_22027; // @[Mux.scala 27:72]
  wire  _T_21625 = bht_rd_addr_hashed_f == 8'h6d; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_109; // @[Reg.scala 27:20]
  wire [1:0] _T_22028 = _T_21625 ? bht_bank_rd_data_out_1_109 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22283 = _T_22282 | _T_22028; // @[Mux.scala 27:72]
  wire  _T_21627 = bht_rd_addr_hashed_f == 8'h6e; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_110; // @[Reg.scala 27:20]
  wire [1:0] _T_22029 = _T_21627 ? bht_bank_rd_data_out_1_110 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22284 = _T_22283 | _T_22029; // @[Mux.scala 27:72]
  wire  _T_21629 = bht_rd_addr_hashed_f == 8'h6f; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_111; // @[Reg.scala 27:20]
  wire [1:0] _T_22030 = _T_21629 ? bht_bank_rd_data_out_1_111 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22285 = _T_22284 | _T_22030; // @[Mux.scala 27:72]
  wire  _T_21631 = bht_rd_addr_hashed_f == 8'h70; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_112; // @[Reg.scala 27:20]
  wire [1:0] _T_22031 = _T_21631 ? bht_bank_rd_data_out_1_112 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22286 = _T_22285 | _T_22031; // @[Mux.scala 27:72]
  wire  _T_21633 = bht_rd_addr_hashed_f == 8'h71; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_113; // @[Reg.scala 27:20]
  wire [1:0] _T_22032 = _T_21633 ? bht_bank_rd_data_out_1_113 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22287 = _T_22286 | _T_22032; // @[Mux.scala 27:72]
  wire  _T_21635 = bht_rd_addr_hashed_f == 8'h72; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_114; // @[Reg.scala 27:20]
  wire [1:0] _T_22033 = _T_21635 ? bht_bank_rd_data_out_1_114 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22288 = _T_22287 | _T_22033; // @[Mux.scala 27:72]
  wire  _T_21637 = bht_rd_addr_hashed_f == 8'h73; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_115; // @[Reg.scala 27:20]
  wire [1:0] _T_22034 = _T_21637 ? bht_bank_rd_data_out_1_115 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22289 = _T_22288 | _T_22034; // @[Mux.scala 27:72]
  wire  _T_21639 = bht_rd_addr_hashed_f == 8'h74; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_116; // @[Reg.scala 27:20]
  wire [1:0] _T_22035 = _T_21639 ? bht_bank_rd_data_out_1_116 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22290 = _T_22289 | _T_22035; // @[Mux.scala 27:72]
  wire  _T_21641 = bht_rd_addr_hashed_f == 8'h75; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_117; // @[Reg.scala 27:20]
  wire [1:0] _T_22036 = _T_21641 ? bht_bank_rd_data_out_1_117 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22291 = _T_22290 | _T_22036; // @[Mux.scala 27:72]
  wire  _T_21643 = bht_rd_addr_hashed_f == 8'h76; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_118; // @[Reg.scala 27:20]
  wire [1:0] _T_22037 = _T_21643 ? bht_bank_rd_data_out_1_118 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22292 = _T_22291 | _T_22037; // @[Mux.scala 27:72]
  wire  _T_21645 = bht_rd_addr_hashed_f == 8'h77; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_119; // @[Reg.scala 27:20]
  wire [1:0] _T_22038 = _T_21645 ? bht_bank_rd_data_out_1_119 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22293 = _T_22292 | _T_22038; // @[Mux.scala 27:72]
  wire  _T_21647 = bht_rd_addr_hashed_f == 8'h78; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_120; // @[Reg.scala 27:20]
  wire [1:0] _T_22039 = _T_21647 ? bht_bank_rd_data_out_1_120 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22294 = _T_22293 | _T_22039; // @[Mux.scala 27:72]
  wire  _T_21649 = bht_rd_addr_hashed_f == 8'h79; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_121; // @[Reg.scala 27:20]
  wire [1:0] _T_22040 = _T_21649 ? bht_bank_rd_data_out_1_121 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22295 = _T_22294 | _T_22040; // @[Mux.scala 27:72]
  wire  _T_21651 = bht_rd_addr_hashed_f == 8'h7a; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_122; // @[Reg.scala 27:20]
  wire [1:0] _T_22041 = _T_21651 ? bht_bank_rd_data_out_1_122 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22296 = _T_22295 | _T_22041; // @[Mux.scala 27:72]
  wire  _T_21653 = bht_rd_addr_hashed_f == 8'h7b; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_123; // @[Reg.scala 27:20]
  wire [1:0] _T_22042 = _T_21653 ? bht_bank_rd_data_out_1_123 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22297 = _T_22296 | _T_22042; // @[Mux.scala 27:72]
  wire  _T_21655 = bht_rd_addr_hashed_f == 8'h7c; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_124; // @[Reg.scala 27:20]
  wire [1:0] _T_22043 = _T_21655 ? bht_bank_rd_data_out_1_124 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22298 = _T_22297 | _T_22043; // @[Mux.scala 27:72]
  wire  _T_21657 = bht_rd_addr_hashed_f == 8'h7d; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_125; // @[Reg.scala 27:20]
  wire [1:0] _T_22044 = _T_21657 ? bht_bank_rd_data_out_1_125 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22299 = _T_22298 | _T_22044; // @[Mux.scala 27:72]
  wire  _T_21659 = bht_rd_addr_hashed_f == 8'h7e; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_126; // @[Reg.scala 27:20]
  wire [1:0] _T_22045 = _T_21659 ? bht_bank_rd_data_out_1_126 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22300 = _T_22299 | _T_22045; // @[Mux.scala 27:72]
  wire  _T_21661 = bht_rd_addr_hashed_f == 8'h7f; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_127; // @[Reg.scala 27:20]
  wire [1:0] _T_22046 = _T_21661 ? bht_bank_rd_data_out_1_127 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22301 = _T_22300 | _T_22046; // @[Mux.scala 27:72]
  wire  _T_21663 = bht_rd_addr_hashed_f == 8'h80; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_128; // @[Reg.scala 27:20]
  wire [1:0] _T_22047 = _T_21663 ? bht_bank_rd_data_out_1_128 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22302 = _T_22301 | _T_22047; // @[Mux.scala 27:72]
  wire  _T_21665 = bht_rd_addr_hashed_f == 8'h81; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_129; // @[Reg.scala 27:20]
  wire [1:0] _T_22048 = _T_21665 ? bht_bank_rd_data_out_1_129 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22303 = _T_22302 | _T_22048; // @[Mux.scala 27:72]
  wire  _T_21667 = bht_rd_addr_hashed_f == 8'h82; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_130; // @[Reg.scala 27:20]
  wire [1:0] _T_22049 = _T_21667 ? bht_bank_rd_data_out_1_130 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22304 = _T_22303 | _T_22049; // @[Mux.scala 27:72]
  wire  _T_21669 = bht_rd_addr_hashed_f == 8'h83; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_131; // @[Reg.scala 27:20]
  wire [1:0] _T_22050 = _T_21669 ? bht_bank_rd_data_out_1_131 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22305 = _T_22304 | _T_22050; // @[Mux.scala 27:72]
  wire  _T_21671 = bht_rd_addr_hashed_f == 8'h84; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_132; // @[Reg.scala 27:20]
  wire [1:0] _T_22051 = _T_21671 ? bht_bank_rd_data_out_1_132 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22306 = _T_22305 | _T_22051; // @[Mux.scala 27:72]
  wire  _T_21673 = bht_rd_addr_hashed_f == 8'h85; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_133; // @[Reg.scala 27:20]
  wire [1:0] _T_22052 = _T_21673 ? bht_bank_rd_data_out_1_133 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22307 = _T_22306 | _T_22052; // @[Mux.scala 27:72]
  wire  _T_21675 = bht_rd_addr_hashed_f == 8'h86; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_134; // @[Reg.scala 27:20]
  wire [1:0] _T_22053 = _T_21675 ? bht_bank_rd_data_out_1_134 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22308 = _T_22307 | _T_22053; // @[Mux.scala 27:72]
  wire  _T_21677 = bht_rd_addr_hashed_f == 8'h87; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_135; // @[Reg.scala 27:20]
  wire [1:0] _T_22054 = _T_21677 ? bht_bank_rd_data_out_1_135 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22309 = _T_22308 | _T_22054; // @[Mux.scala 27:72]
  wire  _T_21679 = bht_rd_addr_hashed_f == 8'h88; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_136; // @[Reg.scala 27:20]
  wire [1:0] _T_22055 = _T_21679 ? bht_bank_rd_data_out_1_136 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22310 = _T_22309 | _T_22055; // @[Mux.scala 27:72]
  wire  _T_21681 = bht_rd_addr_hashed_f == 8'h89; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_137; // @[Reg.scala 27:20]
  wire [1:0] _T_22056 = _T_21681 ? bht_bank_rd_data_out_1_137 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22311 = _T_22310 | _T_22056; // @[Mux.scala 27:72]
  wire  _T_21683 = bht_rd_addr_hashed_f == 8'h8a; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_138; // @[Reg.scala 27:20]
  wire [1:0] _T_22057 = _T_21683 ? bht_bank_rd_data_out_1_138 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22312 = _T_22311 | _T_22057; // @[Mux.scala 27:72]
  wire  _T_21685 = bht_rd_addr_hashed_f == 8'h8b; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_139; // @[Reg.scala 27:20]
  wire [1:0] _T_22058 = _T_21685 ? bht_bank_rd_data_out_1_139 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22313 = _T_22312 | _T_22058; // @[Mux.scala 27:72]
  wire  _T_21687 = bht_rd_addr_hashed_f == 8'h8c; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_140; // @[Reg.scala 27:20]
  wire [1:0] _T_22059 = _T_21687 ? bht_bank_rd_data_out_1_140 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22314 = _T_22313 | _T_22059; // @[Mux.scala 27:72]
  wire  _T_21689 = bht_rd_addr_hashed_f == 8'h8d; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_141; // @[Reg.scala 27:20]
  wire [1:0] _T_22060 = _T_21689 ? bht_bank_rd_data_out_1_141 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22315 = _T_22314 | _T_22060; // @[Mux.scala 27:72]
  wire  _T_21691 = bht_rd_addr_hashed_f == 8'h8e; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_142; // @[Reg.scala 27:20]
  wire [1:0] _T_22061 = _T_21691 ? bht_bank_rd_data_out_1_142 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22316 = _T_22315 | _T_22061; // @[Mux.scala 27:72]
  wire  _T_21693 = bht_rd_addr_hashed_f == 8'h8f; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_143; // @[Reg.scala 27:20]
  wire [1:0] _T_22062 = _T_21693 ? bht_bank_rd_data_out_1_143 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22317 = _T_22316 | _T_22062; // @[Mux.scala 27:72]
  wire  _T_21695 = bht_rd_addr_hashed_f == 8'h90; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_144; // @[Reg.scala 27:20]
  wire [1:0] _T_22063 = _T_21695 ? bht_bank_rd_data_out_1_144 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22318 = _T_22317 | _T_22063; // @[Mux.scala 27:72]
  wire  _T_21697 = bht_rd_addr_hashed_f == 8'h91; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_145; // @[Reg.scala 27:20]
  wire [1:0] _T_22064 = _T_21697 ? bht_bank_rd_data_out_1_145 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22319 = _T_22318 | _T_22064; // @[Mux.scala 27:72]
  wire  _T_21699 = bht_rd_addr_hashed_f == 8'h92; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_146; // @[Reg.scala 27:20]
  wire [1:0] _T_22065 = _T_21699 ? bht_bank_rd_data_out_1_146 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22320 = _T_22319 | _T_22065; // @[Mux.scala 27:72]
  wire  _T_21701 = bht_rd_addr_hashed_f == 8'h93; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_147; // @[Reg.scala 27:20]
  wire [1:0] _T_22066 = _T_21701 ? bht_bank_rd_data_out_1_147 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22321 = _T_22320 | _T_22066; // @[Mux.scala 27:72]
  wire  _T_21703 = bht_rd_addr_hashed_f == 8'h94; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_148; // @[Reg.scala 27:20]
  wire [1:0] _T_22067 = _T_21703 ? bht_bank_rd_data_out_1_148 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22322 = _T_22321 | _T_22067; // @[Mux.scala 27:72]
  wire  _T_21705 = bht_rd_addr_hashed_f == 8'h95; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_149; // @[Reg.scala 27:20]
  wire [1:0] _T_22068 = _T_21705 ? bht_bank_rd_data_out_1_149 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22323 = _T_22322 | _T_22068; // @[Mux.scala 27:72]
  wire  _T_21707 = bht_rd_addr_hashed_f == 8'h96; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_150; // @[Reg.scala 27:20]
  wire [1:0] _T_22069 = _T_21707 ? bht_bank_rd_data_out_1_150 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22324 = _T_22323 | _T_22069; // @[Mux.scala 27:72]
  wire  _T_21709 = bht_rd_addr_hashed_f == 8'h97; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_151; // @[Reg.scala 27:20]
  wire [1:0] _T_22070 = _T_21709 ? bht_bank_rd_data_out_1_151 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22325 = _T_22324 | _T_22070; // @[Mux.scala 27:72]
  wire  _T_21711 = bht_rd_addr_hashed_f == 8'h98; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_152; // @[Reg.scala 27:20]
  wire [1:0] _T_22071 = _T_21711 ? bht_bank_rd_data_out_1_152 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22326 = _T_22325 | _T_22071; // @[Mux.scala 27:72]
  wire  _T_21713 = bht_rd_addr_hashed_f == 8'h99; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_153; // @[Reg.scala 27:20]
  wire [1:0] _T_22072 = _T_21713 ? bht_bank_rd_data_out_1_153 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22327 = _T_22326 | _T_22072; // @[Mux.scala 27:72]
  wire  _T_21715 = bht_rd_addr_hashed_f == 8'h9a; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_154; // @[Reg.scala 27:20]
  wire [1:0] _T_22073 = _T_21715 ? bht_bank_rd_data_out_1_154 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22328 = _T_22327 | _T_22073; // @[Mux.scala 27:72]
  wire  _T_21717 = bht_rd_addr_hashed_f == 8'h9b; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_155; // @[Reg.scala 27:20]
  wire [1:0] _T_22074 = _T_21717 ? bht_bank_rd_data_out_1_155 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22329 = _T_22328 | _T_22074; // @[Mux.scala 27:72]
  wire  _T_21719 = bht_rd_addr_hashed_f == 8'h9c; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_156; // @[Reg.scala 27:20]
  wire [1:0] _T_22075 = _T_21719 ? bht_bank_rd_data_out_1_156 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22330 = _T_22329 | _T_22075; // @[Mux.scala 27:72]
  wire  _T_21721 = bht_rd_addr_hashed_f == 8'h9d; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_157; // @[Reg.scala 27:20]
  wire [1:0] _T_22076 = _T_21721 ? bht_bank_rd_data_out_1_157 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22331 = _T_22330 | _T_22076; // @[Mux.scala 27:72]
  wire  _T_21723 = bht_rd_addr_hashed_f == 8'h9e; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_158; // @[Reg.scala 27:20]
  wire [1:0] _T_22077 = _T_21723 ? bht_bank_rd_data_out_1_158 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22332 = _T_22331 | _T_22077; // @[Mux.scala 27:72]
  wire  _T_21725 = bht_rd_addr_hashed_f == 8'h9f; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_159; // @[Reg.scala 27:20]
  wire [1:0] _T_22078 = _T_21725 ? bht_bank_rd_data_out_1_159 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22333 = _T_22332 | _T_22078; // @[Mux.scala 27:72]
  wire  _T_21727 = bht_rd_addr_hashed_f == 8'ha0; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_160; // @[Reg.scala 27:20]
  wire [1:0] _T_22079 = _T_21727 ? bht_bank_rd_data_out_1_160 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22334 = _T_22333 | _T_22079; // @[Mux.scala 27:72]
  wire  _T_21729 = bht_rd_addr_hashed_f == 8'ha1; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_161; // @[Reg.scala 27:20]
  wire [1:0] _T_22080 = _T_21729 ? bht_bank_rd_data_out_1_161 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22335 = _T_22334 | _T_22080; // @[Mux.scala 27:72]
  wire  _T_21731 = bht_rd_addr_hashed_f == 8'ha2; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_162; // @[Reg.scala 27:20]
  wire [1:0] _T_22081 = _T_21731 ? bht_bank_rd_data_out_1_162 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22336 = _T_22335 | _T_22081; // @[Mux.scala 27:72]
  wire  _T_21733 = bht_rd_addr_hashed_f == 8'ha3; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_163; // @[Reg.scala 27:20]
  wire [1:0] _T_22082 = _T_21733 ? bht_bank_rd_data_out_1_163 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22337 = _T_22336 | _T_22082; // @[Mux.scala 27:72]
  wire  _T_21735 = bht_rd_addr_hashed_f == 8'ha4; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_164; // @[Reg.scala 27:20]
  wire [1:0] _T_22083 = _T_21735 ? bht_bank_rd_data_out_1_164 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22338 = _T_22337 | _T_22083; // @[Mux.scala 27:72]
  wire  _T_21737 = bht_rd_addr_hashed_f == 8'ha5; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_165; // @[Reg.scala 27:20]
  wire [1:0] _T_22084 = _T_21737 ? bht_bank_rd_data_out_1_165 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22339 = _T_22338 | _T_22084; // @[Mux.scala 27:72]
  wire  _T_21739 = bht_rd_addr_hashed_f == 8'ha6; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_166; // @[Reg.scala 27:20]
  wire [1:0] _T_22085 = _T_21739 ? bht_bank_rd_data_out_1_166 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22340 = _T_22339 | _T_22085; // @[Mux.scala 27:72]
  wire  _T_21741 = bht_rd_addr_hashed_f == 8'ha7; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_167; // @[Reg.scala 27:20]
  wire [1:0] _T_22086 = _T_21741 ? bht_bank_rd_data_out_1_167 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22341 = _T_22340 | _T_22086; // @[Mux.scala 27:72]
  wire  _T_21743 = bht_rd_addr_hashed_f == 8'ha8; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_168; // @[Reg.scala 27:20]
  wire [1:0] _T_22087 = _T_21743 ? bht_bank_rd_data_out_1_168 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22342 = _T_22341 | _T_22087; // @[Mux.scala 27:72]
  wire  _T_21745 = bht_rd_addr_hashed_f == 8'ha9; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_169; // @[Reg.scala 27:20]
  wire [1:0] _T_22088 = _T_21745 ? bht_bank_rd_data_out_1_169 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22343 = _T_22342 | _T_22088; // @[Mux.scala 27:72]
  wire  _T_21747 = bht_rd_addr_hashed_f == 8'haa; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_170; // @[Reg.scala 27:20]
  wire [1:0] _T_22089 = _T_21747 ? bht_bank_rd_data_out_1_170 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22344 = _T_22343 | _T_22089; // @[Mux.scala 27:72]
  wire  _T_21749 = bht_rd_addr_hashed_f == 8'hab; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_171; // @[Reg.scala 27:20]
  wire [1:0] _T_22090 = _T_21749 ? bht_bank_rd_data_out_1_171 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22345 = _T_22344 | _T_22090; // @[Mux.scala 27:72]
  wire  _T_21751 = bht_rd_addr_hashed_f == 8'hac; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_172; // @[Reg.scala 27:20]
  wire [1:0] _T_22091 = _T_21751 ? bht_bank_rd_data_out_1_172 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22346 = _T_22345 | _T_22091; // @[Mux.scala 27:72]
  wire  _T_21753 = bht_rd_addr_hashed_f == 8'had; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_173; // @[Reg.scala 27:20]
  wire [1:0] _T_22092 = _T_21753 ? bht_bank_rd_data_out_1_173 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22347 = _T_22346 | _T_22092; // @[Mux.scala 27:72]
  wire  _T_21755 = bht_rd_addr_hashed_f == 8'hae; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_174; // @[Reg.scala 27:20]
  wire [1:0] _T_22093 = _T_21755 ? bht_bank_rd_data_out_1_174 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22348 = _T_22347 | _T_22093; // @[Mux.scala 27:72]
  wire  _T_21757 = bht_rd_addr_hashed_f == 8'haf; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_175; // @[Reg.scala 27:20]
  wire [1:0] _T_22094 = _T_21757 ? bht_bank_rd_data_out_1_175 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22349 = _T_22348 | _T_22094; // @[Mux.scala 27:72]
  wire  _T_21759 = bht_rd_addr_hashed_f == 8'hb0; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_176; // @[Reg.scala 27:20]
  wire [1:0] _T_22095 = _T_21759 ? bht_bank_rd_data_out_1_176 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22350 = _T_22349 | _T_22095; // @[Mux.scala 27:72]
  wire  _T_21761 = bht_rd_addr_hashed_f == 8'hb1; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_177; // @[Reg.scala 27:20]
  wire [1:0] _T_22096 = _T_21761 ? bht_bank_rd_data_out_1_177 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22351 = _T_22350 | _T_22096; // @[Mux.scala 27:72]
  wire  _T_21763 = bht_rd_addr_hashed_f == 8'hb2; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_178; // @[Reg.scala 27:20]
  wire [1:0] _T_22097 = _T_21763 ? bht_bank_rd_data_out_1_178 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22352 = _T_22351 | _T_22097; // @[Mux.scala 27:72]
  wire  _T_21765 = bht_rd_addr_hashed_f == 8'hb3; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_179; // @[Reg.scala 27:20]
  wire [1:0] _T_22098 = _T_21765 ? bht_bank_rd_data_out_1_179 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22353 = _T_22352 | _T_22098; // @[Mux.scala 27:72]
  wire  _T_21767 = bht_rd_addr_hashed_f == 8'hb4; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_180; // @[Reg.scala 27:20]
  wire [1:0] _T_22099 = _T_21767 ? bht_bank_rd_data_out_1_180 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22354 = _T_22353 | _T_22099; // @[Mux.scala 27:72]
  wire  _T_21769 = bht_rd_addr_hashed_f == 8'hb5; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_181; // @[Reg.scala 27:20]
  wire [1:0] _T_22100 = _T_21769 ? bht_bank_rd_data_out_1_181 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22355 = _T_22354 | _T_22100; // @[Mux.scala 27:72]
  wire  _T_21771 = bht_rd_addr_hashed_f == 8'hb6; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_182; // @[Reg.scala 27:20]
  wire [1:0] _T_22101 = _T_21771 ? bht_bank_rd_data_out_1_182 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22356 = _T_22355 | _T_22101; // @[Mux.scala 27:72]
  wire  _T_21773 = bht_rd_addr_hashed_f == 8'hb7; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_183; // @[Reg.scala 27:20]
  wire [1:0] _T_22102 = _T_21773 ? bht_bank_rd_data_out_1_183 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22357 = _T_22356 | _T_22102; // @[Mux.scala 27:72]
  wire  _T_21775 = bht_rd_addr_hashed_f == 8'hb8; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_184; // @[Reg.scala 27:20]
  wire [1:0] _T_22103 = _T_21775 ? bht_bank_rd_data_out_1_184 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22358 = _T_22357 | _T_22103; // @[Mux.scala 27:72]
  wire  _T_21777 = bht_rd_addr_hashed_f == 8'hb9; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_185; // @[Reg.scala 27:20]
  wire [1:0] _T_22104 = _T_21777 ? bht_bank_rd_data_out_1_185 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22359 = _T_22358 | _T_22104; // @[Mux.scala 27:72]
  wire  _T_21779 = bht_rd_addr_hashed_f == 8'hba; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_186; // @[Reg.scala 27:20]
  wire [1:0] _T_22105 = _T_21779 ? bht_bank_rd_data_out_1_186 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22360 = _T_22359 | _T_22105; // @[Mux.scala 27:72]
  wire  _T_21781 = bht_rd_addr_hashed_f == 8'hbb; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_187; // @[Reg.scala 27:20]
  wire [1:0] _T_22106 = _T_21781 ? bht_bank_rd_data_out_1_187 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22361 = _T_22360 | _T_22106; // @[Mux.scala 27:72]
  wire  _T_21783 = bht_rd_addr_hashed_f == 8'hbc; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_188; // @[Reg.scala 27:20]
  wire [1:0] _T_22107 = _T_21783 ? bht_bank_rd_data_out_1_188 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22362 = _T_22361 | _T_22107; // @[Mux.scala 27:72]
  wire  _T_21785 = bht_rd_addr_hashed_f == 8'hbd; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_189; // @[Reg.scala 27:20]
  wire [1:0] _T_22108 = _T_21785 ? bht_bank_rd_data_out_1_189 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22363 = _T_22362 | _T_22108; // @[Mux.scala 27:72]
  wire  _T_21787 = bht_rd_addr_hashed_f == 8'hbe; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_190; // @[Reg.scala 27:20]
  wire [1:0] _T_22109 = _T_21787 ? bht_bank_rd_data_out_1_190 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22364 = _T_22363 | _T_22109; // @[Mux.scala 27:72]
  wire  _T_21789 = bht_rd_addr_hashed_f == 8'hbf; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_191; // @[Reg.scala 27:20]
  wire [1:0] _T_22110 = _T_21789 ? bht_bank_rd_data_out_1_191 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22365 = _T_22364 | _T_22110; // @[Mux.scala 27:72]
  wire  _T_21791 = bht_rd_addr_hashed_f == 8'hc0; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_192; // @[Reg.scala 27:20]
  wire [1:0] _T_22111 = _T_21791 ? bht_bank_rd_data_out_1_192 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22366 = _T_22365 | _T_22111; // @[Mux.scala 27:72]
  wire  _T_21793 = bht_rd_addr_hashed_f == 8'hc1; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_193; // @[Reg.scala 27:20]
  wire [1:0] _T_22112 = _T_21793 ? bht_bank_rd_data_out_1_193 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22367 = _T_22366 | _T_22112; // @[Mux.scala 27:72]
  wire  _T_21795 = bht_rd_addr_hashed_f == 8'hc2; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_194; // @[Reg.scala 27:20]
  wire [1:0] _T_22113 = _T_21795 ? bht_bank_rd_data_out_1_194 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22368 = _T_22367 | _T_22113; // @[Mux.scala 27:72]
  wire  _T_21797 = bht_rd_addr_hashed_f == 8'hc3; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_195; // @[Reg.scala 27:20]
  wire [1:0] _T_22114 = _T_21797 ? bht_bank_rd_data_out_1_195 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22369 = _T_22368 | _T_22114; // @[Mux.scala 27:72]
  wire  _T_21799 = bht_rd_addr_hashed_f == 8'hc4; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_196; // @[Reg.scala 27:20]
  wire [1:0] _T_22115 = _T_21799 ? bht_bank_rd_data_out_1_196 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22370 = _T_22369 | _T_22115; // @[Mux.scala 27:72]
  wire  _T_21801 = bht_rd_addr_hashed_f == 8'hc5; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_197; // @[Reg.scala 27:20]
  wire [1:0] _T_22116 = _T_21801 ? bht_bank_rd_data_out_1_197 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22371 = _T_22370 | _T_22116; // @[Mux.scala 27:72]
  wire  _T_21803 = bht_rd_addr_hashed_f == 8'hc6; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_198; // @[Reg.scala 27:20]
  wire [1:0] _T_22117 = _T_21803 ? bht_bank_rd_data_out_1_198 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22372 = _T_22371 | _T_22117; // @[Mux.scala 27:72]
  wire  _T_21805 = bht_rd_addr_hashed_f == 8'hc7; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_199; // @[Reg.scala 27:20]
  wire [1:0] _T_22118 = _T_21805 ? bht_bank_rd_data_out_1_199 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22373 = _T_22372 | _T_22118; // @[Mux.scala 27:72]
  wire  _T_21807 = bht_rd_addr_hashed_f == 8'hc8; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_200; // @[Reg.scala 27:20]
  wire [1:0] _T_22119 = _T_21807 ? bht_bank_rd_data_out_1_200 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22374 = _T_22373 | _T_22119; // @[Mux.scala 27:72]
  wire  _T_21809 = bht_rd_addr_hashed_f == 8'hc9; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_201; // @[Reg.scala 27:20]
  wire [1:0] _T_22120 = _T_21809 ? bht_bank_rd_data_out_1_201 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22375 = _T_22374 | _T_22120; // @[Mux.scala 27:72]
  wire  _T_21811 = bht_rd_addr_hashed_f == 8'hca; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_202; // @[Reg.scala 27:20]
  wire [1:0] _T_22121 = _T_21811 ? bht_bank_rd_data_out_1_202 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22376 = _T_22375 | _T_22121; // @[Mux.scala 27:72]
  wire  _T_21813 = bht_rd_addr_hashed_f == 8'hcb; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_203; // @[Reg.scala 27:20]
  wire [1:0] _T_22122 = _T_21813 ? bht_bank_rd_data_out_1_203 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22377 = _T_22376 | _T_22122; // @[Mux.scala 27:72]
  wire  _T_21815 = bht_rd_addr_hashed_f == 8'hcc; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_204; // @[Reg.scala 27:20]
  wire [1:0] _T_22123 = _T_21815 ? bht_bank_rd_data_out_1_204 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22378 = _T_22377 | _T_22123; // @[Mux.scala 27:72]
  wire  _T_21817 = bht_rd_addr_hashed_f == 8'hcd; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_205; // @[Reg.scala 27:20]
  wire [1:0] _T_22124 = _T_21817 ? bht_bank_rd_data_out_1_205 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22379 = _T_22378 | _T_22124; // @[Mux.scala 27:72]
  wire  _T_21819 = bht_rd_addr_hashed_f == 8'hce; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_206; // @[Reg.scala 27:20]
  wire [1:0] _T_22125 = _T_21819 ? bht_bank_rd_data_out_1_206 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22380 = _T_22379 | _T_22125; // @[Mux.scala 27:72]
  wire  _T_21821 = bht_rd_addr_hashed_f == 8'hcf; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_207; // @[Reg.scala 27:20]
  wire [1:0] _T_22126 = _T_21821 ? bht_bank_rd_data_out_1_207 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22381 = _T_22380 | _T_22126; // @[Mux.scala 27:72]
  wire  _T_21823 = bht_rd_addr_hashed_f == 8'hd0; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_208; // @[Reg.scala 27:20]
  wire [1:0] _T_22127 = _T_21823 ? bht_bank_rd_data_out_1_208 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22382 = _T_22381 | _T_22127; // @[Mux.scala 27:72]
  wire  _T_21825 = bht_rd_addr_hashed_f == 8'hd1; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_209; // @[Reg.scala 27:20]
  wire [1:0] _T_22128 = _T_21825 ? bht_bank_rd_data_out_1_209 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22383 = _T_22382 | _T_22128; // @[Mux.scala 27:72]
  wire  _T_21827 = bht_rd_addr_hashed_f == 8'hd2; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_210; // @[Reg.scala 27:20]
  wire [1:0] _T_22129 = _T_21827 ? bht_bank_rd_data_out_1_210 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22384 = _T_22383 | _T_22129; // @[Mux.scala 27:72]
  wire  _T_21829 = bht_rd_addr_hashed_f == 8'hd3; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_211; // @[Reg.scala 27:20]
  wire [1:0] _T_22130 = _T_21829 ? bht_bank_rd_data_out_1_211 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22385 = _T_22384 | _T_22130; // @[Mux.scala 27:72]
  wire  _T_21831 = bht_rd_addr_hashed_f == 8'hd4; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_212; // @[Reg.scala 27:20]
  wire [1:0] _T_22131 = _T_21831 ? bht_bank_rd_data_out_1_212 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22386 = _T_22385 | _T_22131; // @[Mux.scala 27:72]
  wire  _T_21833 = bht_rd_addr_hashed_f == 8'hd5; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_213; // @[Reg.scala 27:20]
  wire [1:0] _T_22132 = _T_21833 ? bht_bank_rd_data_out_1_213 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22387 = _T_22386 | _T_22132; // @[Mux.scala 27:72]
  wire  _T_21835 = bht_rd_addr_hashed_f == 8'hd6; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_214; // @[Reg.scala 27:20]
  wire [1:0] _T_22133 = _T_21835 ? bht_bank_rd_data_out_1_214 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22388 = _T_22387 | _T_22133; // @[Mux.scala 27:72]
  wire  _T_21837 = bht_rd_addr_hashed_f == 8'hd7; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_215; // @[Reg.scala 27:20]
  wire [1:0] _T_22134 = _T_21837 ? bht_bank_rd_data_out_1_215 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22389 = _T_22388 | _T_22134; // @[Mux.scala 27:72]
  wire  _T_21839 = bht_rd_addr_hashed_f == 8'hd8; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_216; // @[Reg.scala 27:20]
  wire [1:0] _T_22135 = _T_21839 ? bht_bank_rd_data_out_1_216 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22390 = _T_22389 | _T_22135; // @[Mux.scala 27:72]
  wire  _T_21841 = bht_rd_addr_hashed_f == 8'hd9; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_217; // @[Reg.scala 27:20]
  wire [1:0] _T_22136 = _T_21841 ? bht_bank_rd_data_out_1_217 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22391 = _T_22390 | _T_22136; // @[Mux.scala 27:72]
  wire  _T_21843 = bht_rd_addr_hashed_f == 8'hda; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_218; // @[Reg.scala 27:20]
  wire [1:0] _T_22137 = _T_21843 ? bht_bank_rd_data_out_1_218 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22392 = _T_22391 | _T_22137; // @[Mux.scala 27:72]
  wire  _T_21845 = bht_rd_addr_hashed_f == 8'hdb; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_219; // @[Reg.scala 27:20]
  wire [1:0] _T_22138 = _T_21845 ? bht_bank_rd_data_out_1_219 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22393 = _T_22392 | _T_22138; // @[Mux.scala 27:72]
  wire  _T_21847 = bht_rd_addr_hashed_f == 8'hdc; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_220; // @[Reg.scala 27:20]
  wire [1:0] _T_22139 = _T_21847 ? bht_bank_rd_data_out_1_220 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22394 = _T_22393 | _T_22139; // @[Mux.scala 27:72]
  wire  _T_21849 = bht_rd_addr_hashed_f == 8'hdd; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_221; // @[Reg.scala 27:20]
  wire [1:0] _T_22140 = _T_21849 ? bht_bank_rd_data_out_1_221 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22395 = _T_22394 | _T_22140; // @[Mux.scala 27:72]
  wire  _T_21851 = bht_rd_addr_hashed_f == 8'hde; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_222; // @[Reg.scala 27:20]
  wire [1:0] _T_22141 = _T_21851 ? bht_bank_rd_data_out_1_222 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22396 = _T_22395 | _T_22141; // @[Mux.scala 27:72]
  wire  _T_21853 = bht_rd_addr_hashed_f == 8'hdf; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_223; // @[Reg.scala 27:20]
  wire [1:0] _T_22142 = _T_21853 ? bht_bank_rd_data_out_1_223 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22397 = _T_22396 | _T_22142; // @[Mux.scala 27:72]
  wire  _T_21855 = bht_rd_addr_hashed_f == 8'he0; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_224; // @[Reg.scala 27:20]
  wire [1:0] _T_22143 = _T_21855 ? bht_bank_rd_data_out_1_224 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22398 = _T_22397 | _T_22143; // @[Mux.scala 27:72]
  wire  _T_21857 = bht_rd_addr_hashed_f == 8'he1; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_225; // @[Reg.scala 27:20]
  wire [1:0] _T_22144 = _T_21857 ? bht_bank_rd_data_out_1_225 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22399 = _T_22398 | _T_22144; // @[Mux.scala 27:72]
  wire  _T_21859 = bht_rd_addr_hashed_f == 8'he2; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_226; // @[Reg.scala 27:20]
  wire [1:0] _T_22145 = _T_21859 ? bht_bank_rd_data_out_1_226 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22400 = _T_22399 | _T_22145; // @[Mux.scala 27:72]
  wire  _T_21861 = bht_rd_addr_hashed_f == 8'he3; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_227; // @[Reg.scala 27:20]
  wire [1:0] _T_22146 = _T_21861 ? bht_bank_rd_data_out_1_227 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22401 = _T_22400 | _T_22146; // @[Mux.scala 27:72]
  wire  _T_21863 = bht_rd_addr_hashed_f == 8'he4; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_228; // @[Reg.scala 27:20]
  wire [1:0] _T_22147 = _T_21863 ? bht_bank_rd_data_out_1_228 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22402 = _T_22401 | _T_22147; // @[Mux.scala 27:72]
  wire  _T_21865 = bht_rd_addr_hashed_f == 8'he5; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_229; // @[Reg.scala 27:20]
  wire [1:0] _T_22148 = _T_21865 ? bht_bank_rd_data_out_1_229 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22403 = _T_22402 | _T_22148; // @[Mux.scala 27:72]
  wire  _T_21867 = bht_rd_addr_hashed_f == 8'he6; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_230; // @[Reg.scala 27:20]
  wire [1:0] _T_22149 = _T_21867 ? bht_bank_rd_data_out_1_230 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22404 = _T_22403 | _T_22149; // @[Mux.scala 27:72]
  wire  _T_21869 = bht_rd_addr_hashed_f == 8'he7; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_231; // @[Reg.scala 27:20]
  wire [1:0] _T_22150 = _T_21869 ? bht_bank_rd_data_out_1_231 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22405 = _T_22404 | _T_22150; // @[Mux.scala 27:72]
  wire  _T_21871 = bht_rd_addr_hashed_f == 8'he8; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_232; // @[Reg.scala 27:20]
  wire [1:0] _T_22151 = _T_21871 ? bht_bank_rd_data_out_1_232 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22406 = _T_22405 | _T_22151; // @[Mux.scala 27:72]
  wire  _T_21873 = bht_rd_addr_hashed_f == 8'he9; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_233; // @[Reg.scala 27:20]
  wire [1:0] _T_22152 = _T_21873 ? bht_bank_rd_data_out_1_233 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22407 = _T_22406 | _T_22152; // @[Mux.scala 27:72]
  wire  _T_21875 = bht_rd_addr_hashed_f == 8'hea; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_234; // @[Reg.scala 27:20]
  wire [1:0] _T_22153 = _T_21875 ? bht_bank_rd_data_out_1_234 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22408 = _T_22407 | _T_22153; // @[Mux.scala 27:72]
  wire  _T_21877 = bht_rd_addr_hashed_f == 8'heb; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_235; // @[Reg.scala 27:20]
  wire [1:0] _T_22154 = _T_21877 ? bht_bank_rd_data_out_1_235 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22409 = _T_22408 | _T_22154; // @[Mux.scala 27:72]
  wire  _T_21879 = bht_rd_addr_hashed_f == 8'hec; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_236; // @[Reg.scala 27:20]
  wire [1:0] _T_22155 = _T_21879 ? bht_bank_rd_data_out_1_236 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22410 = _T_22409 | _T_22155; // @[Mux.scala 27:72]
  wire  _T_21881 = bht_rd_addr_hashed_f == 8'hed; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_237; // @[Reg.scala 27:20]
  wire [1:0] _T_22156 = _T_21881 ? bht_bank_rd_data_out_1_237 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22411 = _T_22410 | _T_22156; // @[Mux.scala 27:72]
  wire  _T_21883 = bht_rd_addr_hashed_f == 8'hee; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_238; // @[Reg.scala 27:20]
  wire [1:0] _T_22157 = _T_21883 ? bht_bank_rd_data_out_1_238 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22412 = _T_22411 | _T_22157; // @[Mux.scala 27:72]
  wire  _T_21885 = bht_rd_addr_hashed_f == 8'hef; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_239; // @[Reg.scala 27:20]
  wire [1:0] _T_22158 = _T_21885 ? bht_bank_rd_data_out_1_239 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22413 = _T_22412 | _T_22158; // @[Mux.scala 27:72]
  wire  _T_21887 = bht_rd_addr_hashed_f == 8'hf0; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_240; // @[Reg.scala 27:20]
  wire [1:0] _T_22159 = _T_21887 ? bht_bank_rd_data_out_1_240 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22414 = _T_22413 | _T_22159; // @[Mux.scala 27:72]
  wire  _T_21889 = bht_rd_addr_hashed_f == 8'hf1; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_241; // @[Reg.scala 27:20]
  wire [1:0] _T_22160 = _T_21889 ? bht_bank_rd_data_out_1_241 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22415 = _T_22414 | _T_22160; // @[Mux.scala 27:72]
  wire  _T_21891 = bht_rd_addr_hashed_f == 8'hf2; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_242; // @[Reg.scala 27:20]
  wire [1:0] _T_22161 = _T_21891 ? bht_bank_rd_data_out_1_242 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22416 = _T_22415 | _T_22161; // @[Mux.scala 27:72]
  wire  _T_21893 = bht_rd_addr_hashed_f == 8'hf3; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_243; // @[Reg.scala 27:20]
  wire [1:0] _T_22162 = _T_21893 ? bht_bank_rd_data_out_1_243 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22417 = _T_22416 | _T_22162; // @[Mux.scala 27:72]
  wire  _T_21895 = bht_rd_addr_hashed_f == 8'hf4; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_244; // @[Reg.scala 27:20]
  wire [1:0] _T_22163 = _T_21895 ? bht_bank_rd_data_out_1_244 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22418 = _T_22417 | _T_22163; // @[Mux.scala 27:72]
  wire  _T_21897 = bht_rd_addr_hashed_f == 8'hf5; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_245; // @[Reg.scala 27:20]
  wire [1:0] _T_22164 = _T_21897 ? bht_bank_rd_data_out_1_245 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22419 = _T_22418 | _T_22164; // @[Mux.scala 27:72]
  wire  _T_21899 = bht_rd_addr_hashed_f == 8'hf6; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_246; // @[Reg.scala 27:20]
  wire [1:0] _T_22165 = _T_21899 ? bht_bank_rd_data_out_1_246 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22420 = _T_22419 | _T_22165; // @[Mux.scala 27:72]
  wire  _T_21901 = bht_rd_addr_hashed_f == 8'hf7; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_247; // @[Reg.scala 27:20]
  wire [1:0] _T_22166 = _T_21901 ? bht_bank_rd_data_out_1_247 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22421 = _T_22420 | _T_22166; // @[Mux.scala 27:72]
  wire  _T_21903 = bht_rd_addr_hashed_f == 8'hf8; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_248; // @[Reg.scala 27:20]
  wire [1:0] _T_22167 = _T_21903 ? bht_bank_rd_data_out_1_248 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22422 = _T_22421 | _T_22167; // @[Mux.scala 27:72]
  wire  _T_21905 = bht_rd_addr_hashed_f == 8'hf9; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_249; // @[Reg.scala 27:20]
  wire [1:0] _T_22168 = _T_21905 ? bht_bank_rd_data_out_1_249 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22423 = _T_22422 | _T_22168; // @[Mux.scala 27:72]
  wire  _T_21907 = bht_rd_addr_hashed_f == 8'hfa; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_250; // @[Reg.scala 27:20]
  wire [1:0] _T_22169 = _T_21907 ? bht_bank_rd_data_out_1_250 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22424 = _T_22423 | _T_22169; // @[Mux.scala 27:72]
  wire  _T_21909 = bht_rd_addr_hashed_f == 8'hfb; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_251; // @[Reg.scala 27:20]
  wire [1:0] _T_22170 = _T_21909 ? bht_bank_rd_data_out_1_251 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22425 = _T_22424 | _T_22170; // @[Mux.scala 27:72]
  wire  _T_21911 = bht_rd_addr_hashed_f == 8'hfc; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_252; // @[Reg.scala 27:20]
  wire [1:0] _T_22171 = _T_21911 ? bht_bank_rd_data_out_1_252 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22426 = _T_22425 | _T_22171; // @[Mux.scala 27:72]
  wire  _T_21913 = bht_rd_addr_hashed_f == 8'hfd; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_253; // @[Reg.scala 27:20]
  wire [1:0] _T_22172 = _T_21913 ? bht_bank_rd_data_out_1_253 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22427 = _T_22426 | _T_22172; // @[Mux.scala 27:72]
  wire  _T_21915 = bht_rd_addr_hashed_f == 8'hfe; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_254; // @[Reg.scala 27:20]
  wire [1:0] _T_22173 = _T_21915 ? bht_bank_rd_data_out_1_254 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22428 = _T_22427 | _T_22173; // @[Mux.scala 27:72]
  wire  _T_21917 = bht_rd_addr_hashed_f == 8'hff; // @[el2_ifu_bp_ctl.scala 467:79]
  reg [1:0] bht_bank_rd_data_out_1_255; // @[Reg.scala 27:20]
  wire [1:0] _T_22174 = _T_21917 ? bht_bank_rd_data_out_1_255 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] bht_bank1_rd_data_f = _T_22428 | _T_22174; // @[Mux.scala 27:72]
  wire [1:0] _T_259 = _T_143 ? bht_bank1_rd_data_f : 2'h0; // @[Mux.scala 27:72]
  wire [9:0] _T_572 = {btb_rd_addr_p1_f,2'h0}; // @[Cat.scala 29:58]
  wire [7:0] bht_rd_addr_hashed_p1_f = _T_572[9:2] ^ fghr; // @[el2_lib.scala 194:35]
  wire  _T_22431 = bht_rd_addr_hashed_p1_f == 8'h0; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_0; // @[Reg.scala 27:20]
  wire [1:0] _T_22943 = _T_22431 ? bht_bank_rd_data_out_0_0 : 2'h0; // @[Mux.scala 27:72]
  wire  _T_22433 = bht_rd_addr_hashed_p1_f == 8'h1; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_1; // @[Reg.scala 27:20]
  wire [1:0] _T_22944 = _T_22433 ? bht_bank_rd_data_out_0_1 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23199 = _T_22943 | _T_22944; // @[Mux.scala 27:72]
  wire  _T_22435 = bht_rd_addr_hashed_p1_f == 8'h2; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_2; // @[Reg.scala 27:20]
  wire [1:0] _T_22945 = _T_22435 ? bht_bank_rd_data_out_0_2 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23200 = _T_23199 | _T_22945; // @[Mux.scala 27:72]
  wire  _T_22437 = bht_rd_addr_hashed_p1_f == 8'h3; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_3; // @[Reg.scala 27:20]
  wire [1:0] _T_22946 = _T_22437 ? bht_bank_rd_data_out_0_3 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23201 = _T_23200 | _T_22946; // @[Mux.scala 27:72]
  wire  _T_22439 = bht_rd_addr_hashed_p1_f == 8'h4; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_4; // @[Reg.scala 27:20]
  wire [1:0] _T_22947 = _T_22439 ? bht_bank_rd_data_out_0_4 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23202 = _T_23201 | _T_22947; // @[Mux.scala 27:72]
  wire  _T_22441 = bht_rd_addr_hashed_p1_f == 8'h5; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_5; // @[Reg.scala 27:20]
  wire [1:0] _T_22948 = _T_22441 ? bht_bank_rd_data_out_0_5 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23203 = _T_23202 | _T_22948; // @[Mux.scala 27:72]
  wire  _T_22443 = bht_rd_addr_hashed_p1_f == 8'h6; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_6; // @[Reg.scala 27:20]
  wire [1:0] _T_22949 = _T_22443 ? bht_bank_rd_data_out_0_6 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23204 = _T_23203 | _T_22949; // @[Mux.scala 27:72]
  wire  _T_22445 = bht_rd_addr_hashed_p1_f == 8'h7; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_7; // @[Reg.scala 27:20]
  wire [1:0] _T_22950 = _T_22445 ? bht_bank_rd_data_out_0_7 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23205 = _T_23204 | _T_22950; // @[Mux.scala 27:72]
  wire  _T_22447 = bht_rd_addr_hashed_p1_f == 8'h8; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_8; // @[Reg.scala 27:20]
  wire [1:0] _T_22951 = _T_22447 ? bht_bank_rd_data_out_0_8 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23206 = _T_23205 | _T_22951; // @[Mux.scala 27:72]
  wire  _T_22449 = bht_rd_addr_hashed_p1_f == 8'h9; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_9; // @[Reg.scala 27:20]
  wire [1:0] _T_22952 = _T_22449 ? bht_bank_rd_data_out_0_9 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23207 = _T_23206 | _T_22952; // @[Mux.scala 27:72]
  wire  _T_22451 = bht_rd_addr_hashed_p1_f == 8'ha; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_10; // @[Reg.scala 27:20]
  wire [1:0] _T_22953 = _T_22451 ? bht_bank_rd_data_out_0_10 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23208 = _T_23207 | _T_22953; // @[Mux.scala 27:72]
  wire  _T_22453 = bht_rd_addr_hashed_p1_f == 8'hb; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_11; // @[Reg.scala 27:20]
  wire [1:0] _T_22954 = _T_22453 ? bht_bank_rd_data_out_0_11 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23209 = _T_23208 | _T_22954; // @[Mux.scala 27:72]
  wire  _T_22455 = bht_rd_addr_hashed_p1_f == 8'hc; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_12; // @[Reg.scala 27:20]
  wire [1:0] _T_22955 = _T_22455 ? bht_bank_rd_data_out_0_12 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23210 = _T_23209 | _T_22955; // @[Mux.scala 27:72]
  wire  _T_22457 = bht_rd_addr_hashed_p1_f == 8'hd; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_13; // @[Reg.scala 27:20]
  wire [1:0] _T_22956 = _T_22457 ? bht_bank_rd_data_out_0_13 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23211 = _T_23210 | _T_22956; // @[Mux.scala 27:72]
  wire  _T_22459 = bht_rd_addr_hashed_p1_f == 8'he; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_14; // @[Reg.scala 27:20]
  wire [1:0] _T_22957 = _T_22459 ? bht_bank_rd_data_out_0_14 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23212 = _T_23211 | _T_22957; // @[Mux.scala 27:72]
  wire  _T_22461 = bht_rd_addr_hashed_p1_f == 8'hf; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_15; // @[Reg.scala 27:20]
  wire [1:0] _T_22958 = _T_22461 ? bht_bank_rd_data_out_0_15 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23213 = _T_23212 | _T_22958; // @[Mux.scala 27:72]
  wire  _T_22463 = bht_rd_addr_hashed_p1_f == 8'h10; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_16; // @[Reg.scala 27:20]
  wire [1:0] _T_22959 = _T_22463 ? bht_bank_rd_data_out_0_16 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23214 = _T_23213 | _T_22959; // @[Mux.scala 27:72]
  wire  _T_22465 = bht_rd_addr_hashed_p1_f == 8'h11; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_17; // @[Reg.scala 27:20]
  wire [1:0] _T_22960 = _T_22465 ? bht_bank_rd_data_out_0_17 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23215 = _T_23214 | _T_22960; // @[Mux.scala 27:72]
  wire  _T_22467 = bht_rd_addr_hashed_p1_f == 8'h12; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_18; // @[Reg.scala 27:20]
  wire [1:0] _T_22961 = _T_22467 ? bht_bank_rd_data_out_0_18 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23216 = _T_23215 | _T_22961; // @[Mux.scala 27:72]
  wire  _T_22469 = bht_rd_addr_hashed_p1_f == 8'h13; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_19; // @[Reg.scala 27:20]
  wire [1:0] _T_22962 = _T_22469 ? bht_bank_rd_data_out_0_19 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23217 = _T_23216 | _T_22962; // @[Mux.scala 27:72]
  wire  _T_22471 = bht_rd_addr_hashed_p1_f == 8'h14; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_20; // @[Reg.scala 27:20]
  wire [1:0] _T_22963 = _T_22471 ? bht_bank_rd_data_out_0_20 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23218 = _T_23217 | _T_22963; // @[Mux.scala 27:72]
  wire  _T_22473 = bht_rd_addr_hashed_p1_f == 8'h15; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_21; // @[Reg.scala 27:20]
  wire [1:0] _T_22964 = _T_22473 ? bht_bank_rd_data_out_0_21 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23219 = _T_23218 | _T_22964; // @[Mux.scala 27:72]
  wire  _T_22475 = bht_rd_addr_hashed_p1_f == 8'h16; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_22; // @[Reg.scala 27:20]
  wire [1:0] _T_22965 = _T_22475 ? bht_bank_rd_data_out_0_22 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23220 = _T_23219 | _T_22965; // @[Mux.scala 27:72]
  wire  _T_22477 = bht_rd_addr_hashed_p1_f == 8'h17; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_23; // @[Reg.scala 27:20]
  wire [1:0] _T_22966 = _T_22477 ? bht_bank_rd_data_out_0_23 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23221 = _T_23220 | _T_22966; // @[Mux.scala 27:72]
  wire  _T_22479 = bht_rd_addr_hashed_p1_f == 8'h18; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_24; // @[Reg.scala 27:20]
  wire [1:0] _T_22967 = _T_22479 ? bht_bank_rd_data_out_0_24 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23222 = _T_23221 | _T_22967; // @[Mux.scala 27:72]
  wire  _T_22481 = bht_rd_addr_hashed_p1_f == 8'h19; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_25; // @[Reg.scala 27:20]
  wire [1:0] _T_22968 = _T_22481 ? bht_bank_rd_data_out_0_25 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23223 = _T_23222 | _T_22968; // @[Mux.scala 27:72]
  wire  _T_22483 = bht_rd_addr_hashed_p1_f == 8'h1a; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_26; // @[Reg.scala 27:20]
  wire [1:0] _T_22969 = _T_22483 ? bht_bank_rd_data_out_0_26 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23224 = _T_23223 | _T_22969; // @[Mux.scala 27:72]
  wire  _T_22485 = bht_rd_addr_hashed_p1_f == 8'h1b; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_27; // @[Reg.scala 27:20]
  wire [1:0] _T_22970 = _T_22485 ? bht_bank_rd_data_out_0_27 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23225 = _T_23224 | _T_22970; // @[Mux.scala 27:72]
  wire  _T_22487 = bht_rd_addr_hashed_p1_f == 8'h1c; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_28; // @[Reg.scala 27:20]
  wire [1:0] _T_22971 = _T_22487 ? bht_bank_rd_data_out_0_28 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23226 = _T_23225 | _T_22971; // @[Mux.scala 27:72]
  wire  _T_22489 = bht_rd_addr_hashed_p1_f == 8'h1d; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_29; // @[Reg.scala 27:20]
  wire [1:0] _T_22972 = _T_22489 ? bht_bank_rd_data_out_0_29 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23227 = _T_23226 | _T_22972; // @[Mux.scala 27:72]
  wire  _T_22491 = bht_rd_addr_hashed_p1_f == 8'h1e; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_30; // @[Reg.scala 27:20]
  wire [1:0] _T_22973 = _T_22491 ? bht_bank_rd_data_out_0_30 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23228 = _T_23227 | _T_22973; // @[Mux.scala 27:72]
  wire  _T_22493 = bht_rd_addr_hashed_p1_f == 8'h1f; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_31; // @[Reg.scala 27:20]
  wire [1:0] _T_22974 = _T_22493 ? bht_bank_rd_data_out_0_31 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23229 = _T_23228 | _T_22974; // @[Mux.scala 27:72]
  wire  _T_22495 = bht_rd_addr_hashed_p1_f == 8'h20; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_32; // @[Reg.scala 27:20]
  wire [1:0] _T_22975 = _T_22495 ? bht_bank_rd_data_out_0_32 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23230 = _T_23229 | _T_22975; // @[Mux.scala 27:72]
  wire  _T_22497 = bht_rd_addr_hashed_p1_f == 8'h21; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_33; // @[Reg.scala 27:20]
  wire [1:0] _T_22976 = _T_22497 ? bht_bank_rd_data_out_0_33 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23231 = _T_23230 | _T_22976; // @[Mux.scala 27:72]
  wire  _T_22499 = bht_rd_addr_hashed_p1_f == 8'h22; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_34; // @[Reg.scala 27:20]
  wire [1:0] _T_22977 = _T_22499 ? bht_bank_rd_data_out_0_34 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23232 = _T_23231 | _T_22977; // @[Mux.scala 27:72]
  wire  _T_22501 = bht_rd_addr_hashed_p1_f == 8'h23; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_35; // @[Reg.scala 27:20]
  wire [1:0] _T_22978 = _T_22501 ? bht_bank_rd_data_out_0_35 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23233 = _T_23232 | _T_22978; // @[Mux.scala 27:72]
  wire  _T_22503 = bht_rd_addr_hashed_p1_f == 8'h24; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_36; // @[Reg.scala 27:20]
  wire [1:0] _T_22979 = _T_22503 ? bht_bank_rd_data_out_0_36 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23234 = _T_23233 | _T_22979; // @[Mux.scala 27:72]
  wire  _T_22505 = bht_rd_addr_hashed_p1_f == 8'h25; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_37; // @[Reg.scala 27:20]
  wire [1:0] _T_22980 = _T_22505 ? bht_bank_rd_data_out_0_37 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23235 = _T_23234 | _T_22980; // @[Mux.scala 27:72]
  wire  _T_22507 = bht_rd_addr_hashed_p1_f == 8'h26; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_38; // @[Reg.scala 27:20]
  wire [1:0] _T_22981 = _T_22507 ? bht_bank_rd_data_out_0_38 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23236 = _T_23235 | _T_22981; // @[Mux.scala 27:72]
  wire  _T_22509 = bht_rd_addr_hashed_p1_f == 8'h27; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_39; // @[Reg.scala 27:20]
  wire [1:0] _T_22982 = _T_22509 ? bht_bank_rd_data_out_0_39 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23237 = _T_23236 | _T_22982; // @[Mux.scala 27:72]
  wire  _T_22511 = bht_rd_addr_hashed_p1_f == 8'h28; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_40; // @[Reg.scala 27:20]
  wire [1:0] _T_22983 = _T_22511 ? bht_bank_rd_data_out_0_40 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23238 = _T_23237 | _T_22983; // @[Mux.scala 27:72]
  wire  _T_22513 = bht_rd_addr_hashed_p1_f == 8'h29; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_41; // @[Reg.scala 27:20]
  wire [1:0] _T_22984 = _T_22513 ? bht_bank_rd_data_out_0_41 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23239 = _T_23238 | _T_22984; // @[Mux.scala 27:72]
  wire  _T_22515 = bht_rd_addr_hashed_p1_f == 8'h2a; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_42; // @[Reg.scala 27:20]
  wire [1:0] _T_22985 = _T_22515 ? bht_bank_rd_data_out_0_42 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23240 = _T_23239 | _T_22985; // @[Mux.scala 27:72]
  wire  _T_22517 = bht_rd_addr_hashed_p1_f == 8'h2b; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_43; // @[Reg.scala 27:20]
  wire [1:0] _T_22986 = _T_22517 ? bht_bank_rd_data_out_0_43 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23241 = _T_23240 | _T_22986; // @[Mux.scala 27:72]
  wire  _T_22519 = bht_rd_addr_hashed_p1_f == 8'h2c; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_44; // @[Reg.scala 27:20]
  wire [1:0] _T_22987 = _T_22519 ? bht_bank_rd_data_out_0_44 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23242 = _T_23241 | _T_22987; // @[Mux.scala 27:72]
  wire  _T_22521 = bht_rd_addr_hashed_p1_f == 8'h2d; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_45; // @[Reg.scala 27:20]
  wire [1:0] _T_22988 = _T_22521 ? bht_bank_rd_data_out_0_45 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23243 = _T_23242 | _T_22988; // @[Mux.scala 27:72]
  wire  _T_22523 = bht_rd_addr_hashed_p1_f == 8'h2e; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_46; // @[Reg.scala 27:20]
  wire [1:0] _T_22989 = _T_22523 ? bht_bank_rd_data_out_0_46 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23244 = _T_23243 | _T_22989; // @[Mux.scala 27:72]
  wire  _T_22525 = bht_rd_addr_hashed_p1_f == 8'h2f; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_47; // @[Reg.scala 27:20]
  wire [1:0] _T_22990 = _T_22525 ? bht_bank_rd_data_out_0_47 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23245 = _T_23244 | _T_22990; // @[Mux.scala 27:72]
  wire  _T_22527 = bht_rd_addr_hashed_p1_f == 8'h30; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_48; // @[Reg.scala 27:20]
  wire [1:0] _T_22991 = _T_22527 ? bht_bank_rd_data_out_0_48 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23246 = _T_23245 | _T_22991; // @[Mux.scala 27:72]
  wire  _T_22529 = bht_rd_addr_hashed_p1_f == 8'h31; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_49; // @[Reg.scala 27:20]
  wire [1:0] _T_22992 = _T_22529 ? bht_bank_rd_data_out_0_49 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23247 = _T_23246 | _T_22992; // @[Mux.scala 27:72]
  wire  _T_22531 = bht_rd_addr_hashed_p1_f == 8'h32; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_50; // @[Reg.scala 27:20]
  wire [1:0] _T_22993 = _T_22531 ? bht_bank_rd_data_out_0_50 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23248 = _T_23247 | _T_22993; // @[Mux.scala 27:72]
  wire  _T_22533 = bht_rd_addr_hashed_p1_f == 8'h33; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_51; // @[Reg.scala 27:20]
  wire [1:0] _T_22994 = _T_22533 ? bht_bank_rd_data_out_0_51 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23249 = _T_23248 | _T_22994; // @[Mux.scala 27:72]
  wire  _T_22535 = bht_rd_addr_hashed_p1_f == 8'h34; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_52; // @[Reg.scala 27:20]
  wire [1:0] _T_22995 = _T_22535 ? bht_bank_rd_data_out_0_52 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23250 = _T_23249 | _T_22995; // @[Mux.scala 27:72]
  wire  _T_22537 = bht_rd_addr_hashed_p1_f == 8'h35; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_53; // @[Reg.scala 27:20]
  wire [1:0] _T_22996 = _T_22537 ? bht_bank_rd_data_out_0_53 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23251 = _T_23250 | _T_22996; // @[Mux.scala 27:72]
  wire  _T_22539 = bht_rd_addr_hashed_p1_f == 8'h36; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_54; // @[Reg.scala 27:20]
  wire [1:0] _T_22997 = _T_22539 ? bht_bank_rd_data_out_0_54 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23252 = _T_23251 | _T_22997; // @[Mux.scala 27:72]
  wire  _T_22541 = bht_rd_addr_hashed_p1_f == 8'h37; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_55; // @[Reg.scala 27:20]
  wire [1:0] _T_22998 = _T_22541 ? bht_bank_rd_data_out_0_55 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23253 = _T_23252 | _T_22998; // @[Mux.scala 27:72]
  wire  _T_22543 = bht_rd_addr_hashed_p1_f == 8'h38; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_56; // @[Reg.scala 27:20]
  wire [1:0] _T_22999 = _T_22543 ? bht_bank_rd_data_out_0_56 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23254 = _T_23253 | _T_22999; // @[Mux.scala 27:72]
  wire  _T_22545 = bht_rd_addr_hashed_p1_f == 8'h39; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_57; // @[Reg.scala 27:20]
  wire [1:0] _T_23000 = _T_22545 ? bht_bank_rd_data_out_0_57 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23255 = _T_23254 | _T_23000; // @[Mux.scala 27:72]
  wire  _T_22547 = bht_rd_addr_hashed_p1_f == 8'h3a; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_58; // @[Reg.scala 27:20]
  wire [1:0] _T_23001 = _T_22547 ? bht_bank_rd_data_out_0_58 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23256 = _T_23255 | _T_23001; // @[Mux.scala 27:72]
  wire  _T_22549 = bht_rd_addr_hashed_p1_f == 8'h3b; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_59; // @[Reg.scala 27:20]
  wire [1:0] _T_23002 = _T_22549 ? bht_bank_rd_data_out_0_59 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23257 = _T_23256 | _T_23002; // @[Mux.scala 27:72]
  wire  _T_22551 = bht_rd_addr_hashed_p1_f == 8'h3c; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_60; // @[Reg.scala 27:20]
  wire [1:0] _T_23003 = _T_22551 ? bht_bank_rd_data_out_0_60 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23258 = _T_23257 | _T_23003; // @[Mux.scala 27:72]
  wire  _T_22553 = bht_rd_addr_hashed_p1_f == 8'h3d; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_61; // @[Reg.scala 27:20]
  wire [1:0] _T_23004 = _T_22553 ? bht_bank_rd_data_out_0_61 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23259 = _T_23258 | _T_23004; // @[Mux.scala 27:72]
  wire  _T_22555 = bht_rd_addr_hashed_p1_f == 8'h3e; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_62; // @[Reg.scala 27:20]
  wire [1:0] _T_23005 = _T_22555 ? bht_bank_rd_data_out_0_62 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23260 = _T_23259 | _T_23005; // @[Mux.scala 27:72]
  wire  _T_22557 = bht_rd_addr_hashed_p1_f == 8'h3f; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_63; // @[Reg.scala 27:20]
  wire [1:0] _T_23006 = _T_22557 ? bht_bank_rd_data_out_0_63 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23261 = _T_23260 | _T_23006; // @[Mux.scala 27:72]
  wire  _T_22559 = bht_rd_addr_hashed_p1_f == 8'h40; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_64; // @[Reg.scala 27:20]
  wire [1:0] _T_23007 = _T_22559 ? bht_bank_rd_data_out_0_64 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23262 = _T_23261 | _T_23007; // @[Mux.scala 27:72]
  wire  _T_22561 = bht_rd_addr_hashed_p1_f == 8'h41; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_65; // @[Reg.scala 27:20]
  wire [1:0] _T_23008 = _T_22561 ? bht_bank_rd_data_out_0_65 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23263 = _T_23262 | _T_23008; // @[Mux.scala 27:72]
  wire  _T_22563 = bht_rd_addr_hashed_p1_f == 8'h42; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_66; // @[Reg.scala 27:20]
  wire [1:0] _T_23009 = _T_22563 ? bht_bank_rd_data_out_0_66 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23264 = _T_23263 | _T_23009; // @[Mux.scala 27:72]
  wire  _T_22565 = bht_rd_addr_hashed_p1_f == 8'h43; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_67; // @[Reg.scala 27:20]
  wire [1:0] _T_23010 = _T_22565 ? bht_bank_rd_data_out_0_67 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23265 = _T_23264 | _T_23010; // @[Mux.scala 27:72]
  wire  _T_22567 = bht_rd_addr_hashed_p1_f == 8'h44; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_68; // @[Reg.scala 27:20]
  wire [1:0] _T_23011 = _T_22567 ? bht_bank_rd_data_out_0_68 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23266 = _T_23265 | _T_23011; // @[Mux.scala 27:72]
  wire  _T_22569 = bht_rd_addr_hashed_p1_f == 8'h45; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_69; // @[Reg.scala 27:20]
  wire [1:0] _T_23012 = _T_22569 ? bht_bank_rd_data_out_0_69 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23267 = _T_23266 | _T_23012; // @[Mux.scala 27:72]
  wire  _T_22571 = bht_rd_addr_hashed_p1_f == 8'h46; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_70; // @[Reg.scala 27:20]
  wire [1:0] _T_23013 = _T_22571 ? bht_bank_rd_data_out_0_70 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23268 = _T_23267 | _T_23013; // @[Mux.scala 27:72]
  wire  _T_22573 = bht_rd_addr_hashed_p1_f == 8'h47; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_71; // @[Reg.scala 27:20]
  wire [1:0] _T_23014 = _T_22573 ? bht_bank_rd_data_out_0_71 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23269 = _T_23268 | _T_23014; // @[Mux.scala 27:72]
  wire  _T_22575 = bht_rd_addr_hashed_p1_f == 8'h48; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_72; // @[Reg.scala 27:20]
  wire [1:0] _T_23015 = _T_22575 ? bht_bank_rd_data_out_0_72 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23270 = _T_23269 | _T_23015; // @[Mux.scala 27:72]
  wire  _T_22577 = bht_rd_addr_hashed_p1_f == 8'h49; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_73; // @[Reg.scala 27:20]
  wire [1:0] _T_23016 = _T_22577 ? bht_bank_rd_data_out_0_73 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23271 = _T_23270 | _T_23016; // @[Mux.scala 27:72]
  wire  _T_22579 = bht_rd_addr_hashed_p1_f == 8'h4a; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_74; // @[Reg.scala 27:20]
  wire [1:0] _T_23017 = _T_22579 ? bht_bank_rd_data_out_0_74 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23272 = _T_23271 | _T_23017; // @[Mux.scala 27:72]
  wire  _T_22581 = bht_rd_addr_hashed_p1_f == 8'h4b; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_75; // @[Reg.scala 27:20]
  wire [1:0] _T_23018 = _T_22581 ? bht_bank_rd_data_out_0_75 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23273 = _T_23272 | _T_23018; // @[Mux.scala 27:72]
  wire  _T_22583 = bht_rd_addr_hashed_p1_f == 8'h4c; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_76; // @[Reg.scala 27:20]
  wire [1:0] _T_23019 = _T_22583 ? bht_bank_rd_data_out_0_76 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23274 = _T_23273 | _T_23019; // @[Mux.scala 27:72]
  wire  _T_22585 = bht_rd_addr_hashed_p1_f == 8'h4d; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_77; // @[Reg.scala 27:20]
  wire [1:0] _T_23020 = _T_22585 ? bht_bank_rd_data_out_0_77 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23275 = _T_23274 | _T_23020; // @[Mux.scala 27:72]
  wire  _T_22587 = bht_rd_addr_hashed_p1_f == 8'h4e; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_78; // @[Reg.scala 27:20]
  wire [1:0] _T_23021 = _T_22587 ? bht_bank_rd_data_out_0_78 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23276 = _T_23275 | _T_23021; // @[Mux.scala 27:72]
  wire  _T_22589 = bht_rd_addr_hashed_p1_f == 8'h4f; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_79; // @[Reg.scala 27:20]
  wire [1:0] _T_23022 = _T_22589 ? bht_bank_rd_data_out_0_79 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23277 = _T_23276 | _T_23022; // @[Mux.scala 27:72]
  wire  _T_22591 = bht_rd_addr_hashed_p1_f == 8'h50; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_80; // @[Reg.scala 27:20]
  wire [1:0] _T_23023 = _T_22591 ? bht_bank_rd_data_out_0_80 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23278 = _T_23277 | _T_23023; // @[Mux.scala 27:72]
  wire  _T_22593 = bht_rd_addr_hashed_p1_f == 8'h51; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_81; // @[Reg.scala 27:20]
  wire [1:0] _T_23024 = _T_22593 ? bht_bank_rd_data_out_0_81 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23279 = _T_23278 | _T_23024; // @[Mux.scala 27:72]
  wire  _T_22595 = bht_rd_addr_hashed_p1_f == 8'h52; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_82; // @[Reg.scala 27:20]
  wire [1:0] _T_23025 = _T_22595 ? bht_bank_rd_data_out_0_82 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23280 = _T_23279 | _T_23025; // @[Mux.scala 27:72]
  wire  _T_22597 = bht_rd_addr_hashed_p1_f == 8'h53; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_83; // @[Reg.scala 27:20]
  wire [1:0] _T_23026 = _T_22597 ? bht_bank_rd_data_out_0_83 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23281 = _T_23280 | _T_23026; // @[Mux.scala 27:72]
  wire  _T_22599 = bht_rd_addr_hashed_p1_f == 8'h54; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_84; // @[Reg.scala 27:20]
  wire [1:0] _T_23027 = _T_22599 ? bht_bank_rd_data_out_0_84 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23282 = _T_23281 | _T_23027; // @[Mux.scala 27:72]
  wire  _T_22601 = bht_rd_addr_hashed_p1_f == 8'h55; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_85; // @[Reg.scala 27:20]
  wire [1:0] _T_23028 = _T_22601 ? bht_bank_rd_data_out_0_85 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23283 = _T_23282 | _T_23028; // @[Mux.scala 27:72]
  wire  _T_22603 = bht_rd_addr_hashed_p1_f == 8'h56; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_86; // @[Reg.scala 27:20]
  wire [1:0] _T_23029 = _T_22603 ? bht_bank_rd_data_out_0_86 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23284 = _T_23283 | _T_23029; // @[Mux.scala 27:72]
  wire  _T_22605 = bht_rd_addr_hashed_p1_f == 8'h57; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_87; // @[Reg.scala 27:20]
  wire [1:0] _T_23030 = _T_22605 ? bht_bank_rd_data_out_0_87 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23285 = _T_23284 | _T_23030; // @[Mux.scala 27:72]
  wire  _T_22607 = bht_rd_addr_hashed_p1_f == 8'h58; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_88; // @[Reg.scala 27:20]
  wire [1:0] _T_23031 = _T_22607 ? bht_bank_rd_data_out_0_88 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23286 = _T_23285 | _T_23031; // @[Mux.scala 27:72]
  wire  _T_22609 = bht_rd_addr_hashed_p1_f == 8'h59; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_89; // @[Reg.scala 27:20]
  wire [1:0] _T_23032 = _T_22609 ? bht_bank_rd_data_out_0_89 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23287 = _T_23286 | _T_23032; // @[Mux.scala 27:72]
  wire  _T_22611 = bht_rd_addr_hashed_p1_f == 8'h5a; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_90; // @[Reg.scala 27:20]
  wire [1:0] _T_23033 = _T_22611 ? bht_bank_rd_data_out_0_90 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23288 = _T_23287 | _T_23033; // @[Mux.scala 27:72]
  wire  _T_22613 = bht_rd_addr_hashed_p1_f == 8'h5b; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_91; // @[Reg.scala 27:20]
  wire [1:0] _T_23034 = _T_22613 ? bht_bank_rd_data_out_0_91 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23289 = _T_23288 | _T_23034; // @[Mux.scala 27:72]
  wire  _T_22615 = bht_rd_addr_hashed_p1_f == 8'h5c; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_92; // @[Reg.scala 27:20]
  wire [1:0] _T_23035 = _T_22615 ? bht_bank_rd_data_out_0_92 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23290 = _T_23289 | _T_23035; // @[Mux.scala 27:72]
  wire  _T_22617 = bht_rd_addr_hashed_p1_f == 8'h5d; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_93; // @[Reg.scala 27:20]
  wire [1:0] _T_23036 = _T_22617 ? bht_bank_rd_data_out_0_93 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23291 = _T_23290 | _T_23036; // @[Mux.scala 27:72]
  wire  _T_22619 = bht_rd_addr_hashed_p1_f == 8'h5e; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_94; // @[Reg.scala 27:20]
  wire [1:0] _T_23037 = _T_22619 ? bht_bank_rd_data_out_0_94 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23292 = _T_23291 | _T_23037; // @[Mux.scala 27:72]
  wire  _T_22621 = bht_rd_addr_hashed_p1_f == 8'h5f; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_95; // @[Reg.scala 27:20]
  wire [1:0] _T_23038 = _T_22621 ? bht_bank_rd_data_out_0_95 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23293 = _T_23292 | _T_23038; // @[Mux.scala 27:72]
  wire  _T_22623 = bht_rd_addr_hashed_p1_f == 8'h60; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_96; // @[Reg.scala 27:20]
  wire [1:0] _T_23039 = _T_22623 ? bht_bank_rd_data_out_0_96 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23294 = _T_23293 | _T_23039; // @[Mux.scala 27:72]
  wire  _T_22625 = bht_rd_addr_hashed_p1_f == 8'h61; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_97; // @[Reg.scala 27:20]
  wire [1:0] _T_23040 = _T_22625 ? bht_bank_rd_data_out_0_97 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23295 = _T_23294 | _T_23040; // @[Mux.scala 27:72]
  wire  _T_22627 = bht_rd_addr_hashed_p1_f == 8'h62; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_98; // @[Reg.scala 27:20]
  wire [1:0] _T_23041 = _T_22627 ? bht_bank_rd_data_out_0_98 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23296 = _T_23295 | _T_23041; // @[Mux.scala 27:72]
  wire  _T_22629 = bht_rd_addr_hashed_p1_f == 8'h63; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_99; // @[Reg.scala 27:20]
  wire [1:0] _T_23042 = _T_22629 ? bht_bank_rd_data_out_0_99 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23297 = _T_23296 | _T_23042; // @[Mux.scala 27:72]
  wire  _T_22631 = bht_rd_addr_hashed_p1_f == 8'h64; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_100; // @[Reg.scala 27:20]
  wire [1:0] _T_23043 = _T_22631 ? bht_bank_rd_data_out_0_100 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23298 = _T_23297 | _T_23043; // @[Mux.scala 27:72]
  wire  _T_22633 = bht_rd_addr_hashed_p1_f == 8'h65; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_101; // @[Reg.scala 27:20]
  wire [1:0] _T_23044 = _T_22633 ? bht_bank_rd_data_out_0_101 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23299 = _T_23298 | _T_23044; // @[Mux.scala 27:72]
  wire  _T_22635 = bht_rd_addr_hashed_p1_f == 8'h66; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_102; // @[Reg.scala 27:20]
  wire [1:0] _T_23045 = _T_22635 ? bht_bank_rd_data_out_0_102 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23300 = _T_23299 | _T_23045; // @[Mux.scala 27:72]
  wire  _T_22637 = bht_rd_addr_hashed_p1_f == 8'h67; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_103; // @[Reg.scala 27:20]
  wire [1:0] _T_23046 = _T_22637 ? bht_bank_rd_data_out_0_103 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23301 = _T_23300 | _T_23046; // @[Mux.scala 27:72]
  wire  _T_22639 = bht_rd_addr_hashed_p1_f == 8'h68; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_104; // @[Reg.scala 27:20]
  wire [1:0] _T_23047 = _T_22639 ? bht_bank_rd_data_out_0_104 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23302 = _T_23301 | _T_23047; // @[Mux.scala 27:72]
  wire  _T_22641 = bht_rd_addr_hashed_p1_f == 8'h69; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_105; // @[Reg.scala 27:20]
  wire [1:0] _T_23048 = _T_22641 ? bht_bank_rd_data_out_0_105 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23303 = _T_23302 | _T_23048; // @[Mux.scala 27:72]
  wire  _T_22643 = bht_rd_addr_hashed_p1_f == 8'h6a; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_106; // @[Reg.scala 27:20]
  wire [1:0] _T_23049 = _T_22643 ? bht_bank_rd_data_out_0_106 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23304 = _T_23303 | _T_23049; // @[Mux.scala 27:72]
  wire  _T_22645 = bht_rd_addr_hashed_p1_f == 8'h6b; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_107; // @[Reg.scala 27:20]
  wire [1:0] _T_23050 = _T_22645 ? bht_bank_rd_data_out_0_107 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23305 = _T_23304 | _T_23050; // @[Mux.scala 27:72]
  wire  _T_22647 = bht_rd_addr_hashed_p1_f == 8'h6c; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_108; // @[Reg.scala 27:20]
  wire [1:0] _T_23051 = _T_22647 ? bht_bank_rd_data_out_0_108 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23306 = _T_23305 | _T_23051; // @[Mux.scala 27:72]
  wire  _T_22649 = bht_rd_addr_hashed_p1_f == 8'h6d; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_109; // @[Reg.scala 27:20]
  wire [1:0] _T_23052 = _T_22649 ? bht_bank_rd_data_out_0_109 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23307 = _T_23306 | _T_23052; // @[Mux.scala 27:72]
  wire  _T_22651 = bht_rd_addr_hashed_p1_f == 8'h6e; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_110; // @[Reg.scala 27:20]
  wire [1:0] _T_23053 = _T_22651 ? bht_bank_rd_data_out_0_110 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23308 = _T_23307 | _T_23053; // @[Mux.scala 27:72]
  wire  _T_22653 = bht_rd_addr_hashed_p1_f == 8'h6f; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_111; // @[Reg.scala 27:20]
  wire [1:0] _T_23054 = _T_22653 ? bht_bank_rd_data_out_0_111 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23309 = _T_23308 | _T_23054; // @[Mux.scala 27:72]
  wire  _T_22655 = bht_rd_addr_hashed_p1_f == 8'h70; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_112; // @[Reg.scala 27:20]
  wire [1:0] _T_23055 = _T_22655 ? bht_bank_rd_data_out_0_112 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23310 = _T_23309 | _T_23055; // @[Mux.scala 27:72]
  wire  _T_22657 = bht_rd_addr_hashed_p1_f == 8'h71; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_113; // @[Reg.scala 27:20]
  wire [1:0] _T_23056 = _T_22657 ? bht_bank_rd_data_out_0_113 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23311 = _T_23310 | _T_23056; // @[Mux.scala 27:72]
  wire  _T_22659 = bht_rd_addr_hashed_p1_f == 8'h72; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_114; // @[Reg.scala 27:20]
  wire [1:0] _T_23057 = _T_22659 ? bht_bank_rd_data_out_0_114 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23312 = _T_23311 | _T_23057; // @[Mux.scala 27:72]
  wire  _T_22661 = bht_rd_addr_hashed_p1_f == 8'h73; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_115; // @[Reg.scala 27:20]
  wire [1:0] _T_23058 = _T_22661 ? bht_bank_rd_data_out_0_115 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23313 = _T_23312 | _T_23058; // @[Mux.scala 27:72]
  wire  _T_22663 = bht_rd_addr_hashed_p1_f == 8'h74; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_116; // @[Reg.scala 27:20]
  wire [1:0] _T_23059 = _T_22663 ? bht_bank_rd_data_out_0_116 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23314 = _T_23313 | _T_23059; // @[Mux.scala 27:72]
  wire  _T_22665 = bht_rd_addr_hashed_p1_f == 8'h75; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_117; // @[Reg.scala 27:20]
  wire [1:0] _T_23060 = _T_22665 ? bht_bank_rd_data_out_0_117 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23315 = _T_23314 | _T_23060; // @[Mux.scala 27:72]
  wire  _T_22667 = bht_rd_addr_hashed_p1_f == 8'h76; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_118; // @[Reg.scala 27:20]
  wire [1:0] _T_23061 = _T_22667 ? bht_bank_rd_data_out_0_118 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23316 = _T_23315 | _T_23061; // @[Mux.scala 27:72]
  wire  _T_22669 = bht_rd_addr_hashed_p1_f == 8'h77; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_119; // @[Reg.scala 27:20]
  wire [1:0] _T_23062 = _T_22669 ? bht_bank_rd_data_out_0_119 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23317 = _T_23316 | _T_23062; // @[Mux.scala 27:72]
  wire  _T_22671 = bht_rd_addr_hashed_p1_f == 8'h78; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_120; // @[Reg.scala 27:20]
  wire [1:0] _T_23063 = _T_22671 ? bht_bank_rd_data_out_0_120 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23318 = _T_23317 | _T_23063; // @[Mux.scala 27:72]
  wire  _T_22673 = bht_rd_addr_hashed_p1_f == 8'h79; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_121; // @[Reg.scala 27:20]
  wire [1:0] _T_23064 = _T_22673 ? bht_bank_rd_data_out_0_121 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23319 = _T_23318 | _T_23064; // @[Mux.scala 27:72]
  wire  _T_22675 = bht_rd_addr_hashed_p1_f == 8'h7a; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_122; // @[Reg.scala 27:20]
  wire [1:0] _T_23065 = _T_22675 ? bht_bank_rd_data_out_0_122 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23320 = _T_23319 | _T_23065; // @[Mux.scala 27:72]
  wire  _T_22677 = bht_rd_addr_hashed_p1_f == 8'h7b; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_123; // @[Reg.scala 27:20]
  wire [1:0] _T_23066 = _T_22677 ? bht_bank_rd_data_out_0_123 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23321 = _T_23320 | _T_23066; // @[Mux.scala 27:72]
  wire  _T_22679 = bht_rd_addr_hashed_p1_f == 8'h7c; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_124; // @[Reg.scala 27:20]
  wire [1:0] _T_23067 = _T_22679 ? bht_bank_rd_data_out_0_124 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23322 = _T_23321 | _T_23067; // @[Mux.scala 27:72]
  wire  _T_22681 = bht_rd_addr_hashed_p1_f == 8'h7d; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_125; // @[Reg.scala 27:20]
  wire [1:0] _T_23068 = _T_22681 ? bht_bank_rd_data_out_0_125 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23323 = _T_23322 | _T_23068; // @[Mux.scala 27:72]
  wire  _T_22683 = bht_rd_addr_hashed_p1_f == 8'h7e; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_126; // @[Reg.scala 27:20]
  wire [1:0] _T_23069 = _T_22683 ? bht_bank_rd_data_out_0_126 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23324 = _T_23323 | _T_23069; // @[Mux.scala 27:72]
  wire  _T_22685 = bht_rd_addr_hashed_p1_f == 8'h7f; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_127; // @[Reg.scala 27:20]
  wire [1:0] _T_23070 = _T_22685 ? bht_bank_rd_data_out_0_127 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23325 = _T_23324 | _T_23070; // @[Mux.scala 27:72]
  wire  _T_22687 = bht_rd_addr_hashed_p1_f == 8'h80; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_128; // @[Reg.scala 27:20]
  wire [1:0] _T_23071 = _T_22687 ? bht_bank_rd_data_out_0_128 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23326 = _T_23325 | _T_23071; // @[Mux.scala 27:72]
  wire  _T_22689 = bht_rd_addr_hashed_p1_f == 8'h81; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_129; // @[Reg.scala 27:20]
  wire [1:0] _T_23072 = _T_22689 ? bht_bank_rd_data_out_0_129 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23327 = _T_23326 | _T_23072; // @[Mux.scala 27:72]
  wire  _T_22691 = bht_rd_addr_hashed_p1_f == 8'h82; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_130; // @[Reg.scala 27:20]
  wire [1:0] _T_23073 = _T_22691 ? bht_bank_rd_data_out_0_130 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23328 = _T_23327 | _T_23073; // @[Mux.scala 27:72]
  wire  _T_22693 = bht_rd_addr_hashed_p1_f == 8'h83; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_131; // @[Reg.scala 27:20]
  wire [1:0] _T_23074 = _T_22693 ? bht_bank_rd_data_out_0_131 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23329 = _T_23328 | _T_23074; // @[Mux.scala 27:72]
  wire  _T_22695 = bht_rd_addr_hashed_p1_f == 8'h84; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_132; // @[Reg.scala 27:20]
  wire [1:0] _T_23075 = _T_22695 ? bht_bank_rd_data_out_0_132 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23330 = _T_23329 | _T_23075; // @[Mux.scala 27:72]
  wire  _T_22697 = bht_rd_addr_hashed_p1_f == 8'h85; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_133; // @[Reg.scala 27:20]
  wire [1:0] _T_23076 = _T_22697 ? bht_bank_rd_data_out_0_133 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23331 = _T_23330 | _T_23076; // @[Mux.scala 27:72]
  wire  _T_22699 = bht_rd_addr_hashed_p1_f == 8'h86; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_134; // @[Reg.scala 27:20]
  wire [1:0] _T_23077 = _T_22699 ? bht_bank_rd_data_out_0_134 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23332 = _T_23331 | _T_23077; // @[Mux.scala 27:72]
  wire  _T_22701 = bht_rd_addr_hashed_p1_f == 8'h87; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_135; // @[Reg.scala 27:20]
  wire [1:0] _T_23078 = _T_22701 ? bht_bank_rd_data_out_0_135 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23333 = _T_23332 | _T_23078; // @[Mux.scala 27:72]
  wire  _T_22703 = bht_rd_addr_hashed_p1_f == 8'h88; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_136; // @[Reg.scala 27:20]
  wire [1:0] _T_23079 = _T_22703 ? bht_bank_rd_data_out_0_136 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23334 = _T_23333 | _T_23079; // @[Mux.scala 27:72]
  wire  _T_22705 = bht_rd_addr_hashed_p1_f == 8'h89; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_137; // @[Reg.scala 27:20]
  wire [1:0] _T_23080 = _T_22705 ? bht_bank_rd_data_out_0_137 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23335 = _T_23334 | _T_23080; // @[Mux.scala 27:72]
  wire  _T_22707 = bht_rd_addr_hashed_p1_f == 8'h8a; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_138; // @[Reg.scala 27:20]
  wire [1:0] _T_23081 = _T_22707 ? bht_bank_rd_data_out_0_138 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23336 = _T_23335 | _T_23081; // @[Mux.scala 27:72]
  wire  _T_22709 = bht_rd_addr_hashed_p1_f == 8'h8b; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_139; // @[Reg.scala 27:20]
  wire [1:0] _T_23082 = _T_22709 ? bht_bank_rd_data_out_0_139 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23337 = _T_23336 | _T_23082; // @[Mux.scala 27:72]
  wire  _T_22711 = bht_rd_addr_hashed_p1_f == 8'h8c; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_140; // @[Reg.scala 27:20]
  wire [1:0] _T_23083 = _T_22711 ? bht_bank_rd_data_out_0_140 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23338 = _T_23337 | _T_23083; // @[Mux.scala 27:72]
  wire  _T_22713 = bht_rd_addr_hashed_p1_f == 8'h8d; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_141; // @[Reg.scala 27:20]
  wire [1:0] _T_23084 = _T_22713 ? bht_bank_rd_data_out_0_141 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23339 = _T_23338 | _T_23084; // @[Mux.scala 27:72]
  wire  _T_22715 = bht_rd_addr_hashed_p1_f == 8'h8e; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_142; // @[Reg.scala 27:20]
  wire [1:0] _T_23085 = _T_22715 ? bht_bank_rd_data_out_0_142 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23340 = _T_23339 | _T_23085; // @[Mux.scala 27:72]
  wire  _T_22717 = bht_rd_addr_hashed_p1_f == 8'h8f; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_143; // @[Reg.scala 27:20]
  wire [1:0] _T_23086 = _T_22717 ? bht_bank_rd_data_out_0_143 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23341 = _T_23340 | _T_23086; // @[Mux.scala 27:72]
  wire  _T_22719 = bht_rd_addr_hashed_p1_f == 8'h90; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_144; // @[Reg.scala 27:20]
  wire [1:0] _T_23087 = _T_22719 ? bht_bank_rd_data_out_0_144 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23342 = _T_23341 | _T_23087; // @[Mux.scala 27:72]
  wire  _T_22721 = bht_rd_addr_hashed_p1_f == 8'h91; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_145; // @[Reg.scala 27:20]
  wire [1:0] _T_23088 = _T_22721 ? bht_bank_rd_data_out_0_145 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23343 = _T_23342 | _T_23088; // @[Mux.scala 27:72]
  wire  _T_22723 = bht_rd_addr_hashed_p1_f == 8'h92; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_146; // @[Reg.scala 27:20]
  wire [1:0] _T_23089 = _T_22723 ? bht_bank_rd_data_out_0_146 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23344 = _T_23343 | _T_23089; // @[Mux.scala 27:72]
  wire  _T_22725 = bht_rd_addr_hashed_p1_f == 8'h93; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_147; // @[Reg.scala 27:20]
  wire [1:0] _T_23090 = _T_22725 ? bht_bank_rd_data_out_0_147 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23345 = _T_23344 | _T_23090; // @[Mux.scala 27:72]
  wire  _T_22727 = bht_rd_addr_hashed_p1_f == 8'h94; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_148; // @[Reg.scala 27:20]
  wire [1:0] _T_23091 = _T_22727 ? bht_bank_rd_data_out_0_148 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23346 = _T_23345 | _T_23091; // @[Mux.scala 27:72]
  wire  _T_22729 = bht_rd_addr_hashed_p1_f == 8'h95; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_149; // @[Reg.scala 27:20]
  wire [1:0] _T_23092 = _T_22729 ? bht_bank_rd_data_out_0_149 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23347 = _T_23346 | _T_23092; // @[Mux.scala 27:72]
  wire  _T_22731 = bht_rd_addr_hashed_p1_f == 8'h96; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_150; // @[Reg.scala 27:20]
  wire [1:0] _T_23093 = _T_22731 ? bht_bank_rd_data_out_0_150 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23348 = _T_23347 | _T_23093; // @[Mux.scala 27:72]
  wire  _T_22733 = bht_rd_addr_hashed_p1_f == 8'h97; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_151; // @[Reg.scala 27:20]
  wire [1:0] _T_23094 = _T_22733 ? bht_bank_rd_data_out_0_151 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23349 = _T_23348 | _T_23094; // @[Mux.scala 27:72]
  wire  _T_22735 = bht_rd_addr_hashed_p1_f == 8'h98; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_152; // @[Reg.scala 27:20]
  wire [1:0] _T_23095 = _T_22735 ? bht_bank_rd_data_out_0_152 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23350 = _T_23349 | _T_23095; // @[Mux.scala 27:72]
  wire  _T_22737 = bht_rd_addr_hashed_p1_f == 8'h99; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_153; // @[Reg.scala 27:20]
  wire [1:0] _T_23096 = _T_22737 ? bht_bank_rd_data_out_0_153 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23351 = _T_23350 | _T_23096; // @[Mux.scala 27:72]
  wire  _T_22739 = bht_rd_addr_hashed_p1_f == 8'h9a; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_154; // @[Reg.scala 27:20]
  wire [1:0] _T_23097 = _T_22739 ? bht_bank_rd_data_out_0_154 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23352 = _T_23351 | _T_23097; // @[Mux.scala 27:72]
  wire  _T_22741 = bht_rd_addr_hashed_p1_f == 8'h9b; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_155; // @[Reg.scala 27:20]
  wire [1:0] _T_23098 = _T_22741 ? bht_bank_rd_data_out_0_155 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23353 = _T_23352 | _T_23098; // @[Mux.scala 27:72]
  wire  _T_22743 = bht_rd_addr_hashed_p1_f == 8'h9c; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_156; // @[Reg.scala 27:20]
  wire [1:0] _T_23099 = _T_22743 ? bht_bank_rd_data_out_0_156 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23354 = _T_23353 | _T_23099; // @[Mux.scala 27:72]
  wire  _T_22745 = bht_rd_addr_hashed_p1_f == 8'h9d; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_157; // @[Reg.scala 27:20]
  wire [1:0] _T_23100 = _T_22745 ? bht_bank_rd_data_out_0_157 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23355 = _T_23354 | _T_23100; // @[Mux.scala 27:72]
  wire  _T_22747 = bht_rd_addr_hashed_p1_f == 8'h9e; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_158; // @[Reg.scala 27:20]
  wire [1:0] _T_23101 = _T_22747 ? bht_bank_rd_data_out_0_158 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23356 = _T_23355 | _T_23101; // @[Mux.scala 27:72]
  wire  _T_22749 = bht_rd_addr_hashed_p1_f == 8'h9f; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_159; // @[Reg.scala 27:20]
  wire [1:0] _T_23102 = _T_22749 ? bht_bank_rd_data_out_0_159 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23357 = _T_23356 | _T_23102; // @[Mux.scala 27:72]
  wire  _T_22751 = bht_rd_addr_hashed_p1_f == 8'ha0; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_160; // @[Reg.scala 27:20]
  wire [1:0] _T_23103 = _T_22751 ? bht_bank_rd_data_out_0_160 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23358 = _T_23357 | _T_23103; // @[Mux.scala 27:72]
  wire  _T_22753 = bht_rd_addr_hashed_p1_f == 8'ha1; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_161; // @[Reg.scala 27:20]
  wire [1:0] _T_23104 = _T_22753 ? bht_bank_rd_data_out_0_161 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23359 = _T_23358 | _T_23104; // @[Mux.scala 27:72]
  wire  _T_22755 = bht_rd_addr_hashed_p1_f == 8'ha2; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_162; // @[Reg.scala 27:20]
  wire [1:0] _T_23105 = _T_22755 ? bht_bank_rd_data_out_0_162 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23360 = _T_23359 | _T_23105; // @[Mux.scala 27:72]
  wire  _T_22757 = bht_rd_addr_hashed_p1_f == 8'ha3; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_163; // @[Reg.scala 27:20]
  wire [1:0] _T_23106 = _T_22757 ? bht_bank_rd_data_out_0_163 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23361 = _T_23360 | _T_23106; // @[Mux.scala 27:72]
  wire  _T_22759 = bht_rd_addr_hashed_p1_f == 8'ha4; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_164; // @[Reg.scala 27:20]
  wire [1:0] _T_23107 = _T_22759 ? bht_bank_rd_data_out_0_164 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23362 = _T_23361 | _T_23107; // @[Mux.scala 27:72]
  wire  _T_22761 = bht_rd_addr_hashed_p1_f == 8'ha5; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_165; // @[Reg.scala 27:20]
  wire [1:0] _T_23108 = _T_22761 ? bht_bank_rd_data_out_0_165 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23363 = _T_23362 | _T_23108; // @[Mux.scala 27:72]
  wire  _T_22763 = bht_rd_addr_hashed_p1_f == 8'ha6; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_166; // @[Reg.scala 27:20]
  wire [1:0] _T_23109 = _T_22763 ? bht_bank_rd_data_out_0_166 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23364 = _T_23363 | _T_23109; // @[Mux.scala 27:72]
  wire  _T_22765 = bht_rd_addr_hashed_p1_f == 8'ha7; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_167; // @[Reg.scala 27:20]
  wire [1:0] _T_23110 = _T_22765 ? bht_bank_rd_data_out_0_167 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23365 = _T_23364 | _T_23110; // @[Mux.scala 27:72]
  wire  _T_22767 = bht_rd_addr_hashed_p1_f == 8'ha8; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_168; // @[Reg.scala 27:20]
  wire [1:0] _T_23111 = _T_22767 ? bht_bank_rd_data_out_0_168 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23366 = _T_23365 | _T_23111; // @[Mux.scala 27:72]
  wire  _T_22769 = bht_rd_addr_hashed_p1_f == 8'ha9; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_169; // @[Reg.scala 27:20]
  wire [1:0] _T_23112 = _T_22769 ? bht_bank_rd_data_out_0_169 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23367 = _T_23366 | _T_23112; // @[Mux.scala 27:72]
  wire  _T_22771 = bht_rd_addr_hashed_p1_f == 8'haa; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_170; // @[Reg.scala 27:20]
  wire [1:0] _T_23113 = _T_22771 ? bht_bank_rd_data_out_0_170 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23368 = _T_23367 | _T_23113; // @[Mux.scala 27:72]
  wire  _T_22773 = bht_rd_addr_hashed_p1_f == 8'hab; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_171; // @[Reg.scala 27:20]
  wire [1:0] _T_23114 = _T_22773 ? bht_bank_rd_data_out_0_171 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23369 = _T_23368 | _T_23114; // @[Mux.scala 27:72]
  wire  _T_22775 = bht_rd_addr_hashed_p1_f == 8'hac; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_172; // @[Reg.scala 27:20]
  wire [1:0] _T_23115 = _T_22775 ? bht_bank_rd_data_out_0_172 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23370 = _T_23369 | _T_23115; // @[Mux.scala 27:72]
  wire  _T_22777 = bht_rd_addr_hashed_p1_f == 8'had; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_173; // @[Reg.scala 27:20]
  wire [1:0] _T_23116 = _T_22777 ? bht_bank_rd_data_out_0_173 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23371 = _T_23370 | _T_23116; // @[Mux.scala 27:72]
  wire  _T_22779 = bht_rd_addr_hashed_p1_f == 8'hae; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_174; // @[Reg.scala 27:20]
  wire [1:0] _T_23117 = _T_22779 ? bht_bank_rd_data_out_0_174 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23372 = _T_23371 | _T_23117; // @[Mux.scala 27:72]
  wire  _T_22781 = bht_rd_addr_hashed_p1_f == 8'haf; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_175; // @[Reg.scala 27:20]
  wire [1:0] _T_23118 = _T_22781 ? bht_bank_rd_data_out_0_175 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23373 = _T_23372 | _T_23118; // @[Mux.scala 27:72]
  wire  _T_22783 = bht_rd_addr_hashed_p1_f == 8'hb0; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_176; // @[Reg.scala 27:20]
  wire [1:0] _T_23119 = _T_22783 ? bht_bank_rd_data_out_0_176 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23374 = _T_23373 | _T_23119; // @[Mux.scala 27:72]
  wire  _T_22785 = bht_rd_addr_hashed_p1_f == 8'hb1; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_177; // @[Reg.scala 27:20]
  wire [1:0] _T_23120 = _T_22785 ? bht_bank_rd_data_out_0_177 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23375 = _T_23374 | _T_23120; // @[Mux.scala 27:72]
  wire  _T_22787 = bht_rd_addr_hashed_p1_f == 8'hb2; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_178; // @[Reg.scala 27:20]
  wire [1:0] _T_23121 = _T_22787 ? bht_bank_rd_data_out_0_178 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23376 = _T_23375 | _T_23121; // @[Mux.scala 27:72]
  wire  _T_22789 = bht_rd_addr_hashed_p1_f == 8'hb3; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_179; // @[Reg.scala 27:20]
  wire [1:0] _T_23122 = _T_22789 ? bht_bank_rd_data_out_0_179 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23377 = _T_23376 | _T_23122; // @[Mux.scala 27:72]
  wire  _T_22791 = bht_rd_addr_hashed_p1_f == 8'hb4; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_180; // @[Reg.scala 27:20]
  wire [1:0] _T_23123 = _T_22791 ? bht_bank_rd_data_out_0_180 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23378 = _T_23377 | _T_23123; // @[Mux.scala 27:72]
  wire  _T_22793 = bht_rd_addr_hashed_p1_f == 8'hb5; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_181; // @[Reg.scala 27:20]
  wire [1:0] _T_23124 = _T_22793 ? bht_bank_rd_data_out_0_181 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23379 = _T_23378 | _T_23124; // @[Mux.scala 27:72]
  wire  _T_22795 = bht_rd_addr_hashed_p1_f == 8'hb6; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_182; // @[Reg.scala 27:20]
  wire [1:0] _T_23125 = _T_22795 ? bht_bank_rd_data_out_0_182 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23380 = _T_23379 | _T_23125; // @[Mux.scala 27:72]
  wire  _T_22797 = bht_rd_addr_hashed_p1_f == 8'hb7; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_183; // @[Reg.scala 27:20]
  wire [1:0] _T_23126 = _T_22797 ? bht_bank_rd_data_out_0_183 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23381 = _T_23380 | _T_23126; // @[Mux.scala 27:72]
  wire  _T_22799 = bht_rd_addr_hashed_p1_f == 8'hb8; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_184; // @[Reg.scala 27:20]
  wire [1:0] _T_23127 = _T_22799 ? bht_bank_rd_data_out_0_184 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23382 = _T_23381 | _T_23127; // @[Mux.scala 27:72]
  wire  _T_22801 = bht_rd_addr_hashed_p1_f == 8'hb9; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_185; // @[Reg.scala 27:20]
  wire [1:0] _T_23128 = _T_22801 ? bht_bank_rd_data_out_0_185 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23383 = _T_23382 | _T_23128; // @[Mux.scala 27:72]
  wire  _T_22803 = bht_rd_addr_hashed_p1_f == 8'hba; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_186; // @[Reg.scala 27:20]
  wire [1:0] _T_23129 = _T_22803 ? bht_bank_rd_data_out_0_186 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23384 = _T_23383 | _T_23129; // @[Mux.scala 27:72]
  wire  _T_22805 = bht_rd_addr_hashed_p1_f == 8'hbb; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_187; // @[Reg.scala 27:20]
  wire [1:0] _T_23130 = _T_22805 ? bht_bank_rd_data_out_0_187 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23385 = _T_23384 | _T_23130; // @[Mux.scala 27:72]
  wire  _T_22807 = bht_rd_addr_hashed_p1_f == 8'hbc; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_188; // @[Reg.scala 27:20]
  wire [1:0] _T_23131 = _T_22807 ? bht_bank_rd_data_out_0_188 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23386 = _T_23385 | _T_23131; // @[Mux.scala 27:72]
  wire  _T_22809 = bht_rd_addr_hashed_p1_f == 8'hbd; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_189; // @[Reg.scala 27:20]
  wire [1:0] _T_23132 = _T_22809 ? bht_bank_rd_data_out_0_189 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23387 = _T_23386 | _T_23132; // @[Mux.scala 27:72]
  wire  _T_22811 = bht_rd_addr_hashed_p1_f == 8'hbe; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_190; // @[Reg.scala 27:20]
  wire [1:0] _T_23133 = _T_22811 ? bht_bank_rd_data_out_0_190 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23388 = _T_23387 | _T_23133; // @[Mux.scala 27:72]
  wire  _T_22813 = bht_rd_addr_hashed_p1_f == 8'hbf; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_191; // @[Reg.scala 27:20]
  wire [1:0] _T_23134 = _T_22813 ? bht_bank_rd_data_out_0_191 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23389 = _T_23388 | _T_23134; // @[Mux.scala 27:72]
  wire  _T_22815 = bht_rd_addr_hashed_p1_f == 8'hc0; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_192; // @[Reg.scala 27:20]
  wire [1:0] _T_23135 = _T_22815 ? bht_bank_rd_data_out_0_192 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23390 = _T_23389 | _T_23135; // @[Mux.scala 27:72]
  wire  _T_22817 = bht_rd_addr_hashed_p1_f == 8'hc1; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_193; // @[Reg.scala 27:20]
  wire [1:0] _T_23136 = _T_22817 ? bht_bank_rd_data_out_0_193 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23391 = _T_23390 | _T_23136; // @[Mux.scala 27:72]
  wire  _T_22819 = bht_rd_addr_hashed_p1_f == 8'hc2; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_194; // @[Reg.scala 27:20]
  wire [1:0] _T_23137 = _T_22819 ? bht_bank_rd_data_out_0_194 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23392 = _T_23391 | _T_23137; // @[Mux.scala 27:72]
  wire  _T_22821 = bht_rd_addr_hashed_p1_f == 8'hc3; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_195; // @[Reg.scala 27:20]
  wire [1:0] _T_23138 = _T_22821 ? bht_bank_rd_data_out_0_195 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23393 = _T_23392 | _T_23138; // @[Mux.scala 27:72]
  wire  _T_22823 = bht_rd_addr_hashed_p1_f == 8'hc4; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_196; // @[Reg.scala 27:20]
  wire [1:0] _T_23139 = _T_22823 ? bht_bank_rd_data_out_0_196 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23394 = _T_23393 | _T_23139; // @[Mux.scala 27:72]
  wire  _T_22825 = bht_rd_addr_hashed_p1_f == 8'hc5; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_197; // @[Reg.scala 27:20]
  wire [1:0] _T_23140 = _T_22825 ? bht_bank_rd_data_out_0_197 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23395 = _T_23394 | _T_23140; // @[Mux.scala 27:72]
  wire  _T_22827 = bht_rd_addr_hashed_p1_f == 8'hc6; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_198; // @[Reg.scala 27:20]
  wire [1:0] _T_23141 = _T_22827 ? bht_bank_rd_data_out_0_198 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23396 = _T_23395 | _T_23141; // @[Mux.scala 27:72]
  wire  _T_22829 = bht_rd_addr_hashed_p1_f == 8'hc7; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_199; // @[Reg.scala 27:20]
  wire [1:0] _T_23142 = _T_22829 ? bht_bank_rd_data_out_0_199 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23397 = _T_23396 | _T_23142; // @[Mux.scala 27:72]
  wire  _T_22831 = bht_rd_addr_hashed_p1_f == 8'hc8; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_200; // @[Reg.scala 27:20]
  wire [1:0] _T_23143 = _T_22831 ? bht_bank_rd_data_out_0_200 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23398 = _T_23397 | _T_23143; // @[Mux.scala 27:72]
  wire  _T_22833 = bht_rd_addr_hashed_p1_f == 8'hc9; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_201; // @[Reg.scala 27:20]
  wire [1:0] _T_23144 = _T_22833 ? bht_bank_rd_data_out_0_201 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23399 = _T_23398 | _T_23144; // @[Mux.scala 27:72]
  wire  _T_22835 = bht_rd_addr_hashed_p1_f == 8'hca; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_202; // @[Reg.scala 27:20]
  wire [1:0] _T_23145 = _T_22835 ? bht_bank_rd_data_out_0_202 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23400 = _T_23399 | _T_23145; // @[Mux.scala 27:72]
  wire  _T_22837 = bht_rd_addr_hashed_p1_f == 8'hcb; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_203; // @[Reg.scala 27:20]
  wire [1:0] _T_23146 = _T_22837 ? bht_bank_rd_data_out_0_203 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23401 = _T_23400 | _T_23146; // @[Mux.scala 27:72]
  wire  _T_22839 = bht_rd_addr_hashed_p1_f == 8'hcc; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_204; // @[Reg.scala 27:20]
  wire [1:0] _T_23147 = _T_22839 ? bht_bank_rd_data_out_0_204 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23402 = _T_23401 | _T_23147; // @[Mux.scala 27:72]
  wire  _T_22841 = bht_rd_addr_hashed_p1_f == 8'hcd; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_205; // @[Reg.scala 27:20]
  wire [1:0] _T_23148 = _T_22841 ? bht_bank_rd_data_out_0_205 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23403 = _T_23402 | _T_23148; // @[Mux.scala 27:72]
  wire  _T_22843 = bht_rd_addr_hashed_p1_f == 8'hce; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_206; // @[Reg.scala 27:20]
  wire [1:0] _T_23149 = _T_22843 ? bht_bank_rd_data_out_0_206 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23404 = _T_23403 | _T_23149; // @[Mux.scala 27:72]
  wire  _T_22845 = bht_rd_addr_hashed_p1_f == 8'hcf; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_207; // @[Reg.scala 27:20]
  wire [1:0] _T_23150 = _T_22845 ? bht_bank_rd_data_out_0_207 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23405 = _T_23404 | _T_23150; // @[Mux.scala 27:72]
  wire  _T_22847 = bht_rd_addr_hashed_p1_f == 8'hd0; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_208; // @[Reg.scala 27:20]
  wire [1:0] _T_23151 = _T_22847 ? bht_bank_rd_data_out_0_208 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23406 = _T_23405 | _T_23151; // @[Mux.scala 27:72]
  wire  _T_22849 = bht_rd_addr_hashed_p1_f == 8'hd1; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_209; // @[Reg.scala 27:20]
  wire [1:0] _T_23152 = _T_22849 ? bht_bank_rd_data_out_0_209 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23407 = _T_23406 | _T_23152; // @[Mux.scala 27:72]
  wire  _T_22851 = bht_rd_addr_hashed_p1_f == 8'hd2; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_210; // @[Reg.scala 27:20]
  wire [1:0] _T_23153 = _T_22851 ? bht_bank_rd_data_out_0_210 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23408 = _T_23407 | _T_23153; // @[Mux.scala 27:72]
  wire  _T_22853 = bht_rd_addr_hashed_p1_f == 8'hd3; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_211; // @[Reg.scala 27:20]
  wire [1:0] _T_23154 = _T_22853 ? bht_bank_rd_data_out_0_211 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23409 = _T_23408 | _T_23154; // @[Mux.scala 27:72]
  wire  _T_22855 = bht_rd_addr_hashed_p1_f == 8'hd4; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_212; // @[Reg.scala 27:20]
  wire [1:0] _T_23155 = _T_22855 ? bht_bank_rd_data_out_0_212 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23410 = _T_23409 | _T_23155; // @[Mux.scala 27:72]
  wire  _T_22857 = bht_rd_addr_hashed_p1_f == 8'hd5; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_213; // @[Reg.scala 27:20]
  wire [1:0] _T_23156 = _T_22857 ? bht_bank_rd_data_out_0_213 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23411 = _T_23410 | _T_23156; // @[Mux.scala 27:72]
  wire  _T_22859 = bht_rd_addr_hashed_p1_f == 8'hd6; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_214; // @[Reg.scala 27:20]
  wire [1:0] _T_23157 = _T_22859 ? bht_bank_rd_data_out_0_214 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23412 = _T_23411 | _T_23157; // @[Mux.scala 27:72]
  wire  _T_22861 = bht_rd_addr_hashed_p1_f == 8'hd7; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_215; // @[Reg.scala 27:20]
  wire [1:0] _T_23158 = _T_22861 ? bht_bank_rd_data_out_0_215 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23413 = _T_23412 | _T_23158; // @[Mux.scala 27:72]
  wire  _T_22863 = bht_rd_addr_hashed_p1_f == 8'hd8; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_216; // @[Reg.scala 27:20]
  wire [1:0] _T_23159 = _T_22863 ? bht_bank_rd_data_out_0_216 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23414 = _T_23413 | _T_23159; // @[Mux.scala 27:72]
  wire  _T_22865 = bht_rd_addr_hashed_p1_f == 8'hd9; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_217; // @[Reg.scala 27:20]
  wire [1:0] _T_23160 = _T_22865 ? bht_bank_rd_data_out_0_217 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23415 = _T_23414 | _T_23160; // @[Mux.scala 27:72]
  wire  _T_22867 = bht_rd_addr_hashed_p1_f == 8'hda; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_218; // @[Reg.scala 27:20]
  wire [1:0] _T_23161 = _T_22867 ? bht_bank_rd_data_out_0_218 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23416 = _T_23415 | _T_23161; // @[Mux.scala 27:72]
  wire  _T_22869 = bht_rd_addr_hashed_p1_f == 8'hdb; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_219; // @[Reg.scala 27:20]
  wire [1:0] _T_23162 = _T_22869 ? bht_bank_rd_data_out_0_219 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23417 = _T_23416 | _T_23162; // @[Mux.scala 27:72]
  wire  _T_22871 = bht_rd_addr_hashed_p1_f == 8'hdc; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_220; // @[Reg.scala 27:20]
  wire [1:0] _T_23163 = _T_22871 ? bht_bank_rd_data_out_0_220 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23418 = _T_23417 | _T_23163; // @[Mux.scala 27:72]
  wire  _T_22873 = bht_rd_addr_hashed_p1_f == 8'hdd; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_221; // @[Reg.scala 27:20]
  wire [1:0] _T_23164 = _T_22873 ? bht_bank_rd_data_out_0_221 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23419 = _T_23418 | _T_23164; // @[Mux.scala 27:72]
  wire  _T_22875 = bht_rd_addr_hashed_p1_f == 8'hde; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_222; // @[Reg.scala 27:20]
  wire [1:0] _T_23165 = _T_22875 ? bht_bank_rd_data_out_0_222 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23420 = _T_23419 | _T_23165; // @[Mux.scala 27:72]
  wire  _T_22877 = bht_rd_addr_hashed_p1_f == 8'hdf; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_223; // @[Reg.scala 27:20]
  wire [1:0] _T_23166 = _T_22877 ? bht_bank_rd_data_out_0_223 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23421 = _T_23420 | _T_23166; // @[Mux.scala 27:72]
  wire  _T_22879 = bht_rd_addr_hashed_p1_f == 8'he0; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_224; // @[Reg.scala 27:20]
  wire [1:0] _T_23167 = _T_22879 ? bht_bank_rd_data_out_0_224 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23422 = _T_23421 | _T_23167; // @[Mux.scala 27:72]
  wire  _T_22881 = bht_rd_addr_hashed_p1_f == 8'he1; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_225; // @[Reg.scala 27:20]
  wire [1:0] _T_23168 = _T_22881 ? bht_bank_rd_data_out_0_225 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23423 = _T_23422 | _T_23168; // @[Mux.scala 27:72]
  wire  _T_22883 = bht_rd_addr_hashed_p1_f == 8'he2; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_226; // @[Reg.scala 27:20]
  wire [1:0] _T_23169 = _T_22883 ? bht_bank_rd_data_out_0_226 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23424 = _T_23423 | _T_23169; // @[Mux.scala 27:72]
  wire  _T_22885 = bht_rd_addr_hashed_p1_f == 8'he3; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_227; // @[Reg.scala 27:20]
  wire [1:0] _T_23170 = _T_22885 ? bht_bank_rd_data_out_0_227 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23425 = _T_23424 | _T_23170; // @[Mux.scala 27:72]
  wire  _T_22887 = bht_rd_addr_hashed_p1_f == 8'he4; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_228; // @[Reg.scala 27:20]
  wire [1:0] _T_23171 = _T_22887 ? bht_bank_rd_data_out_0_228 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23426 = _T_23425 | _T_23171; // @[Mux.scala 27:72]
  wire  _T_22889 = bht_rd_addr_hashed_p1_f == 8'he5; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_229; // @[Reg.scala 27:20]
  wire [1:0] _T_23172 = _T_22889 ? bht_bank_rd_data_out_0_229 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23427 = _T_23426 | _T_23172; // @[Mux.scala 27:72]
  wire  _T_22891 = bht_rd_addr_hashed_p1_f == 8'he6; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_230; // @[Reg.scala 27:20]
  wire [1:0] _T_23173 = _T_22891 ? bht_bank_rd_data_out_0_230 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23428 = _T_23427 | _T_23173; // @[Mux.scala 27:72]
  wire  _T_22893 = bht_rd_addr_hashed_p1_f == 8'he7; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_231; // @[Reg.scala 27:20]
  wire [1:0] _T_23174 = _T_22893 ? bht_bank_rd_data_out_0_231 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23429 = _T_23428 | _T_23174; // @[Mux.scala 27:72]
  wire  _T_22895 = bht_rd_addr_hashed_p1_f == 8'he8; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_232; // @[Reg.scala 27:20]
  wire [1:0] _T_23175 = _T_22895 ? bht_bank_rd_data_out_0_232 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23430 = _T_23429 | _T_23175; // @[Mux.scala 27:72]
  wire  _T_22897 = bht_rd_addr_hashed_p1_f == 8'he9; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_233; // @[Reg.scala 27:20]
  wire [1:0] _T_23176 = _T_22897 ? bht_bank_rd_data_out_0_233 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23431 = _T_23430 | _T_23176; // @[Mux.scala 27:72]
  wire  _T_22899 = bht_rd_addr_hashed_p1_f == 8'hea; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_234; // @[Reg.scala 27:20]
  wire [1:0] _T_23177 = _T_22899 ? bht_bank_rd_data_out_0_234 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23432 = _T_23431 | _T_23177; // @[Mux.scala 27:72]
  wire  _T_22901 = bht_rd_addr_hashed_p1_f == 8'heb; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_235; // @[Reg.scala 27:20]
  wire [1:0] _T_23178 = _T_22901 ? bht_bank_rd_data_out_0_235 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23433 = _T_23432 | _T_23178; // @[Mux.scala 27:72]
  wire  _T_22903 = bht_rd_addr_hashed_p1_f == 8'hec; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_236; // @[Reg.scala 27:20]
  wire [1:0] _T_23179 = _T_22903 ? bht_bank_rd_data_out_0_236 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23434 = _T_23433 | _T_23179; // @[Mux.scala 27:72]
  wire  _T_22905 = bht_rd_addr_hashed_p1_f == 8'hed; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_237; // @[Reg.scala 27:20]
  wire [1:0] _T_23180 = _T_22905 ? bht_bank_rd_data_out_0_237 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23435 = _T_23434 | _T_23180; // @[Mux.scala 27:72]
  wire  _T_22907 = bht_rd_addr_hashed_p1_f == 8'hee; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_238; // @[Reg.scala 27:20]
  wire [1:0] _T_23181 = _T_22907 ? bht_bank_rd_data_out_0_238 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23436 = _T_23435 | _T_23181; // @[Mux.scala 27:72]
  wire  _T_22909 = bht_rd_addr_hashed_p1_f == 8'hef; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_239; // @[Reg.scala 27:20]
  wire [1:0] _T_23182 = _T_22909 ? bht_bank_rd_data_out_0_239 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23437 = _T_23436 | _T_23182; // @[Mux.scala 27:72]
  wire  _T_22911 = bht_rd_addr_hashed_p1_f == 8'hf0; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_240; // @[Reg.scala 27:20]
  wire [1:0] _T_23183 = _T_22911 ? bht_bank_rd_data_out_0_240 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23438 = _T_23437 | _T_23183; // @[Mux.scala 27:72]
  wire  _T_22913 = bht_rd_addr_hashed_p1_f == 8'hf1; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_241; // @[Reg.scala 27:20]
  wire [1:0] _T_23184 = _T_22913 ? bht_bank_rd_data_out_0_241 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23439 = _T_23438 | _T_23184; // @[Mux.scala 27:72]
  wire  _T_22915 = bht_rd_addr_hashed_p1_f == 8'hf2; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_242; // @[Reg.scala 27:20]
  wire [1:0] _T_23185 = _T_22915 ? bht_bank_rd_data_out_0_242 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23440 = _T_23439 | _T_23185; // @[Mux.scala 27:72]
  wire  _T_22917 = bht_rd_addr_hashed_p1_f == 8'hf3; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_243; // @[Reg.scala 27:20]
  wire [1:0] _T_23186 = _T_22917 ? bht_bank_rd_data_out_0_243 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23441 = _T_23440 | _T_23186; // @[Mux.scala 27:72]
  wire  _T_22919 = bht_rd_addr_hashed_p1_f == 8'hf4; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_244; // @[Reg.scala 27:20]
  wire [1:0] _T_23187 = _T_22919 ? bht_bank_rd_data_out_0_244 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23442 = _T_23441 | _T_23187; // @[Mux.scala 27:72]
  wire  _T_22921 = bht_rd_addr_hashed_p1_f == 8'hf5; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_245; // @[Reg.scala 27:20]
  wire [1:0] _T_23188 = _T_22921 ? bht_bank_rd_data_out_0_245 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23443 = _T_23442 | _T_23188; // @[Mux.scala 27:72]
  wire  _T_22923 = bht_rd_addr_hashed_p1_f == 8'hf6; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_246; // @[Reg.scala 27:20]
  wire [1:0] _T_23189 = _T_22923 ? bht_bank_rd_data_out_0_246 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23444 = _T_23443 | _T_23189; // @[Mux.scala 27:72]
  wire  _T_22925 = bht_rd_addr_hashed_p1_f == 8'hf7; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_247; // @[Reg.scala 27:20]
  wire [1:0] _T_23190 = _T_22925 ? bht_bank_rd_data_out_0_247 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23445 = _T_23444 | _T_23190; // @[Mux.scala 27:72]
  wire  _T_22927 = bht_rd_addr_hashed_p1_f == 8'hf8; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_248; // @[Reg.scala 27:20]
  wire [1:0] _T_23191 = _T_22927 ? bht_bank_rd_data_out_0_248 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23446 = _T_23445 | _T_23191; // @[Mux.scala 27:72]
  wire  _T_22929 = bht_rd_addr_hashed_p1_f == 8'hf9; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_249; // @[Reg.scala 27:20]
  wire [1:0] _T_23192 = _T_22929 ? bht_bank_rd_data_out_0_249 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23447 = _T_23446 | _T_23192; // @[Mux.scala 27:72]
  wire  _T_22931 = bht_rd_addr_hashed_p1_f == 8'hfa; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_250; // @[Reg.scala 27:20]
  wire [1:0] _T_23193 = _T_22931 ? bht_bank_rd_data_out_0_250 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23448 = _T_23447 | _T_23193; // @[Mux.scala 27:72]
  wire  _T_22933 = bht_rd_addr_hashed_p1_f == 8'hfb; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_251; // @[Reg.scala 27:20]
  wire [1:0] _T_23194 = _T_22933 ? bht_bank_rd_data_out_0_251 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23449 = _T_23448 | _T_23194; // @[Mux.scala 27:72]
  wire  _T_22935 = bht_rd_addr_hashed_p1_f == 8'hfc; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_252; // @[Reg.scala 27:20]
  wire [1:0] _T_23195 = _T_22935 ? bht_bank_rd_data_out_0_252 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23450 = _T_23449 | _T_23195; // @[Mux.scala 27:72]
  wire  _T_22937 = bht_rd_addr_hashed_p1_f == 8'hfd; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_253; // @[Reg.scala 27:20]
  wire [1:0] _T_23196 = _T_22937 ? bht_bank_rd_data_out_0_253 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23451 = _T_23450 | _T_23196; // @[Mux.scala 27:72]
  wire  _T_22939 = bht_rd_addr_hashed_p1_f == 8'hfe; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_254; // @[Reg.scala 27:20]
  wire [1:0] _T_23197 = _T_22939 ? bht_bank_rd_data_out_0_254 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23452 = _T_23451 | _T_23197; // @[Mux.scala 27:72]
  wire  _T_22941 = bht_rd_addr_hashed_p1_f == 8'hff; // @[el2_ifu_bp_ctl.scala 468:85]
  reg [1:0] bht_bank_rd_data_out_0_255; // @[Reg.scala 27:20]
  wire [1:0] _T_23198 = _T_22941 ? bht_bank_rd_data_out_0_255 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] bht_bank0_rd_data_p1_f = _T_23452 | _T_23198; // @[Mux.scala 27:72]
  wire [1:0] _T_260 = io_ifc_fetch_addr_f[0] ? bht_bank0_rd_data_p1_f : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] bht_vbank1_rd_data_f = _T_259 | _T_260; // @[Mux.scala 27:72]
  wire  _T_264 = bht_force_taken_f[1] | bht_vbank1_rd_data_f[1]; // @[el2_ifu_bp_ctl.scala 293:42]
  wire [1:0] wayhit_f = tag_match_way0_expanded_f | tag_match_way1_expanded_f; // @[el2_ifu_bp_ctl.scala 167:44]
  wire [1:0] _T_158 = _T_143 ? wayhit_f : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] wayhit_p1_f = tag_match_way0_expanded_p1_f | tag_match_way1_expanded_p1_f; // @[el2_ifu_bp_ctl.scala 169:50]
  wire [1:0] _T_157 = {wayhit_p1_f[0],wayhit_f[1]}; // @[Cat.scala 29:58]
  wire [1:0] _T_159 = io_ifc_fetch_addr_f[0] ? _T_157 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_160 = _T_158 | _T_159; // @[Mux.scala 27:72]
  wire  eoc_near = &io_ifc_fetch_addr_f[4:2]; // @[el2_ifu_bp_ctl.scala 253:64]
  wire  _T_218 = ~eoc_near; // @[el2_ifu_bp_ctl.scala 256:15]
  wire [1:0] _T_220 = ~io_ifc_fetch_addr_f[1:0]; // @[el2_ifu_bp_ctl.scala 256:28]
  wire  _T_221 = |_T_220; // @[el2_ifu_bp_ctl.scala 256:58]
  wire  eoc_mask = _T_218 | _T_221; // @[el2_ifu_bp_ctl.scala 256:25]
  wire [1:0] _T_162 = {eoc_mask,1'h1}; // @[Cat.scala 29:58]
  wire [1:0] vwayhit_f = _T_160 & _T_162; // @[el2_ifu_bp_ctl.scala 215:71]
  wire  _T_266 = _T_264 & vwayhit_f[1]; // @[el2_ifu_bp_ctl.scala 293:69]
  wire [1:0] _T_20895 = _T_21407 ? bht_bank_rd_data_out_0_0 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20896 = _T_21409 ? bht_bank_rd_data_out_0_1 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21151 = _T_20895 | _T_20896; // @[Mux.scala 27:72]
  wire [1:0] _T_20897 = _T_21411 ? bht_bank_rd_data_out_0_2 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21152 = _T_21151 | _T_20897; // @[Mux.scala 27:72]
  wire [1:0] _T_20898 = _T_21413 ? bht_bank_rd_data_out_0_3 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21153 = _T_21152 | _T_20898; // @[Mux.scala 27:72]
  wire [1:0] _T_20899 = _T_21415 ? bht_bank_rd_data_out_0_4 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21154 = _T_21153 | _T_20899; // @[Mux.scala 27:72]
  wire [1:0] _T_20900 = _T_21417 ? bht_bank_rd_data_out_0_5 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21155 = _T_21154 | _T_20900; // @[Mux.scala 27:72]
  wire [1:0] _T_20901 = _T_21419 ? bht_bank_rd_data_out_0_6 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21156 = _T_21155 | _T_20901; // @[Mux.scala 27:72]
  wire [1:0] _T_20902 = _T_21421 ? bht_bank_rd_data_out_0_7 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21157 = _T_21156 | _T_20902; // @[Mux.scala 27:72]
  wire [1:0] _T_20903 = _T_21423 ? bht_bank_rd_data_out_0_8 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21158 = _T_21157 | _T_20903; // @[Mux.scala 27:72]
  wire [1:0] _T_20904 = _T_21425 ? bht_bank_rd_data_out_0_9 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21159 = _T_21158 | _T_20904; // @[Mux.scala 27:72]
  wire [1:0] _T_20905 = _T_21427 ? bht_bank_rd_data_out_0_10 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21160 = _T_21159 | _T_20905; // @[Mux.scala 27:72]
  wire [1:0] _T_20906 = _T_21429 ? bht_bank_rd_data_out_0_11 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21161 = _T_21160 | _T_20906; // @[Mux.scala 27:72]
  wire [1:0] _T_20907 = _T_21431 ? bht_bank_rd_data_out_0_12 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21162 = _T_21161 | _T_20907; // @[Mux.scala 27:72]
  wire [1:0] _T_20908 = _T_21433 ? bht_bank_rd_data_out_0_13 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21163 = _T_21162 | _T_20908; // @[Mux.scala 27:72]
  wire [1:0] _T_20909 = _T_21435 ? bht_bank_rd_data_out_0_14 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21164 = _T_21163 | _T_20909; // @[Mux.scala 27:72]
  wire [1:0] _T_20910 = _T_21437 ? bht_bank_rd_data_out_0_15 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21165 = _T_21164 | _T_20910; // @[Mux.scala 27:72]
  wire [1:0] _T_20911 = _T_21439 ? bht_bank_rd_data_out_0_16 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21166 = _T_21165 | _T_20911; // @[Mux.scala 27:72]
  wire [1:0] _T_20912 = _T_21441 ? bht_bank_rd_data_out_0_17 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21167 = _T_21166 | _T_20912; // @[Mux.scala 27:72]
  wire [1:0] _T_20913 = _T_21443 ? bht_bank_rd_data_out_0_18 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21168 = _T_21167 | _T_20913; // @[Mux.scala 27:72]
  wire [1:0] _T_20914 = _T_21445 ? bht_bank_rd_data_out_0_19 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21169 = _T_21168 | _T_20914; // @[Mux.scala 27:72]
  wire [1:0] _T_20915 = _T_21447 ? bht_bank_rd_data_out_0_20 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21170 = _T_21169 | _T_20915; // @[Mux.scala 27:72]
  wire [1:0] _T_20916 = _T_21449 ? bht_bank_rd_data_out_0_21 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21171 = _T_21170 | _T_20916; // @[Mux.scala 27:72]
  wire [1:0] _T_20917 = _T_21451 ? bht_bank_rd_data_out_0_22 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21172 = _T_21171 | _T_20917; // @[Mux.scala 27:72]
  wire [1:0] _T_20918 = _T_21453 ? bht_bank_rd_data_out_0_23 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21173 = _T_21172 | _T_20918; // @[Mux.scala 27:72]
  wire [1:0] _T_20919 = _T_21455 ? bht_bank_rd_data_out_0_24 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21174 = _T_21173 | _T_20919; // @[Mux.scala 27:72]
  wire [1:0] _T_20920 = _T_21457 ? bht_bank_rd_data_out_0_25 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21175 = _T_21174 | _T_20920; // @[Mux.scala 27:72]
  wire [1:0] _T_20921 = _T_21459 ? bht_bank_rd_data_out_0_26 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21176 = _T_21175 | _T_20921; // @[Mux.scala 27:72]
  wire [1:0] _T_20922 = _T_21461 ? bht_bank_rd_data_out_0_27 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21177 = _T_21176 | _T_20922; // @[Mux.scala 27:72]
  wire [1:0] _T_20923 = _T_21463 ? bht_bank_rd_data_out_0_28 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21178 = _T_21177 | _T_20923; // @[Mux.scala 27:72]
  wire [1:0] _T_20924 = _T_21465 ? bht_bank_rd_data_out_0_29 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21179 = _T_21178 | _T_20924; // @[Mux.scala 27:72]
  wire [1:0] _T_20925 = _T_21467 ? bht_bank_rd_data_out_0_30 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21180 = _T_21179 | _T_20925; // @[Mux.scala 27:72]
  wire [1:0] _T_20926 = _T_21469 ? bht_bank_rd_data_out_0_31 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21181 = _T_21180 | _T_20926; // @[Mux.scala 27:72]
  wire [1:0] _T_20927 = _T_21471 ? bht_bank_rd_data_out_0_32 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21182 = _T_21181 | _T_20927; // @[Mux.scala 27:72]
  wire [1:0] _T_20928 = _T_21473 ? bht_bank_rd_data_out_0_33 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21183 = _T_21182 | _T_20928; // @[Mux.scala 27:72]
  wire [1:0] _T_20929 = _T_21475 ? bht_bank_rd_data_out_0_34 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21184 = _T_21183 | _T_20929; // @[Mux.scala 27:72]
  wire [1:0] _T_20930 = _T_21477 ? bht_bank_rd_data_out_0_35 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21185 = _T_21184 | _T_20930; // @[Mux.scala 27:72]
  wire [1:0] _T_20931 = _T_21479 ? bht_bank_rd_data_out_0_36 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21186 = _T_21185 | _T_20931; // @[Mux.scala 27:72]
  wire [1:0] _T_20932 = _T_21481 ? bht_bank_rd_data_out_0_37 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21187 = _T_21186 | _T_20932; // @[Mux.scala 27:72]
  wire [1:0] _T_20933 = _T_21483 ? bht_bank_rd_data_out_0_38 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21188 = _T_21187 | _T_20933; // @[Mux.scala 27:72]
  wire [1:0] _T_20934 = _T_21485 ? bht_bank_rd_data_out_0_39 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21189 = _T_21188 | _T_20934; // @[Mux.scala 27:72]
  wire [1:0] _T_20935 = _T_21487 ? bht_bank_rd_data_out_0_40 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21190 = _T_21189 | _T_20935; // @[Mux.scala 27:72]
  wire [1:0] _T_20936 = _T_21489 ? bht_bank_rd_data_out_0_41 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21191 = _T_21190 | _T_20936; // @[Mux.scala 27:72]
  wire [1:0] _T_20937 = _T_21491 ? bht_bank_rd_data_out_0_42 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21192 = _T_21191 | _T_20937; // @[Mux.scala 27:72]
  wire [1:0] _T_20938 = _T_21493 ? bht_bank_rd_data_out_0_43 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21193 = _T_21192 | _T_20938; // @[Mux.scala 27:72]
  wire [1:0] _T_20939 = _T_21495 ? bht_bank_rd_data_out_0_44 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21194 = _T_21193 | _T_20939; // @[Mux.scala 27:72]
  wire [1:0] _T_20940 = _T_21497 ? bht_bank_rd_data_out_0_45 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21195 = _T_21194 | _T_20940; // @[Mux.scala 27:72]
  wire [1:0] _T_20941 = _T_21499 ? bht_bank_rd_data_out_0_46 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21196 = _T_21195 | _T_20941; // @[Mux.scala 27:72]
  wire [1:0] _T_20942 = _T_21501 ? bht_bank_rd_data_out_0_47 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21197 = _T_21196 | _T_20942; // @[Mux.scala 27:72]
  wire [1:0] _T_20943 = _T_21503 ? bht_bank_rd_data_out_0_48 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21198 = _T_21197 | _T_20943; // @[Mux.scala 27:72]
  wire [1:0] _T_20944 = _T_21505 ? bht_bank_rd_data_out_0_49 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21199 = _T_21198 | _T_20944; // @[Mux.scala 27:72]
  wire [1:0] _T_20945 = _T_21507 ? bht_bank_rd_data_out_0_50 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21200 = _T_21199 | _T_20945; // @[Mux.scala 27:72]
  wire [1:0] _T_20946 = _T_21509 ? bht_bank_rd_data_out_0_51 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21201 = _T_21200 | _T_20946; // @[Mux.scala 27:72]
  wire [1:0] _T_20947 = _T_21511 ? bht_bank_rd_data_out_0_52 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21202 = _T_21201 | _T_20947; // @[Mux.scala 27:72]
  wire [1:0] _T_20948 = _T_21513 ? bht_bank_rd_data_out_0_53 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21203 = _T_21202 | _T_20948; // @[Mux.scala 27:72]
  wire [1:0] _T_20949 = _T_21515 ? bht_bank_rd_data_out_0_54 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21204 = _T_21203 | _T_20949; // @[Mux.scala 27:72]
  wire [1:0] _T_20950 = _T_21517 ? bht_bank_rd_data_out_0_55 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21205 = _T_21204 | _T_20950; // @[Mux.scala 27:72]
  wire [1:0] _T_20951 = _T_21519 ? bht_bank_rd_data_out_0_56 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21206 = _T_21205 | _T_20951; // @[Mux.scala 27:72]
  wire [1:0] _T_20952 = _T_21521 ? bht_bank_rd_data_out_0_57 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21207 = _T_21206 | _T_20952; // @[Mux.scala 27:72]
  wire [1:0] _T_20953 = _T_21523 ? bht_bank_rd_data_out_0_58 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21208 = _T_21207 | _T_20953; // @[Mux.scala 27:72]
  wire [1:0] _T_20954 = _T_21525 ? bht_bank_rd_data_out_0_59 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21209 = _T_21208 | _T_20954; // @[Mux.scala 27:72]
  wire [1:0] _T_20955 = _T_21527 ? bht_bank_rd_data_out_0_60 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21210 = _T_21209 | _T_20955; // @[Mux.scala 27:72]
  wire [1:0] _T_20956 = _T_21529 ? bht_bank_rd_data_out_0_61 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21211 = _T_21210 | _T_20956; // @[Mux.scala 27:72]
  wire [1:0] _T_20957 = _T_21531 ? bht_bank_rd_data_out_0_62 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21212 = _T_21211 | _T_20957; // @[Mux.scala 27:72]
  wire [1:0] _T_20958 = _T_21533 ? bht_bank_rd_data_out_0_63 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21213 = _T_21212 | _T_20958; // @[Mux.scala 27:72]
  wire [1:0] _T_20959 = _T_21535 ? bht_bank_rd_data_out_0_64 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21214 = _T_21213 | _T_20959; // @[Mux.scala 27:72]
  wire [1:0] _T_20960 = _T_21537 ? bht_bank_rd_data_out_0_65 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21215 = _T_21214 | _T_20960; // @[Mux.scala 27:72]
  wire [1:0] _T_20961 = _T_21539 ? bht_bank_rd_data_out_0_66 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21216 = _T_21215 | _T_20961; // @[Mux.scala 27:72]
  wire [1:0] _T_20962 = _T_21541 ? bht_bank_rd_data_out_0_67 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21217 = _T_21216 | _T_20962; // @[Mux.scala 27:72]
  wire [1:0] _T_20963 = _T_21543 ? bht_bank_rd_data_out_0_68 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21218 = _T_21217 | _T_20963; // @[Mux.scala 27:72]
  wire [1:0] _T_20964 = _T_21545 ? bht_bank_rd_data_out_0_69 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21219 = _T_21218 | _T_20964; // @[Mux.scala 27:72]
  wire [1:0] _T_20965 = _T_21547 ? bht_bank_rd_data_out_0_70 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21220 = _T_21219 | _T_20965; // @[Mux.scala 27:72]
  wire [1:0] _T_20966 = _T_21549 ? bht_bank_rd_data_out_0_71 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21221 = _T_21220 | _T_20966; // @[Mux.scala 27:72]
  wire [1:0] _T_20967 = _T_21551 ? bht_bank_rd_data_out_0_72 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21222 = _T_21221 | _T_20967; // @[Mux.scala 27:72]
  wire [1:0] _T_20968 = _T_21553 ? bht_bank_rd_data_out_0_73 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21223 = _T_21222 | _T_20968; // @[Mux.scala 27:72]
  wire [1:0] _T_20969 = _T_21555 ? bht_bank_rd_data_out_0_74 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21224 = _T_21223 | _T_20969; // @[Mux.scala 27:72]
  wire [1:0] _T_20970 = _T_21557 ? bht_bank_rd_data_out_0_75 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21225 = _T_21224 | _T_20970; // @[Mux.scala 27:72]
  wire [1:0] _T_20971 = _T_21559 ? bht_bank_rd_data_out_0_76 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21226 = _T_21225 | _T_20971; // @[Mux.scala 27:72]
  wire [1:0] _T_20972 = _T_21561 ? bht_bank_rd_data_out_0_77 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21227 = _T_21226 | _T_20972; // @[Mux.scala 27:72]
  wire [1:0] _T_20973 = _T_21563 ? bht_bank_rd_data_out_0_78 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21228 = _T_21227 | _T_20973; // @[Mux.scala 27:72]
  wire [1:0] _T_20974 = _T_21565 ? bht_bank_rd_data_out_0_79 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21229 = _T_21228 | _T_20974; // @[Mux.scala 27:72]
  wire [1:0] _T_20975 = _T_21567 ? bht_bank_rd_data_out_0_80 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21230 = _T_21229 | _T_20975; // @[Mux.scala 27:72]
  wire [1:0] _T_20976 = _T_21569 ? bht_bank_rd_data_out_0_81 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21231 = _T_21230 | _T_20976; // @[Mux.scala 27:72]
  wire [1:0] _T_20977 = _T_21571 ? bht_bank_rd_data_out_0_82 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21232 = _T_21231 | _T_20977; // @[Mux.scala 27:72]
  wire [1:0] _T_20978 = _T_21573 ? bht_bank_rd_data_out_0_83 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21233 = _T_21232 | _T_20978; // @[Mux.scala 27:72]
  wire [1:0] _T_20979 = _T_21575 ? bht_bank_rd_data_out_0_84 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21234 = _T_21233 | _T_20979; // @[Mux.scala 27:72]
  wire [1:0] _T_20980 = _T_21577 ? bht_bank_rd_data_out_0_85 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21235 = _T_21234 | _T_20980; // @[Mux.scala 27:72]
  wire [1:0] _T_20981 = _T_21579 ? bht_bank_rd_data_out_0_86 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21236 = _T_21235 | _T_20981; // @[Mux.scala 27:72]
  wire [1:0] _T_20982 = _T_21581 ? bht_bank_rd_data_out_0_87 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21237 = _T_21236 | _T_20982; // @[Mux.scala 27:72]
  wire [1:0] _T_20983 = _T_21583 ? bht_bank_rd_data_out_0_88 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21238 = _T_21237 | _T_20983; // @[Mux.scala 27:72]
  wire [1:0] _T_20984 = _T_21585 ? bht_bank_rd_data_out_0_89 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21239 = _T_21238 | _T_20984; // @[Mux.scala 27:72]
  wire [1:0] _T_20985 = _T_21587 ? bht_bank_rd_data_out_0_90 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21240 = _T_21239 | _T_20985; // @[Mux.scala 27:72]
  wire [1:0] _T_20986 = _T_21589 ? bht_bank_rd_data_out_0_91 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21241 = _T_21240 | _T_20986; // @[Mux.scala 27:72]
  wire [1:0] _T_20987 = _T_21591 ? bht_bank_rd_data_out_0_92 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21242 = _T_21241 | _T_20987; // @[Mux.scala 27:72]
  wire [1:0] _T_20988 = _T_21593 ? bht_bank_rd_data_out_0_93 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21243 = _T_21242 | _T_20988; // @[Mux.scala 27:72]
  wire [1:0] _T_20989 = _T_21595 ? bht_bank_rd_data_out_0_94 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21244 = _T_21243 | _T_20989; // @[Mux.scala 27:72]
  wire [1:0] _T_20990 = _T_21597 ? bht_bank_rd_data_out_0_95 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21245 = _T_21244 | _T_20990; // @[Mux.scala 27:72]
  wire [1:0] _T_20991 = _T_21599 ? bht_bank_rd_data_out_0_96 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21246 = _T_21245 | _T_20991; // @[Mux.scala 27:72]
  wire [1:0] _T_20992 = _T_21601 ? bht_bank_rd_data_out_0_97 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21247 = _T_21246 | _T_20992; // @[Mux.scala 27:72]
  wire [1:0] _T_20993 = _T_21603 ? bht_bank_rd_data_out_0_98 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21248 = _T_21247 | _T_20993; // @[Mux.scala 27:72]
  wire [1:0] _T_20994 = _T_21605 ? bht_bank_rd_data_out_0_99 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21249 = _T_21248 | _T_20994; // @[Mux.scala 27:72]
  wire [1:0] _T_20995 = _T_21607 ? bht_bank_rd_data_out_0_100 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21250 = _T_21249 | _T_20995; // @[Mux.scala 27:72]
  wire [1:0] _T_20996 = _T_21609 ? bht_bank_rd_data_out_0_101 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21251 = _T_21250 | _T_20996; // @[Mux.scala 27:72]
  wire [1:0] _T_20997 = _T_21611 ? bht_bank_rd_data_out_0_102 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21252 = _T_21251 | _T_20997; // @[Mux.scala 27:72]
  wire [1:0] _T_20998 = _T_21613 ? bht_bank_rd_data_out_0_103 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21253 = _T_21252 | _T_20998; // @[Mux.scala 27:72]
  wire [1:0] _T_20999 = _T_21615 ? bht_bank_rd_data_out_0_104 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21254 = _T_21253 | _T_20999; // @[Mux.scala 27:72]
  wire [1:0] _T_21000 = _T_21617 ? bht_bank_rd_data_out_0_105 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21255 = _T_21254 | _T_21000; // @[Mux.scala 27:72]
  wire [1:0] _T_21001 = _T_21619 ? bht_bank_rd_data_out_0_106 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21256 = _T_21255 | _T_21001; // @[Mux.scala 27:72]
  wire [1:0] _T_21002 = _T_21621 ? bht_bank_rd_data_out_0_107 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21257 = _T_21256 | _T_21002; // @[Mux.scala 27:72]
  wire [1:0] _T_21003 = _T_21623 ? bht_bank_rd_data_out_0_108 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21258 = _T_21257 | _T_21003; // @[Mux.scala 27:72]
  wire [1:0] _T_21004 = _T_21625 ? bht_bank_rd_data_out_0_109 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21259 = _T_21258 | _T_21004; // @[Mux.scala 27:72]
  wire [1:0] _T_21005 = _T_21627 ? bht_bank_rd_data_out_0_110 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21260 = _T_21259 | _T_21005; // @[Mux.scala 27:72]
  wire [1:0] _T_21006 = _T_21629 ? bht_bank_rd_data_out_0_111 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21261 = _T_21260 | _T_21006; // @[Mux.scala 27:72]
  wire [1:0] _T_21007 = _T_21631 ? bht_bank_rd_data_out_0_112 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21262 = _T_21261 | _T_21007; // @[Mux.scala 27:72]
  wire [1:0] _T_21008 = _T_21633 ? bht_bank_rd_data_out_0_113 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21263 = _T_21262 | _T_21008; // @[Mux.scala 27:72]
  wire [1:0] _T_21009 = _T_21635 ? bht_bank_rd_data_out_0_114 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21264 = _T_21263 | _T_21009; // @[Mux.scala 27:72]
  wire [1:0] _T_21010 = _T_21637 ? bht_bank_rd_data_out_0_115 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21265 = _T_21264 | _T_21010; // @[Mux.scala 27:72]
  wire [1:0] _T_21011 = _T_21639 ? bht_bank_rd_data_out_0_116 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21266 = _T_21265 | _T_21011; // @[Mux.scala 27:72]
  wire [1:0] _T_21012 = _T_21641 ? bht_bank_rd_data_out_0_117 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21267 = _T_21266 | _T_21012; // @[Mux.scala 27:72]
  wire [1:0] _T_21013 = _T_21643 ? bht_bank_rd_data_out_0_118 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21268 = _T_21267 | _T_21013; // @[Mux.scala 27:72]
  wire [1:0] _T_21014 = _T_21645 ? bht_bank_rd_data_out_0_119 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21269 = _T_21268 | _T_21014; // @[Mux.scala 27:72]
  wire [1:0] _T_21015 = _T_21647 ? bht_bank_rd_data_out_0_120 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21270 = _T_21269 | _T_21015; // @[Mux.scala 27:72]
  wire [1:0] _T_21016 = _T_21649 ? bht_bank_rd_data_out_0_121 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21271 = _T_21270 | _T_21016; // @[Mux.scala 27:72]
  wire [1:0] _T_21017 = _T_21651 ? bht_bank_rd_data_out_0_122 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21272 = _T_21271 | _T_21017; // @[Mux.scala 27:72]
  wire [1:0] _T_21018 = _T_21653 ? bht_bank_rd_data_out_0_123 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21273 = _T_21272 | _T_21018; // @[Mux.scala 27:72]
  wire [1:0] _T_21019 = _T_21655 ? bht_bank_rd_data_out_0_124 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21274 = _T_21273 | _T_21019; // @[Mux.scala 27:72]
  wire [1:0] _T_21020 = _T_21657 ? bht_bank_rd_data_out_0_125 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21275 = _T_21274 | _T_21020; // @[Mux.scala 27:72]
  wire [1:0] _T_21021 = _T_21659 ? bht_bank_rd_data_out_0_126 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21276 = _T_21275 | _T_21021; // @[Mux.scala 27:72]
  wire [1:0] _T_21022 = _T_21661 ? bht_bank_rd_data_out_0_127 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21277 = _T_21276 | _T_21022; // @[Mux.scala 27:72]
  wire [1:0] _T_21023 = _T_21663 ? bht_bank_rd_data_out_0_128 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21278 = _T_21277 | _T_21023; // @[Mux.scala 27:72]
  wire [1:0] _T_21024 = _T_21665 ? bht_bank_rd_data_out_0_129 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21279 = _T_21278 | _T_21024; // @[Mux.scala 27:72]
  wire [1:0] _T_21025 = _T_21667 ? bht_bank_rd_data_out_0_130 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21280 = _T_21279 | _T_21025; // @[Mux.scala 27:72]
  wire [1:0] _T_21026 = _T_21669 ? bht_bank_rd_data_out_0_131 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21281 = _T_21280 | _T_21026; // @[Mux.scala 27:72]
  wire [1:0] _T_21027 = _T_21671 ? bht_bank_rd_data_out_0_132 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21282 = _T_21281 | _T_21027; // @[Mux.scala 27:72]
  wire [1:0] _T_21028 = _T_21673 ? bht_bank_rd_data_out_0_133 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21283 = _T_21282 | _T_21028; // @[Mux.scala 27:72]
  wire [1:0] _T_21029 = _T_21675 ? bht_bank_rd_data_out_0_134 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21284 = _T_21283 | _T_21029; // @[Mux.scala 27:72]
  wire [1:0] _T_21030 = _T_21677 ? bht_bank_rd_data_out_0_135 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21285 = _T_21284 | _T_21030; // @[Mux.scala 27:72]
  wire [1:0] _T_21031 = _T_21679 ? bht_bank_rd_data_out_0_136 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21286 = _T_21285 | _T_21031; // @[Mux.scala 27:72]
  wire [1:0] _T_21032 = _T_21681 ? bht_bank_rd_data_out_0_137 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21287 = _T_21286 | _T_21032; // @[Mux.scala 27:72]
  wire [1:0] _T_21033 = _T_21683 ? bht_bank_rd_data_out_0_138 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21288 = _T_21287 | _T_21033; // @[Mux.scala 27:72]
  wire [1:0] _T_21034 = _T_21685 ? bht_bank_rd_data_out_0_139 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21289 = _T_21288 | _T_21034; // @[Mux.scala 27:72]
  wire [1:0] _T_21035 = _T_21687 ? bht_bank_rd_data_out_0_140 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21290 = _T_21289 | _T_21035; // @[Mux.scala 27:72]
  wire [1:0] _T_21036 = _T_21689 ? bht_bank_rd_data_out_0_141 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21291 = _T_21290 | _T_21036; // @[Mux.scala 27:72]
  wire [1:0] _T_21037 = _T_21691 ? bht_bank_rd_data_out_0_142 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21292 = _T_21291 | _T_21037; // @[Mux.scala 27:72]
  wire [1:0] _T_21038 = _T_21693 ? bht_bank_rd_data_out_0_143 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21293 = _T_21292 | _T_21038; // @[Mux.scala 27:72]
  wire [1:0] _T_21039 = _T_21695 ? bht_bank_rd_data_out_0_144 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21294 = _T_21293 | _T_21039; // @[Mux.scala 27:72]
  wire [1:0] _T_21040 = _T_21697 ? bht_bank_rd_data_out_0_145 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21295 = _T_21294 | _T_21040; // @[Mux.scala 27:72]
  wire [1:0] _T_21041 = _T_21699 ? bht_bank_rd_data_out_0_146 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21296 = _T_21295 | _T_21041; // @[Mux.scala 27:72]
  wire [1:0] _T_21042 = _T_21701 ? bht_bank_rd_data_out_0_147 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21297 = _T_21296 | _T_21042; // @[Mux.scala 27:72]
  wire [1:0] _T_21043 = _T_21703 ? bht_bank_rd_data_out_0_148 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21298 = _T_21297 | _T_21043; // @[Mux.scala 27:72]
  wire [1:0] _T_21044 = _T_21705 ? bht_bank_rd_data_out_0_149 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21299 = _T_21298 | _T_21044; // @[Mux.scala 27:72]
  wire [1:0] _T_21045 = _T_21707 ? bht_bank_rd_data_out_0_150 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21300 = _T_21299 | _T_21045; // @[Mux.scala 27:72]
  wire [1:0] _T_21046 = _T_21709 ? bht_bank_rd_data_out_0_151 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21301 = _T_21300 | _T_21046; // @[Mux.scala 27:72]
  wire [1:0] _T_21047 = _T_21711 ? bht_bank_rd_data_out_0_152 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21302 = _T_21301 | _T_21047; // @[Mux.scala 27:72]
  wire [1:0] _T_21048 = _T_21713 ? bht_bank_rd_data_out_0_153 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21303 = _T_21302 | _T_21048; // @[Mux.scala 27:72]
  wire [1:0] _T_21049 = _T_21715 ? bht_bank_rd_data_out_0_154 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21304 = _T_21303 | _T_21049; // @[Mux.scala 27:72]
  wire [1:0] _T_21050 = _T_21717 ? bht_bank_rd_data_out_0_155 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21305 = _T_21304 | _T_21050; // @[Mux.scala 27:72]
  wire [1:0] _T_21051 = _T_21719 ? bht_bank_rd_data_out_0_156 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21306 = _T_21305 | _T_21051; // @[Mux.scala 27:72]
  wire [1:0] _T_21052 = _T_21721 ? bht_bank_rd_data_out_0_157 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21307 = _T_21306 | _T_21052; // @[Mux.scala 27:72]
  wire [1:0] _T_21053 = _T_21723 ? bht_bank_rd_data_out_0_158 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21308 = _T_21307 | _T_21053; // @[Mux.scala 27:72]
  wire [1:0] _T_21054 = _T_21725 ? bht_bank_rd_data_out_0_159 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21309 = _T_21308 | _T_21054; // @[Mux.scala 27:72]
  wire [1:0] _T_21055 = _T_21727 ? bht_bank_rd_data_out_0_160 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21310 = _T_21309 | _T_21055; // @[Mux.scala 27:72]
  wire [1:0] _T_21056 = _T_21729 ? bht_bank_rd_data_out_0_161 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21311 = _T_21310 | _T_21056; // @[Mux.scala 27:72]
  wire [1:0] _T_21057 = _T_21731 ? bht_bank_rd_data_out_0_162 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21312 = _T_21311 | _T_21057; // @[Mux.scala 27:72]
  wire [1:0] _T_21058 = _T_21733 ? bht_bank_rd_data_out_0_163 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21313 = _T_21312 | _T_21058; // @[Mux.scala 27:72]
  wire [1:0] _T_21059 = _T_21735 ? bht_bank_rd_data_out_0_164 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21314 = _T_21313 | _T_21059; // @[Mux.scala 27:72]
  wire [1:0] _T_21060 = _T_21737 ? bht_bank_rd_data_out_0_165 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21315 = _T_21314 | _T_21060; // @[Mux.scala 27:72]
  wire [1:0] _T_21061 = _T_21739 ? bht_bank_rd_data_out_0_166 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21316 = _T_21315 | _T_21061; // @[Mux.scala 27:72]
  wire [1:0] _T_21062 = _T_21741 ? bht_bank_rd_data_out_0_167 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21317 = _T_21316 | _T_21062; // @[Mux.scala 27:72]
  wire [1:0] _T_21063 = _T_21743 ? bht_bank_rd_data_out_0_168 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21318 = _T_21317 | _T_21063; // @[Mux.scala 27:72]
  wire [1:0] _T_21064 = _T_21745 ? bht_bank_rd_data_out_0_169 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21319 = _T_21318 | _T_21064; // @[Mux.scala 27:72]
  wire [1:0] _T_21065 = _T_21747 ? bht_bank_rd_data_out_0_170 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21320 = _T_21319 | _T_21065; // @[Mux.scala 27:72]
  wire [1:0] _T_21066 = _T_21749 ? bht_bank_rd_data_out_0_171 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21321 = _T_21320 | _T_21066; // @[Mux.scala 27:72]
  wire [1:0] _T_21067 = _T_21751 ? bht_bank_rd_data_out_0_172 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21322 = _T_21321 | _T_21067; // @[Mux.scala 27:72]
  wire [1:0] _T_21068 = _T_21753 ? bht_bank_rd_data_out_0_173 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21323 = _T_21322 | _T_21068; // @[Mux.scala 27:72]
  wire [1:0] _T_21069 = _T_21755 ? bht_bank_rd_data_out_0_174 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21324 = _T_21323 | _T_21069; // @[Mux.scala 27:72]
  wire [1:0] _T_21070 = _T_21757 ? bht_bank_rd_data_out_0_175 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21325 = _T_21324 | _T_21070; // @[Mux.scala 27:72]
  wire [1:0] _T_21071 = _T_21759 ? bht_bank_rd_data_out_0_176 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21326 = _T_21325 | _T_21071; // @[Mux.scala 27:72]
  wire [1:0] _T_21072 = _T_21761 ? bht_bank_rd_data_out_0_177 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21327 = _T_21326 | _T_21072; // @[Mux.scala 27:72]
  wire [1:0] _T_21073 = _T_21763 ? bht_bank_rd_data_out_0_178 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21328 = _T_21327 | _T_21073; // @[Mux.scala 27:72]
  wire [1:0] _T_21074 = _T_21765 ? bht_bank_rd_data_out_0_179 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21329 = _T_21328 | _T_21074; // @[Mux.scala 27:72]
  wire [1:0] _T_21075 = _T_21767 ? bht_bank_rd_data_out_0_180 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21330 = _T_21329 | _T_21075; // @[Mux.scala 27:72]
  wire [1:0] _T_21076 = _T_21769 ? bht_bank_rd_data_out_0_181 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21331 = _T_21330 | _T_21076; // @[Mux.scala 27:72]
  wire [1:0] _T_21077 = _T_21771 ? bht_bank_rd_data_out_0_182 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21332 = _T_21331 | _T_21077; // @[Mux.scala 27:72]
  wire [1:0] _T_21078 = _T_21773 ? bht_bank_rd_data_out_0_183 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21333 = _T_21332 | _T_21078; // @[Mux.scala 27:72]
  wire [1:0] _T_21079 = _T_21775 ? bht_bank_rd_data_out_0_184 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21334 = _T_21333 | _T_21079; // @[Mux.scala 27:72]
  wire [1:0] _T_21080 = _T_21777 ? bht_bank_rd_data_out_0_185 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21335 = _T_21334 | _T_21080; // @[Mux.scala 27:72]
  wire [1:0] _T_21081 = _T_21779 ? bht_bank_rd_data_out_0_186 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21336 = _T_21335 | _T_21081; // @[Mux.scala 27:72]
  wire [1:0] _T_21082 = _T_21781 ? bht_bank_rd_data_out_0_187 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21337 = _T_21336 | _T_21082; // @[Mux.scala 27:72]
  wire [1:0] _T_21083 = _T_21783 ? bht_bank_rd_data_out_0_188 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21338 = _T_21337 | _T_21083; // @[Mux.scala 27:72]
  wire [1:0] _T_21084 = _T_21785 ? bht_bank_rd_data_out_0_189 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21339 = _T_21338 | _T_21084; // @[Mux.scala 27:72]
  wire [1:0] _T_21085 = _T_21787 ? bht_bank_rd_data_out_0_190 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21340 = _T_21339 | _T_21085; // @[Mux.scala 27:72]
  wire [1:0] _T_21086 = _T_21789 ? bht_bank_rd_data_out_0_191 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21341 = _T_21340 | _T_21086; // @[Mux.scala 27:72]
  wire [1:0] _T_21087 = _T_21791 ? bht_bank_rd_data_out_0_192 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21342 = _T_21341 | _T_21087; // @[Mux.scala 27:72]
  wire [1:0] _T_21088 = _T_21793 ? bht_bank_rd_data_out_0_193 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21343 = _T_21342 | _T_21088; // @[Mux.scala 27:72]
  wire [1:0] _T_21089 = _T_21795 ? bht_bank_rd_data_out_0_194 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21344 = _T_21343 | _T_21089; // @[Mux.scala 27:72]
  wire [1:0] _T_21090 = _T_21797 ? bht_bank_rd_data_out_0_195 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21345 = _T_21344 | _T_21090; // @[Mux.scala 27:72]
  wire [1:0] _T_21091 = _T_21799 ? bht_bank_rd_data_out_0_196 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21346 = _T_21345 | _T_21091; // @[Mux.scala 27:72]
  wire [1:0] _T_21092 = _T_21801 ? bht_bank_rd_data_out_0_197 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21347 = _T_21346 | _T_21092; // @[Mux.scala 27:72]
  wire [1:0] _T_21093 = _T_21803 ? bht_bank_rd_data_out_0_198 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21348 = _T_21347 | _T_21093; // @[Mux.scala 27:72]
  wire [1:0] _T_21094 = _T_21805 ? bht_bank_rd_data_out_0_199 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21349 = _T_21348 | _T_21094; // @[Mux.scala 27:72]
  wire [1:0] _T_21095 = _T_21807 ? bht_bank_rd_data_out_0_200 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21350 = _T_21349 | _T_21095; // @[Mux.scala 27:72]
  wire [1:0] _T_21096 = _T_21809 ? bht_bank_rd_data_out_0_201 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21351 = _T_21350 | _T_21096; // @[Mux.scala 27:72]
  wire [1:0] _T_21097 = _T_21811 ? bht_bank_rd_data_out_0_202 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21352 = _T_21351 | _T_21097; // @[Mux.scala 27:72]
  wire [1:0] _T_21098 = _T_21813 ? bht_bank_rd_data_out_0_203 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21353 = _T_21352 | _T_21098; // @[Mux.scala 27:72]
  wire [1:0] _T_21099 = _T_21815 ? bht_bank_rd_data_out_0_204 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21354 = _T_21353 | _T_21099; // @[Mux.scala 27:72]
  wire [1:0] _T_21100 = _T_21817 ? bht_bank_rd_data_out_0_205 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21355 = _T_21354 | _T_21100; // @[Mux.scala 27:72]
  wire [1:0] _T_21101 = _T_21819 ? bht_bank_rd_data_out_0_206 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21356 = _T_21355 | _T_21101; // @[Mux.scala 27:72]
  wire [1:0] _T_21102 = _T_21821 ? bht_bank_rd_data_out_0_207 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21357 = _T_21356 | _T_21102; // @[Mux.scala 27:72]
  wire [1:0] _T_21103 = _T_21823 ? bht_bank_rd_data_out_0_208 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21358 = _T_21357 | _T_21103; // @[Mux.scala 27:72]
  wire [1:0] _T_21104 = _T_21825 ? bht_bank_rd_data_out_0_209 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21359 = _T_21358 | _T_21104; // @[Mux.scala 27:72]
  wire [1:0] _T_21105 = _T_21827 ? bht_bank_rd_data_out_0_210 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21360 = _T_21359 | _T_21105; // @[Mux.scala 27:72]
  wire [1:0] _T_21106 = _T_21829 ? bht_bank_rd_data_out_0_211 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21361 = _T_21360 | _T_21106; // @[Mux.scala 27:72]
  wire [1:0] _T_21107 = _T_21831 ? bht_bank_rd_data_out_0_212 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21362 = _T_21361 | _T_21107; // @[Mux.scala 27:72]
  wire [1:0] _T_21108 = _T_21833 ? bht_bank_rd_data_out_0_213 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21363 = _T_21362 | _T_21108; // @[Mux.scala 27:72]
  wire [1:0] _T_21109 = _T_21835 ? bht_bank_rd_data_out_0_214 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21364 = _T_21363 | _T_21109; // @[Mux.scala 27:72]
  wire [1:0] _T_21110 = _T_21837 ? bht_bank_rd_data_out_0_215 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21365 = _T_21364 | _T_21110; // @[Mux.scala 27:72]
  wire [1:0] _T_21111 = _T_21839 ? bht_bank_rd_data_out_0_216 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21366 = _T_21365 | _T_21111; // @[Mux.scala 27:72]
  wire [1:0] _T_21112 = _T_21841 ? bht_bank_rd_data_out_0_217 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21367 = _T_21366 | _T_21112; // @[Mux.scala 27:72]
  wire [1:0] _T_21113 = _T_21843 ? bht_bank_rd_data_out_0_218 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21368 = _T_21367 | _T_21113; // @[Mux.scala 27:72]
  wire [1:0] _T_21114 = _T_21845 ? bht_bank_rd_data_out_0_219 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21369 = _T_21368 | _T_21114; // @[Mux.scala 27:72]
  wire [1:0] _T_21115 = _T_21847 ? bht_bank_rd_data_out_0_220 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21370 = _T_21369 | _T_21115; // @[Mux.scala 27:72]
  wire [1:0] _T_21116 = _T_21849 ? bht_bank_rd_data_out_0_221 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21371 = _T_21370 | _T_21116; // @[Mux.scala 27:72]
  wire [1:0] _T_21117 = _T_21851 ? bht_bank_rd_data_out_0_222 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21372 = _T_21371 | _T_21117; // @[Mux.scala 27:72]
  wire [1:0] _T_21118 = _T_21853 ? bht_bank_rd_data_out_0_223 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21373 = _T_21372 | _T_21118; // @[Mux.scala 27:72]
  wire [1:0] _T_21119 = _T_21855 ? bht_bank_rd_data_out_0_224 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21374 = _T_21373 | _T_21119; // @[Mux.scala 27:72]
  wire [1:0] _T_21120 = _T_21857 ? bht_bank_rd_data_out_0_225 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21375 = _T_21374 | _T_21120; // @[Mux.scala 27:72]
  wire [1:0] _T_21121 = _T_21859 ? bht_bank_rd_data_out_0_226 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21376 = _T_21375 | _T_21121; // @[Mux.scala 27:72]
  wire [1:0] _T_21122 = _T_21861 ? bht_bank_rd_data_out_0_227 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21377 = _T_21376 | _T_21122; // @[Mux.scala 27:72]
  wire [1:0] _T_21123 = _T_21863 ? bht_bank_rd_data_out_0_228 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21378 = _T_21377 | _T_21123; // @[Mux.scala 27:72]
  wire [1:0] _T_21124 = _T_21865 ? bht_bank_rd_data_out_0_229 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21379 = _T_21378 | _T_21124; // @[Mux.scala 27:72]
  wire [1:0] _T_21125 = _T_21867 ? bht_bank_rd_data_out_0_230 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21380 = _T_21379 | _T_21125; // @[Mux.scala 27:72]
  wire [1:0] _T_21126 = _T_21869 ? bht_bank_rd_data_out_0_231 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21381 = _T_21380 | _T_21126; // @[Mux.scala 27:72]
  wire [1:0] _T_21127 = _T_21871 ? bht_bank_rd_data_out_0_232 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21382 = _T_21381 | _T_21127; // @[Mux.scala 27:72]
  wire [1:0] _T_21128 = _T_21873 ? bht_bank_rd_data_out_0_233 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21383 = _T_21382 | _T_21128; // @[Mux.scala 27:72]
  wire [1:0] _T_21129 = _T_21875 ? bht_bank_rd_data_out_0_234 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21384 = _T_21383 | _T_21129; // @[Mux.scala 27:72]
  wire [1:0] _T_21130 = _T_21877 ? bht_bank_rd_data_out_0_235 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21385 = _T_21384 | _T_21130; // @[Mux.scala 27:72]
  wire [1:0] _T_21131 = _T_21879 ? bht_bank_rd_data_out_0_236 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21386 = _T_21385 | _T_21131; // @[Mux.scala 27:72]
  wire [1:0] _T_21132 = _T_21881 ? bht_bank_rd_data_out_0_237 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21387 = _T_21386 | _T_21132; // @[Mux.scala 27:72]
  wire [1:0] _T_21133 = _T_21883 ? bht_bank_rd_data_out_0_238 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21388 = _T_21387 | _T_21133; // @[Mux.scala 27:72]
  wire [1:0] _T_21134 = _T_21885 ? bht_bank_rd_data_out_0_239 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21389 = _T_21388 | _T_21134; // @[Mux.scala 27:72]
  wire [1:0] _T_21135 = _T_21887 ? bht_bank_rd_data_out_0_240 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21390 = _T_21389 | _T_21135; // @[Mux.scala 27:72]
  wire [1:0] _T_21136 = _T_21889 ? bht_bank_rd_data_out_0_241 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21391 = _T_21390 | _T_21136; // @[Mux.scala 27:72]
  wire [1:0] _T_21137 = _T_21891 ? bht_bank_rd_data_out_0_242 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21392 = _T_21391 | _T_21137; // @[Mux.scala 27:72]
  wire [1:0] _T_21138 = _T_21893 ? bht_bank_rd_data_out_0_243 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21393 = _T_21392 | _T_21138; // @[Mux.scala 27:72]
  wire [1:0] _T_21139 = _T_21895 ? bht_bank_rd_data_out_0_244 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21394 = _T_21393 | _T_21139; // @[Mux.scala 27:72]
  wire [1:0] _T_21140 = _T_21897 ? bht_bank_rd_data_out_0_245 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21395 = _T_21394 | _T_21140; // @[Mux.scala 27:72]
  wire [1:0] _T_21141 = _T_21899 ? bht_bank_rd_data_out_0_246 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21396 = _T_21395 | _T_21141; // @[Mux.scala 27:72]
  wire [1:0] _T_21142 = _T_21901 ? bht_bank_rd_data_out_0_247 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21397 = _T_21396 | _T_21142; // @[Mux.scala 27:72]
  wire [1:0] _T_21143 = _T_21903 ? bht_bank_rd_data_out_0_248 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21398 = _T_21397 | _T_21143; // @[Mux.scala 27:72]
  wire [1:0] _T_21144 = _T_21905 ? bht_bank_rd_data_out_0_249 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21399 = _T_21398 | _T_21144; // @[Mux.scala 27:72]
  wire [1:0] _T_21145 = _T_21907 ? bht_bank_rd_data_out_0_250 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21400 = _T_21399 | _T_21145; // @[Mux.scala 27:72]
  wire [1:0] _T_21146 = _T_21909 ? bht_bank_rd_data_out_0_251 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21401 = _T_21400 | _T_21146; // @[Mux.scala 27:72]
  wire [1:0] _T_21147 = _T_21911 ? bht_bank_rd_data_out_0_252 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21402 = _T_21401 | _T_21147; // @[Mux.scala 27:72]
  wire [1:0] _T_21148 = _T_21913 ? bht_bank_rd_data_out_0_253 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21403 = _T_21402 | _T_21148; // @[Mux.scala 27:72]
  wire [1:0] _T_21149 = _T_21915 ? bht_bank_rd_data_out_0_254 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21404 = _T_21403 | _T_21149; // @[Mux.scala 27:72]
  wire [1:0] _T_21150 = _T_21917 ? bht_bank_rd_data_out_0_255 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] bht_bank0_rd_data_f = _T_21404 | _T_21150; // @[Mux.scala 27:72]
  wire [1:0] _T_251 = _T_143 ? bht_bank0_rd_data_f : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_252 = io_ifc_fetch_addr_f[0] ? bht_bank1_rd_data_f : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] bht_vbank0_rd_data_f = _T_251 | _T_252; // @[Mux.scala 27:72]
  wire  _T_269 = bht_force_taken_f[0] | bht_vbank0_rd_data_f[1]; // @[el2_ifu_bp_ctl.scala 294:45]
  wire  _T_271 = _T_269 & vwayhit_f[0]; // @[el2_ifu_bp_ctl.scala 294:72]
  wire [1:0] bht_dir_f = {_T_266,_T_271}; // @[Cat.scala 29:58]
  wire  _T_14 = ~bht_dir_f[0]; // @[el2_ifu_bp_ctl.scala 108:23]
  wire [1:0] btb_sel_f = {_T_14,bht_dir_f[0]}; // @[Cat.scala 29:58]
  wire [1:0] fetch_start_f = {io_ifc_fetch_addr_f[0],_T_143}; // @[Cat.scala 29:58]
  wire  _T_32 = io_exu_mp_btag == fetch_rd_tag_f; // @[el2_ifu_bp_ctl.scala 126:46]
  wire  _T_33 = _T_32 & exu_mp_valid; // @[el2_ifu_bp_ctl.scala 126:66]
  wire  _T_34 = _T_33 & io_ifc_fetch_req_f; // @[el2_ifu_bp_ctl.scala 126:81]
  wire  _T_35 = io_exu_mp_index == btb_rd_addr_f; // @[el2_ifu_bp_ctl.scala 126:117]
  wire  fetch_mp_collision_f = _T_34 & _T_35; // @[el2_ifu_bp_ctl.scala 126:102]
  wire  _T_36 = io_exu_mp_btag == fetch_rd_tag_p1_f; // @[el2_ifu_bp_ctl.scala 127:49]
  wire  _T_37 = _T_36 & exu_mp_valid; // @[el2_ifu_bp_ctl.scala 127:72]
  wire  _T_38 = _T_37 & io_ifc_fetch_req_f; // @[el2_ifu_bp_ctl.scala 127:87]
  wire  _T_39 = io_exu_mp_index == btb_rd_addr_p1_f; // @[el2_ifu_bp_ctl.scala 127:123]
  wire  fetch_mp_collision_p1_f = _T_38 & _T_39; // @[el2_ifu_bp_ctl.scala 127:108]
  reg  exu_mp_way_f; // @[el2_ifu_bp_ctl.scala 131:55]
  reg  exu_flush_final_d1; // @[el2_ifu_bp_ctl.scala 132:61]
  wire [255:0] mp_wrindex_dec = 256'h1 << io_exu_mp_index; // @[el2_ifu_bp_ctl.scala 203:28]
  wire [255:0] fetch_wrindex_dec = 256'h1 << btb_rd_addr_f; // @[el2_ifu_bp_ctl.scala 206:31]
  wire [255:0] fetch_wrindex_p1_dec = 256'h1 << btb_rd_addr_p1_f; // @[el2_ifu_bp_ctl.scala 209:34]
  wire [255:0] _T_149 = exu_mp_valid ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12]
  wire [255:0] mp_wrlru_b0 = mp_wrindex_dec & _T_149; // @[el2_ifu_bp_ctl.scala 212:36]
  wire  _T_165 = vwayhit_f[0] | vwayhit_f[1]; // @[el2_ifu_bp_ctl.scala 218:42]
  wire  _T_166 = _T_165 & io_ifc_fetch_req_f; // @[el2_ifu_bp_ctl.scala 218:58]
  wire  lru_update_valid_f = _T_166 & _T; // @[el2_ifu_bp_ctl.scala 218:79]
  wire [255:0] _T_169 = lru_update_valid_f ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12]
  wire [255:0] fetch_wrlru_b0 = fetch_wrindex_dec & _T_169; // @[el2_ifu_bp_ctl.scala 220:42]
  wire [255:0] fetch_wrlru_p1_b0 = fetch_wrindex_p1_dec & _T_169; // @[el2_ifu_bp_ctl.scala 221:48]
  wire [255:0] _T_172 = ~mp_wrlru_b0; // @[el2_ifu_bp_ctl.scala 223:25]
  wire [255:0] _T_173 = ~fetch_wrlru_b0; // @[el2_ifu_bp_ctl.scala 223:40]
  wire [255:0] btb_lru_b0_hold = _T_172 & _T_173; // @[el2_ifu_bp_ctl.scala 223:38]
  wire  _T_175 = ~io_exu_mp_pkt_way; // @[el2_ifu_bp_ctl.scala 230:40]
  wire [255:0] _T_178 = _T_175 ? mp_wrlru_b0 : 256'h0; // @[Mux.scala 27:72]
  wire [255:0] _T_179 = tag_match_way0_f ? fetch_wrlru_b0 : 256'h0; // @[Mux.scala 27:72]
  wire [255:0] _T_180 = tag_match_way0_p1_f ? fetch_wrlru_p1_b0 : 256'h0; // @[Mux.scala 27:72]
  wire [255:0] _T_181 = _T_178 | _T_179; // @[Mux.scala 27:72]
  wire [255:0] _T_182 = _T_181 | _T_180; // @[Mux.scala 27:72]
  reg [255:0] btb_lru_b0_f; // @[el2_lib.scala 481:16]
  wire [255:0] _T_184 = btb_lru_b0_hold & btb_lru_b0_f; // @[el2_ifu_bp_ctl.scala 232:102]
  wire [255:0] _T_186 = fetch_wrindex_dec & btb_lru_b0_f; // @[el2_ifu_bp_ctl.scala 235:78]
  wire  _T_187 = |_T_186; // @[el2_ifu_bp_ctl.scala 235:94]
  wire  btb_lru_rd_f = fetch_mp_collision_f ? exu_mp_way_f : _T_187; // @[el2_ifu_bp_ctl.scala 235:25]
  wire [255:0] _T_189 = fetch_wrindex_p1_dec & btb_lru_b0_f; // @[el2_ifu_bp_ctl.scala 237:87]
  wire  _T_190 = |_T_189; // @[el2_ifu_bp_ctl.scala 237:103]
  wire  btb_lru_rd_p1_f = fetch_mp_collision_p1_f ? exu_mp_way_f : _T_190; // @[el2_ifu_bp_ctl.scala 237:28]
  wire [1:0] _T_193 = {btb_lru_rd_f,btb_lru_rd_f}; // @[Cat.scala 29:58]
  wire [1:0] _T_196 = {btb_lru_rd_p1_f,btb_lru_rd_f}; // @[Cat.scala 29:58]
  wire [1:0] _T_197 = _T_143 ? _T_193 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_198 = io_ifc_fetch_addr_f[0] ? _T_196 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] btb_vlru_rd_f = _T_197 | _T_198; // @[Mux.scala 27:72]
  wire [1:0] _T_207 = {tag_match_way1_expanded_p1_f[0],tag_match_way1_expanded_f[1]}; // @[Cat.scala 29:58]
  wire [1:0] _T_208 = _T_143 ? tag_match_way1_expanded_f : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_209 = io_ifc_fetch_addr_f[0] ? _T_207 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] tag_match_vway1_expanded_f = _T_208 | _T_209; // @[Mux.scala 27:72]
  wire [1:0] _T_211 = ~vwayhit_f; // @[el2_ifu_bp_ctl.scala 247:52]
  wire [1:0] _T_212 = _T_211 & btb_vlru_rd_f; // @[el2_ifu_bp_ctl.scala 247:63]
  wire [15:0] _T_229 = btb_sel_f[1] ? btb_vbank1_rd_data_f[16:1] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_230 = btb_sel_f[0] ? btb_vbank0_rd_data_f[16:1] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] btb_sel_data_f = _T_229 | _T_230; // @[Mux.scala 27:72]
  wire [11:0] btb_rd_tgt_f = btb_sel_data_f[15:4]; // @[el2_ifu_bp_ctl.scala 263:36]
  wire  btb_rd_pc4_f = btb_sel_data_f[3]; // @[el2_ifu_bp_ctl.scala 264:36]
  wire  btb_rd_call_f = btb_sel_data_f[1]; // @[el2_ifu_bp_ctl.scala 265:37]
  wire  btb_rd_ret_f = btb_sel_data_f[0]; // @[el2_ifu_bp_ctl.scala 266:36]
  wire [1:0] _T_279 = {bht_vbank1_rd_data_f[1],bht_vbank0_rd_data_f[1]}; // @[Cat.scala 29:58]
  wire [1:0] hist1_raw = bht_force_taken_f | _T_279; // @[el2_ifu_bp_ctl.scala 300:34]
  wire [1:0] _T_233 = vwayhit_f & hist1_raw; // @[el2_ifu_bp_ctl.scala 273:39]
  wire  _T_234 = |_T_233; // @[el2_ifu_bp_ctl.scala 273:52]
  wire  _T_235 = _T_234 & io_ifc_fetch_req_f; // @[el2_ifu_bp_ctl.scala 273:56]
  wire  _T_236 = ~leak_one_f_d1; // @[el2_ifu_bp_ctl.scala 273:79]
  wire  _T_237 = _T_235 & _T_236; // @[el2_ifu_bp_ctl.scala 273:77]
  wire  _T_238 = ~io_dec_tlu_bpred_disable; // @[el2_ifu_bp_ctl.scala 273:96]
  wire  _T_274 = io_ifu_bp_hit_taken_f & btb_sel_f[1]; // @[el2_ifu_bp_ctl.scala 297:51]
  wire  _T_275 = ~io_ifu_bp_hit_taken_f; // @[el2_ifu_bp_ctl.scala 297:69]
  wire  _T_285 = vwayhit_f[1] & btb_vbank1_rd_data_f[4]; // @[el2_ifu_bp_ctl.scala 306:34]
  wire  _T_288 = vwayhit_f[0] & btb_vbank0_rd_data_f[4]; // @[el2_ifu_bp_ctl.scala 307:34]
  wire  _T_291 = ~btb_vbank1_rd_data_f[2]; // @[el2_ifu_bp_ctl.scala 310:37]
  wire  _T_292 = vwayhit_f[1] & _T_291; // @[el2_ifu_bp_ctl.scala 310:35]
  wire  _T_294 = _T_292 & btb_vbank1_rd_data_f[1]; // @[el2_ifu_bp_ctl.scala 310:65]
  wire  _T_297 = ~btb_vbank0_rd_data_f[2]; // @[el2_ifu_bp_ctl.scala 311:37]
  wire  _T_298 = vwayhit_f[0] & _T_297; // @[el2_ifu_bp_ctl.scala 311:35]
  wire  _T_300 = _T_298 & btb_vbank0_rd_data_f[1]; // @[el2_ifu_bp_ctl.scala 311:65]
  wire [1:0] num_valids = vwayhit_f[1] + vwayhit_f[0]; // @[el2_ifu_bp_ctl.scala 314:35]
  wire [1:0] _T_303 = btb_sel_f & bht_dir_f; // @[el2_ifu_bp_ctl.scala 317:28]
  wire  final_h = |_T_303; // @[el2_ifu_bp_ctl.scala 317:41]
  wire  _T_304 = num_valids == 2'h2; // @[el2_ifu_bp_ctl.scala 321:41]
  wire [7:0] _T_308 = {fghr[5:0],1'h0,final_h}; // @[Cat.scala 29:58]
  wire  _T_309 = num_valids == 2'h1; // @[el2_ifu_bp_ctl.scala 322:41]
  wire [7:0] _T_312 = {fghr[6:0],final_h}; // @[Cat.scala 29:58]
  wire  _T_313 = num_valids == 2'h0; // @[el2_ifu_bp_ctl.scala 323:41]
  wire [7:0] _T_316 = _T_304 ? _T_308 : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_317 = _T_309 ? _T_312 : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_318 = _T_313 ? fghr : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_319 = _T_316 | _T_317; // @[Mux.scala 27:72]
  wire [7:0] merged_ghr = _T_319 | _T_318; // @[Mux.scala 27:72]
  wire  _T_322 = ~exu_flush_final_d1; // @[el2_ifu_bp_ctl.scala 332:27]
  wire  _T_323 = _T_322 & io_ifc_fetch_req_f; // @[el2_ifu_bp_ctl.scala 332:47]
  wire  _T_324 = _T_323 & io_ic_hit_f; // @[el2_ifu_bp_ctl.scala 332:70]
  wire  _T_326 = _T_324 & _T_236; // @[el2_ifu_bp_ctl.scala 332:84]
  wire  _T_329 = io_ifc_fetch_req_f & io_ic_hit_f; // @[el2_ifu_bp_ctl.scala 333:70]
  wire  _T_331 = _T_329 & _T_236; // @[el2_ifu_bp_ctl.scala 333:84]
  wire  _T_332 = ~_T_331; // @[el2_ifu_bp_ctl.scala 333:49]
  wire  _T_333 = _T_322 & _T_332; // @[el2_ifu_bp_ctl.scala 333:47]
  wire [7:0] _T_335 = exu_flush_final_d1 ? io_exu_mp_fghr : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_336 = _T_326 ? merged_ghr : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_337 = _T_333 ? fghr : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_338 = _T_335 | _T_336; // @[Mux.scala 27:72]
  wire [1:0] _T_343 = io_dec_tlu_bpred_disable ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [1:0] _T_344 = ~_T_343; // @[el2_ifu_bp_ctl.scala 342:36]
  wire  _T_348 = ~fetch_start_f[0]; // @[el2_ifu_bp_ctl.scala 346:36]
  wire  _T_349 = bht_dir_f[0] & _T_348; // @[el2_ifu_bp_ctl.scala 346:34]
  wire  _T_353 = _T_14 & fetch_start_f[0]; // @[el2_ifu_bp_ctl.scala 346:72]
  wire  _T_354 = _T_349 | _T_353; // @[el2_ifu_bp_ctl.scala 346:55]
  wire  _T_357 = bht_dir_f[0] & fetch_start_f[0]; // @[el2_ifu_bp_ctl.scala 347:34]
  wire  _T_362 = _T_14 & _T_348; // @[el2_ifu_bp_ctl.scala 347:71]
  wire  _T_363 = _T_357 | _T_362; // @[el2_ifu_bp_ctl.scala 347:54]
  wire [1:0] bloc_f = {_T_354,_T_363}; // @[Cat.scala 29:58]
  wire  _T_367 = _T_14 & io_ifc_fetch_addr_f[0]; // @[el2_ifu_bp_ctl.scala 349:35]
  wire  _T_368 = ~btb_rd_pc4_f; // @[el2_ifu_bp_ctl.scala 349:62]
  wire  use_fa_plus = _T_367 & _T_368; // @[el2_ifu_bp_ctl.scala 349:60]
  wire  _T_371 = fetch_start_f[0] & btb_sel_f[0]; // @[el2_ifu_bp_ctl.scala 351:44]
  wire  btb_fg_crossing_f = _T_371 & btb_rd_pc4_f; // @[el2_ifu_bp_ctl.scala 351:59]
  wire  bp_total_branch_offset_f = bloc_f[1] ^ btb_rd_pc4_f; // @[el2_ifu_bp_ctl.scala 352:43]
  wire  _T_375 = io_ifc_fetch_req_f & _T_275; // @[el2_ifu_bp_ctl.scala 354:85]
  reg [29:0] ifc_fetch_adder_prior; // @[el2_lib.scala 481:16]
  wire  _T_380 = ~btb_fg_crossing_f; // @[el2_ifu_bp_ctl.scala 360:32]
  wire  _T_381 = ~use_fa_plus; // @[el2_ifu_bp_ctl.scala 360:53]
  wire  _T_382 = _T_380 & _T_381; // @[el2_ifu_bp_ctl.scala 360:51]
  wire [29:0] _T_385 = use_fa_plus ? fetch_addr_p1_f : 30'h0; // @[Mux.scala 27:72]
  wire [29:0] _T_386 = btb_fg_crossing_f ? ifc_fetch_adder_prior : 30'h0; // @[Mux.scala 27:72]
  wire [29:0] _T_387 = _T_382 ? io_ifc_fetch_addr_f[30:1] : 30'h0; // @[Mux.scala 27:72]
  wire [29:0] _T_388 = _T_385 | _T_386; // @[Mux.scala 27:72]
  wire [29:0] adder_pc_in_f = _T_388 | _T_387; // @[Mux.scala 27:72]
  wire [31:0] _T_392 = {adder_pc_in_f,bp_total_branch_offset_f,1'h0}; // @[Cat.scala 29:58]
  wire [12:0] _T_393 = {btb_rd_tgt_f,1'h0}; // @[Cat.scala 29:58]
  wire [12:0] _T_396 = _T_392[12:1] + _T_393[12:1]; // @[el2_lib.scala 204:31]
  wire [18:0] _T_399 = _T_392[31:13] + 19'h1; // @[el2_lib.scala 205:27]
  wire [18:0] _T_402 = _T_392[31:13] - 19'h1; // @[el2_lib.scala 206:27]
  wire  _T_405 = ~_T_396[12]; // @[el2_lib.scala 208:28]
  wire  _T_406 = _T_393[12] ^ _T_405; // @[el2_lib.scala 208:26]
  wire  _T_409 = ~_T_393[12]; // @[el2_lib.scala 209:20]
  wire  _T_411 = _T_409 & _T_396[12]; // @[el2_lib.scala 209:26]
  wire  _T_415 = _T_393[12] & _T_405; // @[el2_lib.scala 210:26]
  wire [18:0] _T_417 = _T_406 ? _T_392[31:13] : 19'h0; // @[Mux.scala 27:72]
  wire [18:0] _T_418 = _T_411 ? _T_399 : 19'h0; // @[Mux.scala 27:72]
  wire [18:0] _T_419 = _T_415 ? _T_402 : 19'h0; // @[Mux.scala 27:72]
  wire [18:0] _T_420 = _T_417 | _T_418; // @[Mux.scala 27:72]
  wire [18:0] _T_421 = _T_420 | _T_419; // @[Mux.scala 27:72]
  wire [31:0] bp_btb_target_adder_f = {_T_421,_T_396[11:0],1'h0}; // @[Cat.scala 29:58]
  wire  _T_425 = ~btb_rd_call_f; // @[el2_ifu_bp_ctl.scala 369:49]
  wire  _T_426 = btb_rd_ret_f & _T_425; // @[el2_ifu_bp_ctl.scala 369:47]
  reg [31:0] rets_out_0; // @[el2_lib.scala 481:16]
  wire  _T_428 = _T_426 & rets_out_0[0]; // @[el2_ifu_bp_ctl.scala 369:64]
  wire [12:0] _T_439 = {11'h0,_T_368,1'h0}; // @[Cat.scala 29:58]
  wire [12:0] _T_442 = _T_392[12:1] + _T_439[12:1]; // @[el2_lib.scala 204:31]
  wire  _T_451 = ~_T_442[12]; // @[el2_lib.scala 208:28]
  wire  _T_452 = _T_439[12] ^ _T_451; // @[el2_lib.scala 208:26]
  wire  _T_455 = ~_T_439[12]; // @[el2_lib.scala 209:20]
  wire  _T_457 = _T_455 & _T_442[12]; // @[el2_lib.scala 209:26]
  wire  _T_461 = _T_439[12] & _T_451; // @[el2_lib.scala 210:26]
  wire [18:0] _T_463 = _T_452 ? _T_392[31:13] : 19'h0; // @[Mux.scala 27:72]
  wire [18:0] _T_464 = _T_457 ? _T_399 : 19'h0; // @[Mux.scala 27:72]
  wire [18:0] _T_465 = _T_461 ? _T_402 : 19'h0; // @[Mux.scala 27:72]
  wire [18:0] _T_466 = _T_463 | _T_464; // @[Mux.scala 27:72]
  wire [18:0] _T_467 = _T_466 | _T_465; // @[Mux.scala 27:72]
  wire [31:0] bp_rs_call_target_f = {_T_467,_T_442[11:0],1'h0}; // @[Cat.scala 29:58]
  wire  _T_471 = ~btb_rd_ret_f; // @[el2_ifu_bp_ctl.scala 375:33]
  wire  _T_472 = btb_rd_call_f & _T_471; // @[el2_ifu_bp_ctl.scala 375:31]
  wire  rs_push = _T_472 & io_ifu_bp_hit_taken_f; // @[el2_ifu_bp_ctl.scala 375:47]
  wire  rs_pop = _T_426 & io_ifu_bp_hit_taken_f; // @[el2_ifu_bp_ctl.scala 376:46]
  wire  _T_475 = ~rs_push; // @[el2_ifu_bp_ctl.scala 377:17]
  wire  _T_476 = ~rs_pop; // @[el2_ifu_bp_ctl.scala 377:28]
  wire  rs_hold = _T_475 & _T_476; // @[el2_ifu_bp_ctl.scala 377:26]
  wire [31:0] _T_479 = {bp_rs_call_target_f[31:1],1'h1}; // @[Cat.scala 29:58]
  wire [31:0] _T_481 = rs_push ? _T_479 : 32'h0; // @[Mux.scala 27:72]
  reg [31:0] rets_out_1; // @[el2_lib.scala 481:16]
  wire [31:0] _T_482 = rs_pop ? rets_out_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_486 = rs_push ? rets_out_0 : 32'h0; // @[Mux.scala 27:72]
  reg [31:0] rets_out_2; // @[el2_lib.scala 481:16]
  wire [31:0] _T_487 = rs_pop ? rets_out_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_491 = rs_push ? rets_out_1 : 32'h0; // @[Mux.scala 27:72]
  reg [31:0] rets_out_3; // @[el2_lib.scala 481:16]
  wire [31:0] _T_492 = rs_pop ? rets_out_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_496 = rs_push ? rets_out_2 : 32'h0; // @[Mux.scala 27:72]
  reg [31:0] rets_out_4; // @[el2_lib.scala 481:16]
  wire [31:0] _T_497 = rs_pop ? rets_out_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_501 = rs_push ? rets_out_3 : 32'h0; // @[Mux.scala 27:72]
  reg [31:0] rets_out_5; // @[el2_lib.scala 481:16]
  wire [31:0] _T_502 = rs_pop ? rets_out_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_506 = rs_push ? rets_out_4 : 32'h0; // @[Mux.scala 27:72]
  reg [31:0] rets_out_6; // @[el2_lib.scala 481:16]
  wire [31:0] _T_507 = rs_pop ? rets_out_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_511 = rs_push ? rets_out_5 : 32'h0; // @[Mux.scala 27:72]
  reg [31:0] rets_out_7; // @[el2_lib.scala 481:16]
  wire [31:0] _T_512 = rs_pop ? rets_out_7 : 32'h0; // @[Mux.scala 27:72]
  wire  _T_530 = ~dec_tlu_error_wb; // @[el2_ifu_bp_ctl.scala 392:35]
  wire  btb_valid = exu_mp_valid & _T_530; // @[el2_ifu_bp_ctl.scala 392:32]
  wire  _T_531 = io_exu_mp_pkt_pcall | io_exu_mp_pkt_pja; // @[el2_ifu_bp_ctl.scala 396:89]
  wire  _T_532 = io_exu_mp_pkt_pret | io_exu_mp_pkt_pja; // @[el2_ifu_bp_ctl.scala 396:113]
  wire [2:0] _T_534 = {_T_531,_T_532,btb_valid}; // @[Cat.scala 29:58]
  wire [18:0] _T_537 = {io_exu_mp_btag,io_exu_mp_pkt_toffset,io_exu_mp_pkt_pc4,io_exu_mp_pkt_boffset}; // @[Cat.scala 29:58]
  wire  exu_mp_valid_write = exu_mp_valid & io_exu_mp_pkt_ataken; // @[el2_ifu_bp_ctl.scala 397:41]
  wire  _T_539 = _T_175 & exu_mp_valid_write; // @[el2_ifu_bp_ctl.scala 400:39]
  wire  _T_541 = _T_539 & _T_530; // @[el2_ifu_bp_ctl.scala 400:60]
  wire  _T_542 = ~io_dec_tlu_br0_r_pkt_way; // @[el2_ifu_bp_ctl.scala 400:87]
  wire  _T_543 = _T_542 & dec_tlu_error_wb; // @[el2_ifu_bp_ctl.scala 400:104]
  wire  btb_wr_en_way0 = _T_541 | _T_543; // @[el2_ifu_bp_ctl.scala 400:83]
  wire  _T_544 = io_exu_mp_pkt_way & exu_mp_valid_write; // @[el2_ifu_bp_ctl.scala 401:36]
  wire  _T_546 = _T_544 & _T_530; // @[el2_ifu_bp_ctl.scala 401:57]
  wire  _T_547 = io_dec_tlu_br0_r_pkt_way & dec_tlu_error_wb; // @[el2_ifu_bp_ctl.scala 401:98]
  wire  btb_wr_en_way1 = _T_546 | _T_547; // @[el2_ifu_bp_ctl.scala 401:80]
  wire [7:0] btb_wr_addr = dec_tlu_error_wb ? io_exu_i0_br_index_r : io_exu_mp_index; // @[el2_ifu_bp_ctl.scala 404:24]
  wire  middle_of_bank = io_exu_mp_pkt_pc4 ^ io_exu_mp_pkt_boffset; // @[el2_ifu_bp_ctl.scala 405:35]
  wire  _T_549 = ~io_exu_mp_pkt_pcall; // @[el2_ifu_bp_ctl.scala 408:43]
  wire  _T_550 = exu_mp_valid & _T_549; // @[el2_ifu_bp_ctl.scala 408:41]
  wire  _T_551 = ~io_exu_mp_pkt_pret; // @[el2_ifu_bp_ctl.scala 408:58]
  wire  _T_552 = _T_550 & _T_551; // @[el2_ifu_bp_ctl.scala 408:56]
  wire  _T_553 = ~io_exu_mp_pkt_pja; // @[el2_ifu_bp_ctl.scala 408:72]
  wire  _T_554 = _T_552 & _T_553; // @[el2_ifu_bp_ctl.scala 408:70]
  wire [1:0] _T_556 = _T_554 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire  _T_557 = ~middle_of_bank; // @[el2_ifu_bp_ctl.scala 408:106]
  wire [1:0] _T_558 = {middle_of_bank,_T_557}; // @[Cat.scala 29:58]
  wire [1:0] bht_wr_en0 = _T_556 & _T_558; // @[el2_ifu_bp_ctl.scala 408:84]
  wire [1:0] _T_560 = io_dec_tlu_br0_r_pkt_valid ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire  _T_561 = ~io_dec_tlu_br0_r_pkt_middle; // @[el2_ifu_bp_ctl.scala 409:75]
  wire [1:0] _T_562 = {io_dec_tlu_br0_r_pkt_middle,_T_561}; // @[Cat.scala 29:58]
  wire [1:0] bht_wr_en2 = _T_560 & _T_562; // @[el2_ifu_bp_ctl.scala 409:46]
  wire [9:0] _T_563 = {io_exu_mp_index,2'h0}; // @[Cat.scala 29:58]
  wire [7:0] mp_hashed = _T_563[9:2] ^ io_exu_mp_eghr; // @[el2_lib.scala 194:35]
  wire [9:0] _T_566 = {io_exu_i0_br_index_r,2'h0}; // @[Cat.scala 29:58]
  wire [7:0] br0_hashed_wb = _T_566[9:2] ^ io_exu_i0_br_fghr_r; // @[el2_lib.scala 194:35]
  wire  _T_575 = btb_wr_addr == 8'h0; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_578 = btb_wr_addr == 8'h1; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_581 = btb_wr_addr == 8'h2; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_584 = btb_wr_addr == 8'h3; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_587 = btb_wr_addr == 8'h4; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_590 = btb_wr_addr == 8'h5; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_593 = btb_wr_addr == 8'h6; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_596 = btb_wr_addr == 8'h7; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_599 = btb_wr_addr == 8'h8; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_602 = btb_wr_addr == 8'h9; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_605 = btb_wr_addr == 8'ha; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_608 = btb_wr_addr == 8'hb; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_611 = btb_wr_addr == 8'hc; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_614 = btb_wr_addr == 8'hd; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_617 = btb_wr_addr == 8'he; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_620 = btb_wr_addr == 8'hf; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_623 = btb_wr_addr == 8'h10; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_626 = btb_wr_addr == 8'h11; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_629 = btb_wr_addr == 8'h12; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_632 = btb_wr_addr == 8'h13; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_635 = btb_wr_addr == 8'h14; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_638 = btb_wr_addr == 8'h15; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_641 = btb_wr_addr == 8'h16; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_644 = btb_wr_addr == 8'h17; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_647 = btb_wr_addr == 8'h18; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_650 = btb_wr_addr == 8'h19; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_653 = btb_wr_addr == 8'h1a; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_656 = btb_wr_addr == 8'h1b; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_659 = btb_wr_addr == 8'h1c; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_662 = btb_wr_addr == 8'h1d; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_665 = btb_wr_addr == 8'h1e; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_668 = btb_wr_addr == 8'h1f; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_671 = btb_wr_addr == 8'h20; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_674 = btb_wr_addr == 8'h21; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_677 = btb_wr_addr == 8'h22; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_680 = btb_wr_addr == 8'h23; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_683 = btb_wr_addr == 8'h24; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_686 = btb_wr_addr == 8'h25; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_689 = btb_wr_addr == 8'h26; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_692 = btb_wr_addr == 8'h27; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_695 = btb_wr_addr == 8'h28; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_698 = btb_wr_addr == 8'h29; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_701 = btb_wr_addr == 8'h2a; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_704 = btb_wr_addr == 8'h2b; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_707 = btb_wr_addr == 8'h2c; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_710 = btb_wr_addr == 8'h2d; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_713 = btb_wr_addr == 8'h2e; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_716 = btb_wr_addr == 8'h2f; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_719 = btb_wr_addr == 8'h30; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_722 = btb_wr_addr == 8'h31; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_725 = btb_wr_addr == 8'h32; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_728 = btb_wr_addr == 8'h33; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_731 = btb_wr_addr == 8'h34; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_734 = btb_wr_addr == 8'h35; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_737 = btb_wr_addr == 8'h36; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_740 = btb_wr_addr == 8'h37; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_743 = btb_wr_addr == 8'h38; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_746 = btb_wr_addr == 8'h39; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_749 = btb_wr_addr == 8'h3a; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_752 = btb_wr_addr == 8'h3b; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_755 = btb_wr_addr == 8'h3c; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_758 = btb_wr_addr == 8'h3d; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_761 = btb_wr_addr == 8'h3e; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_764 = btb_wr_addr == 8'h3f; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_767 = btb_wr_addr == 8'h40; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_770 = btb_wr_addr == 8'h41; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_773 = btb_wr_addr == 8'h42; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_776 = btb_wr_addr == 8'h43; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_779 = btb_wr_addr == 8'h44; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_782 = btb_wr_addr == 8'h45; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_785 = btb_wr_addr == 8'h46; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_788 = btb_wr_addr == 8'h47; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_791 = btb_wr_addr == 8'h48; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_794 = btb_wr_addr == 8'h49; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_797 = btb_wr_addr == 8'h4a; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_800 = btb_wr_addr == 8'h4b; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_803 = btb_wr_addr == 8'h4c; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_806 = btb_wr_addr == 8'h4d; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_809 = btb_wr_addr == 8'h4e; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_812 = btb_wr_addr == 8'h4f; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_815 = btb_wr_addr == 8'h50; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_818 = btb_wr_addr == 8'h51; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_821 = btb_wr_addr == 8'h52; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_824 = btb_wr_addr == 8'h53; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_827 = btb_wr_addr == 8'h54; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_830 = btb_wr_addr == 8'h55; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_833 = btb_wr_addr == 8'h56; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_836 = btb_wr_addr == 8'h57; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_839 = btb_wr_addr == 8'h58; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_842 = btb_wr_addr == 8'h59; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_845 = btb_wr_addr == 8'h5a; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_848 = btb_wr_addr == 8'h5b; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_851 = btb_wr_addr == 8'h5c; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_854 = btb_wr_addr == 8'h5d; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_857 = btb_wr_addr == 8'h5e; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_860 = btb_wr_addr == 8'h5f; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_863 = btb_wr_addr == 8'h60; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_866 = btb_wr_addr == 8'h61; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_869 = btb_wr_addr == 8'h62; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_872 = btb_wr_addr == 8'h63; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_875 = btb_wr_addr == 8'h64; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_878 = btb_wr_addr == 8'h65; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_881 = btb_wr_addr == 8'h66; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_884 = btb_wr_addr == 8'h67; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_887 = btb_wr_addr == 8'h68; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_890 = btb_wr_addr == 8'h69; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_893 = btb_wr_addr == 8'h6a; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_896 = btb_wr_addr == 8'h6b; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_899 = btb_wr_addr == 8'h6c; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_902 = btb_wr_addr == 8'h6d; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_905 = btb_wr_addr == 8'h6e; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_908 = btb_wr_addr == 8'h6f; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_911 = btb_wr_addr == 8'h70; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_914 = btb_wr_addr == 8'h71; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_917 = btb_wr_addr == 8'h72; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_920 = btb_wr_addr == 8'h73; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_923 = btb_wr_addr == 8'h74; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_926 = btb_wr_addr == 8'h75; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_929 = btb_wr_addr == 8'h76; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_932 = btb_wr_addr == 8'h77; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_935 = btb_wr_addr == 8'h78; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_938 = btb_wr_addr == 8'h79; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_941 = btb_wr_addr == 8'h7a; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_944 = btb_wr_addr == 8'h7b; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_947 = btb_wr_addr == 8'h7c; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_950 = btb_wr_addr == 8'h7d; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_953 = btb_wr_addr == 8'h7e; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_956 = btb_wr_addr == 8'h7f; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_959 = btb_wr_addr == 8'h80; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_962 = btb_wr_addr == 8'h81; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_965 = btb_wr_addr == 8'h82; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_968 = btb_wr_addr == 8'h83; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_971 = btb_wr_addr == 8'h84; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_974 = btb_wr_addr == 8'h85; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_977 = btb_wr_addr == 8'h86; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_980 = btb_wr_addr == 8'h87; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_983 = btb_wr_addr == 8'h88; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_986 = btb_wr_addr == 8'h89; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_989 = btb_wr_addr == 8'h8a; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_992 = btb_wr_addr == 8'h8b; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_995 = btb_wr_addr == 8'h8c; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_998 = btb_wr_addr == 8'h8d; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1001 = btb_wr_addr == 8'h8e; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1004 = btb_wr_addr == 8'h8f; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1007 = btb_wr_addr == 8'h90; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1010 = btb_wr_addr == 8'h91; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1013 = btb_wr_addr == 8'h92; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1016 = btb_wr_addr == 8'h93; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1019 = btb_wr_addr == 8'h94; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1022 = btb_wr_addr == 8'h95; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1025 = btb_wr_addr == 8'h96; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1028 = btb_wr_addr == 8'h97; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1031 = btb_wr_addr == 8'h98; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1034 = btb_wr_addr == 8'h99; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1037 = btb_wr_addr == 8'h9a; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1040 = btb_wr_addr == 8'h9b; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1043 = btb_wr_addr == 8'h9c; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1046 = btb_wr_addr == 8'h9d; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1049 = btb_wr_addr == 8'h9e; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1052 = btb_wr_addr == 8'h9f; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1055 = btb_wr_addr == 8'ha0; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1058 = btb_wr_addr == 8'ha1; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1061 = btb_wr_addr == 8'ha2; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1064 = btb_wr_addr == 8'ha3; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1067 = btb_wr_addr == 8'ha4; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1070 = btb_wr_addr == 8'ha5; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1073 = btb_wr_addr == 8'ha6; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1076 = btb_wr_addr == 8'ha7; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1079 = btb_wr_addr == 8'ha8; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1082 = btb_wr_addr == 8'ha9; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1085 = btb_wr_addr == 8'haa; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1088 = btb_wr_addr == 8'hab; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1091 = btb_wr_addr == 8'hac; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1094 = btb_wr_addr == 8'had; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1097 = btb_wr_addr == 8'hae; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1100 = btb_wr_addr == 8'haf; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1103 = btb_wr_addr == 8'hb0; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1106 = btb_wr_addr == 8'hb1; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1109 = btb_wr_addr == 8'hb2; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1112 = btb_wr_addr == 8'hb3; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1115 = btb_wr_addr == 8'hb4; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1118 = btb_wr_addr == 8'hb5; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1121 = btb_wr_addr == 8'hb6; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1124 = btb_wr_addr == 8'hb7; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1127 = btb_wr_addr == 8'hb8; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1130 = btb_wr_addr == 8'hb9; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1133 = btb_wr_addr == 8'hba; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1136 = btb_wr_addr == 8'hbb; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1139 = btb_wr_addr == 8'hbc; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1142 = btb_wr_addr == 8'hbd; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1145 = btb_wr_addr == 8'hbe; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1148 = btb_wr_addr == 8'hbf; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1151 = btb_wr_addr == 8'hc0; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1154 = btb_wr_addr == 8'hc1; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1157 = btb_wr_addr == 8'hc2; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1160 = btb_wr_addr == 8'hc3; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1163 = btb_wr_addr == 8'hc4; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1166 = btb_wr_addr == 8'hc5; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1169 = btb_wr_addr == 8'hc6; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1172 = btb_wr_addr == 8'hc7; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1175 = btb_wr_addr == 8'hc8; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1178 = btb_wr_addr == 8'hc9; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1181 = btb_wr_addr == 8'hca; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1184 = btb_wr_addr == 8'hcb; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1187 = btb_wr_addr == 8'hcc; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1190 = btb_wr_addr == 8'hcd; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1193 = btb_wr_addr == 8'hce; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1196 = btb_wr_addr == 8'hcf; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1199 = btb_wr_addr == 8'hd0; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1202 = btb_wr_addr == 8'hd1; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1205 = btb_wr_addr == 8'hd2; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1208 = btb_wr_addr == 8'hd3; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1211 = btb_wr_addr == 8'hd4; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1214 = btb_wr_addr == 8'hd5; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1217 = btb_wr_addr == 8'hd6; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1220 = btb_wr_addr == 8'hd7; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1223 = btb_wr_addr == 8'hd8; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1226 = btb_wr_addr == 8'hd9; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1229 = btb_wr_addr == 8'hda; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1232 = btb_wr_addr == 8'hdb; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1235 = btb_wr_addr == 8'hdc; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1238 = btb_wr_addr == 8'hdd; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1241 = btb_wr_addr == 8'hde; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1244 = btb_wr_addr == 8'hdf; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1247 = btb_wr_addr == 8'he0; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1250 = btb_wr_addr == 8'he1; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1253 = btb_wr_addr == 8'he2; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1256 = btb_wr_addr == 8'he3; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1259 = btb_wr_addr == 8'he4; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1262 = btb_wr_addr == 8'he5; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1265 = btb_wr_addr == 8'he6; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1268 = btb_wr_addr == 8'he7; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1271 = btb_wr_addr == 8'he8; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1274 = btb_wr_addr == 8'he9; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1277 = btb_wr_addr == 8'hea; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1280 = btb_wr_addr == 8'heb; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1283 = btb_wr_addr == 8'hec; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1286 = btb_wr_addr == 8'hed; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1289 = btb_wr_addr == 8'hee; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1292 = btb_wr_addr == 8'hef; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1295 = btb_wr_addr == 8'hf0; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1298 = btb_wr_addr == 8'hf1; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1301 = btb_wr_addr == 8'hf2; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1304 = btb_wr_addr == 8'hf3; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1307 = btb_wr_addr == 8'hf4; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1310 = btb_wr_addr == 8'hf5; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1313 = btb_wr_addr == 8'hf6; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1316 = btb_wr_addr == 8'hf7; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1319 = btb_wr_addr == 8'hf8; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1322 = btb_wr_addr == 8'hf9; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1325 = btb_wr_addr == 8'hfa; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1328 = btb_wr_addr == 8'hfb; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1331 = btb_wr_addr == 8'hfc; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1334 = btb_wr_addr == 8'hfd; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1337 = btb_wr_addr == 8'hfe; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_1340 = btb_wr_addr == 8'hff; // @[el2_ifu_bp_ctl.scala 427:95]
  wire  _T_6209 = mp_hashed[7:4] == 4'h0; // @[el2_ifu_bp_ctl.scala 441:109]
  wire  _T_6211 = bht_wr_en0[0] & _T_6209; // @[el2_ifu_bp_ctl.scala 441:44]
  wire  _T_6214 = br0_hashed_wb[7:4] == 4'h0; // @[el2_ifu_bp_ctl.scala 442:109]
  wire  _T_6216 = bht_wr_en2[0] & _T_6214; // @[el2_ifu_bp_ctl.scala 442:44]
  wire  _T_6220 = mp_hashed[7:4] == 4'h1; // @[el2_ifu_bp_ctl.scala 441:109]
  wire  _T_6222 = bht_wr_en0[0] & _T_6220; // @[el2_ifu_bp_ctl.scala 441:44]
  wire  _T_6225 = br0_hashed_wb[7:4] == 4'h1; // @[el2_ifu_bp_ctl.scala 442:109]
  wire  _T_6227 = bht_wr_en2[0] & _T_6225; // @[el2_ifu_bp_ctl.scala 442:44]
  wire  _T_6231 = mp_hashed[7:4] == 4'h2; // @[el2_ifu_bp_ctl.scala 441:109]
  wire  _T_6233 = bht_wr_en0[0] & _T_6231; // @[el2_ifu_bp_ctl.scala 441:44]
  wire  _T_6236 = br0_hashed_wb[7:4] == 4'h2; // @[el2_ifu_bp_ctl.scala 442:109]
  wire  _T_6238 = bht_wr_en2[0] & _T_6236; // @[el2_ifu_bp_ctl.scala 442:44]
  wire  _T_6242 = mp_hashed[7:4] == 4'h3; // @[el2_ifu_bp_ctl.scala 441:109]
  wire  _T_6244 = bht_wr_en0[0] & _T_6242; // @[el2_ifu_bp_ctl.scala 441:44]
  wire  _T_6247 = br0_hashed_wb[7:4] == 4'h3; // @[el2_ifu_bp_ctl.scala 442:109]
  wire  _T_6249 = bht_wr_en2[0] & _T_6247; // @[el2_ifu_bp_ctl.scala 442:44]
  wire  _T_6253 = mp_hashed[7:4] == 4'h4; // @[el2_ifu_bp_ctl.scala 441:109]
  wire  _T_6255 = bht_wr_en0[0] & _T_6253; // @[el2_ifu_bp_ctl.scala 441:44]
  wire  _T_6258 = br0_hashed_wb[7:4] == 4'h4; // @[el2_ifu_bp_ctl.scala 442:109]
  wire  _T_6260 = bht_wr_en2[0] & _T_6258; // @[el2_ifu_bp_ctl.scala 442:44]
  wire  _T_6264 = mp_hashed[7:4] == 4'h5; // @[el2_ifu_bp_ctl.scala 441:109]
  wire  _T_6266 = bht_wr_en0[0] & _T_6264; // @[el2_ifu_bp_ctl.scala 441:44]
  wire  _T_6269 = br0_hashed_wb[7:4] == 4'h5; // @[el2_ifu_bp_ctl.scala 442:109]
  wire  _T_6271 = bht_wr_en2[0] & _T_6269; // @[el2_ifu_bp_ctl.scala 442:44]
  wire  _T_6275 = mp_hashed[7:4] == 4'h6; // @[el2_ifu_bp_ctl.scala 441:109]
  wire  _T_6277 = bht_wr_en0[0] & _T_6275; // @[el2_ifu_bp_ctl.scala 441:44]
  wire  _T_6280 = br0_hashed_wb[7:4] == 4'h6; // @[el2_ifu_bp_ctl.scala 442:109]
  wire  _T_6282 = bht_wr_en2[0] & _T_6280; // @[el2_ifu_bp_ctl.scala 442:44]
  wire  _T_6286 = mp_hashed[7:4] == 4'h7; // @[el2_ifu_bp_ctl.scala 441:109]
  wire  _T_6288 = bht_wr_en0[0] & _T_6286; // @[el2_ifu_bp_ctl.scala 441:44]
  wire  _T_6291 = br0_hashed_wb[7:4] == 4'h7; // @[el2_ifu_bp_ctl.scala 442:109]
  wire  _T_6293 = bht_wr_en2[0] & _T_6291; // @[el2_ifu_bp_ctl.scala 442:44]
  wire  _T_6297 = mp_hashed[7:4] == 4'h8; // @[el2_ifu_bp_ctl.scala 441:109]
  wire  _T_6299 = bht_wr_en0[0] & _T_6297; // @[el2_ifu_bp_ctl.scala 441:44]
  wire  _T_6302 = br0_hashed_wb[7:4] == 4'h8; // @[el2_ifu_bp_ctl.scala 442:109]
  wire  _T_6304 = bht_wr_en2[0] & _T_6302; // @[el2_ifu_bp_ctl.scala 442:44]
  wire  _T_6308 = mp_hashed[7:4] == 4'h9; // @[el2_ifu_bp_ctl.scala 441:109]
  wire  _T_6310 = bht_wr_en0[0] & _T_6308; // @[el2_ifu_bp_ctl.scala 441:44]
  wire  _T_6313 = br0_hashed_wb[7:4] == 4'h9; // @[el2_ifu_bp_ctl.scala 442:109]
  wire  _T_6315 = bht_wr_en2[0] & _T_6313; // @[el2_ifu_bp_ctl.scala 442:44]
  wire  _T_6319 = mp_hashed[7:4] == 4'ha; // @[el2_ifu_bp_ctl.scala 441:109]
  wire  _T_6321 = bht_wr_en0[0] & _T_6319; // @[el2_ifu_bp_ctl.scala 441:44]
  wire  _T_6324 = br0_hashed_wb[7:4] == 4'ha; // @[el2_ifu_bp_ctl.scala 442:109]
  wire  _T_6326 = bht_wr_en2[0] & _T_6324; // @[el2_ifu_bp_ctl.scala 442:44]
  wire  _T_6330 = mp_hashed[7:4] == 4'hb; // @[el2_ifu_bp_ctl.scala 441:109]
  wire  _T_6332 = bht_wr_en0[0] & _T_6330; // @[el2_ifu_bp_ctl.scala 441:44]
  wire  _T_6335 = br0_hashed_wb[7:4] == 4'hb; // @[el2_ifu_bp_ctl.scala 442:109]
  wire  _T_6337 = bht_wr_en2[0] & _T_6335; // @[el2_ifu_bp_ctl.scala 442:44]
  wire  _T_6341 = mp_hashed[7:4] == 4'hc; // @[el2_ifu_bp_ctl.scala 441:109]
  wire  _T_6343 = bht_wr_en0[0] & _T_6341; // @[el2_ifu_bp_ctl.scala 441:44]
  wire  _T_6346 = br0_hashed_wb[7:4] == 4'hc; // @[el2_ifu_bp_ctl.scala 442:109]
  wire  _T_6348 = bht_wr_en2[0] & _T_6346; // @[el2_ifu_bp_ctl.scala 442:44]
  wire  _T_6352 = mp_hashed[7:4] == 4'hd; // @[el2_ifu_bp_ctl.scala 441:109]
  wire  _T_6354 = bht_wr_en0[0] & _T_6352; // @[el2_ifu_bp_ctl.scala 441:44]
  wire  _T_6357 = br0_hashed_wb[7:4] == 4'hd; // @[el2_ifu_bp_ctl.scala 442:109]
  wire  _T_6359 = bht_wr_en2[0] & _T_6357; // @[el2_ifu_bp_ctl.scala 442:44]
  wire  _T_6363 = mp_hashed[7:4] == 4'he; // @[el2_ifu_bp_ctl.scala 441:109]
  wire  _T_6365 = bht_wr_en0[0] & _T_6363; // @[el2_ifu_bp_ctl.scala 441:44]
  wire  _T_6368 = br0_hashed_wb[7:4] == 4'he; // @[el2_ifu_bp_ctl.scala 442:109]
  wire  _T_6370 = bht_wr_en2[0] & _T_6368; // @[el2_ifu_bp_ctl.scala 442:44]
  wire  _T_6374 = mp_hashed[7:4] == 4'hf; // @[el2_ifu_bp_ctl.scala 441:109]
  wire  _T_6376 = bht_wr_en0[0] & _T_6374; // @[el2_ifu_bp_ctl.scala 441:44]
  wire  _T_6379 = br0_hashed_wb[7:4] == 4'hf; // @[el2_ifu_bp_ctl.scala 442:109]
  wire  _T_6381 = bht_wr_en2[0] & _T_6379; // @[el2_ifu_bp_ctl.scala 442:44]
  wire  _T_6387 = bht_wr_en0[1] & _T_6209; // @[el2_ifu_bp_ctl.scala 441:44]
  wire  _T_6392 = bht_wr_en2[1] & _T_6214; // @[el2_ifu_bp_ctl.scala 442:44]
  wire  _T_6398 = bht_wr_en0[1] & _T_6220; // @[el2_ifu_bp_ctl.scala 441:44]
  wire  _T_6403 = bht_wr_en2[1] & _T_6225; // @[el2_ifu_bp_ctl.scala 442:44]
  wire  _T_6409 = bht_wr_en0[1] & _T_6231; // @[el2_ifu_bp_ctl.scala 441:44]
  wire  _T_6414 = bht_wr_en2[1] & _T_6236; // @[el2_ifu_bp_ctl.scala 442:44]
  wire  _T_6420 = bht_wr_en0[1] & _T_6242; // @[el2_ifu_bp_ctl.scala 441:44]
  wire  _T_6425 = bht_wr_en2[1] & _T_6247; // @[el2_ifu_bp_ctl.scala 442:44]
  wire  _T_6431 = bht_wr_en0[1] & _T_6253; // @[el2_ifu_bp_ctl.scala 441:44]
  wire  _T_6436 = bht_wr_en2[1] & _T_6258; // @[el2_ifu_bp_ctl.scala 442:44]
  wire  _T_6442 = bht_wr_en0[1] & _T_6264; // @[el2_ifu_bp_ctl.scala 441:44]
  wire  _T_6447 = bht_wr_en2[1] & _T_6269; // @[el2_ifu_bp_ctl.scala 442:44]
  wire  _T_6453 = bht_wr_en0[1] & _T_6275; // @[el2_ifu_bp_ctl.scala 441:44]
  wire  _T_6458 = bht_wr_en2[1] & _T_6280; // @[el2_ifu_bp_ctl.scala 442:44]
  wire  _T_6464 = bht_wr_en0[1] & _T_6286; // @[el2_ifu_bp_ctl.scala 441:44]
  wire  _T_6469 = bht_wr_en2[1] & _T_6291; // @[el2_ifu_bp_ctl.scala 442:44]
  wire  _T_6475 = bht_wr_en0[1] & _T_6297; // @[el2_ifu_bp_ctl.scala 441:44]
  wire  _T_6480 = bht_wr_en2[1] & _T_6302; // @[el2_ifu_bp_ctl.scala 442:44]
  wire  _T_6486 = bht_wr_en0[1] & _T_6308; // @[el2_ifu_bp_ctl.scala 441:44]
  wire  _T_6491 = bht_wr_en2[1] & _T_6313; // @[el2_ifu_bp_ctl.scala 442:44]
  wire  _T_6497 = bht_wr_en0[1] & _T_6319; // @[el2_ifu_bp_ctl.scala 441:44]
  wire  _T_6502 = bht_wr_en2[1] & _T_6324; // @[el2_ifu_bp_ctl.scala 442:44]
  wire  _T_6508 = bht_wr_en0[1] & _T_6330; // @[el2_ifu_bp_ctl.scala 441:44]
  wire  _T_6513 = bht_wr_en2[1] & _T_6335; // @[el2_ifu_bp_ctl.scala 442:44]
  wire  _T_6519 = bht_wr_en0[1] & _T_6341; // @[el2_ifu_bp_ctl.scala 441:44]
  wire  _T_6524 = bht_wr_en2[1] & _T_6346; // @[el2_ifu_bp_ctl.scala 442:44]
  wire  _T_6530 = bht_wr_en0[1] & _T_6352; // @[el2_ifu_bp_ctl.scala 441:44]
  wire  _T_6535 = bht_wr_en2[1] & _T_6357; // @[el2_ifu_bp_ctl.scala 442:44]
  wire  _T_6541 = bht_wr_en0[1] & _T_6363; // @[el2_ifu_bp_ctl.scala 441:44]
  wire  _T_6546 = bht_wr_en2[1] & _T_6368; // @[el2_ifu_bp_ctl.scala 442:44]
  wire  _T_6552 = bht_wr_en0[1] & _T_6374; // @[el2_ifu_bp_ctl.scala 441:44]
  wire  _T_6557 = bht_wr_en2[1] & _T_6379; // @[el2_ifu_bp_ctl.scala 442:44]
  wire  _T_6561 = br0_hashed_wb[3:0] == 4'h0; // @[el2_ifu_bp_ctl.scala 447:74]
  wire  _T_6562 = bht_wr_en2[0] & _T_6561; // @[el2_ifu_bp_ctl.scala 447:23]
  wire  _T_6565 = _T_6562 & _T_6214; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_6570 = br0_hashed_wb[3:0] == 4'h1; // @[el2_ifu_bp_ctl.scala 447:74]
  wire  _T_6571 = bht_wr_en2[0] & _T_6570; // @[el2_ifu_bp_ctl.scala 447:23]
  wire  _T_6574 = _T_6571 & _T_6214; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_6579 = br0_hashed_wb[3:0] == 4'h2; // @[el2_ifu_bp_ctl.scala 447:74]
  wire  _T_6580 = bht_wr_en2[0] & _T_6579; // @[el2_ifu_bp_ctl.scala 447:23]
  wire  _T_6583 = _T_6580 & _T_6214; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_6588 = br0_hashed_wb[3:0] == 4'h3; // @[el2_ifu_bp_ctl.scala 447:74]
  wire  _T_6589 = bht_wr_en2[0] & _T_6588; // @[el2_ifu_bp_ctl.scala 447:23]
  wire  _T_6592 = _T_6589 & _T_6214; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_6597 = br0_hashed_wb[3:0] == 4'h4; // @[el2_ifu_bp_ctl.scala 447:74]
  wire  _T_6598 = bht_wr_en2[0] & _T_6597; // @[el2_ifu_bp_ctl.scala 447:23]
  wire  _T_6601 = _T_6598 & _T_6214; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_6606 = br0_hashed_wb[3:0] == 4'h5; // @[el2_ifu_bp_ctl.scala 447:74]
  wire  _T_6607 = bht_wr_en2[0] & _T_6606; // @[el2_ifu_bp_ctl.scala 447:23]
  wire  _T_6610 = _T_6607 & _T_6214; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_6615 = br0_hashed_wb[3:0] == 4'h6; // @[el2_ifu_bp_ctl.scala 447:74]
  wire  _T_6616 = bht_wr_en2[0] & _T_6615; // @[el2_ifu_bp_ctl.scala 447:23]
  wire  _T_6619 = _T_6616 & _T_6214; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_6624 = br0_hashed_wb[3:0] == 4'h7; // @[el2_ifu_bp_ctl.scala 447:74]
  wire  _T_6625 = bht_wr_en2[0] & _T_6624; // @[el2_ifu_bp_ctl.scala 447:23]
  wire  _T_6628 = _T_6625 & _T_6214; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_6633 = br0_hashed_wb[3:0] == 4'h8; // @[el2_ifu_bp_ctl.scala 447:74]
  wire  _T_6634 = bht_wr_en2[0] & _T_6633; // @[el2_ifu_bp_ctl.scala 447:23]
  wire  _T_6637 = _T_6634 & _T_6214; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_6642 = br0_hashed_wb[3:0] == 4'h9; // @[el2_ifu_bp_ctl.scala 447:74]
  wire  _T_6643 = bht_wr_en2[0] & _T_6642; // @[el2_ifu_bp_ctl.scala 447:23]
  wire  _T_6646 = _T_6643 & _T_6214; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_6651 = br0_hashed_wb[3:0] == 4'ha; // @[el2_ifu_bp_ctl.scala 447:74]
  wire  _T_6652 = bht_wr_en2[0] & _T_6651; // @[el2_ifu_bp_ctl.scala 447:23]
  wire  _T_6655 = _T_6652 & _T_6214; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_6660 = br0_hashed_wb[3:0] == 4'hb; // @[el2_ifu_bp_ctl.scala 447:74]
  wire  _T_6661 = bht_wr_en2[0] & _T_6660; // @[el2_ifu_bp_ctl.scala 447:23]
  wire  _T_6664 = _T_6661 & _T_6214; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_6669 = br0_hashed_wb[3:0] == 4'hc; // @[el2_ifu_bp_ctl.scala 447:74]
  wire  _T_6670 = bht_wr_en2[0] & _T_6669; // @[el2_ifu_bp_ctl.scala 447:23]
  wire  _T_6673 = _T_6670 & _T_6214; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_6678 = br0_hashed_wb[3:0] == 4'hd; // @[el2_ifu_bp_ctl.scala 447:74]
  wire  _T_6679 = bht_wr_en2[0] & _T_6678; // @[el2_ifu_bp_ctl.scala 447:23]
  wire  _T_6682 = _T_6679 & _T_6214; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_6687 = br0_hashed_wb[3:0] == 4'he; // @[el2_ifu_bp_ctl.scala 447:74]
  wire  _T_6688 = bht_wr_en2[0] & _T_6687; // @[el2_ifu_bp_ctl.scala 447:23]
  wire  _T_6691 = _T_6688 & _T_6214; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_6696 = br0_hashed_wb[3:0] == 4'hf; // @[el2_ifu_bp_ctl.scala 447:74]
  wire  _T_6697 = bht_wr_en2[0] & _T_6696; // @[el2_ifu_bp_ctl.scala 447:23]
  wire  _T_6700 = _T_6697 & _T_6214; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_6709 = _T_6562 & _T_6225; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_6718 = _T_6571 & _T_6225; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_6727 = _T_6580 & _T_6225; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_6736 = _T_6589 & _T_6225; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_6745 = _T_6598 & _T_6225; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_6754 = _T_6607 & _T_6225; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_6763 = _T_6616 & _T_6225; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_6772 = _T_6625 & _T_6225; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_6781 = _T_6634 & _T_6225; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_6790 = _T_6643 & _T_6225; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_6799 = _T_6652 & _T_6225; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_6808 = _T_6661 & _T_6225; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_6817 = _T_6670 & _T_6225; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_6826 = _T_6679 & _T_6225; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_6835 = _T_6688 & _T_6225; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_6844 = _T_6697 & _T_6225; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_6853 = _T_6562 & _T_6236; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_6862 = _T_6571 & _T_6236; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_6871 = _T_6580 & _T_6236; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_6880 = _T_6589 & _T_6236; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_6889 = _T_6598 & _T_6236; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_6898 = _T_6607 & _T_6236; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_6907 = _T_6616 & _T_6236; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_6916 = _T_6625 & _T_6236; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_6925 = _T_6634 & _T_6236; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_6934 = _T_6643 & _T_6236; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_6943 = _T_6652 & _T_6236; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_6952 = _T_6661 & _T_6236; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_6961 = _T_6670 & _T_6236; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_6970 = _T_6679 & _T_6236; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_6979 = _T_6688 & _T_6236; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_6988 = _T_6697 & _T_6236; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_6997 = _T_6562 & _T_6247; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_7006 = _T_6571 & _T_6247; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_7015 = _T_6580 & _T_6247; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_7024 = _T_6589 & _T_6247; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_7033 = _T_6598 & _T_6247; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_7042 = _T_6607 & _T_6247; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_7051 = _T_6616 & _T_6247; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_7060 = _T_6625 & _T_6247; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_7069 = _T_6634 & _T_6247; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_7078 = _T_6643 & _T_6247; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_7087 = _T_6652 & _T_6247; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_7096 = _T_6661 & _T_6247; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_7105 = _T_6670 & _T_6247; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_7114 = _T_6679 & _T_6247; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_7123 = _T_6688 & _T_6247; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_7132 = _T_6697 & _T_6247; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_7141 = _T_6562 & _T_6258; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_7150 = _T_6571 & _T_6258; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_7159 = _T_6580 & _T_6258; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_7168 = _T_6589 & _T_6258; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_7177 = _T_6598 & _T_6258; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_7186 = _T_6607 & _T_6258; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_7195 = _T_6616 & _T_6258; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_7204 = _T_6625 & _T_6258; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_7213 = _T_6634 & _T_6258; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_7222 = _T_6643 & _T_6258; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_7231 = _T_6652 & _T_6258; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_7240 = _T_6661 & _T_6258; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_7249 = _T_6670 & _T_6258; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_7258 = _T_6679 & _T_6258; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_7267 = _T_6688 & _T_6258; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_7276 = _T_6697 & _T_6258; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_7285 = _T_6562 & _T_6269; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_7294 = _T_6571 & _T_6269; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_7303 = _T_6580 & _T_6269; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_7312 = _T_6589 & _T_6269; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_7321 = _T_6598 & _T_6269; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_7330 = _T_6607 & _T_6269; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_7339 = _T_6616 & _T_6269; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_7348 = _T_6625 & _T_6269; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_7357 = _T_6634 & _T_6269; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_7366 = _T_6643 & _T_6269; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_7375 = _T_6652 & _T_6269; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_7384 = _T_6661 & _T_6269; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_7393 = _T_6670 & _T_6269; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_7402 = _T_6679 & _T_6269; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_7411 = _T_6688 & _T_6269; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_7420 = _T_6697 & _T_6269; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_7429 = _T_6562 & _T_6280; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_7438 = _T_6571 & _T_6280; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_7447 = _T_6580 & _T_6280; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_7456 = _T_6589 & _T_6280; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_7465 = _T_6598 & _T_6280; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_7474 = _T_6607 & _T_6280; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_7483 = _T_6616 & _T_6280; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_7492 = _T_6625 & _T_6280; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_7501 = _T_6634 & _T_6280; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_7510 = _T_6643 & _T_6280; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_7519 = _T_6652 & _T_6280; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_7528 = _T_6661 & _T_6280; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_7537 = _T_6670 & _T_6280; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_7546 = _T_6679 & _T_6280; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_7555 = _T_6688 & _T_6280; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_7564 = _T_6697 & _T_6280; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_7573 = _T_6562 & _T_6291; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_7582 = _T_6571 & _T_6291; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_7591 = _T_6580 & _T_6291; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_7600 = _T_6589 & _T_6291; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_7609 = _T_6598 & _T_6291; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_7618 = _T_6607 & _T_6291; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_7627 = _T_6616 & _T_6291; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_7636 = _T_6625 & _T_6291; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_7645 = _T_6634 & _T_6291; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_7654 = _T_6643 & _T_6291; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_7663 = _T_6652 & _T_6291; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_7672 = _T_6661 & _T_6291; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_7681 = _T_6670 & _T_6291; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_7690 = _T_6679 & _T_6291; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_7699 = _T_6688 & _T_6291; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_7708 = _T_6697 & _T_6291; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_7717 = _T_6562 & _T_6302; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_7726 = _T_6571 & _T_6302; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_7735 = _T_6580 & _T_6302; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_7744 = _T_6589 & _T_6302; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_7753 = _T_6598 & _T_6302; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_7762 = _T_6607 & _T_6302; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_7771 = _T_6616 & _T_6302; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_7780 = _T_6625 & _T_6302; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_7789 = _T_6634 & _T_6302; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_7798 = _T_6643 & _T_6302; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_7807 = _T_6652 & _T_6302; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_7816 = _T_6661 & _T_6302; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_7825 = _T_6670 & _T_6302; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_7834 = _T_6679 & _T_6302; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_7843 = _T_6688 & _T_6302; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_7852 = _T_6697 & _T_6302; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_7861 = _T_6562 & _T_6313; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_7870 = _T_6571 & _T_6313; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_7879 = _T_6580 & _T_6313; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_7888 = _T_6589 & _T_6313; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_7897 = _T_6598 & _T_6313; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_7906 = _T_6607 & _T_6313; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_7915 = _T_6616 & _T_6313; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_7924 = _T_6625 & _T_6313; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_7933 = _T_6634 & _T_6313; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_7942 = _T_6643 & _T_6313; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_7951 = _T_6652 & _T_6313; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_7960 = _T_6661 & _T_6313; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_7969 = _T_6670 & _T_6313; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_7978 = _T_6679 & _T_6313; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_7987 = _T_6688 & _T_6313; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_7996 = _T_6697 & _T_6313; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_8005 = _T_6562 & _T_6324; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_8014 = _T_6571 & _T_6324; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_8023 = _T_6580 & _T_6324; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_8032 = _T_6589 & _T_6324; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_8041 = _T_6598 & _T_6324; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_8050 = _T_6607 & _T_6324; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_8059 = _T_6616 & _T_6324; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_8068 = _T_6625 & _T_6324; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_8077 = _T_6634 & _T_6324; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_8086 = _T_6643 & _T_6324; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_8095 = _T_6652 & _T_6324; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_8104 = _T_6661 & _T_6324; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_8113 = _T_6670 & _T_6324; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_8122 = _T_6679 & _T_6324; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_8131 = _T_6688 & _T_6324; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_8140 = _T_6697 & _T_6324; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_8149 = _T_6562 & _T_6335; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_8158 = _T_6571 & _T_6335; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_8167 = _T_6580 & _T_6335; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_8176 = _T_6589 & _T_6335; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_8185 = _T_6598 & _T_6335; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_8194 = _T_6607 & _T_6335; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_8203 = _T_6616 & _T_6335; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_8212 = _T_6625 & _T_6335; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_8221 = _T_6634 & _T_6335; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_8230 = _T_6643 & _T_6335; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_8239 = _T_6652 & _T_6335; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_8248 = _T_6661 & _T_6335; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_8257 = _T_6670 & _T_6335; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_8266 = _T_6679 & _T_6335; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_8275 = _T_6688 & _T_6335; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_8284 = _T_6697 & _T_6335; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_8293 = _T_6562 & _T_6346; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_8302 = _T_6571 & _T_6346; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_8311 = _T_6580 & _T_6346; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_8320 = _T_6589 & _T_6346; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_8329 = _T_6598 & _T_6346; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_8338 = _T_6607 & _T_6346; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_8347 = _T_6616 & _T_6346; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_8356 = _T_6625 & _T_6346; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_8365 = _T_6634 & _T_6346; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_8374 = _T_6643 & _T_6346; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_8383 = _T_6652 & _T_6346; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_8392 = _T_6661 & _T_6346; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_8401 = _T_6670 & _T_6346; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_8410 = _T_6679 & _T_6346; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_8419 = _T_6688 & _T_6346; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_8428 = _T_6697 & _T_6346; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_8437 = _T_6562 & _T_6357; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_8446 = _T_6571 & _T_6357; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_8455 = _T_6580 & _T_6357; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_8464 = _T_6589 & _T_6357; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_8473 = _T_6598 & _T_6357; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_8482 = _T_6607 & _T_6357; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_8491 = _T_6616 & _T_6357; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_8500 = _T_6625 & _T_6357; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_8509 = _T_6634 & _T_6357; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_8518 = _T_6643 & _T_6357; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_8527 = _T_6652 & _T_6357; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_8536 = _T_6661 & _T_6357; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_8545 = _T_6670 & _T_6357; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_8554 = _T_6679 & _T_6357; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_8563 = _T_6688 & _T_6357; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_8572 = _T_6697 & _T_6357; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_8581 = _T_6562 & _T_6368; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_8590 = _T_6571 & _T_6368; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_8599 = _T_6580 & _T_6368; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_8608 = _T_6589 & _T_6368; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_8617 = _T_6598 & _T_6368; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_8626 = _T_6607 & _T_6368; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_8635 = _T_6616 & _T_6368; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_8644 = _T_6625 & _T_6368; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_8653 = _T_6634 & _T_6368; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_8662 = _T_6643 & _T_6368; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_8671 = _T_6652 & _T_6368; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_8680 = _T_6661 & _T_6368; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_8689 = _T_6670 & _T_6368; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_8698 = _T_6679 & _T_6368; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_8707 = _T_6688 & _T_6368; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_8716 = _T_6697 & _T_6368; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_8725 = _T_6562 & _T_6379; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_8734 = _T_6571 & _T_6379; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_8743 = _T_6580 & _T_6379; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_8752 = _T_6589 & _T_6379; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_8761 = _T_6598 & _T_6379; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_8770 = _T_6607 & _T_6379; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_8779 = _T_6616 & _T_6379; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_8788 = _T_6625 & _T_6379; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_8797 = _T_6634 & _T_6379; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_8806 = _T_6643 & _T_6379; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_8815 = _T_6652 & _T_6379; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_8824 = _T_6661 & _T_6379; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_8833 = _T_6670 & _T_6379; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_8842 = _T_6679 & _T_6379; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_8851 = _T_6688 & _T_6379; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_8860 = _T_6697 & _T_6379; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_8866 = bht_wr_en2[1] & _T_6561; // @[el2_ifu_bp_ctl.scala 447:23]
  wire  _T_8869 = _T_8866 & _T_6214; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_8875 = bht_wr_en2[1] & _T_6570; // @[el2_ifu_bp_ctl.scala 447:23]
  wire  _T_8878 = _T_8875 & _T_6214; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_8884 = bht_wr_en2[1] & _T_6579; // @[el2_ifu_bp_ctl.scala 447:23]
  wire  _T_8887 = _T_8884 & _T_6214; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_8893 = bht_wr_en2[1] & _T_6588; // @[el2_ifu_bp_ctl.scala 447:23]
  wire  _T_8896 = _T_8893 & _T_6214; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_8902 = bht_wr_en2[1] & _T_6597; // @[el2_ifu_bp_ctl.scala 447:23]
  wire  _T_8905 = _T_8902 & _T_6214; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_8911 = bht_wr_en2[1] & _T_6606; // @[el2_ifu_bp_ctl.scala 447:23]
  wire  _T_8914 = _T_8911 & _T_6214; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_8920 = bht_wr_en2[1] & _T_6615; // @[el2_ifu_bp_ctl.scala 447:23]
  wire  _T_8923 = _T_8920 & _T_6214; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_8929 = bht_wr_en2[1] & _T_6624; // @[el2_ifu_bp_ctl.scala 447:23]
  wire  _T_8932 = _T_8929 & _T_6214; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_8938 = bht_wr_en2[1] & _T_6633; // @[el2_ifu_bp_ctl.scala 447:23]
  wire  _T_8941 = _T_8938 & _T_6214; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_8947 = bht_wr_en2[1] & _T_6642; // @[el2_ifu_bp_ctl.scala 447:23]
  wire  _T_8950 = _T_8947 & _T_6214; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_8956 = bht_wr_en2[1] & _T_6651; // @[el2_ifu_bp_ctl.scala 447:23]
  wire  _T_8959 = _T_8956 & _T_6214; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_8965 = bht_wr_en2[1] & _T_6660; // @[el2_ifu_bp_ctl.scala 447:23]
  wire  _T_8968 = _T_8965 & _T_6214; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_8974 = bht_wr_en2[1] & _T_6669; // @[el2_ifu_bp_ctl.scala 447:23]
  wire  _T_8977 = _T_8974 & _T_6214; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_8983 = bht_wr_en2[1] & _T_6678; // @[el2_ifu_bp_ctl.scala 447:23]
  wire  _T_8986 = _T_8983 & _T_6214; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_8992 = bht_wr_en2[1] & _T_6687; // @[el2_ifu_bp_ctl.scala 447:23]
  wire  _T_8995 = _T_8992 & _T_6214; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_9001 = bht_wr_en2[1] & _T_6696; // @[el2_ifu_bp_ctl.scala 447:23]
  wire  _T_9004 = _T_9001 & _T_6214; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_9013 = _T_8866 & _T_6225; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_9022 = _T_8875 & _T_6225; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_9031 = _T_8884 & _T_6225; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_9040 = _T_8893 & _T_6225; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_9049 = _T_8902 & _T_6225; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_9058 = _T_8911 & _T_6225; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_9067 = _T_8920 & _T_6225; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_9076 = _T_8929 & _T_6225; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_9085 = _T_8938 & _T_6225; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_9094 = _T_8947 & _T_6225; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_9103 = _T_8956 & _T_6225; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_9112 = _T_8965 & _T_6225; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_9121 = _T_8974 & _T_6225; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_9130 = _T_8983 & _T_6225; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_9139 = _T_8992 & _T_6225; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_9148 = _T_9001 & _T_6225; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_9157 = _T_8866 & _T_6236; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_9166 = _T_8875 & _T_6236; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_9175 = _T_8884 & _T_6236; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_9184 = _T_8893 & _T_6236; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_9193 = _T_8902 & _T_6236; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_9202 = _T_8911 & _T_6236; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_9211 = _T_8920 & _T_6236; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_9220 = _T_8929 & _T_6236; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_9229 = _T_8938 & _T_6236; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_9238 = _T_8947 & _T_6236; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_9247 = _T_8956 & _T_6236; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_9256 = _T_8965 & _T_6236; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_9265 = _T_8974 & _T_6236; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_9274 = _T_8983 & _T_6236; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_9283 = _T_8992 & _T_6236; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_9292 = _T_9001 & _T_6236; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_9301 = _T_8866 & _T_6247; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_9310 = _T_8875 & _T_6247; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_9319 = _T_8884 & _T_6247; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_9328 = _T_8893 & _T_6247; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_9337 = _T_8902 & _T_6247; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_9346 = _T_8911 & _T_6247; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_9355 = _T_8920 & _T_6247; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_9364 = _T_8929 & _T_6247; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_9373 = _T_8938 & _T_6247; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_9382 = _T_8947 & _T_6247; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_9391 = _T_8956 & _T_6247; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_9400 = _T_8965 & _T_6247; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_9409 = _T_8974 & _T_6247; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_9418 = _T_8983 & _T_6247; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_9427 = _T_8992 & _T_6247; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_9436 = _T_9001 & _T_6247; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_9445 = _T_8866 & _T_6258; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_9454 = _T_8875 & _T_6258; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_9463 = _T_8884 & _T_6258; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_9472 = _T_8893 & _T_6258; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_9481 = _T_8902 & _T_6258; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_9490 = _T_8911 & _T_6258; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_9499 = _T_8920 & _T_6258; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_9508 = _T_8929 & _T_6258; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_9517 = _T_8938 & _T_6258; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_9526 = _T_8947 & _T_6258; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_9535 = _T_8956 & _T_6258; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_9544 = _T_8965 & _T_6258; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_9553 = _T_8974 & _T_6258; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_9562 = _T_8983 & _T_6258; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_9571 = _T_8992 & _T_6258; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_9580 = _T_9001 & _T_6258; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_9589 = _T_8866 & _T_6269; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_9598 = _T_8875 & _T_6269; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_9607 = _T_8884 & _T_6269; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_9616 = _T_8893 & _T_6269; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_9625 = _T_8902 & _T_6269; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_9634 = _T_8911 & _T_6269; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_9643 = _T_8920 & _T_6269; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_9652 = _T_8929 & _T_6269; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_9661 = _T_8938 & _T_6269; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_9670 = _T_8947 & _T_6269; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_9679 = _T_8956 & _T_6269; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_9688 = _T_8965 & _T_6269; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_9697 = _T_8974 & _T_6269; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_9706 = _T_8983 & _T_6269; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_9715 = _T_8992 & _T_6269; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_9724 = _T_9001 & _T_6269; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_9733 = _T_8866 & _T_6280; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_9742 = _T_8875 & _T_6280; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_9751 = _T_8884 & _T_6280; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_9760 = _T_8893 & _T_6280; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_9769 = _T_8902 & _T_6280; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_9778 = _T_8911 & _T_6280; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_9787 = _T_8920 & _T_6280; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_9796 = _T_8929 & _T_6280; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_9805 = _T_8938 & _T_6280; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_9814 = _T_8947 & _T_6280; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_9823 = _T_8956 & _T_6280; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_9832 = _T_8965 & _T_6280; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_9841 = _T_8974 & _T_6280; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_9850 = _T_8983 & _T_6280; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_9859 = _T_8992 & _T_6280; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_9868 = _T_9001 & _T_6280; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_9877 = _T_8866 & _T_6291; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_9886 = _T_8875 & _T_6291; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_9895 = _T_8884 & _T_6291; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_9904 = _T_8893 & _T_6291; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_9913 = _T_8902 & _T_6291; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_9922 = _T_8911 & _T_6291; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_9931 = _T_8920 & _T_6291; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_9940 = _T_8929 & _T_6291; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_9949 = _T_8938 & _T_6291; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_9958 = _T_8947 & _T_6291; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_9967 = _T_8956 & _T_6291; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_9976 = _T_8965 & _T_6291; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_9985 = _T_8974 & _T_6291; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_9994 = _T_8983 & _T_6291; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_10003 = _T_8992 & _T_6291; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_10012 = _T_9001 & _T_6291; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_10021 = _T_8866 & _T_6302; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_10030 = _T_8875 & _T_6302; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_10039 = _T_8884 & _T_6302; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_10048 = _T_8893 & _T_6302; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_10057 = _T_8902 & _T_6302; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_10066 = _T_8911 & _T_6302; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_10075 = _T_8920 & _T_6302; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_10084 = _T_8929 & _T_6302; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_10093 = _T_8938 & _T_6302; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_10102 = _T_8947 & _T_6302; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_10111 = _T_8956 & _T_6302; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_10120 = _T_8965 & _T_6302; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_10129 = _T_8974 & _T_6302; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_10138 = _T_8983 & _T_6302; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_10147 = _T_8992 & _T_6302; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_10156 = _T_9001 & _T_6302; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_10165 = _T_8866 & _T_6313; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_10174 = _T_8875 & _T_6313; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_10183 = _T_8884 & _T_6313; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_10192 = _T_8893 & _T_6313; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_10201 = _T_8902 & _T_6313; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_10210 = _T_8911 & _T_6313; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_10219 = _T_8920 & _T_6313; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_10228 = _T_8929 & _T_6313; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_10237 = _T_8938 & _T_6313; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_10246 = _T_8947 & _T_6313; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_10255 = _T_8956 & _T_6313; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_10264 = _T_8965 & _T_6313; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_10273 = _T_8974 & _T_6313; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_10282 = _T_8983 & _T_6313; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_10291 = _T_8992 & _T_6313; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_10300 = _T_9001 & _T_6313; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_10309 = _T_8866 & _T_6324; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_10318 = _T_8875 & _T_6324; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_10327 = _T_8884 & _T_6324; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_10336 = _T_8893 & _T_6324; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_10345 = _T_8902 & _T_6324; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_10354 = _T_8911 & _T_6324; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_10363 = _T_8920 & _T_6324; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_10372 = _T_8929 & _T_6324; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_10381 = _T_8938 & _T_6324; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_10390 = _T_8947 & _T_6324; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_10399 = _T_8956 & _T_6324; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_10408 = _T_8965 & _T_6324; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_10417 = _T_8974 & _T_6324; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_10426 = _T_8983 & _T_6324; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_10435 = _T_8992 & _T_6324; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_10444 = _T_9001 & _T_6324; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_10453 = _T_8866 & _T_6335; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_10462 = _T_8875 & _T_6335; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_10471 = _T_8884 & _T_6335; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_10480 = _T_8893 & _T_6335; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_10489 = _T_8902 & _T_6335; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_10498 = _T_8911 & _T_6335; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_10507 = _T_8920 & _T_6335; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_10516 = _T_8929 & _T_6335; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_10525 = _T_8938 & _T_6335; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_10534 = _T_8947 & _T_6335; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_10543 = _T_8956 & _T_6335; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_10552 = _T_8965 & _T_6335; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_10561 = _T_8974 & _T_6335; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_10570 = _T_8983 & _T_6335; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_10579 = _T_8992 & _T_6335; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_10588 = _T_9001 & _T_6335; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_10597 = _T_8866 & _T_6346; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_10606 = _T_8875 & _T_6346; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_10615 = _T_8884 & _T_6346; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_10624 = _T_8893 & _T_6346; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_10633 = _T_8902 & _T_6346; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_10642 = _T_8911 & _T_6346; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_10651 = _T_8920 & _T_6346; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_10660 = _T_8929 & _T_6346; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_10669 = _T_8938 & _T_6346; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_10678 = _T_8947 & _T_6346; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_10687 = _T_8956 & _T_6346; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_10696 = _T_8965 & _T_6346; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_10705 = _T_8974 & _T_6346; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_10714 = _T_8983 & _T_6346; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_10723 = _T_8992 & _T_6346; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_10732 = _T_9001 & _T_6346; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_10741 = _T_8866 & _T_6357; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_10750 = _T_8875 & _T_6357; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_10759 = _T_8884 & _T_6357; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_10768 = _T_8893 & _T_6357; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_10777 = _T_8902 & _T_6357; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_10786 = _T_8911 & _T_6357; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_10795 = _T_8920 & _T_6357; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_10804 = _T_8929 & _T_6357; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_10813 = _T_8938 & _T_6357; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_10822 = _T_8947 & _T_6357; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_10831 = _T_8956 & _T_6357; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_10840 = _T_8965 & _T_6357; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_10849 = _T_8974 & _T_6357; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_10858 = _T_8983 & _T_6357; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_10867 = _T_8992 & _T_6357; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_10876 = _T_9001 & _T_6357; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_10885 = _T_8866 & _T_6368; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_10894 = _T_8875 & _T_6368; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_10903 = _T_8884 & _T_6368; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_10912 = _T_8893 & _T_6368; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_10921 = _T_8902 & _T_6368; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_10930 = _T_8911 & _T_6368; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_10939 = _T_8920 & _T_6368; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_10948 = _T_8929 & _T_6368; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_10957 = _T_8938 & _T_6368; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_10966 = _T_8947 & _T_6368; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_10975 = _T_8956 & _T_6368; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_10984 = _T_8965 & _T_6368; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_10993 = _T_8974 & _T_6368; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_11002 = _T_8983 & _T_6368; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_11011 = _T_8992 & _T_6368; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_11020 = _T_9001 & _T_6368; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_11029 = _T_8866 & _T_6379; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_11038 = _T_8875 & _T_6379; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_11047 = _T_8884 & _T_6379; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_11056 = _T_8893 & _T_6379; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_11065 = _T_8902 & _T_6379; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_11074 = _T_8911 & _T_6379; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_11083 = _T_8920 & _T_6379; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_11092 = _T_8929 & _T_6379; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_11101 = _T_8938 & _T_6379; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_11110 = _T_8947 & _T_6379; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_11119 = _T_8956 & _T_6379; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_11128 = _T_8965 & _T_6379; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_11137 = _T_8974 & _T_6379; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_11146 = _T_8983 & _T_6379; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_11155 = _T_8992 & _T_6379; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_11164 = _T_9001 & _T_6379; // @[el2_ifu_bp_ctl.scala 447:81]
  wire  _T_11169 = mp_hashed[3:0] == 4'h0; // @[el2_ifu_bp_ctl.scala 455:97]
  wire  _T_11170 = bht_wr_en0[0] & _T_11169; // @[el2_ifu_bp_ctl.scala 455:45]
  wire  _T_11174 = _T_11170 & _T_6209; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_0_0 = _T_11174 | _T_6565; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_11186 = mp_hashed[3:0] == 4'h1; // @[el2_ifu_bp_ctl.scala 455:97]
  wire  _T_11187 = bht_wr_en0[0] & _T_11186; // @[el2_ifu_bp_ctl.scala 455:45]
  wire  _T_11191 = _T_11187 & _T_6209; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_0_1 = _T_11191 | _T_6574; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_11203 = mp_hashed[3:0] == 4'h2; // @[el2_ifu_bp_ctl.scala 455:97]
  wire  _T_11204 = bht_wr_en0[0] & _T_11203; // @[el2_ifu_bp_ctl.scala 455:45]
  wire  _T_11208 = _T_11204 & _T_6209; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_0_2 = _T_11208 | _T_6583; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_11220 = mp_hashed[3:0] == 4'h3; // @[el2_ifu_bp_ctl.scala 455:97]
  wire  _T_11221 = bht_wr_en0[0] & _T_11220; // @[el2_ifu_bp_ctl.scala 455:45]
  wire  _T_11225 = _T_11221 & _T_6209; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_0_3 = _T_11225 | _T_6592; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_11237 = mp_hashed[3:0] == 4'h4; // @[el2_ifu_bp_ctl.scala 455:97]
  wire  _T_11238 = bht_wr_en0[0] & _T_11237; // @[el2_ifu_bp_ctl.scala 455:45]
  wire  _T_11242 = _T_11238 & _T_6209; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_0_4 = _T_11242 | _T_6601; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_11254 = mp_hashed[3:0] == 4'h5; // @[el2_ifu_bp_ctl.scala 455:97]
  wire  _T_11255 = bht_wr_en0[0] & _T_11254; // @[el2_ifu_bp_ctl.scala 455:45]
  wire  _T_11259 = _T_11255 & _T_6209; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_0_5 = _T_11259 | _T_6610; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_11271 = mp_hashed[3:0] == 4'h6; // @[el2_ifu_bp_ctl.scala 455:97]
  wire  _T_11272 = bht_wr_en0[0] & _T_11271; // @[el2_ifu_bp_ctl.scala 455:45]
  wire  _T_11276 = _T_11272 & _T_6209; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_0_6 = _T_11276 | _T_6619; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_11288 = mp_hashed[3:0] == 4'h7; // @[el2_ifu_bp_ctl.scala 455:97]
  wire  _T_11289 = bht_wr_en0[0] & _T_11288; // @[el2_ifu_bp_ctl.scala 455:45]
  wire  _T_11293 = _T_11289 & _T_6209; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_0_7 = _T_11293 | _T_6628; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_11305 = mp_hashed[3:0] == 4'h8; // @[el2_ifu_bp_ctl.scala 455:97]
  wire  _T_11306 = bht_wr_en0[0] & _T_11305; // @[el2_ifu_bp_ctl.scala 455:45]
  wire  _T_11310 = _T_11306 & _T_6209; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_0_8 = _T_11310 | _T_6637; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_11322 = mp_hashed[3:0] == 4'h9; // @[el2_ifu_bp_ctl.scala 455:97]
  wire  _T_11323 = bht_wr_en0[0] & _T_11322; // @[el2_ifu_bp_ctl.scala 455:45]
  wire  _T_11327 = _T_11323 & _T_6209; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_0_9 = _T_11327 | _T_6646; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_11339 = mp_hashed[3:0] == 4'ha; // @[el2_ifu_bp_ctl.scala 455:97]
  wire  _T_11340 = bht_wr_en0[0] & _T_11339; // @[el2_ifu_bp_ctl.scala 455:45]
  wire  _T_11344 = _T_11340 & _T_6209; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_0_10 = _T_11344 | _T_6655; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_11356 = mp_hashed[3:0] == 4'hb; // @[el2_ifu_bp_ctl.scala 455:97]
  wire  _T_11357 = bht_wr_en0[0] & _T_11356; // @[el2_ifu_bp_ctl.scala 455:45]
  wire  _T_11361 = _T_11357 & _T_6209; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_0_11 = _T_11361 | _T_6664; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_11373 = mp_hashed[3:0] == 4'hc; // @[el2_ifu_bp_ctl.scala 455:97]
  wire  _T_11374 = bht_wr_en0[0] & _T_11373; // @[el2_ifu_bp_ctl.scala 455:45]
  wire  _T_11378 = _T_11374 & _T_6209; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_0_12 = _T_11378 | _T_6673; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_11390 = mp_hashed[3:0] == 4'hd; // @[el2_ifu_bp_ctl.scala 455:97]
  wire  _T_11391 = bht_wr_en0[0] & _T_11390; // @[el2_ifu_bp_ctl.scala 455:45]
  wire  _T_11395 = _T_11391 & _T_6209; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_0_13 = _T_11395 | _T_6682; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_11407 = mp_hashed[3:0] == 4'he; // @[el2_ifu_bp_ctl.scala 455:97]
  wire  _T_11408 = bht_wr_en0[0] & _T_11407; // @[el2_ifu_bp_ctl.scala 455:45]
  wire  _T_11412 = _T_11408 & _T_6209; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_0_14 = _T_11412 | _T_6691; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_11424 = mp_hashed[3:0] == 4'hf; // @[el2_ifu_bp_ctl.scala 455:97]
  wire  _T_11425 = bht_wr_en0[0] & _T_11424; // @[el2_ifu_bp_ctl.scala 455:45]
  wire  _T_11429 = _T_11425 & _T_6209; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_0_15 = _T_11429 | _T_6700; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_11446 = _T_11170 & _T_6220; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_1_0 = _T_11446 | _T_6709; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_11463 = _T_11187 & _T_6220; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_1_1 = _T_11463 | _T_6718; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_11480 = _T_11204 & _T_6220; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_1_2 = _T_11480 | _T_6727; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_11497 = _T_11221 & _T_6220; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_1_3 = _T_11497 | _T_6736; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_11514 = _T_11238 & _T_6220; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_1_4 = _T_11514 | _T_6745; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_11531 = _T_11255 & _T_6220; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_1_5 = _T_11531 | _T_6754; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_11548 = _T_11272 & _T_6220; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_1_6 = _T_11548 | _T_6763; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_11565 = _T_11289 & _T_6220; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_1_7 = _T_11565 | _T_6772; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_11582 = _T_11306 & _T_6220; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_1_8 = _T_11582 | _T_6781; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_11599 = _T_11323 & _T_6220; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_1_9 = _T_11599 | _T_6790; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_11616 = _T_11340 & _T_6220; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_1_10 = _T_11616 | _T_6799; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_11633 = _T_11357 & _T_6220; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_1_11 = _T_11633 | _T_6808; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_11650 = _T_11374 & _T_6220; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_1_12 = _T_11650 | _T_6817; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_11667 = _T_11391 & _T_6220; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_1_13 = _T_11667 | _T_6826; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_11684 = _T_11408 & _T_6220; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_1_14 = _T_11684 | _T_6835; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_11701 = _T_11425 & _T_6220; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_1_15 = _T_11701 | _T_6844; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_11718 = _T_11170 & _T_6231; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_2_0 = _T_11718 | _T_6853; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_11735 = _T_11187 & _T_6231; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_2_1 = _T_11735 | _T_6862; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_11752 = _T_11204 & _T_6231; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_2_2 = _T_11752 | _T_6871; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_11769 = _T_11221 & _T_6231; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_2_3 = _T_11769 | _T_6880; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_11786 = _T_11238 & _T_6231; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_2_4 = _T_11786 | _T_6889; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_11803 = _T_11255 & _T_6231; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_2_5 = _T_11803 | _T_6898; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_11820 = _T_11272 & _T_6231; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_2_6 = _T_11820 | _T_6907; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_11837 = _T_11289 & _T_6231; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_2_7 = _T_11837 | _T_6916; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_11854 = _T_11306 & _T_6231; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_2_8 = _T_11854 | _T_6925; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_11871 = _T_11323 & _T_6231; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_2_9 = _T_11871 | _T_6934; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_11888 = _T_11340 & _T_6231; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_2_10 = _T_11888 | _T_6943; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_11905 = _T_11357 & _T_6231; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_2_11 = _T_11905 | _T_6952; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_11922 = _T_11374 & _T_6231; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_2_12 = _T_11922 | _T_6961; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_11939 = _T_11391 & _T_6231; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_2_13 = _T_11939 | _T_6970; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_11956 = _T_11408 & _T_6231; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_2_14 = _T_11956 | _T_6979; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_11973 = _T_11425 & _T_6231; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_2_15 = _T_11973 | _T_6988; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_11990 = _T_11170 & _T_6242; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_3_0 = _T_11990 | _T_6997; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_12007 = _T_11187 & _T_6242; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_3_1 = _T_12007 | _T_7006; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_12024 = _T_11204 & _T_6242; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_3_2 = _T_12024 | _T_7015; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_12041 = _T_11221 & _T_6242; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_3_3 = _T_12041 | _T_7024; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_12058 = _T_11238 & _T_6242; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_3_4 = _T_12058 | _T_7033; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_12075 = _T_11255 & _T_6242; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_3_5 = _T_12075 | _T_7042; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_12092 = _T_11272 & _T_6242; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_3_6 = _T_12092 | _T_7051; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_12109 = _T_11289 & _T_6242; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_3_7 = _T_12109 | _T_7060; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_12126 = _T_11306 & _T_6242; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_3_8 = _T_12126 | _T_7069; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_12143 = _T_11323 & _T_6242; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_3_9 = _T_12143 | _T_7078; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_12160 = _T_11340 & _T_6242; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_3_10 = _T_12160 | _T_7087; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_12177 = _T_11357 & _T_6242; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_3_11 = _T_12177 | _T_7096; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_12194 = _T_11374 & _T_6242; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_3_12 = _T_12194 | _T_7105; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_12211 = _T_11391 & _T_6242; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_3_13 = _T_12211 | _T_7114; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_12228 = _T_11408 & _T_6242; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_3_14 = _T_12228 | _T_7123; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_12245 = _T_11425 & _T_6242; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_3_15 = _T_12245 | _T_7132; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_12262 = _T_11170 & _T_6253; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_4_0 = _T_12262 | _T_7141; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_12279 = _T_11187 & _T_6253; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_4_1 = _T_12279 | _T_7150; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_12296 = _T_11204 & _T_6253; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_4_2 = _T_12296 | _T_7159; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_12313 = _T_11221 & _T_6253; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_4_3 = _T_12313 | _T_7168; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_12330 = _T_11238 & _T_6253; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_4_4 = _T_12330 | _T_7177; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_12347 = _T_11255 & _T_6253; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_4_5 = _T_12347 | _T_7186; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_12364 = _T_11272 & _T_6253; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_4_6 = _T_12364 | _T_7195; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_12381 = _T_11289 & _T_6253; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_4_7 = _T_12381 | _T_7204; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_12398 = _T_11306 & _T_6253; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_4_8 = _T_12398 | _T_7213; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_12415 = _T_11323 & _T_6253; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_4_9 = _T_12415 | _T_7222; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_12432 = _T_11340 & _T_6253; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_4_10 = _T_12432 | _T_7231; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_12449 = _T_11357 & _T_6253; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_4_11 = _T_12449 | _T_7240; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_12466 = _T_11374 & _T_6253; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_4_12 = _T_12466 | _T_7249; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_12483 = _T_11391 & _T_6253; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_4_13 = _T_12483 | _T_7258; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_12500 = _T_11408 & _T_6253; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_4_14 = _T_12500 | _T_7267; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_12517 = _T_11425 & _T_6253; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_4_15 = _T_12517 | _T_7276; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_12534 = _T_11170 & _T_6264; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_5_0 = _T_12534 | _T_7285; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_12551 = _T_11187 & _T_6264; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_5_1 = _T_12551 | _T_7294; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_12568 = _T_11204 & _T_6264; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_5_2 = _T_12568 | _T_7303; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_12585 = _T_11221 & _T_6264; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_5_3 = _T_12585 | _T_7312; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_12602 = _T_11238 & _T_6264; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_5_4 = _T_12602 | _T_7321; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_12619 = _T_11255 & _T_6264; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_5_5 = _T_12619 | _T_7330; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_12636 = _T_11272 & _T_6264; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_5_6 = _T_12636 | _T_7339; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_12653 = _T_11289 & _T_6264; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_5_7 = _T_12653 | _T_7348; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_12670 = _T_11306 & _T_6264; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_5_8 = _T_12670 | _T_7357; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_12687 = _T_11323 & _T_6264; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_5_9 = _T_12687 | _T_7366; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_12704 = _T_11340 & _T_6264; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_5_10 = _T_12704 | _T_7375; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_12721 = _T_11357 & _T_6264; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_5_11 = _T_12721 | _T_7384; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_12738 = _T_11374 & _T_6264; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_5_12 = _T_12738 | _T_7393; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_12755 = _T_11391 & _T_6264; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_5_13 = _T_12755 | _T_7402; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_12772 = _T_11408 & _T_6264; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_5_14 = _T_12772 | _T_7411; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_12789 = _T_11425 & _T_6264; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_5_15 = _T_12789 | _T_7420; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_12806 = _T_11170 & _T_6275; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_6_0 = _T_12806 | _T_7429; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_12823 = _T_11187 & _T_6275; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_6_1 = _T_12823 | _T_7438; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_12840 = _T_11204 & _T_6275; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_6_2 = _T_12840 | _T_7447; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_12857 = _T_11221 & _T_6275; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_6_3 = _T_12857 | _T_7456; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_12874 = _T_11238 & _T_6275; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_6_4 = _T_12874 | _T_7465; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_12891 = _T_11255 & _T_6275; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_6_5 = _T_12891 | _T_7474; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_12908 = _T_11272 & _T_6275; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_6_6 = _T_12908 | _T_7483; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_12925 = _T_11289 & _T_6275; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_6_7 = _T_12925 | _T_7492; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_12942 = _T_11306 & _T_6275; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_6_8 = _T_12942 | _T_7501; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_12959 = _T_11323 & _T_6275; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_6_9 = _T_12959 | _T_7510; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_12976 = _T_11340 & _T_6275; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_6_10 = _T_12976 | _T_7519; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_12993 = _T_11357 & _T_6275; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_6_11 = _T_12993 | _T_7528; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_13010 = _T_11374 & _T_6275; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_6_12 = _T_13010 | _T_7537; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_13027 = _T_11391 & _T_6275; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_6_13 = _T_13027 | _T_7546; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_13044 = _T_11408 & _T_6275; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_6_14 = _T_13044 | _T_7555; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_13061 = _T_11425 & _T_6275; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_6_15 = _T_13061 | _T_7564; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_13078 = _T_11170 & _T_6286; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_7_0 = _T_13078 | _T_7573; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_13095 = _T_11187 & _T_6286; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_7_1 = _T_13095 | _T_7582; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_13112 = _T_11204 & _T_6286; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_7_2 = _T_13112 | _T_7591; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_13129 = _T_11221 & _T_6286; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_7_3 = _T_13129 | _T_7600; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_13146 = _T_11238 & _T_6286; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_7_4 = _T_13146 | _T_7609; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_13163 = _T_11255 & _T_6286; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_7_5 = _T_13163 | _T_7618; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_13180 = _T_11272 & _T_6286; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_7_6 = _T_13180 | _T_7627; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_13197 = _T_11289 & _T_6286; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_7_7 = _T_13197 | _T_7636; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_13214 = _T_11306 & _T_6286; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_7_8 = _T_13214 | _T_7645; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_13231 = _T_11323 & _T_6286; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_7_9 = _T_13231 | _T_7654; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_13248 = _T_11340 & _T_6286; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_7_10 = _T_13248 | _T_7663; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_13265 = _T_11357 & _T_6286; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_7_11 = _T_13265 | _T_7672; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_13282 = _T_11374 & _T_6286; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_7_12 = _T_13282 | _T_7681; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_13299 = _T_11391 & _T_6286; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_7_13 = _T_13299 | _T_7690; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_13316 = _T_11408 & _T_6286; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_7_14 = _T_13316 | _T_7699; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_13333 = _T_11425 & _T_6286; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_7_15 = _T_13333 | _T_7708; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_13350 = _T_11170 & _T_6297; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_8_0 = _T_13350 | _T_7717; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_13367 = _T_11187 & _T_6297; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_8_1 = _T_13367 | _T_7726; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_13384 = _T_11204 & _T_6297; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_8_2 = _T_13384 | _T_7735; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_13401 = _T_11221 & _T_6297; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_8_3 = _T_13401 | _T_7744; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_13418 = _T_11238 & _T_6297; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_8_4 = _T_13418 | _T_7753; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_13435 = _T_11255 & _T_6297; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_8_5 = _T_13435 | _T_7762; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_13452 = _T_11272 & _T_6297; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_8_6 = _T_13452 | _T_7771; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_13469 = _T_11289 & _T_6297; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_8_7 = _T_13469 | _T_7780; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_13486 = _T_11306 & _T_6297; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_8_8 = _T_13486 | _T_7789; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_13503 = _T_11323 & _T_6297; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_8_9 = _T_13503 | _T_7798; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_13520 = _T_11340 & _T_6297; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_8_10 = _T_13520 | _T_7807; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_13537 = _T_11357 & _T_6297; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_8_11 = _T_13537 | _T_7816; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_13554 = _T_11374 & _T_6297; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_8_12 = _T_13554 | _T_7825; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_13571 = _T_11391 & _T_6297; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_8_13 = _T_13571 | _T_7834; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_13588 = _T_11408 & _T_6297; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_8_14 = _T_13588 | _T_7843; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_13605 = _T_11425 & _T_6297; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_8_15 = _T_13605 | _T_7852; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_13622 = _T_11170 & _T_6308; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_9_0 = _T_13622 | _T_7861; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_13639 = _T_11187 & _T_6308; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_9_1 = _T_13639 | _T_7870; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_13656 = _T_11204 & _T_6308; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_9_2 = _T_13656 | _T_7879; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_13673 = _T_11221 & _T_6308; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_9_3 = _T_13673 | _T_7888; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_13690 = _T_11238 & _T_6308; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_9_4 = _T_13690 | _T_7897; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_13707 = _T_11255 & _T_6308; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_9_5 = _T_13707 | _T_7906; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_13724 = _T_11272 & _T_6308; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_9_6 = _T_13724 | _T_7915; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_13741 = _T_11289 & _T_6308; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_9_7 = _T_13741 | _T_7924; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_13758 = _T_11306 & _T_6308; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_9_8 = _T_13758 | _T_7933; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_13775 = _T_11323 & _T_6308; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_9_9 = _T_13775 | _T_7942; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_13792 = _T_11340 & _T_6308; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_9_10 = _T_13792 | _T_7951; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_13809 = _T_11357 & _T_6308; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_9_11 = _T_13809 | _T_7960; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_13826 = _T_11374 & _T_6308; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_9_12 = _T_13826 | _T_7969; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_13843 = _T_11391 & _T_6308; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_9_13 = _T_13843 | _T_7978; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_13860 = _T_11408 & _T_6308; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_9_14 = _T_13860 | _T_7987; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_13877 = _T_11425 & _T_6308; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_9_15 = _T_13877 | _T_7996; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_13894 = _T_11170 & _T_6319; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_10_0 = _T_13894 | _T_8005; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_13911 = _T_11187 & _T_6319; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_10_1 = _T_13911 | _T_8014; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_13928 = _T_11204 & _T_6319; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_10_2 = _T_13928 | _T_8023; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_13945 = _T_11221 & _T_6319; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_10_3 = _T_13945 | _T_8032; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_13962 = _T_11238 & _T_6319; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_10_4 = _T_13962 | _T_8041; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_13979 = _T_11255 & _T_6319; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_10_5 = _T_13979 | _T_8050; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_13996 = _T_11272 & _T_6319; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_10_6 = _T_13996 | _T_8059; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_14013 = _T_11289 & _T_6319; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_10_7 = _T_14013 | _T_8068; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_14030 = _T_11306 & _T_6319; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_10_8 = _T_14030 | _T_8077; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_14047 = _T_11323 & _T_6319; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_10_9 = _T_14047 | _T_8086; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_14064 = _T_11340 & _T_6319; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_10_10 = _T_14064 | _T_8095; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_14081 = _T_11357 & _T_6319; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_10_11 = _T_14081 | _T_8104; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_14098 = _T_11374 & _T_6319; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_10_12 = _T_14098 | _T_8113; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_14115 = _T_11391 & _T_6319; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_10_13 = _T_14115 | _T_8122; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_14132 = _T_11408 & _T_6319; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_10_14 = _T_14132 | _T_8131; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_14149 = _T_11425 & _T_6319; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_10_15 = _T_14149 | _T_8140; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_14166 = _T_11170 & _T_6330; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_11_0 = _T_14166 | _T_8149; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_14183 = _T_11187 & _T_6330; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_11_1 = _T_14183 | _T_8158; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_14200 = _T_11204 & _T_6330; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_11_2 = _T_14200 | _T_8167; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_14217 = _T_11221 & _T_6330; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_11_3 = _T_14217 | _T_8176; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_14234 = _T_11238 & _T_6330; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_11_4 = _T_14234 | _T_8185; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_14251 = _T_11255 & _T_6330; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_11_5 = _T_14251 | _T_8194; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_14268 = _T_11272 & _T_6330; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_11_6 = _T_14268 | _T_8203; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_14285 = _T_11289 & _T_6330; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_11_7 = _T_14285 | _T_8212; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_14302 = _T_11306 & _T_6330; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_11_8 = _T_14302 | _T_8221; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_14319 = _T_11323 & _T_6330; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_11_9 = _T_14319 | _T_8230; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_14336 = _T_11340 & _T_6330; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_11_10 = _T_14336 | _T_8239; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_14353 = _T_11357 & _T_6330; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_11_11 = _T_14353 | _T_8248; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_14370 = _T_11374 & _T_6330; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_11_12 = _T_14370 | _T_8257; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_14387 = _T_11391 & _T_6330; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_11_13 = _T_14387 | _T_8266; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_14404 = _T_11408 & _T_6330; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_11_14 = _T_14404 | _T_8275; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_14421 = _T_11425 & _T_6330; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_11_15 = _T_14421 | _T_8284; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_14438 = _T_11170 & _T_6341; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_12_0 = _T_14438 | _T_8293; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_14455 = _T_11187 & _T_6341; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_12_1 = _T_14455 | _T_8302; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_14472 = _T_11204 & _T_6341; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_12_2 = _T_14472 | _T_8311; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_14489 = _T_11221 & _T_6341; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_12_3 = _T_14489 | _T_8320; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_14506 = _T_11238 & _T_6341; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_12_4 = _T_14506 | _T_8329; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_14523 = _T_11255 & _T_6341; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_12_5 = _T_14523 | _T_8338; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_14540 = _T_11272 & _T_6341; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_12_6 = _T_14540 | _T_8347; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_14557 = _T_11289 & _T_6341; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_12_7 = _T_14557 | _T_8356; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_14574 = _T_11306 & _T_6341; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_12_8 = _T_14574 | _T_8365; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_14591 = _T_11323 & _T_6341; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_12_9 = _T_14591 | _T_8374; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_14608 = _T_11340 & _T_6341; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_12_10 = _T_14608 | _T_8383; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_14625 = _T_11357 & _T_6341; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_12_11 = _T_14625 | _T_8392; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_14642 = _T_11374 & _T_6341; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_12_12 = _T_14642 | _T_8401; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_14659 = _T_11391 & _T_6341; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_12_13 = _T_14659 | _T_8410; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_14676 = _T_11408 & _T_6341; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_12_14 = _T_14676 | _T_8419; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_14693 = _T_11425 & _T_6341; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_12_15 = _T_14693 | _T_8428; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_14710 = _T_11170 & _T_6352; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_13_0 = _T_14710 | _T_8437; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_14727 = _T_11187 & _T_6352; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_13_1 = _T_14727 | _T_8446; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_14744 = _T_11204 & _T_6352; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_13_2 = _T_14744 | _T_8455; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_14761 = _T_11221 & _T_6352; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_13_3 = _T_14761 | _T_8464; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_14778 = _T_11238 & _T_6352; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_13_4 = _T_14778 | _T_8473; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_14795 = _T_11255 & _T_6352; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_13_5 = _T_14795 | _T_8482; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_14812 = _T_11272 & _T_6352; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_13_6 = _T_14812 | _T_8491; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_14829 = _T_11289 & _T_6352; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_13_7 = _T_14829 | _T_8500; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_14846 = _T_11306 & _T_6352; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_13_8 = _T_14846 | _T_8509; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_14863 = _T_11323 & _T_6352; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_13_9 = _T_14863 | _T_8518; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_14880 = _T_11340 & _T_6352; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_13_10 = _T_14880 | _T_8527; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_14897 = _T_11357 & _T_6352; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_13_11 = _T_14897 | _T_8536; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_14914 = _T_11374 & _T_6352; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_13_12 = _T_14914 | _T_8545; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_14931 = _T_11391 & _T_6352; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_13_13 = _T_14931 | _T_8554; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_14948 = _T_11408 & _T_6352; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_13_14 = _T_14948 | _T_8563; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_14965 = _T_11425 & _T_6352; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_13_15 = _T_14965 | _T_8572; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_14982 = _T_11170 & _T_6363; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_14_0 = _T_14982 | _T_8581; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_14999 = _T_11187 & _T_6363; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_14_1 = _T_14999 | _T_8590; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_15016 = _T_11204 & _T_6363; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_14_2 = _T_15016 | _T_8599; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_15033 = _T_11221 & _T_6363; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_14_3 = _T_15033 | _T_8608; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_15050 = _T_11238 & _T_6363; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_14_4 = _T_15050 | _T_8617; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_15067 = _T_11255 & _T_6363; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_14_5 = _T_15067 | _T_8626; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_15084 = _T_11272 & _T_6363; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_14_6 = _T_15084 | _T_8635; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_15101 = _T_11289 & _T_6363; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_14_7 = _T_15101 | _T_8644; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_15118 = _T_11306 & _T_6363; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_14_8 = _T_15118 | _T_8653; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_15135 = _T_11323 & _T_6363; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_14_9 = _T_15135 | _T_8662; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_15152 = _T_11340 & _T_6363; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_14_10 = _T_15152 | _T_8671; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_15169 = _T_11357 & _T_6363; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_14_11 = _T_15169 | _T_8680; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_15186 = _T_11374 & _T_6363; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_14_12 = _T_15186 | _T_8689; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_15203 = _T_11391 & _T_6363; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_14_13 = _T_15203 | _T_8698; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_15220 = _T_11408 & _T_6363; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_14_14 = _T_15220 | _T_8707; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_15237 = _T_11425 & _T_6363; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_14_15 = _T_15237 | _T_8716; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_15254 = _T_11170 & _T_6374; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_15_0 = _T_15254 | _T_8725; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_15271 = _T_11187 & _T_6374; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_15_1 = _T_15271 | _T_8734; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_15288 = _T_11204 & _T_6374; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_15_2 = _T_15288 | _T_8743; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_15305 = _T_11221 & _T_6374; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_15_3 = _T_15305 | _T_8752; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_15322 = _T_11238 & _T_6374; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_15_4 = _T_15322 | _T_8761; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_15339 = _T_11255 & _T_6374; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_15_5 = _T_15339 | _T_8770; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_15356 = _T_11272 & _T_6374; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_15_6 = _T_15356 | _T_8779; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_15373 = _T_11289 & _T_6374; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_15_7 = _T_15373 | _T_8788; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_15390 = _T_11306 & _T_6374; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_15_8 = _T_15390 | _T_8797; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_15407 = _T_11323 & _T_6374; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_15_9 = _T_15407 | _T_8806; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_15424 = _T_11340 & _T_6374; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_15_10 = _T_15424 | _T_8815; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_15441 = _T_11357 & _T_6374; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_15_11 = _T_15441 | _T_8824; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_15458 = _T_11374 & _T_6374; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_15_12 = _T_15458 | _T_8833; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_15475 = _T_11391 & _T_6374; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_15_13 = _T_15475 | _T_8842; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_15492 = _T_11408 & _T_6374; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_15_14 = _T_15492 | _T_8851; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_15509 = _T_11425 & _T_6374; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_0_15_15 = _T_15509 | _T_8860; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_15522 = bht_wr_en0[1] & _T_11169; // @[el2_ifu_bp_ctl.scala 455:45]
  wire  _T_15526 = _T_15522 & _T_6209; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_0_0 = _T_15526 | _T_8869; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_15539 = bht_wr_en0[1] & _T_11186; // @[el2_ifu_bp_ctl.scala 455:45]
  wire  _T_15543 = _T_15539 & _T_6209; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_0_1 = _T_15543 | _T_8878; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_15556 = bht_wr_en0[1] & _T_11203; // @[el2_ifu_bp_ctl.scala 455:45]
  wire  _T_15560 = _T_15556 & _T_6209; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_0_2 = _T_15560 | _T_8887; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_15573 = bht_wr_en0[1] & _T_11220; // @[el2_ifu_bp_ctl.scala 455:45]
  wire  _T_15577 = _T_15573 & _T_6209; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_0_3 = _T_15577 | _T_8896; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_15590 = bht_wr_en0[1] & _T_11237; // @[el2_ifu_bp_ctl.scala 455:45]
  wire  _T_15594 = _T_15590 & _T_6209; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_0_4 = _T_15594 | _T_8905; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_15607 = bht_wr_en0[1] & _T_11254; // @[el2_ifu_bp_ctl.scala 455:45]
  wire  _T_15611 = _T_15607 & _T_6209; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_0_5 = _T_15611 | _T_8914; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_15624 = bht_wr_en0[1] & _T_11271; // @[el2_ifu_bp_ctl.scala 455:45]
  wire  _T_15628 = _T_15624 & _T_6209; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_0_6 = _T_15628 | _T_8923; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_15641 = bht_wr_en0[1] & _T_11288; // @[el2_ifu_bp_ctl.scala 455:45]
  wire  _T_15645 = _T_15641 & _T_6209; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_0_7 = _T_15645 | _T_8932; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_15658 = bht_wr_en0[1] & _T_11305; // @[el2_ifu_bp_ctl.scala 455:45]
  wire  _T_15662 = _T_15658 & _T_6209; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_0_8 = _T_15662 | _T_8941; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_15675 = bht_wr_en0[1] & _T_11322; // @[el2_ifu_bp_ctl.scala 455:45]
  wire  _T_15679 = _T_15675 & _T_6209; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_0_9 = _T_15679 | _T_8950; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_15692 = bht_wr_en0[1] & _T_11339; // @[el2_ifu_bp_ctl.scala 455:45]
  wire  _T_15696 = _T_15692 & _T_6209; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_0_10 = _T_15696 | _T_8959; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_15709 = bht_wr_en0[1] & _T_11356; // @[el2_ifu_bp_ctl.scala 455:45]
  wire  _T_15713 = _T_15709 & _T_6209; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_0_11 = _T_15713 | _T_8968; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_15726 = bht_wr_en0[1] & _T_11373; // @[el2_ifu_bp_ctl.scala 455:45]
  wire  _T_15730 = _T_15726 & _T_6209; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_0_12 = _T_15730 | _T_8977; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_15743 = bht_wr_en0[1] & _T_11390; // @[el2_ifu_bp_ctl.scala 455:45]
  wire  _T_15747 = _T_15743 & _T_6209; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_0_13 = _T_15747 | _T_8986; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_15760 = bht_wr_en0[1] & _T_11407; // @[el2_ifu_bp_ctl.scala 455:45]
  wire  _T_15764 = _T_15760 & _T_6209; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_0_14 = _T_15764 | _T_8995; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_15777 = bht_wr_en0[1] & _T_11424; // @[el2_ifu_bp_ctl.scala 455:45]
  wire  _T_15781 = _T_15777 & _T_6209; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_0_15 = _T_15781 | _T_9004; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_15798 = _T_15522 & _T_6220; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_1_0 = _T_15798 | _T_9013; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_15815 = _T_15539 & _T_6220; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_1_1 = _T_15815 | _T_9022; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_15832 = _T_15556 & _T_6220; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_1_2 = _T_15832 | _T_9031; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_15849 = _T_15573 & _T_6220; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_1_3 = _T_15849 | _T_9040; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_15866 = _T_15590 & _T_6220; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_1_4 = _T_15866 | _T_9049; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_15883 = _T_15607 & _T_6220; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_1_5 = _T_15883 | _T_9058; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_15900 = _T_15624 & _T_6220; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_1_6 = _T_15900 | _T_9067; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_15917 = _T_15641 & _T_6220; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_1_7 = _T_15917 | _T_9076; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_15934 = _T_15658 & _T_6220; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_1_8 = _T_15934 | _T_9085; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_15951 = _T_15675 & _T_6220; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_1_9 = _T_15951 | _T_9094; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_15968 = _T_15692 & _T_6220; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_1_10 = _T_15968 | _T_9103; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_15985 = _T_15709 & _T_6220; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_1_11 = _T_15985 | _T_9112; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_16002 = _T_15726 & _T_6220; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_1_12 = _T_16002 | _T_9121; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_16019 = _T_15743 & _T_6220; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_1_13 = _T_16019 | _T_9130; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_16036 = _T_15760 & _T_6220; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_1_14 = _T_16036 | _T_9139; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_16053 = _T_15777 & _T_6220; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_1_15 = _T_16053 | _T_9148; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_16070 = _T_15522 & _T_6231; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_2_0 = _T_16070 | _T_9157; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_16087 = _T_15539 & _T_6231; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_2_1 = _T_16087 | _T_9166; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_16104 = _T_15556 & _T_6231; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_2_2 = _T_16104 | _T_9175; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_16121 = _T_15573 & _T_6231; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_2_3 = _T_16121 | _T_9184; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_16138 = _T_15590 & _T_6231; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_2_4 = _T_16138 | _T_9193; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_16155 = _T_15607 & _T_6231; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_2_5 = _T_16155 | _T_9202; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_16172 = _T_15624 & _T_6231; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_2_6 = _T_16172 | _T_9211; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_16189 = _T_15641 & _T_6231; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_2_7 = _T_16189 | _T_9220; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_16206 = _T_15658 & _T_6231; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_2_8 = _T_16206 | _T_9229; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_16223 = _T_15675 & _T_6231; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_2_9 = _T_16223 | _T_9238; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_16240 = _T_15692 & _T_6231; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_2_10 = _T_16240 | _T_9247; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_16257 = _T_15709 & _T_6231; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_2_11 = _T_16257 | _T_9256; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_16274 = _T_15726 & _T_6231; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_2_12 = _T_16274 | _T_9265; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_16291 = _T_15743 & _T_6231; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_2_13 = _T_16291 | _T_9274; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_16308 = _T_15760 & _T_6231; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_2_14 = _T_16308 | _T_9283; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_16325 = _T_15777 & _T_6231; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_2_15 = _T_16325 | _T_9292; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_16342 = _T_15522 & _T_6242; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_3_0 = _T_16342 | _T_9301; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_16359 = _T_15539 & _T_6242; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_3_1 = _T_16359 | _T_9310; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_16376 = _T_15556 & _T_6242; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_3_2 = _T_16376 | _T_9319; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_16393 = _T_15573 & _T_6242; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_3_3 = _T_16393 | _T_9328; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_16410 = _T_15590 & _T_6242; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_3_4 = _T_16410 | _T_9337; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_16427 = _T_15607 & _T_6242; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_3_5 = _T_16427 | _T_9346; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_16444 = _T_15624 & _T_6242; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_3_6 = _T_16444 | _T_9355; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_16461 = _T_15641 & _T_6242; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_3_7 = _T_16461 | _T_9364; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_16478 = _T_15658 & _T_6242; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_3_8 = _T_16478 | _T_9373; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_16495 = _T_15675 & _T_6242; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_3_9 = _T_16495 | _T_9382; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_16512 = _T_15692 & _T_6242; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_3_10 = _T_16512 | _T_9391; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_16529 = _T_15709 & _T_6242; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_3_11 = _T_16529 | _T_9400; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_16546 = _T_15726 & _T_6242; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_3_12 = _T_16546 | _T_9409; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_16563 = _T_15743 & _T_6242; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_3_13 = _T_16563 | _T_9418; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_16580 = _T_15760 & _T_6242; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_3_14 = _T_16580 | _T_9427; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_16597 = _T_15777 & _T_6242; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_3_15 = _T_16597 | _T_9436; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_16614 = _T_15522 & _T_6253; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_4_0 = _T_16614 | _T_9445; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_16631 = _T_15539 & _T_6253; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_4_1 = _T_16631 | _T_9454; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_16648 = _T_15556 & _T_6253; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_4_2 = _T_16648 | _T_9463; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_16665 = _T_15573 & _T_6253; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_4_3 = _T_16665 | _T_9472; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_16682 = _T_15590 & _T_6253; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_4_4 = _T_16682 | _T_9481; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_16699 = _T_15607 & _T_6253; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_4_5 = _T_16699 | _T_9490; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_16716 = _T_15624 & _T_6253; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_4_6 = _T_16716 | _T_9499; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_16733 = _T_15641 & _T_6253; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_4_7 = _T_16733 | _T_9508; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_16750 = _T_15658 & _T_6253; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_4_8 = _T_16750 | _T_9517; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_16767 = _T_15675 & _T_6253; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_4_9 = _T_16767 | _T_9526; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_16784 = _T_15692 & _T_6253; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_4_10 = _T_16784 | _T_9535; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_16801 = _T_15709 & _T_6253; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_4_11 = _T_16801 | _T_9544; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_16818 = _T_15726 & _T_6253; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_4_12 = _T_16818 | _T_9553; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_16835 = _T_15743 & _T_6253; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_4_13 = _T_16835 | _T_9562; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_16852 = _T_15760 & _T_6253; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_4_14 = _T_16852 | _T_9571; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_16869 = _T_15777 & _T_6253; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_4_15 = _T_16869 | _T_9580; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_16886 = _T_15522 & _T_6264; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_5_0 = _T_16886 | _T_9589; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_16903 = _T_15539 & _T_6264; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_5_1 = _T_16903 | _T_9598; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_16920 = _T_15556 & _T_6264; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_5_2 = _T_16920 | _T_9607; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_16937 = _T_15573 & _T_6264; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_5_3 = _T_16937 | _T_9616; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_16954 = _T_15590 & _T_6264; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_5_4 = _T_16954 | _T_9625; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_16971 = _T_15607 & _T_6264; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_5_5 = _T_16971 | _T_9634; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_16988 = _T_15624 & _T_6264; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_5_6 = _T_16988 | _T_9643; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_17005 = _T_15641 & _T_6264; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_5_7 = _T_17005 | _T_9652; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_17022 = _T_15658 & _T_6264; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_5_8 = _T_17022 | _T_9661; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_17039 = _T_15675 & _T_6264; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_5_9 = _T_17039 | _T_9670; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_17056 = _T_15692 & _T_6264; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_5_10 = _T_17056 | _T_9679; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_17073 = _T_15709 & _T_6264; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_5_11 = _T_17073 | _T_9688; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_17090 = _T_15726 & _T_6264; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_5_12 = _T_17090 | _T_9697; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_17107 = _T_15743 & _T_6264; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_5_13 = _T_17107 | _T_9706; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_17124 = _T_15760 & _T_6264; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_5_14 = _T_17124 | _T_9715; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_17141 = _T_15777 & _T_6264; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_5_15 = _T_17141 | _T_9724; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_17158 = _T_15522 & _T_6275; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_6_0 = _T_17158 | _T_9733; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_17175 = _T_15539 & _T_6275; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_6_1 = _T_17175 | _T_9742; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_17192 = _T_15556 & _T_6275; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_6_2 = _T_17192 | _T_9751; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_17209 = _T_15573 & _T_6275; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_6_3 = _T_17209 | _T_9760; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_17226 = _T_15590 & _T_6275; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_6_4 = _T_17226 | _T_9769; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_17243 = _T_15607 & _T_6275; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_6_5 = _T_17243 | _T_9778; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_17260 = _T_15624 & _T_6275; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_6_6 = _T_17260 | _T_9787; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_17277 = _T_15641 & _T_6275; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_6_7 = _T_17277 | _T_9796; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_17294 = _T_15658 & _T_6275; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_6_8 = _T_17294 | _T_9805; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_17311 = _T_15675 & _T_6275; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_6_9 = _T_17311 | _T_9814; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_17328 = _T_15692 & _T_6275; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_6_10 = _T_17328 | _T_9823; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_17345 = _T_15709 & _T_6275; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_6_11 = _T_17345 | _T_9832; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_17362 = _T_15726 & _T_6275; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_6_12 = _T_17362 | _T_9841; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_17379 = _T_15743 & _T_6275; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_6_13 = _T_17379 | _T_9850; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_17396 = _T_15760 & _T_6275; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_6_14 = _T_17396 | _T_9859; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_17413 = _T_15777 & _T_6275; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_6_15 = _T_17413 | _T_9868; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_17430 = _T_15522 & _T_6286; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_7_0 = _T_17430 | _T_9877; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_17447 = _T_15539 & _T_6286; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_7_1 = _T_17447 | _T_9886; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_17464 = _T_15556 & _T_6286; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_7_2 = _T_17464 | _T_9895; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_17481 = _T_15573 & _T_6286; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_7_3 = _T_17481 | _T_9904; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_17498 = _T_15590 & _T_6286; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_7_4 = _T_17498 | _T_9913; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_17515 = _T_15607 & _T_6286; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_7_5 = _T_17515 | _T_9922; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_17532 = _T_15624 & _T_6286; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_7_6 = _T_17532 | _T_9931; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_17549 = _T_15641 & _T_6286; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_7_7 = _T_17549 | _T_9940; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_17566 = _T_15658 & _T_6286; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_7_8 = _T_17566 | _T_9949; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_17583 = _T_15675 & _T_6286; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_7_9 = _T_17583 | _T_9958; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_17600 = _T_15692 & _T_6286; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_7_10 = _T_17600 | _T_9967; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_17617 = _T_15709 & _T_6286; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_7_11 = _T_17617 | _T_9976; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_17634 = _T_15726 & _T_6286; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_7_12 = _T_17634 | _T_9985; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_17651 = _T_15743 & _T_6286; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_7_13 = _T_17651 | _T_9994; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_17668 = _T_15760 & _T_6286; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_7_14 = _T_17668 | _T_10003; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_17685 = _T_15777 & _T_6286; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_7_15 = _T_17685 | _T_10012; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_17702 = _T_15522 & _T_6297; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_8_0 = _T_17702 | _T_10021; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_17719 = _T_15539 & _T_6297; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_8_1 = _T_17719 | _T_10030; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_17736 = _T_15556 & _T_6297; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_8_2 = _T_17736 | _T_10039; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_17753 = _T_15573 & _T_6297; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_8_3 = _T_17753 | _T_10048; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_17770 = _T_15590 & _T_6297; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_8_4 = _T_17770 | _T_10057; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_17787 = _T_15607 & _T_6297; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_8_5 = _T_17787 | _T_10066; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_17804 = _T_15624 & _T_6297; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_8_6 = _T_17804 | _T_10075; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_17821 = _T_15641 & _T_6297; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_8_7 = _T_17821 | _T_10084; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_17838 = _T_15658 & _T_6297; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_8_8 = _T_17838 | _T_10093; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_17855 = _T_15675 & _T_6297; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_8_9 = _T_17855 | _T_10102; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_17872 = _T_15692 & _T_6297; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_8_10 = _T_17872 | _T_10111; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_17889 = _T_15709 & _T_6297; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_8_11 = _T_17889 | _T_10120; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_17906 = _T_15726 & _T_6297; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_8_12 = _T_17906 | _T_10129; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_17923 = _T_15743 & _T_6297; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_8_13 = _T_17923 | _T_10138; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_17940 = _T_15760 & _T_6297; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_8_14 = _T_17940 | _T_10147; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_17957 = _T_15777 & _T_6297; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_8_15 = _T_17957 | _T_10156; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_17974 = _T_15522 & _T_6308; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_9_0 = _T_17974 | _T_10165; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_17991 = _T_15539 & _T_6308; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_9_1 = _T_17991 | _T_10174; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_18008 = _T_15556 & _T_6308; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_9_2 = _T_18008 | _T_10183; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_18025 = _T_15573 & _T_6308; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_9_3 = _T_18025 | _T_10192; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_18042 = _T_15590 & _T_6308; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_9_4 = _T_18042 | _T_10201; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_18059 = _T_15607 & _T_6308; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_9_5 = _T_18059 | _T_10210; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_18076 = _T_15624 & _T_6308; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_9_6 = _T_18076 | _T_10219; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_18093 = _T_15641 & _T_6308; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_9_7 = _T_18093 | _T_10228; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_18110 = _T_15658 & _T_6308; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_9_8 = _T_18110 | _T_10237; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_18127 = _T_15675 & _T_6308; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_9_9 = _T_18127 | _T_10246; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_18144 = _T_15692 & _T_6308; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_9_10 = _T_18144 | _T_10255; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_18161 = _T_15709 & _T_6308; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_9_11 = _T_18161 | _T_10264; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_18178 = _T_15726 & _T_6308; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_9_12 = _T_18178 | _T_10273; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_18195 = _T_15743 & _T_6308; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_9_13 = _T_18195 | _T_10282; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_18212 = _T_15760 & _T_6308; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_9_14 = _T_18212 | _T_10291; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_18229 = _T_15777 & _T_6308; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_9_15 = _T_18229 | _T_10300; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_18246 = _T_15522 & _T_6319; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_10_0 = _T_18246 | _T_10309; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_18263 = _T_15539 & _T_6319; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_10_1 = _T_18263 | _T_10318; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_18280 = _T_15556 & _T_6319; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_10_2 = _T_18280 | _T_10327; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_18297 = _T_15573 & _T_6319; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_10_3 = _T_18297 | _T_10336; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_18314 = _T_15590 & _T_6319; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_10_4 = _T_18314 | _T_10345; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_18331 = _T_15607 & _T_6319; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_10_5 = _T_18331 | _T_10354; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_18348 = _T_15624 & _T_6319; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_10_6 = _T_18348 | _T_10363; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_18365 = _T_15641 & _T_6319; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_10_7 = _T_18365 | _T_10372; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_18382 = _T_15658 & _T_6319; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_10_8 = _T_18382 | _T_10381; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_18399 = _T_15675 & _T_6319; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_10_9 = _T_18399 | _T_10390; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_18416 = _T_15692 & _T_6319; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_10_10 = _T_18416 | _T_10399; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_18433 = _T_15709 & _T_6319; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_10_11 = _T_18433 | _T_10408; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_18450 = _T_15726 & _T_6319; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_10_12 = _T_18450 | _T_10417; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_18467 = _T_15743 & _T_6319; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_10_13 = _T_18467 | _T_10426; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_18484 = _T_15760 & _T_6319; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_10_14 = _T_18484 | _T_10435; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_18501 = _T_15777 & _T_6319; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_10_15 = _T_18501 | _T_10444; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_18518 = _T_15522 & _T_6330; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_11_0 = _T_18518 | _T_10453; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_18535 = _T_15539 & _T_6330; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_11_1 = _T_18535 | _T_10462; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_18552 = _T_15556 & _T_6330; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_11_2 = _T_18552 | _T_10471; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_18569 = _T_15573 & _T_6330; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_11_3 = _T_18569 | _T_10480; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_18586 = _T_15590 & _T_6330; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_11_4 = _T_18586 | _T_10489; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_18603 = _T_15607 & _T_6330; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_11_5 = _T_18603 | _T_10498; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_18620 = _T_15624 & _T_6330; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_11_6 = _T_18620 | _T_10507; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_18637 = _T_15641 & _T_6330; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_11_7 = _T_18637 | _T_10516; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_18654 = _T_15658 & _T_6330; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_11_8 = _T_18654 | _T_10525; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_18671 = _T_15675 & _T_6330; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_11_9 = _T_18671 | _T_10534; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_18688 = _T_15692 & _T_6330; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_11_10 = _T_18688 | _T_10543; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_18705 = _T_15709 & _T_6330; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_11_11 = _T_18705 | _T_10552; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_18722 = _T_15726 & _T_6330; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_11_12 = _T_18722 | _T_10561; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_18739 = _T_15743 & _T_6330; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_11_13 = _T_18739 | _T_10570; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_18756 = _T_15760 & _T_6330; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_11_14 = _T_18756 | _T_10579; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_18773 = _T_15777 & _T_6330; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_11_15 = _T_18773 | _T_10588; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_18790 = _T_15522 & _T_6341; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_12_0 = _T_18790 | _T_10597; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_18807 = _T_15539 & _T_6341; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_12_1 = _T_18807 | _T_10606; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_18824 = _T_15556 & _T_6341; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_12_2 = _T_18824 | _T_10615; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_18841 = _T_15573 & _T_6341; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_12_3 = _T_18841 | _T_10624; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_18858 = _T_15590 & _T_6341; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_12_4 = _T_18858 | _T_10633; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_18875 = _T_15607 & _T_6341; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_12_5 = _T_18875 | _T_10642; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_18892 = _T_15624 & _T_6341; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_12_6 = _T_18892 | _T_10651; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_18909 = _T_15641 & _T_6341; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_12_7 = _T_18909 | _T_10660; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_18926 = _T_15658 & _T_6341; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_12_8 = _T_18926 | _T_10669; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_18943 = _T_15675 & _T_6341; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_12_9 = _T_18943 | _T_10678; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_18960 = _T_15692 & _T_6341; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_12_10 = _T_18960 | _T_10687; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_18977 = _T_15709 & _T_6341; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_12_11 = _T_18977 | _T_10696; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_18994 = _T_15726 & _T_6341; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_12_12 = _T_18994 | _T_10705; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_19011 = _T_15743 & _T_6341; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_12_13 = _T_19011 | _T_10714; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_19028 = _T_15760 & _T_6341; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_12_14 = _T_19028 | _T_10723; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_19045 = _T_15777 & _T_6341; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_12_15 = _T_19045 | _T_10732; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_19062 = _T_15522 & _T_6352; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_13_0 = _T_19062 | _T_10741; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_19079 = _T_15539 & _T_6352; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_13_1 = _T_19079 | _T_10750; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_19096 = _T_15556 & _T_6352; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_13_2 = _T_19096 | _T_10759; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_19113 = _T_15573 & _T_6352; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_13_3 = _T_19113 | _T_10768; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_19130 = _T_15590 & _T_6352; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_13_4 = _T_19130 | _T_10777; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_19147 = _T_15607 & _T_6352; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_13_5 = _T_19147 | _T_10786; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_19164 = _T_15624 & _T_6352; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_13_6 = _T_19164 | _T_10795; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_19181 = _T_15641 & _T_6352; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_13_7 = _T_19181 | _T_10804; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_19198 = _T_15658 & _T_6352; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_13_8 = _T_19198 | _T_10813; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_19215 = _T_15675 & _T_6352; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_13_9 = _T_19215 | _T_10822; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_19232 = _T_15692 & _T_6352; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_13_10 = _T_19232 | _T_10831; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_19249 = _T_15709 & _T_6352; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_13_11 = _T_19249 | _T_10840; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_19266 = _T_15726 & _T_6352; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_13_12 = _T_19266 | _T_10849; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_19283 = _T_15743 & _T_6352; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_13_13 = _T_19283 | _T_10858; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_19300 = _T_15760 & _T_6352; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_13_14 = _T_19300 | _T_10867; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_19317 = _T_15777 & _T_6352; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_13_15 = _T_19317 | _T_10876; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_19334 = _T_15522 & _T_6363; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_14_0 = _T_19334 | _T_10885; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_19351 = _T_15539 & _T_6363; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_14_1 = _T_19351 | _T_10894; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_19368 = _T_15556 & _T_6363; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_14_2 = _T_19368 | _T_10903; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_19385 = _T_15573 & _T_6363; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_14_3 = _T_19385 | _T_10912; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_19402 = _T_15590 & _T_6363; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_14_4 = _T_19402 | _T_10921; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_19419 = _T_15607 & _T_6363; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_14_5 = _T_19419 | _T_10930; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_19436 = _T_15624 & _T_6363; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_14_6 = _T_19436 | _T_10939; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_19453 = _T_15641 & _T_6363; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_14_7 = _T_19453 | _T_10948; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_19470 = _T_15658 & _T_6363; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_14_8 = _T_19470 | _T_10957; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_19487 = _T_15675 & _T_6363; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_14_9 = _T_19487 | _T_10966; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_19504 = _T_15692 & _T_6363; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_14_10 = _T_19504 | _T_10975; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_19521 = _T_15709 & _T_6363; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_14_11 = _T_19521 | _T_10984; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_19538 = _T_15726 & _T_6363; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_14_12 = _T_19538 | _T_10993; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_19555 = _T_15743 & _T_6363; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_14_13 = _T_19555 | _T_11002; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_19572 = _T_15760 & _T_6363; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_14_14 = _T_19572 | _T_11011; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_19589 = _T_15777 & _T_6363; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_14_15 = _T_19589 | _T_11020; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_19606 = _T_15522 & _T_6374; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_15_0 = _T_19606 | _T_11029; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_19623 = _T_15539 & _T_6374; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_15_1 = _T_19623 | _T_11038; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_19640 = _T_15556 & _T_6374; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_15_2 = _T_19640 | _T_11047; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_19657 = _T_15573 & _T_6374; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_15_3 = _T_19657 | _T_11056; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_19674 = _T_15590 & _T_6374; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_15_4 = _T_19674 | _T_11065; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_19691 = _T_15607 & _T_6374; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_15_5 = _T_19691 | _T_11074; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_19708 = _T_15624 & _T_6374; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_15_6 = _T_19708 | _T_11083; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_19725 = _T_15641 & _T_6374; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_15_7 = _T_19725 | _T_11092; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_19742 = _T_15658 & _T_6374; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_15_8 = _T_19742 | _T_11101; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_19759 = _T_15675 & _T_6374; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_15_9 = _T_19759 | _T_11110; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_19776 = _T_15692 & _T_6374; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_15_10 = _T_19776 | _T_11119; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_19793 = _T_15709 & _T_6374; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_15_11 = _T_19793 | _T_11128; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_19810 = _T_15726 & _T_6374; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_15_12 = _T_19810 | _T_11137; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_19827 = _T_15743 & _T_6374; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_15_13 = _T_19827 | _T_11146; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_19844 = _T_15760 & _T_6374; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_15_14 = _T_19844 | _T_11155; // @[el2_ifu_bp_ctl.scala 455:223]
  wire  _T_19861 = _T_15777 & _T_6374; // @[el2_ifu_bp_ctl.scala 455:110]
  wire  bht_bank_sel_1_15_15 = _T_19861 | _T_11164; // @[el2_ifu_bp_ctl.scala 455:223]
  rvclkhdr rvclkhdr ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_io_l1clk),
    .io_clk(rvclkhdr_io_clk),
    .io_en(rvclkhdr_io_en),
    .io_scan_mode(rvclkhdr_io_scan_mode)
  );
  rvclkhdr rvclkhdr_1 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_1_io_l1clk),
    .io_clk(rvclkhdr_1_io_clk),
    .io_en(rvclkhdr_1_io_en),
    .io_scan_mode(rvclkhdr_1_io_scan_mode)
  );
  rvclkhdr rvclkhdr_2 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_2_io_l1clk),
    .io_clk(rvclkhdr_2_io_clk),
    .io_en(rvclkhdr_2_io_en),
    .io_scan_mode(rvclkhdr_2_io_scan_mode)
  );
  rvclkhdr rvclkhdr_3 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_3_io_l1clk),
    .io_clk(rvclkhdr_3_io_clk),
    .io_en(rvclkhdr_3_io_en),
    .io_scan_mode(rvclkhdr_3_io_scan_mode)
  );
  rvclkhdr rvclkhdr_4 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_4_io_l1clk),
    .io_clk(rvclkhdr_4_io_clk),
    .io_en(rvclkhdr_4_io_en),
    .io_scan_mode(rvclkhdr_4_io_scan_mode)
  );
  rvclkhdr rvclkhdr_5 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_5_io_l1clk),
    .io_clk(rvclkhdr_5_io_clk),
    .io_en(rvclkhdr_5_io_en),
    .io_scan_mode(rvclkhdr_5_io_scan_mode)
  );
  rvclkhdr rvclkhdr_6 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_6_io_l1clk),
    .io_clk(rvclkhdr_6_io_clk),
    .io_en(rvclkhdr_6_io_en),
    .io_scan_mode(rvclkhdr_6_io_scan_mode)
  );
  rvclkhdr rvclkhdr_7 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_7_io_l1clk),
    .io_clk(rvclkhdr_7_io_clk),
    .io_en(rvclkhdr_7_io_en),
    .io_scan_mode(rvclkhdr_7_io_scan_mode)
  );
  rvclkhdr rvclkhdr_8 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_8_io_l1clk),
    .io_clk(rvclkhdr_8_io_clk),
    .io_en(rvclkhdr_8_io_en),
    .io_scan_mode(rvclkhdr_8_io_scan_mode)
  );
  rvclkhdr rvclkhdr_9 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_9_io_l1clk),
    .io_clk(rvclkhdr_9_io_clk),
    .io_en(rvclkhdr_9_io_en),
    .io_scan_mode(rvclkhdr_9_io_scan_mode)
  );
  rvclkhdr rvclkhdr_10 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_10_io_l1clk),
    .io_clk(rvclkhdr_10_io_clk),
    .io_en(rvclkhdr_10_io_en),
    .io_scan_mode(rvclkhdr_10_io_scan_mode)
  );
  rvclkhdr rvclkhdr_11 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_11_io_l1clk),
    .io_clk(rvclkhdr_11_io_clk),
    .io_en(rvclkhdr_11_io_en),
    .io_scan_mode(rvclkhdr_11_io_scan_mode)
  );
  rvclkhdr rvclkhdr_12 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_12_io_l1clk),
    .io_clk(rvclkhdr_12_io_clk),
    .io_en(rvclkhdr_12_io_en),
    .io_scan_mode(rvclkhdr_12_io_scan_mode)
  );
  rvclkhdr rvclkhdr_13 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_13_io_l1clk),
    .io_clk(rvclkhdr_13_io_clk),
    .io_en(rvclkhdr_13_io_en),
    .io_scan_mode(rvclkhdr_13_io_scan_mode)
  );
  rvclkhdr rvclkhdr_14 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_14_io_l1clk),
    .io_clk(rvclkhdr_14_io_clk),
    .io_en(rvclkhdr_14_io_en),
    .io_scan_mode(rvclkhdr_14_io_scan_mode)
  );
  rvclkhdr rvclkhdr_15 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_15_io_l1clk),
    .io_clk(rvclkhdr_15_io_clk),
    .io_en(rvclkhdr_15_io_en),
    .io_scan_mode(rvclkhdr_15_io_scan_mode)
  );
  rvclkhdr rvclkhdr_16 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_16_io_l1clk),
    .io_clk(rvclkhdr_16_io_clk),
    .io_en(rvclkhdr_16_io_en),
    .io_scan_mode(rvclkhdr_16_io_scan_mode)
  );
  rvclkhdr rvclkhdr_17 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_17_io_l1clk),
    .io_clk(rvclkhdr_17_io_clk),
    .io_en(rvclkhdr_17_io_en),
    .io_scan_mode(rvclkhdr_17_io_scan_mode)
  );
  rvclkhdr rvclkhdr_18 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_18_io_l1clk),
    .io_clk(rvclkhdr_18_io_clk),
    .io_en(rvclkhdr_18_io_en),
    .io_scan_mode(rvclkhdr_18_io_scan_mode)
  );
  rvclkhdr rvclkhdr_19 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_19_io_l1clk),
    .io_clk(rvclkhdr_19_io_clk),
    .io_en(rvclkhdr_19_io_en),
    .io_scan_mode(rvclkhdr_19_io_scan_mode)
  );
  rvclkhdr rvclkhdr_20 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_20_io_l1clk),
    .io_clk(rvclkhdr_20_io_clk),
    .io_en(rvclkhdr_20_io_en),
    .io_scan_mode(rvclkhdr_20_io_scan_mode)
  );
  rvclkhdr rvclkhdr_21 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_21_io_l1clk),
    .io_clk(rvclkhdr_21_io_clk),
    .io_en(rvclkhdr_21_io_en),
    .io_scan_mode(rvclkhdr_21_io_scan_mode)
  );
  rvclkhdr rvclkhdr_22 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_22_io_l1clk),
    .io_clk(rvclkhdr_22_io_clk),
    .io_en(rvclkhdr_22_io_en),
    .io_scan_mode(rvclkhdr_22_io_scan_mode)
  );
  rvclkhdr rvclkhdr_23 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_23_io_l1clk),
    .io_clk(rvclkhdr_23_io_clk),
    .io_en(rvclkhdr_23_io_en),
    .io_scan_mode(rvclkhdr_23_io_scan_mode)
  );
  rvclkhdr rvclkhdr_24 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_24_io_l1clk),
    .io_clk(rvclkhdr_24_io_clk),
    .io_en(rvclkhdr_24_io_en),
    .io_scan_mode(rvclkhdr_24_io_scan_mode)
  );
  rvclkhdr rvclkhdr_25 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_25_io_l1clk),
    .io_clk(rvclkhdr_25_io_clk),
    .io_en(rvclkhdr_25_io_en),
    .io_scan_mode(rvclkhdr_25_io_scan_mode)
  );
  rvclkhdr rvclkhdr_26 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_26_io_l1clk),
    .io_clk(rvclkhdr_26_io_clk),
    .io_en(rvclkhdr_26_io_en),
    .io_scan_mode(rvclkhdr_26_io_scan_mode)
  );
  rvclkhdr rvclkhdr_27 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_27_io_l1clk),
    .io_clk(rvclkhdr_27_io_clk),
    .io_en(rvclkhdr_27_io_en),
    .io_scan_mode(rvclkhdr_27_io_scan_mode)
  );
  rvclkhdr rvclkhdr_28 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_28_io_l1clk),
    .io_clk(rvclkhdr_28_io_clk),
    .io_en(rvclkhdr_28_io_en),
    .io_scan_mode(rvclkhdr_28_io_scan_mode)
  );
  rvclkhdr rvclkhdr_29 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_29_io_l1clk),
    .io_clk(rvclkhdr_29_io_clk),
    .io_en(rvclkhdr_29_io_en),
    .io_scan_mode(rvclkhdr_29_io_scan_mode)
  );
  rvclkhdr rvclkhdr_30 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_30_io_l1clk),
    .io_clk(rvclkhdr_30_io_clk),
    .io_en(rvclkhdr_30_io_en),
    .io_scan_mode(rvclkhdr_30_io_scan_mode)
  );
  rvclkhdr rvclkhdr_31 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_31_io_l1clk),
    .io_clk(rvclkhdr_31_io_clk),
    .io_en(rvclkhdr_31_io_en),
    .io_scan_mode(rvclkhdr_31_io_scan_mode)
  );
  rvclkhdr rvclkhdr_32 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_32_io_l1clk),
    .io_clk(rvclkhdr_32_io_clk),
    .io_en(rvclkhdr_32_io_en),
    .io_scan_mode(rvclkhdr_32_io_scan_mode)
  );
  rvclkhdr rvclkhdr_33 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_33_io_l1clk),
    .io_clk(rvclkhdr_33_io_clk),
    .io_en(rvclkhdr_33_io_en),
    .io_scan_mode(rvclkhdr_33_io_scan_mode)
  );
  rvclkhdr rvclkhdr_34 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_34_io_l1clk),
    .io_clk(rvclkhdr_34_io_clk),
    .io_en(rvclkhdr_34_io_en),
    .io_scan_mode(rvclkhdr_34_io_scan_mode)
  );
  rvclkhdr rvclkhdr_35 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_35_io_l1clk),
    .io_clk(rvclkhdr_35_io_clk),
    .io_en(rvclkhdr_35_io_en),
    .io_scan_mode(rvclkhdr_35_io_scan_mode)
  );
  rvclkhdr rvclkhdr_36 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_36_io_l1clk),
    .io_clk(rvclkhdr_36_io_clk),
    .io_en(rvclkhdr_36_io_en),
    .io_scan_mode(rvclkhdr_36_io_scan_mode)
  );
  rvclkhdr rvclkhdr_37 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_37_io_l1clk),
    .io_clk(rvclkhdr_37_io_clk),
    .io_en(rvclkhdr_37_io_en),
    .io_scan_mode(rvclkhdr_37_io_scan_mode)
  );
  rvclkhdr rvclkhdr_38 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_38_io_l1clk),
    .io_clk(rvclkhdr_38_io_clk),
    .io_en(rvclkhdr_38_io_en),
    .io_scan_mode(rvclkhdr_38_io_scan_mode)
  );
  rvclkhdr rvclkhdr_39 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_39_io_l1clk),
    .io_clk(rvclkhdr_39_io_clk),
    .io_en(rvclkhdr_39_io_en),
    .io_scan_mode(rvclkhdr_39_io_scan_mode)
  );
  rvclkhdr rvclkhdr_40 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_40_io_l1clk),
    .io_clk(rvclkhdr_40_io_clk),
    .io_en(rvclkhdr_40_io_en),
    .io_scan_mode(rvclkhdr_40_io_scan_mode)
  );
  rvclkhdr rvclkhdr_41 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_41_io_l1clk),
    .io_clk(rvclkhdr_41_io_clk),
    .io_en(rvclkhdr_41_io_en),
    .io_scan_mode(rvclkhdr_41_io_scan_mode)
  );
  rvclkhdr rvclkhdr_42 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_42_io_l1clk),
    .io_clk(rvclkhdr_42_io_clk),
    .io_en(rvclkhdr_42_io_en),
    .io_scan_mode(rvclkhdr_42_io_scan_mode)
  );
  rvclkhdr rvclkhdr_43 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_43_io_l1clk),
    .io_clk(rvclkhdr_43_io_clk),
    .io_en(rvclkhdr_43_io_en),
    .io_scan_mode(rvclkhdr_43_io_scan_mode)
  );
  rvclkhdr rvclkhdr_44 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_44_io_l1clk),
    .io_clk(rvclkhdr_44_io_clk),
    .io_en(rvclkhdr_44_io_en),
    .io_scan_mode(rvclkhdr_44_io_scan_mode)
  );
  rvclkhdr rvclkhdr_45 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_45_io_l1clk),
    .io_clk(rvclkhdr_45_io_clk),
    .io_en(rvclkhdr_45_io_en),
    .io_scan_mode(rvclkhdr_45_io_scan_mode)
  );
  rvclkhdr rvclkhdr_46 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_46_io_l1clk),
    .io_clk(rvclkhdr_46_io_clk),
    .io_en(rvclkhdr_46_io_en),
    .io_scan_mode(rvclkhdr_46_io_scan_mode)
  );
  rvclkhdr rvclkhdr_47 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_47_io_l1clk),
    .io_clk(rvclkhdr_47_io_clk),
    .io_en(rvclkhdr_47_io_en),
    .io_scan_mode(rvclkhdr_47_io_scan_mode)
  );
  rvclkhdr rvclkhdr_48 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_48_io_l1clk),
    .io_clk(rvclkhdr_48_io_clk),
    .io_en(rvclkhdr_48_io_en),
    .io_scan_mode(rvclkhdr_48_io_scan_mode)
  );
  rvclkhdr rvclkhdr_49 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_49_io_l1clk),
    .io_clk(rvclkhdr_49_io_clk),
    .io_en(rvclkhdr_49_io_en),
    .io_scan_mode(rvclkhdr_49_io_scan_mode)
  );
  rvclkhdr rvclkhdr_50 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_50_io_l1clk),
    .io_clk(rvclkhdr_50_io_clk),
    .io_en(rvclkhdr_50_io_en),
    .io_scan_mode(rvclkhdr_50_io_scan_mode)
  );
  rvclkhdr rvclkhdr_51 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_51_io_l1clk),
    .io_clk(rvclkhdr_51_io_clk),
    .io_en(rvclkhdr_51_io_en),
    .io_scan_mode(rvclkhdr_51_io_scan_mode)
  );
  rvclkhdr rvclkhdr_52 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_52_io_l1clk),
    .io_clk(rvclkhdr_52_io_clk),
    .io_en(rvclkhdr_52_io_en),
    .io_scan_mode(rvclkhdr_52_io_scan_mode)
  );
  rvclkhdr rvclkhdr_53 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_53_io_l1clk),
    .io_clk(rvclkhdr_53_io_clk),
    .io_en(rvclkhdr_53_io_en),
    .io_scan_mode(rvclkhdr_53_io_scan_mode)
  );
  rvclkhdr rvclkhdr_54 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_54_io_l1clk),
    .io_clk(rvclkhdr_54_io_clk),
    .io_en(rvclkhdr_54_io_en),
    .io_scan_mode(rvclkhdr_54_io_scan_mode)
  );
  rvclkhdr rvclkhdr_55 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_55_io_l1clk),
    .io_clk(rvclkhdr_55_io_clk),
    .io_en(rvclkhdr_55_io_en),
    .io_scan_mode(rvclkhdr_55_io_scan_mode)
  );
  rvclkhdr rvclkhdr_56 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_56_io_l1clk),
    .io_clk(rvclkhdr_56_io_clk),
    .io_en(rvclkhdr_56_io_en),
    .io_scan_mode(rvclkhdr_56_io_scan_mode)
  );
  rvclkhdr rvclkhdr_57 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_57_io_l1clk),
    .io_clk(rvclkhdr_57_io_clk),
    .io_en(rvclkhdr_57_io_en),
    .io_scan_mode(rvclkhdr_57_io_scan_mode)
  );
  rvclkhdr rvclkhdr_58 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_58_io_l1clk),
    .io_clk(rvclkhdr_58_io_clk),
    .io_en(rvclkhdr_58_io_en),
    .io_scan_mode(rvclkhdr_58_io_scan_mode)
  );
  rvclkhdr rvclkhdr_59 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_59_io_l1clk),
    .io_clk(rvclkhdr_59_io_clk),
    .io_en(rvclkhdr_59_io_en),
    .io_scan_mode(rvclkhdr_59_io_scan_mode)
  );
  rvclkhdr rvclkhdr_60 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_60_io_l1clk),
    .io_clk(rvclkhdr_60_io_clk),
    .io_en(rvclkhdr_60_io_en),
    .io_scan_mode(rvclkhdr_60_io_scan_mode)
  );
  rvclkhdr rvclkhdr_61 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_61_io_l1clk),
    .io_clk(rvclkhdr_61_io_clk),
    .io_en(rvclkhdr_61_io_en),
    .io_scan_mode(rvclkhdr_61_io_scan_mode)
  );
  rvclkhdr rvclkhdr_62 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_62_io_l1clk),
    .io_clk(rvclkhdr_62_io_clk),
    .io_en(rvclkhdr_62_io_en),
    .io_scan_mode(rvclkhdr_62_io_scan_mode)
  );
  rvclkhdr rvclkhdr_63 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_63_io_l1clk),
    .io_clk(rvclkhdr_63_io_clk),
    .io_en(rvclkhdr_63_io_en),
    .io_scan_mode(rvclkhdr_63_io_scan_mode)
  );
  rvclkhdr rvclkhdr_64 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_64_io_l1clk),
    .io_clk(rvclkhdr_64_io_clk),
    .io_en(rvclkhdr_64_io_en),
    .io_scan_mode(rvclkhdr_64_io_scan_mode)
  );
  rvclkhdr rvclkhdr_65 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_65_io_l1clk),
    .io_clk(rvclkhdr_65_io_clk),
    .io_en(rvclkhdr_65_io_en),
    .io_scan_mode(rvclkhdr_65_io_scan_mode)
  );
  rvclkhdr rvclkhdr_66 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_66_io_l1clk),
    .io_clk(rvclkhdr_66_io_clk),
    .io_en(rvclkhdr_66_io_en),
    .io_scan_mode(rvclkhdr_66_io_scan_mode)
  );
  rvclkhdr rvclkhdr_67 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_67_io_l1clk),
    .io_clk(rvclkhdr_67_io_clk),
    .io_en(rvclkhdr_67_io_en),
    .io_scan_mode(rvclkhdr_67_io_scan_mode)
  );
  rvclkhdr rvclkhdr_68 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_68_io_l1clk),
    .io_clk(rvclkhdr_68_io_clk),
    .io_en(rvclkhdr_68_io_en),
    .io_scan_mode(rvclkhdr_68_io_scan_mode)
  );
  rvclkhdr rvclkhdr_69 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_69_io_l1clk),
    .io_clk(rvclkhdr_69_io_clk),
    .io_en(rvclkhdr_69_io_en),
    .io_scan_mode(rvclkhdr_69_io_scan_mode)
  );
  rvclkhdr rvclkhdr_70 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_70_io_l1clk),
    .io_clk(rvclkhdr_70_io_clk),
    .io_en(rvclkhdr_70_io_en),
    .io_scan_mode(rvclkhdr_70_io_scan_mode)
  );
  rvclkhdr rvclkhdr_71 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_71_io_l1clk),
    .io_clk(rvclkhdr_71_io_clk),
    .io_en(rvclkhdr_71_io_en),
    .io_scan_mode(rvclkhdr_71_io_scan_mode)
  );
  rvclkhdr rvclkhdr_72 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_72_io_l1clk),
    .io_clk(rvclkhdr_72_io_clk),
    .io_en(rvclkhdr_72_io_en),
    .io_scan_mode(rvclkhdr_72_io_scan_mode)
  );
  rvclkhdr rvclkhdr_73 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_73_io_l1clk),
    .io_clk(rvclkhdr_73_io_clk),
    .io_en(rvclkhdr_73_io_en),
    .io_scan_mode(rvclkhdr_73_io_scan_mode)
  );
  rvclkhdr rvclkhdr_74 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_74_io_l1clk),
    .io_clk(rvclkhdr_74_io_clk),
    .io_en(rvclkhdr_74_io_en),
    .io_scan_mode(rvclkhdr_74_io_scan_mode)
  );
  rvclkhdr rvclkhdr_75 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_75_io_l1clk),
    .io_clk(rvclkhdr_75_io_clk),
    .io_en(rvclkhdr_75_io_en),
    .io_scan_mode(rvclkhdr_75_io_scan_mode)
  );
  rvclkhdr rvclkhdr_76 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_76_io_l1clk),
    .io_clk(rvclkhdr_76_io_clk),
    .io_en(rvclkhdr_76_io_en),
    .io_scan_mode(rvclkhdr_76_io_scan_mode)
  );
  rvclkhdr rvclkhdr_77 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_77_io_l1clk),
    .io_clk(rvclkhdr_77_io_clk),
    .io_en(rvclkhdr_77_io_en),
    .io_scan_mode(rvclkhdr_77_io_scan_mode)
  );
  rvclkhdr rvclkhdr_78 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_78_io_l1clk),
    .io_clk(rvclkhdr_78_io_clk),
    .io_en(rvclkhdr_78_io_en),
    .io_scan_mode(rvclkhdr_78_io_scan_mode)
  );
  rvclkhdr rvclkhdr_79 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_79_io_l1clk),
    .io_clk(rvclkhdr_79_io_clk),
    .io_en(rvclkhdr_79_io_en),
    .io_scan_mode(rvclkhdr_79_io_scan_mode)
  );
  rvclkhdr rvclkhdr_80 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_80_io_l1clk),
    .io_clk(rvclkhdr_80_io_clk),
    .io_en(rvclkhdr_80_io_en),
    .io_scan_mode(rvclkhdr_80_io_scan_mode)
  );
  rvclkhdr rvclkhdr_81 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_81_io_l1clk),
    .io_clk(rvclkhdr_81_io_clk),
    .io_en(rvclkhdr_81_io_en),
    .io_scan_mode(rvclkhdr_81_io_scan_mode)
  );
  rvclkhdr rvclkhdr_82 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_82_io_l1clk),
    .io_clk(rvclkhdr_82_io_clk),
    .io_en(rvclkhdr_82_io_en),
    .io_scan_mode(rvclkhdr_82_io_scan_mode)
  );
  rvclkhdr rvclkhdr_83 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_83_io_l1clk),
    .io_clk(rvclkhdr_83_io_clk),
    .io_en(rvclkhdr_83_io_en),
    .io_scan_mode(rvclkhdr_83_io_scan_mode)
  );
  rvclkhdr rvclkhdr_84 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_84_io_l1clk),
    .io_clk(rvclkhdr_84_io_clk),
    .io_en(rvclkhdr_84_io_en),
    .io_scan_mode(rvclkhdr_84_io_scan_mode)
  );
  rvclkhdr rvclkhdr_85 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_85_io_l1clk),
    .io_clk(rvclkhdr_85_io_clk),
    .io_en(rvclkhdr_85_io_en),
    .io_scan_mode(rvclkhdr_85_io_scan_mode)
  );
  rvclkhdr rvclkhdr_86 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_86_io_l1clk),
    .io_clk(rvclkhdr_86_io_clk),
    .io_en(rvclkhdr_86_io_en),
    .io_scan_mode(rvclkhdr_86_io_scan_mode)
  );
  rvclkhdr rvclkhdr_87 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_87_io_l1clk),
    .io_clk(rvclkhdr_87_io_clk),
    .io_en(rvclkhdr_87_io_en),
    .io_scan_mode(rvclkhdr_87_io_scan_mode)
  );
  rvclkhdr rvclkhdr_88 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_88_io_l1clk),
    .io_clk(rvclkhdr_88_io_clk),
    .io_en(rvclkhdr_88_io_en),
    .io_scan_mode(rvclkhdr_88_io_scan_mode)
  );
  rvclkhdr rvclkhdr_89 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_89_io_l1clk),
    .io_clk(rvclkhdr_89_io_clk),
    .io_en(rvclkhdr_89_io_en),
    .io_scan_mode(rvclkhdr_89_io_scan_mode)
  );
  rvclkhdr rvclkhdr_90 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_90_io_l1clk),
    .io_clk(rvclkhdr_90_io_clk),
    .io_en(rvclkhdr_90_io_en),
    .io_scan_mode(rvclkhdr_90_io_scan_mode)
  );
  rvclkhdr rvclkhdr_91 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_91_io_l1clk),
    .io_clk(rvclkhdr_91_io_clk),
    .io_en(rvclkhdr_91_io_en),
    .io_scan_mode(rvclkhdr_91_io_scan_mode)
  );
  rvclkhdr rvclkhdr_92 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_92_io_l1clk),
    .io_clk(rvclkhdr_92_io_clk),
    .io_en(rvclkhdr_92_io_en),
    .io_scan_mode(rvclkhdr_92_io_scan_mode)
  );
  rvclkhdr rvclkhdr_93 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_93_io_l1clk),
    .io_clk(rvclkhdr_93_io_clk),
    .io_en(rvclkhdr_93_io_en),
    .io_scan_mode(rvclkhdr_93_io_scan_mode)
  );
  rvclkhdr rvclkhdr_94 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_94_io_l1clk),
    .io_clk(rvclkhdr_94_io_clk),
    .io_en(rvclkhdr_94_io_en),
    .io_scan_mode(rvclkhdr_94_io_scan_mode)
  );
  rvclkhdr rvclkhdr_95 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_95_io_l1clk),
    .io_clk(rvclkhdr_95_io_clk),
    .io_en(rvclkhdr_95_io_en),
    .io_scan_mode(rvclkhdr_95_io_scan_mode)
  );
  rvclkhdr rvclkhdr_96 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_96_io_l1clk),
    .io_clk(rvclkhdr_96_io_clk),
    .io_en(rvclkhdr_96_io_en),
    .io_scan_mode(rvclkhdr_96_io_scan_mode)
  );
  rvclkhdr rvclkhdr_97 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_97_io_l1clk),
    .io_clk(rvclkhdr_97_io_clk),
    .io_en(rvclkhdr_97_io_en),
    .io_scan_mode(rvclkhdr_97_io_scan_mode)
  );
  rvclkhdr rvclkhdr_98 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_98_io_l1clk),
    .io_clk(rvclkhdr_98_io_clk),
    .io_en(rvclkhdr_98_io_en),
    .io_scan_mode(rvclkhdr_98_io_scan_mode)
  );
  rvclkhdr rvclkhdr_99 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_99_io_l1clk),
    .io_clk(rvclkhdr_99_io_clk),
    .io_en(rvclkhdr_99_io_en),
    .io_scan_mode(rvclkhdr_99_io_scan_mode)
  );
  rvclkhdr rvclkhdr_100 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_100_io_l1clk),
    .io_clk(rvclkhdr_100_io_clk),
    .io_en(rvclkhdr_100_io_en),
    .io_scan_mode(rvclkhdr_100_io_scan_mode)
  );
  rvclkhdr rvclkhdr_101 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_101_io_l1clk),
    .io_clk(rvclkhdr_101_io_clk),
    .io_en(rvclkhdr_101_io_en),
    .io_scan_mode(rvclkhdr_101_io_scan_mode)
  );
  rvclkhdr rvclkhdr_102 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_102_io_l1clk),
    .io_clk(rvclkhdr_102_io_clk),
    .io_en(rvclkhdr_102_io_en),
    .io_scan_mode(rvclkhdr_102_io_scan_mode)
  );
  rvclkhdr rvclkhdr_103 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_103_io_l1clk),
    .io_clk(rvclkhdr_103_io_clk),
    .io_en(rvclkhdr_103_io_en),
    .io_scan_mode(rvclkhdr_103_io_scan_mode)
  );
  rvclkhdr rvclkhdr_104 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_104_io_l1clk),
    .io_clk(rvclkhdr_104_io_clk),
    .io_en(rvclkhdr_104_io_en),
    .io_scan_mode(rvclkhdr_104_io_scan_mode)
  );
  rvclkhdr rvclkhdr_105 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_105_io_l1clk),
    .io_clk(rvclkhdr_105_io_clk),
    .io_en(rvclkhdr_105_io_en),
    .io_scan_mode(rvclkhdr_105_io_scan_mode)
  );
  rvclkhdr rvclkhdr_106 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_106_io_l1clk),
    .io_clk(rvclkhdr_106_io_clk),
    .io_en(rvclkhdr_106_io_en),
    .io_scan_mode(rvclkhdr_106_io_scan_mode)
  );
  rvclkhdr rvclkhdr_107 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_107_io_l1clk),
    .io_clk(rvclkhdr_107_io_clk),
    .io_en(rvclkhdr_107_io_en),
    .io_scan_mode(rvclkhdr_107_io_scan_mode)
  );
  rvclkhdr rvclkhdr_108 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_108_io_l1clk),
    .io_clk(rvclkhdr_108_io_clk),
    .io_en(rvclkhdr_108_io_en),
    .io_scan_mode(rvclkhdr_108_io_scan_mode)
  );
  rvclkhdr rvclkhdr_109 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_109_io_l1clk),
    .io_clk(rvclkhdr_109_io_clk),
    .io_en(rvclkhdr_109_io_en),
    .io_scan_mode(rvclkhdr_109_io_scan_mode)
  );
  rvclkhdr rvclkhdr_110 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_110_io_l1clk),
    .io_clk(rvclkhdr_110_io_clk),
    .io_en(rvclkhdr_110_io_en),
    .io_scan_mode(rvclkhdr_110_io_scan_mode)
  );
  rvclkhdr rvclkhdr_111 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_111_io_l1clk),
    .io_clk(rvclkhdr_111_io_clk),
    .io_en(rvclkhdr_111_io_en),
    .io_scan_mode(rvclkhdr_111_io_scan_mode)
  );
  rvclkhdr rvclkhdr_112 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_112_io_l1clk),
    .io_clk(rvclkhdr_112_io_clk),
    .io_en(rvclkhdr_112_io_en),
    .io_scan_mode(rvclkhdr_112_io_scan_mode)
  );
  rvclkhdr rvclkhdr_113 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_113_io_l1clk),
    .io_clk(rvclkhdr_113_io_clk),
    .io_en(rvclkhdr_113_io_en),
    .io_scan_mode(rvclkhdr_113_io_scan_mode)
  );
  rvclkhdr rvclkhdr_114 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_114_io_l1clk),
    .io_clk(rvclkhdr_114_io_clk),
    .io_en(rvclkhdr_114_io_en),
    .io_scan_mode(rvclkhdr_114_io_scan_mode)
  );
  rvclkhdr rvclkhdr_115 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_115_io_l1clk),
    .io_clk(rvclkhdr_115_io_clk),
    .io_en(rvclkhdr_115_io_en),
    .io_scan_mode(rvclkhdr_115_io_scan_mode)
  );
  rvclkhdr rvclkhdr_116 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_116_io_l1clk),
    .io_clk(rvclkhdr_116_io_clk),
    .io_en(rvclkhdr_116_io_en),
    .io_scan_mode(rvclkhdr_116_io_scan_mode)
  );
  rvclkhdr rvclkhdr_117 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_117_io_l1clk),
    .io_clk(rvclkhdr_117_io_clk),
    .io_en(rvclkhdr_117_io_en),
    .io_scan_mode(rvclkhdr_117_io_scan_mode)
  );
  rvclkhdr rvclkhdr_118 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_118_io_l1clk),
    .io_clk(rvclkhdr_118_io_clk),
    .io_en(rvclkhdr_118_io_en),
    .io_scan_mode(rvclkhdr_118_io_scan_mode)
  );
  rvclkhdr rvclkhdr_119 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_119_io_l1clk),
    .io_clk(rvclkhdr_119_io_clk),
    .io_en(rvclkhdr_119_io_en),
    .io_scan_mode(rvclkhdr_119_io_scan_mode)
  );
  rvclkhdr rvclkhdr_120 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_120_io_l1clk),
    .io_clk(rvclkhdr_120_io_clk),
    .io_en(rvclkhdr_120_io_en),
    .io_scan_mode(rvclkhdr_120_io_scan_mode)
  );
  rvclkhdr rvclkhdr_121 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_121_io_l1clk),
    .io_clk(rvclkhdr_121_io_clk),
    .io_en(rvclkhdr_121_io_en),
    .io_scan_mode(rvclkhdr_121_io_scan_mode)
  );
  rvclkhdr rvclkhdr_122 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_122_io_l1clk),
    .io_clk(rvclkhdr_122_io_clk),
    .io_en(rvclkhdr_122_io_en),
    .io_scan_mode(rvclkhdr_122_io_scan_mode)
  );
  rvclkhdr rvclkhdr_123 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_123_io_l1clk),
    .io_clk(rvclkhdr_123_io_clk),
    .io_en(rvclkhdr_123_io_en),
    .io_scan_mode(rvclkhdr_123_io_scan_mode)
  );
  rvclkhdr rvclkhdr_124 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_124_io_l1clk),
    .io_clk(rvclkhdr_124_io_clk),
    .io_en(rvclkhdr_124_io_en),
    .io_scan_mode(rvclkhdr_124_io_scan_mode)
  );
  rvclkhdr rvclkhdr_125 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_125_io_l1clk),
    .io_clk(rvclkhdr_125_io_clk),
    .io_en(rvclkhdr_125_io_en),
    .io_scan_mode(rvclkhdr_125_io_scan_mode)
  );
  rvclkhdr rvclkhdr_126 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_126_io_l1clk),
    .io_clk(rvclkhdr_126_io_clk),
    .io_en(rvclkhdr_126_io_en),
    .io_scan_mode(rvclkhdr_126_io_scan_mode)
  );
  rvclkhdr rvclkhdr_127 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_127_io_l1clk),
    .io_clk(rvclkhdr_127_io_clk),
    .io_en(rvclkhdr_127_io_en),
    .io_scan_mode(rvclkhdr_127_io_scan_mode)
  );
  rvclkhdr rvclkhdr_128 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_128_io_l1clk),
    .io_clk(rvclkhdr_128_io_clk),
    .io_en(rvclkhdr_128_io_en),
    .io_scan_mode(rvclkhdr_128_io_scan_mode)
  );
  rvclkhdr rvclkhdr_129 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_129_io_l1clk),
    .io_clk(rvclkhdr_129_io_clk),
    .io_en(rvclkhdr_129_io_en),
    .io_scan_mode(rvclkhdr_129_io_scan_mode)
  );
  rvclkhdr rvclkhdr_130 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_130_io_l1clk),
    .io_clk(rvclkhdr_130_io_clk),
    .io_en(rvclkhdr_130_io_en),
    .io_scan_mode(rvclkhdr_130_io_scan_mode)
  );
  rvclkhdr rvclkhdr_131 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_131_io_l1clk),
    .io_clk(rvclkhdr_131_io_clk),
    .io_en(rvclkhdr_131_io_en),
    .io_scan_mode(rvclkhdr_131_io_scan_mode)
  );
  rvclkhdr rvclkhdr_132 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_132_io_l1clk),
    .io_clk(rvclkhdr_132_io_clk),
    .io_en(rvclkhdr_132_io_en),
    .io_scan_mode(rvclkhdr_132_io_scan_mode)
  );
  rvclkhdr rvclkhdr_133 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_133_io_l1clk),
    .io_clk(rvclkhdr_133_io_clk),
    .io_en(rvclkhdr_133_io_en),
    .io_scan_mode(rvclkhdr_133_io_scan_mode)
  );
  rvclkhdr rvclkhdr_134 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_134_io_l1clk),
    .io_clk(rvclkhdr_134_io_clk),
    .io_en(rvclkhdr_134_io_en),
    .io_scan_mode(rvclkhdr_134_io_scan_mode)
  );
  rvclkhdr rvclkhdr_135 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_135_io_l1clk),
    .io_clk(rvclkhdr_135_io_clk),
    .io_en(rvclkhdr_135_io_en),
    .io_scan_mode(rvclkhdr_135_io_scan_mode)
  );
  rvclkhdr rvclkhdr_136 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_136_io_l1clk),
    .io_clk(rvclkhdr_136_io_clk),
    .io_en(rvclkhdr_136_io_en),
    .io_scan_mode(rvclkhdr_136_io_scan_mode)
  );
  rvclkhdr rvclkhdr_137 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_137_io_l1clk),
    .io_clk(rvclkhdr_137_io_clk),
    .io_en(rvclkhdr_137_io_en),
    .io_scan_mode(rvclkhdr_137_io_scan_mode)
  );
  rvclkhdr rvclkhdr_138 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_138_io_l1clk),
    .io_clk(rvclkhdr_138_io_clk),
    .io_en(rvclkhdr_138_io_en),
    .io_scan_mode(rvclkhdr_138_io_scan_mode)
  );
  rvclkhdr rvclkhdr_139 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_139_io_l1clk),
    .io_clk(rvclkhdr_139_io_clk),
    .io_en(rvclkhdr_139_io_en),
    .io_scan_mode(rvclkhdr_139_io_scan_mode)
  );
  rvclkhdr rvclkhdr_140 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_140_io_l1clk),
    .io_clk(rvclkhdr_140_io_clk),
    .io_en(rvclkhdr_140_io_en),
    .io_scan_mode(rvclkhdr_140_io_scan_mode)
  );
  rvclkhdr rvclkhdr_141 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_141_io_l1clk),
    .io_clk(rvclkhdr_141_io_clk),
    .io_en(rvclkhdr_141_io_en),
    .io_scan_mode(rvclkhdr_141_io_scan_mode)
  );
  rvclkhdr rvclkhdr_142 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_142_io_l1clk),
    .io_clk(rvclkhdr_142_io_clk),
    .io_en(rvclkhdr_142_io_en),
    .io_scan_mode(rvclkhdr_142_io_scan_mode)
  );
  rvclkhdr rvclkhdr_143 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_143_io_l1clk),
    .io_clk(rvclkhdr_143_io_clk),
    .io_en(rvclkhdr_143_io_en),
    .io_scan_mode(rvclkhdr_143_io_scan_mode)
  );
  rvclkhdr rvclkhdr_144 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_144_io_l1clk),
    .io_clk(rvclkhdr_144_io_clk),
    .io_en(rvclkhdr_144_io_en),
    .io_scan_mode(rvclkhdr_144_io_scan_mode)
  );
  rvclkhdr rvclkhdr_145 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_145_io_l1clk),
    .io_clk(rvclkhdr_145_io_clk),
    .io_en(rvclkhdr_145_io_en),
    .io_scan_mode(rvclkhdr_145_io_scan_mode)
  );
  rvclkhdr rvclkhdr_146 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_146_io_l1clk),
    .io_clk(rvclkhdr_146_io_clk),
    .io_en(rvclkhdr_146_io_en),
    .io_scan_mode(rvclkhdr_146_io_scan_mode)
  );
  rvclkhdr rvclkhdr_147 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_147_io_l1clk),
    .io_clk(rvclkhdr_147_io_clk),
    .io_en(rvclkhdr_147_io_en),
    .io_scan_mode(rvclkhdr_147_io_scan_mode)
  );
  rvclkhdr rvclkhdr_148 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_148_io_l1clk),
    .io_clk(rvclkhdr_148_io_clk),
    .io_en(rvclkhdr_148_io_en),
    .io_scan_mode(rvclkhdr_148_io_scan_mode)
  );
  rvclkhdr rvclkhdr_149 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_149_io_l1clk),
    .io_clk(rvclkhdr_149_io_clk),
    .io_en(rvclkhdr_149_io_en),
    .io_scan_mode(rvclkhdr_149_io_scan_mode)
  );
  rvclkhdr rvclkhdr_150 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_150_io_l1clk),
    .io_clk(rvclkhdr_150_io_clk),
    .io_en(rvclkhdr_150_io_en),
    .io_scan_mode(rvclkhdr_150_io_scan_mode)
  );
  rvclkhdr rvclkhdr_151 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_151_io_l1clk),
    .io_clk(rvclkhdr_151_io_clk),
    .io_en(rvclkhdr_151_io_en),
    .io_scan_mode(rvclkhdr_151_io_scan_mode)
  );
  rvclkhdr rvclkhdr_152 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_152_io_l1clk),
    .io_clk(rvclkhdr_152_io_clk),
    .io_en(rvclkhdr_152_io_en),
    .io_scan_mode(rvclkhdr_152_io_scan_mode)
  );
  rvclkhdr rvclkhdr_153 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_153_io_l1clk),
    .io_clk(rvclkhdr_153_io_clk),
    .io_en(rvclkhdr_153_io_en),
    .io_scan_mode(rvclkhdr_153_io_scan_mode)
  );
  rvclkhdr rvclkhdr_154 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_154_io_l1clk),
    .io_clk(rvclkhdr_154_io_clk),
    .io_en(rvclkhdr_154_io_en),
    .io_scan_mode(rvclkhdr_154_io_scan_mode)
  );
  rvclkhdr rvclkhdr_155 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_155_io_l1clk),
    .io_clk(rvclkhdr_155_io_clk),
    .io_en(rvclkhdr_155_io_en),
    .io_scan_mode(rvclkhdr_155_io_scan_mode)
  );
  rvclkhdr rvclkhdr_156 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_156_io_l1clk),
    .io_clk(rvclkhdr_156_io_clk),
    .io_en(rvclkhdr_156_io_en),
    .io_scan_mode(rvclkhdr_156_io_scan_mode)
  );
  rvclkhdr rvclkhdr_157 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_157_io_l1clk),
    .io_clk(rvclkhdr_157_io_clk),
    .io_en(rvclkhdr_157_io_en),
    .io_scan_mode(rvclkhdr_157_io_scan_mode)
  );
  rvclkhdr rvclkhdr_158 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_158_io_l1clk),
    .io_clk(rvclkhdr_158_io_clk),
    .io_en(rvclkhdr_158_io_en),
    .io_scan_mode(rvclkhdr_158_io_scan_mode)
  );
  rvclkhdr rvclkhdr_159 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_159_io_l1clk),
    .io_clk(rvclkhdr_159_io_clk),
    .io_en(rvclkhdr_159_io_en),
    .io_scan_mode(rvclkhdr_159_io_scan_mode)
  );
  rvclkhdr rvclkhdr_160 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_160_io_l1clk),
    .io_clk(rvclkhdr_160_io_clk),
    .io_en(rvclkhdr_160_io_en),
    .io_scan_mode(rvclkhdr_160_io_scan_mode)
  );
  rvclkhdr rvclkhdr_161 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_161_io_l1clk),
    .io_clk(rvclkhdr_161_io_clk),
    .io_en(rvclkhdr_161_io_en),
    .io_scan_mode(rvclkhdr_161_io_scan_mode)
  );
  rvclkhdr rvclkhdr_162 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_162_io_l1clk),
    .io_clk(rvclkhdr_162_io_clk),
    .io_en(rvclkhdr_162_io_en),
    .io_scan_mode(rvclkhdr_162_io_scan_mode)
  );
  rvclkhdr rvclkhdr_163 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_163_io_l1clk),
    .io_clk(rvclkhdr_163_io_clk),
    .io_en(rvclkhdr_163_io_en),
    .io_scan_mode(rvclkhdr_163_io_scan_mode)
  );
  rvclkhdr rvclkhdr_164 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_164_io_l1clk),
    .io_clk(rvclkhdr_164_io_clk),
    .io_en(rvclkhdr_164_io_en),
    .io_scan_mode(rvclkhdr_164_io_scan_mode)
  );
  rvclkhdr rvclkhdr_165 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_165_io_l1clk),
    .io_clk(rvclkhdr_165_io_clk),
    .io_en(rvclkhdr_165_io_en),
    .io_scan_mode(rvclkhdr_165_io_scan_mode)
  );
  rvclkhdr rvclkhdr_166 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_166_io_l1clk),
    .io_clk(rvclkhdr_166_io_clk),
    .io_en(rvclkhdr_166_io_en),
    .io_scan_mode(rvclkhdr_166_io_scan_mode)
  );
  rvclkhdr rvclkhdr_167 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_167_io_l1clk),
    .io_clk(rvclkhdr_167_io_clk),
    .io_en(rvclkhdr_167_io_en),
    .io_scan_mode(rvclkhdr_167_io_scan_mode)
  );
  rvclkhdr rvclkhdr_168 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_168_io_l1clk),
    .io_clk(rvclkhdr_168_io_clk),
    .io_en(rvclkhdr_168_io_en),
    .io_scan_mode(rvclkhdr_168_io_scan_mode)
  );
  rvclkhdr rvclkhdr_169 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_169_io_l1clk),
    .io_clk(rvclkhdr_169_io_clk),
    .io_en(rvclkhdr_169_io_en),
    .io_scan_mode(rvclkhdr_169_io_scan_mode)
  );
  rvclkhdr rvclkhdr_170 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_170_io_l1clk),
    .io_clk(rvclkhdr_170_io_clk),
    .io_en(rvclkhdr_170_io_en),
    .io_scan_mode(rvclkhdr_170_io_scan_mode)
  );
  rvclkhdr rvclkhdr_171 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_171_io_l1clk),
    .io_clk(rvclkhdr_171_io_clk),
    .io_en(rvclkhdr_171_io_en),
    .io_scan_mode(rvclkhdr_171_io_scan_mode)
  );
  rvclkhdr rvclkhdr_172 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_172_io_l1clk),
    .io_clk(rvclkhdr_172_io_clk),
    .io_en(rvclkhdr_172_io_en),
    .io_scan_mode(rvclkhdr_172_io_scan_mode)
  );
  rvclkhdr rvclkhdr_173 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_173_io_l1clk),
    .io_clk(rvclkhdr_173_io_clk),
    .io_en(rvclkhdr_173_io_en),
    .io_scan_mode(rvclkhdr_173_io_scan_mode)
  );
  rvclkhdr rvclkhdr_174 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_174_io_l1clk),
    .io_clk(rvclkhdr_174_io_clk),
    .io_en(rvclkhdr_174_io_en),
    .io_scan_mode(rvclkhdr_174_io_scan_mode)
  );
  rvclkhdr rvclkhdr_175 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_175_io_l1clk),
    .io_clk(rvclkhdr_175_io_clk),
    .io_en(rvclkhdr_175_io_en),
    .io_scan_mode(rvclkhdr_175_io_scan_mode)
  );
  rvclkhdr rvclkhdr_176 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_176_io_l1clk),
    .io_clk(rvclkhdr_176_io_clk),
    .io_en(rvclkhdr_176_io_en),
    .io_scan_mode(rvclkhdr_176_io_scan_mode)
  );
  rvclkhdr rvclkhdr_177 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_177_io_l1clk),
    .io_clk(rvclkhdr_177_io_clk),
    .io_en(rvclkhdr_177_io_en),
    .io_scan_mode(rvclkhdr_177_io_scan_mode)
  );
  rvclkhdr rvclkhdr_178 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_178_io_l1clk),
    .io_clk(rvclkhdr_178_io_clk),
    .io_en(rvclkhdr_178_io_en),
    .io_scan_mode(rvclkhdr_178_io_scan_mode)
  );
  rvclkhdr rvclkhdr_179 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_179_io_l1clk),
    .io_clk(rvclkhdr_179_io_clk),
    .io_en(rvclkhdr_179_io_en),
    .io_scan_mode(rvclkhdr_179_io_scan_mode)
  );
  rvclkhdr rvclkhdr_180 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_180_io_l1clk),
    .io_clk(rvclkhdr_180_io_clk),
    .io_en(rvclkhdr_180_io_en),
    .io_scan_mode(rvclkhdr_180_io_scan_mode)
  );
  rvclkhdr rvclkhdr_181 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_181_io_l1clk),
    .io_clk(rvclkhdr_181_io_clk),
    .io_en(rvclkhdr_181_io_en),
    .io_scan_mode(rvclkhdr_181_io_scan_mode)
  );
  rvclkhdr rvclkhdr_182 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_182_io_l1clk),
    .io_clk(rvclkhdr_182_io_clk),
    .io_en(rvclkhdr_182_io_en),
    .io_scan_mode(rvclkhdr_182_io_scan_mode)
  );
  rvclkhdr rvclkhdr_183 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_183_io_l1clk),
    .io_clk(rvclkhdr_183_io_clk),
    .io_en(rvclkhdr_183_io_en),
    .io_scan_mode(rvclkhdr_183_io_scan_mode)
  );
  rvclkhdr rvclkhdr_184 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_184_io_l1clk),
    .io_clk(rvclkhdr_184_io_clk),
    .io_en(rvclkhdr_184_io_en),
    .io_scan_mode(rvclkhdr_184_io_scan_mode)
  );
  rvclkhdr rvclkhdr_185 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_185_io_l1clk),
    .io_clk(rvclkhdr_185_io_clk),
    .io_en(rvclkhdr_185_io_en),
    .io_scan_mode(rvclkhdr_185_io_scan_mode)
  );
  rvclkhdr rvclkhdr_186 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_186_io_l1clk),
    .io_clk(rvclkhdr_186_io_clk),
    .io_en(rvclkhdr_186_io_en),
    .io_scan_mode(rvclkhdr_186_io_scan_mode)
  );
  rvclkhdr rvclkhdr_187 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_187_io_l1clk),
    .io_clk(rvclkhdr_187_io_clk),
    .io_en(rvclkhdr_187_io_en),
    .io_scan_mode(rvclkhdr_187_io_scan_mode)
  );
  rvclkhdr rvclkhdr_188 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_188_io_l1clk),
    .io_clk(rvclkhdr_188_io_clk),
    .io_en(rvclkhdr_188_io_en),
    .io_scan_mode(rvclkhdr_188_io_scan_mode)
  );
  rvclkhdr rvclkhdr_189 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_189_io_l1clk),
    .io_clk(rvclkhdr_189_io_clk),
    .io_en(rvclkhdr_189_io_en),
    .io_scan_mode(rvclkhdr_189_io_scan_mode)
  );
  rvclkhdr rvclkhdr_190 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_190_io_l1clk),
    .io_clk(rvclkhdr_190_io_clk),
    .io_en(rvclkhdr_190_io_en),
    .io_scan_mode(rvclkhdr_190_io_scan_mode)
  );
  rvclkhdr rvclkhdr_191 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_191_io_l1clk),
    .io_clk(rvclkhdr_191_io_clk),
    .io_en(rvclkhdr_191_io_en),
    .io_scan_mode(rvclkhdr_191_io_scan_mode)
  );
  rvclkhdr rvclkhdr_192 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_192_io_l1clk),
    .io_clk(rvclkhdr_192_io_clk),
    .io_en(rvclkhdr_192_io_en),
    .io_scan_mode(rvclkhdr_192_io_scan_mode)
  );
  rvclkhdr rvclkhdr_193 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_193_io_l1clk),
    .io_clk(rvclkhdr_193_io_clk),
    .io_en(rvclkhdr_193_io_en),
    .io_scan_mode(rvclkhdr_193_io_scan_mode)
  );
  rvclkhdr rvclkhdr_194 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_194_io_l1clk),
    .io_clk(rvclkhdr_194_io_clk),
    .io_en(rvclkhdr_194_io_en),
    .io_scan_mode(rvclkhdr_194_io_scan_mode)
  );
  rvclkhdr rvclkhdr_195 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_195_io_l1clk),
    .io_clk(rvclkhdr_195_io_clk),
    .io_en(rvclkhdr_195_io_en),
    .io_scan_mode(rvclkhdr_195_io_scan_mode)
  );
  rvclkhdr rvclkhdr_196 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_196_io_l1clk),
    .io_clk(rvclkhdr_196_io_clk),
    .io_en(rvclkhdr_196_io_en),
    .io_scan_mode(rvclkhdr_196_io_scan_mode)
  );
  rvclkhdr rvclkhdr_197 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_197_io_l1clk),
    .io_clk(rvclkhdr_197_io_clk),
    .io_en(rvclkhdr_197_io_en),
    .io_scan_mode(rvclkhdr_197_io_scan_mode)
  );
  rvclkhdr rvclkhdr_198 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_198_io_l1clk),
    .io_clk(rvclkhdr_198_io_clk),
    .io_en(rvclkhdr_198_io_en),
    .io_scan_mode(rvclkhdr_198_io_scan_mode)
  );
  rvclkhdr rvclkhdr_199 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_199_io_l1clk),
    .io_clk(rvclkhdr_199_io_clk),
    .io_en(rvclkhdr_199_io_en),
    .io_scan_mode(rvclkhdr_199_io_scan_mode)
  );
  rvclkhdr rvclkhdr_200 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_200_io_l1clk),
    .io_clk(rvclkhdr_200_io_clk),
    .io_en(rvclkhdr_200_io_en),
    .io_scan_mode(rvclkhdr_200_io_scan_mode)
  );
  rvclkhdr rvclkhdr_201 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_201_io_l1clk),
    .io_clk(rvclkhdr_201_io_clk),
    .io_en(rvclkhdr_201_io_en),
    .io_scan_mode(rvclkhdr_201_io_scan_mode)
  );
  rvclkhdr rvclkhdr_202 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_202_io_l1clk),
    .io_clk(rvclkhdr_202_io_clk),
    .io_en(rvclkhdr_202_io_en),
    .io_scan_mode(rvclkhdr_202_io_scan_mode)
  );
  rvclkhdr rvclkhdr_203 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_203_io_l1clk),
    .io_clk(rvclkhdr_203_io_clk),
    .io_en(rvclkhdr_203_io_en),
    .io_scan_mode(rvclkhdr_203_io_scan_mode)
  );
  rvclkhdr rvclkhdr_204 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_204_io_l1clk),
    .io_clk(rvclkhdr_204_io_clk),
    .io_en(rvclkhdr_204_io_en),
    .io_scan_mode(rvclkhdr_204_io_scan_mode)
  );
  rvclkhdr rvclkhdr_205 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_205_io_l1clk),
    .io_clk(rvclkhdr_205_io_clk),
    .io_en(rvclkhdr_205_io_en),
    .io_scan_mode(rvclkhdr_205_io_scan_mode)
  );
  rvclkhdr rvclkhdr_206 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_206_io_l1clk),
    .io_clk(rvclkhdr_206_io_clk),
    .io_en(rvclkhdr_206_io_en),
    .io_scan_mode(rvclkhdr_206_io_scan_mode)
  );
  rvclkhdr rvclkhdr_207 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_207_io_l1clk),
    .io_clk(rvclkhdr_207_io_clk),
    .io_en(rvclkhdr_207_io_en),
    .io_scan_mode(rvclkhdr_207_io_scan_mode)
  );
  rvclkhdr rvclkhdr_208 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_208_io_l1clk),
    .io_clk(rvclkhdr_208_io_clk),
    .io_en(rvclkhdr_208_io_en),
    .io_scan_mode(rvclkhdr_208_io_scan_mode)
  );
  rvclkhdr rvclkhdr_209 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_209_io_l1clk),
    .io_clk(rvclkhdr_209_io_clk),
    .io_en(rvclkhdr_209_io_en),
    .io_scan_mode(rvclkhdr_209_io_scan_mode)
  );
  rvclkhdr rvclkhdr_210 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_210_io_l1clk),
    .io_clk(rvclkhdr_210_io_clk),
    .io_en(rvclkhdr_210_io_en),
    .io_scan_mode(rvclkhdr_210_io_scan_mode)
  );
  rvclkhdr rvclkhdr_211 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_211_io_l1clk),
    .io_clk(rvclkhdr_211_io_clk),
    .io_en(rvclkhdr_211_io_en),
    .io_scan_mode(rvclkhdr_211_io_scan_mode)
  );
  rvclkhdr rvclkhdr_212 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_212_io_l1clk),
    .io_clk(rvclkhdr_212_io_clk),
    .io_en(rvclkhdr_212_io_en),
    .io_scan_mode(rvclkhdr_212_io_scan_mode)
  );
  rvclkhdr rvclkhdr_213 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_213_io_l1clk),
    .io_clk(rvclkhdr_213_io_clk),
    .io_en(rvclkhdr_213_io_en),
    .io_scan_mode(rvclkhdr_213_io_scan_mode)
  );
  rvclkhdr rvclkhdr_214 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_214_io_l1clk),
    .io_clk(rvclkhdr_214_io_clk),
    .io_en(rvclkhdr_214_io_en),
    .io_scan_mode(rvclkhdr_214_io_scan_mode)
  );
  rvclkhdr rvclkhdr_215 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_215_io_l1clk),
    .io_clk(rvclkhdr_215_io_clk),
    .io_en(rvclkhdr_215_io_en),
    .io_scan_mode(rvclkhdr_215_io_scan_mode)
  );
  rvclkhdr rvclkhdr_216 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_216_io_l1clk),
    .io_clk(rvclkhdr_216_io_clk),
    .io_en(rvclkhdr_216_io_en),
    .io_scan_mode(rvclkhdr_216_io_scan_mode)
  );
  rvclkhdr rvclkhdr_217 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_217_io_l1clk),
    .io_clk(rvclkhdr_217_io_clk),
    .io_en(rvclkhdr_217_io_en),
    .io_scan_mode(rvclkhdr_217_io_scan_mode)
  );
  rvclkhdr rvclkhdr_218 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_218_io_l1clk),
    .io_clk(rvclkhdr_218_io_clk),
    .io_en(rvclkhdr_218_io_en),
    .io_scan_mode(rvclkhdr_218_io_scan_mode)
  );
  rvclkhdr rvclkhdr_219 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_219_io_l1clk),
    .io_clk(rvclkhdr_219_io_clk),
    .io_en(rvclkhdr_219_io_en),
    .io_scan_mode(rvclkhdr_219_io_scan_mode)
  );
  rvclkhdr rvclkhdr_220 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_220_io_l1clk),
    .io_clk(rvclkhdr_220_io_clk),
    .io_en(rvclkhdr_220_io_en),
    .io_scan_mode(rvclkhdr_220_io_scan_mode)
  );
  rvclkhdr rvclkhdr_221 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_221_io_l1clk),
    .io_clk(rvclkhdr_221_io_clk),
    .io_en(rvclkhdr_221_io_en),
    .io_scan_mode(rvclkhdr_221_io_scan_mode)
  );
  rvclkhdr rvclkhdr_222 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_222_io_l1clk),
    .io_clk(rvclkhdr_222_io_clk),
    .io_en(rvclkhdr_222_io_en),
    .io_scan_mode(rvclkhdr_222_io_scan_mode)
  );
  rvclkhdr rvclkhdr_223 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_223_io_l1clk),
    .io_clk(rvclkhdr_223_io_clk),
    .io_en(rvclkhdr_223_io_en),
    .io_scan_mode(rvclkhdr_223_io_scan_mode)
  );
  rvclkhdr rvclkhdr_224 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_224_io_l1clk),
    .io_clk(rvclkhdr_224_io_clk),
    .io_en(rvclkhdr_224_io_en),
    .io_scan_mode(rvclkhdr_224_io_scan_mode)
  );
  rvclkhdr rvclkhdr_225 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_225_io_l1clk),
    .io_clk(rvclkhdr_225_io_clk),
    .io_en(rvclkhdr_225_io_en),
    .io_scan_mode(rvclkhdr_225_io_scan_mode)
  );
  rvclkhdr rvclkhdr_226 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_226_io_l1clk),
    .io_clk(rvclkhdr_226_io_clk),
    .io_en(rvclkhdr_226_io_en),
    .io_scan_mode(rvclkhdr_226_io_scan_mode)
  );
  rvclkhdr rvclkhdr_227 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_227_io_l1clk),
    .io_clk(rvclkhdr_227_io_clk),
    .io_en(rvclkhdr_227_io_en),
    .io_scan_mode(rvclkhdr_227_io_scan_mode)
  );
  rvclkhdr rvclkhdr_228 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_228_io_l1clk),
    .io_clk(rvclkhdr_228_io_clk),
    .io_en(rvclkhdr_228_io_en),
    .io_scan_mode(rvclkhdr_228_io_scan_mode)
  );
  rvclkhdr rvclkhdr_229 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_229_io_l1clk),
    .io_clk(rvclkhdr_229_io_clk),
    .io_en(rvclkhdr_229_io_en),
    .io_scan_mode(rvclkhdr_229_io_scan_mode)
  );
  rvclkhdr rvclkhdr_230 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_230_io_l1clk),
    .io_clk(rvclkhdr_230_io_clk),
    .io_en(rvclkhdr_230_io_en),
    .io_scan_mode(rvclkhdr_230_io_scan_mode)
  );
  rvclkhdr rvclkhdr_231 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_231_io_l1clk),
    .io_clk(rvclkhdr_231_io_clk),
    .io_en(rvclkhdr_231_io_en),
    .io_scan_mode(rvclkhdr_231_io_scan_mode)
  );
  rvclkhdr rvclkhdr_232 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_232_io_l1clk),
    .io_clk(rvclkhdr_232_io_clk),
    .io_en(rvclkhdr_232_io_en),
    .io_scan_mode(rvclkhdr_232_io_scan_mode)
  );
  rvclkhdr rvclkhdr_233 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_233_io_l1clk),
    .io_clk(rvclkhdr_233_io_clk),
    .io_en(rvclkhdr_233_io_en),
    .io_scan_mode(rvclkhdr_233_io_scan_mode)
  );
  rvclkhdr rvclkhdr_234 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_234_io_l1clk),
    .io_clk(rvclkhdr_234_io_clk),
    .io_en(rvclkhdr_234_io_en),
    .io_scan_mode(rvclkhdr_234_io_scan_mode)
  );
  rvclkhdr rvclkhdr_235 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_235_io_l1clk),
    .io_clk(rvclkhdr_235_io_clk),
    .io_en(rvclkhdr_235_io_en),
    .io_scan_mode(rvclkhdr_235_io_scan_mode)
  );
  rvclkhdr rvclkhdr_236 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_236_io_l1clk),
    .io_clk(rvclkhdr_236_io_clk),
    .io_en(rvclkhdr_236_io_en),
    .io_scan_mode(rvclkhdr_236_io_scan_mode)
  );
  rvclkhdr rvclkhdr_237 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_237_io_l1clk),
    .io_clk(rvclkhdr_237_io_clk),
    .io_en(rvclkhdr_237_io_en),
    .io_scan_mode(rvclkhdr_237_io_scan_mode)
  );
  rvclkhdr rvclkhdr_238 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_238_io_l1clk),
    .io_clk(rvclkhdr_238_io_clk),
    .io_en(rvclkhdr_238_io_en),
    .io_scan_mode(rvclkhdr_238_io_scan_mode)
  );
  rvclkhdr rvclkhdr_239 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_239_io_l1clk),
    .io_clk(rvclkhdr_239_io_clk),
    .io_en(rvclkhdr_239_io_en),
    .io_scan_mode(rvclkhdr_239_io_scan_mode)
  );
  rvclkhdr rvclkhdr_240 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_240_io_l1clk),
    .io_clk(rvclkhdr_240_io_clk),
    .io_en(rvclkhdr_240_io_en),
    .io_scan_mode(rvclkhdr_240_io_scan_mode)
  );
  rvclkhdr rvclkhdr_241 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_241_io_l1clk),
    .io_clk(rvclkhdr_241_io_clk),
    .io_en(rvclkhdr_241_io_en),
    .io_scan_mode(rvclkhdr_241_io_scan_mode)
  );
  rvclkhdr rvclkhdr_242 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_242_io_l1clk),
    .io_clk(rvclkhdr_242_io_clk),
    .io_en(rvclkhdr_242_io_en),
    .io_scan_mode(rvclkhdr_242_io_scan_mode)
  );
  rvclkhdr rvclkhdr_243 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_243_io_l1clk),
    .io_clk(rvclkhdr_243_io_clk),
    .io_en(rvclkhdr_243_io_en),
    .io_scan_mode(rvclkhdr_243_io_scan_mode)
  );
  rvclkhdr rvclkhdr_244 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_244_io_l1clk),
    .io_clk(rvclkhdr_244_io_clk),
    .io_en(rvclkhdr_244_io_en),
    .io_scan_mode(rvclkhdr_244_io_scan_mode)
  );
  rvclkhdr rvclkhdr_245 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_245_io_l1clk),
    .io_clk(rvclkhdr_245_io_clk),
    .io_en(rvclkhdr_245_io_en),
    .io_scan_mode(rvclkhdr_245_io_scan_mode)
  );
  rvclkhdr rvclkhdr_246 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_246_io_l1clk),
    .io_clk(rvclkhdr_246_io_clk),
    .io_en(rvclkhdr_246_io_en),
    .io_scan_mode(rvclkhdr_246_io_scan_mode)
  );
  rvclkhdr rvclkhdr_247 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_247_io_l1clk),
    .io_clk(rvclkhdr_247_io_clk),
    .io_en(rvclkhdr_247_io_en),
    .io_scan_mode(rvclkhdr_247_io_scan_mode)
  );
  rvclkhdr rvclkhdr_248 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_248_io_l1clk),
    .io_clk(rvclkhdr_248_io_clk),
    .io_en(rvclkhdr_248_io_en),
    .io_scan_mode(rvclkhdr_248_io_scan_mode)
  );
  rvclkhdr rvclkhdr_249 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_249_io_l1clk),
    .io_clk(rvclkhdr_249_io_clk),
    .io_en(rvclkhdr_249_io_en),
    .io_scan_mode(rvclkhdr_249_io_scan_mode)
  );
  rvclkhdr rvclkhdr_250 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_250_io_l1clk),
    .io_clk(rvclkhdr_250_io_clk),
    .io_en(rvclkhdr_250_io_en),
    .io_scan_mode(rvclkhdr_250_io_scan_mode)
  );
  rvclkhdr rvclkhdr_251 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_251_io_l1clk),
    .io_clk(rvclkhdr_251_io_clk),
    .io_en(rvclkhdr_251_io_en),
    .io_scan_mode(rvclkhdr_251_io_scan_mode)
  );
  rvclkhdr rvclkhdr_252 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_252_io_l1clk),
    .io_clk(rvclkhdr_252_io_clk),
    .io_en(rvclkhdr_252_io_en),
    .io_scan_mode(rvclkhdr_252_io_scan_mode)
  );
  rvclkhdr rvclkhdr_253 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_253_io_l1clk),
    .io_clk(rvclkhdr_253_io_clk),
    .io_en(rvclkhdr_253_io_en),
    .io_scan_mode(rvclkhdr_253_io_scan_mode)
  );
  rvclkhdr rvclkhdr_254 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_254_io_l1clk),
    .io_clk(rvclkhdr_254_io_clk),
    .io_en(rvclkhdr_254_io_en),
    .io_scan_mode(rvclkhdr_254_io_scan_mode)
  );
  rvclkhdr rvclkhdr_255 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_255_io_l1clk),
    .io_clk(rvclkhdr_255_io_clk),
    .io_en(rvclkhdr_255_io_en),
    .io_scan_mode(rvclkhdr_255_io_scan_mode)
  );
  rvclkhdr rvclkhdr_256 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_256_io_l1clk),
    .io_clk(rvclkhdr_256_io_clk),
    .io_en(rvclkhdr_256_io_en),
    .io_scan_mode(rvclkhdr_256_io_scan_mode)
  );
  rvclkhdr rvclkhdr_257 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_257_io_l1clk),
    .io_clk(rvclkhdr_257_io_clk),
    .io_en(rvclkhdr_257_io_en),
    .io_scan_mode(rvclkhdr_257_io_scan_mode)
  );
  rvclkhdr rvclkhdr_258 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_258_io_l1clk),
    .io_clk(rvclkhdr_258_io_clk),
    .io_en(rvclkhdr_258_io_en),
    .io_scan_mode(rvclkhdr_258_io_scan_mode)
  );
  rvclkhdr rvclkhdr_259 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_259_io_l1clk),
    .io_clk(rvclkhdr_259_io_clk),
    .io_en(rvclkhdr_259_io_en),
    .io_scan_mode(rvclkhdr_259_io_scan_mode)
  );
  rvclkhdr rvclkhdr_260 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_260_io_l1clk),
    .io_clk(rvclkhdr_260_io_clk),
    .io_en(rvclkhdr_260_io_en),
    .io_scan_mode(rvclkhdr_260_io_scan_mode)
  );
  rvclkhdr rvclkhdr_261 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_261_io_l1clk),
    .io_clk(rvclkhdr_261_io_clk),
    .io_en(rvclkhdr_261_io_en),
    .io_scan_mode(rvclkhdr_261_io_scan_mode)
  );
  rvclkhdr rvclkhdr_262 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_262_io_l1clk),
    .io_clk(rvclkhdr_262_io_clk),
    .io_en(rvclkhdr_262_io_en),
    .io_scan_mode(rvclkhdr_262_io_scan_mode)
  );
  rvclkhdr rvclkhdr_263 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_263_io_l1clk),
    .io_clk(rvclkhdr_263_io_clk),
    .io_en(rvclkhdr_263_io_en),
    .io_scan_mode(rvclkhdr_263_io_scan_mode)
  );
  rvclkhdr rvclkhdr_264 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_264_io_l1clk),
    .io_clk(rvclkhdr_264_io_clk),
    .io_en(rvclkhdr_264_io_en),
    .io_scan_mode(rvclkhdr_264_io_scan_mode)
  );
  rvclkhdr rvclkhdr_265 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_265_io_l1clk),
    .io_clk(rvclkhdr_265_io_clk),
    .io_en(rvclkhdr_265_io_en),
    .io_scan_mode(rvclkhdr_265_io_scan_mode)
  );
  rvclkhdr rvclkhdr_266 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_266_io_l1clk),
    .io_clk(rvclkhdr_266_io_clk),
    .io_en(rvclkhdr_266_io_en),
    .io_scan_mode(rvclkhdr_266_io_scan_mode)
  );
  rvclkhdr rvclkhdr_267 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_267_io_l1clk),
    .io_clk(rvclkhdr_267_io_clk),
    .io_en(rvclkhdr_267_io_en),
    .io_scan_mode(rvclkhdr_267_io_scan_mode)
  );
  rvclkhdr rvclkhdr_268 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_268_io_l1clk),
    .io_clk(rvclkhdr_268_io_clk),
    .io_en(rvclkhdr_268_io_en),
    .io_scan_mode(rvclkhdr_268_io_scan_mode)
  );
  rvclkhdr rvclkhdr_269 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_269_io_l1clk),
    .io_clk(rvclkhdr_269_io_clk),
    .io_en(rvclkhdr_269_io_en),
    .io_scan_mode(rvclkhdr_269_io_scan_mode)
  );
  rvclkhdr rvclkhdr_270 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_270_io_l1clk),
    .io_clk(rvclkhdr_270_io_clk),
    .io_en(rvclkhdr_270_io_en),
    .io_scan_mode(rvclkhdr_270_io_scan_mode)
  );
  rvclkhdr rvclkhdr_271 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_271_io_l1clk),
    .io_clk(rvclkhdr_271_io_clk),
    .io_en(rvclkhdr_271_io_en),
    .io_scan_mode(rvclkhdr_271_io_scan_mode)
  );
  rvclkhdr rvclkhdr_272 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_272_io_l1clk),
    .io_clk(rvclkhdr_272_io_clk),
    .io_en(rvclkhdr_272_io_en),
    .io_scan_mode(rvclkhdr_272_io_scan_mode)
  );
  rvclkhdr rvclkhdr_273 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_273_io_l1clk),
    .io_clk(rvclkhdr_273_io_clk),
    .io_en(rvclkhdr_273_io_en),
    .io_scan_mode(rvclkhdr_273_io_scan_mode)
  );
  rvclkhdr rvclkhdr_274 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_274_io_l1clk),
    .io_clk(rvclkhdr_274_io_clk),
    .io_en(rvclkhdr_274_io_en),
    .io_scan_mode(rvclkhdr_274_io_scan_mode)
  );
  rvclkhdr rvclkhdr_275 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_275_io_l1clk),
    .io_clk(rvclkhdr_275_io_clk),
    .io_en(rvclkhdr_275_io_en),
    .io_scan_mode(rvclkhdr_275_io_scan_mode)
  );
  rvclkhdr rvclkhdr_276 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_276_io_l1clk),
    .io_clk(rvclkhdr_276_io_clk),
    .io_en(rvclkhdr_276_io_en),
    .io_scan_mode(rvclkhdr_276_io_scan_mode)
  );
  rvclkhdr rvclkhdr_277 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_277_io_l1clk),
    .io_clk(rvclkhdr_277_io_clk),
    .io_en(rvclkhdr_277_io_en),
    .io_scan_mode(rvclkhdr_277_io_scan_mode)
  );
  rvclkhdr rvclkhdr_278 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_278_io_l1clk),
    .io_clk(rvclkhdr_278_io_clk),
    .io_en(rvclkhdr_278_io_en),
    .io_scan_mode(rvclkhdr_278_io_scan_mode)
  );
  rvclkhdr rvclkhdr_279 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_279_io_l1clk),
    .io_clk(rvclkhdr_279_io_clk),
    .io_en(rvclkhdr_279_io_en),
    .io_scan_mode(rvclkhdr_279_io_scan_mode)
  );
  rvclkhdr rvclkhdr_280 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_280_io_l1clk),
    .io_clk(rvclkhdr_280_io_clk),
    .io_en(rvclkhdr_280_io_en),
    .io_scan_mode(rvclkhdr_280_io_scan_mode)
  );
  rvclkhdr rvclkhdr_281 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_281_io_l1clk),
    .io_clk(rvclkhdr_281_io_clk),
    .io_en(rvclkhdr_281_io_en),
    .io_scan_mode(rvclkhdr_281_io_scan_mode)
  );
  rvclkhdr rvclkhdr_282 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_282_io_l1clk),
    .io_clk(rvclkhdr_282_io_clk),
    .io_en(rvclkhdr_282_io_en),
    .io_scan_mode(rvclkhdr_282_io_scan_mode)
  );
  rvclkhdr rvclkhdr_283 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_283_io_l1clk),
    .io_clk(rvclkhdr_283_io_clk),
    .io_en(rvclkhdr_283_io_en),
    .io_scan_mode(rvclkhdr_283_io_scan_mode)
  );
  rvclkhdr rvclkhdr_284 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_284_io_l1clk),
    .io_clk(rvclkhdr_284_io_clk),
    .io_en(rvclkhdr_284_io_en),
    .io_scan_mode(rvclkhdr_284_io_scan_mode)
  );
  rvclkhdr rvclkhdr_285 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_285_io_l1clk),
    .io_clk(rvclkhdr_285_io_clk),
    .io_en(rvclkhdr_285_io_en),
    .io_scan_mode(rvclkhdr_285_io_scan_mode)
  );
  rvclkhdr rvclkhdr_286 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_286_io_l1clk),
    .io_clk(rvclkhdr_286_io_clk),
    .io_en(rvclkhdr_286_io_en),
    .io_scan_mode(rvclkhdr_286_io_scan_mode)
  );
  rvclkhdr rvclkhdr_287 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_287_io_l1clk),
    .io_clk(rvclkhdr_287_io_clk),
    .io_en(rvclkhdr_287_io_en),
    .io_scan_mode(rvclkhdr_287_io_scan_mode)
  );
  rvclkhdr rvclkhdr_288 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_288_io_l1clk),
    .io_clk(rvclkhdr_288_io_clk),
    .io_en(rvclkhdr_288_io_en),
    .io_scan_mode(rvclkhdr_288_io_scan_mode)
  );
  rvclkhdr rvclkhdr_289 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_289_io_l1clk),
    .io_clk(rvclkhdr_289_io_clk),
    .io_en(rvclkhdr_289_io_en),
    .io_scan_mode(rvclkhdr_289_io_scan_mode)
  );
  rvclkhdr rvclkhdr_290 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_290_io_l1clk),
    .io_clk(rvclkhdr_290_io_clk),
    .io_en(rvclkhdr_290_io_en),
    .io_scan_mode(rvclkhdr_290_io_scan_mode)
  );
  rvclkhdr rvclkhdr_291 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_291_io_l1clk),
    .io_clk(rvclkhdr_291_io_clk),
    .io_en(rvclkhdr_291_io_en),
    .io_scan_mode(rvclkhdr_291_io_scan_mode)
  );
  rvclkhdr rvclkhdr_292 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_292_io_l1clk),
    .io_clk(rvclkhdr_292_io_clk),
    .io_en(rvclkhdr_292_io_en),
    .io_scan_mode(rvclkhdr_292_io_scan_mode)
  );
  rvclkhdr rvclkhdr_293 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_293_io_l1clk),
    .io_clk(rvclkhdr_293_io_clk),
    .io_en(rvclkhdr_293_io_en),
    .io_scan_mode(rvclkhdr_293_io_scan_mode)
  );
  rvclkhdr rvclkhdr_294 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_294_io_l1clk),
    .io_clk(rvclkhdr_294_io_clk),
    .io_en(rvclkhdr_294_io_en),
    .io_scan_mode(rvclkhdr_294_io_scan_mode)
  );
  rvclkhdr rvclkhdr_295 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_295_io_l1clk),
    .io_clk(rvclkhdr_295_io_clk),
    .io_en(rvclkhdr_295_io_en),
    .io_scan_mode(rvclkhdr_295_io_scan_mode)
  );
  rvclkhdr rvclkhdr_296 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_296_io_l1clk),
    .io_clk(rvclkhdr_296_io_clk),
    .io_en(rvclkhdr_296_io_en),
    .io_scan_mode(rvclkhdr_296_io_scan_mode)
  );
  rvclkhdr rvclkhdr_297 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_297_io_l1clk),
    .io_clk(rvclkhdr_297_io_clk),
    .io_en(rvclkhdr_297_io_en),
    .io_scan_mode(rvclkhdr_297_io_scan_mode)
  );
  rvclkhdr rvclkhdr_298 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_298_io_l1clk),
    .io_clk(rvclkhdr_298_io_clk),
    .io_en(rvclkhdr_298_io_en),
    .io_scan_mode(rvclkhdr_298_io_scan_mode)
  );
  rvclkhdr rvclkhdr_299 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_299_io_l1clk),
    .io_clk(rvclkhdr_299_io_clk),
    .io_en(rvclkhdr_299_io_en),
    .io_scan_mode(rvclkhdr_299_io_scan_mode)
  );
  rvclkhdr rvclkhdr_300 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_300_io_l1clk),
    .io_clk(rvclkhdr_300_io_clk),
    .io_en(rvclkhdr_300_io_en),
    .io_scan_mode(rvclkhdr_300_io_scan_mode)
  );
  rvclkhdr rvclkhdr_301 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_301_io_l1clk),
    .io_clk(rvclkhdr_301_io_clk),
    .io_en(rvclkhdr_301_io_en),
    .io_scan_mode(rvclkhdr_301_io_scan_mode)
  );
  rvclkhdr rvclkhdr_302 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_302_io_l1clk),
    .io_clk(rvclkhdr_302_io_clk),
    .io_en(rvclkhdr_302_io_en),
    .io_scan_mode(rvclkhdr_302_io_scan_mode)
  );
  rvclkhdr rvclkhdr_303 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_303_io_l1clk),
    .io_clk(rvclkhdr_303_io_clk),
    .io_en(rvclkhdr_303_io_en),
    .io_scan_mode(rvclkhdr_303_io_scan_mode)
  );
  rvclkhdr rvclkhdr_304 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_304_io_l1clk),
    .io_clk(rvclkhdr_304_io_clk),
    .io_en(rvclkhdr_304_io_en),
    .io_scan_mode(rvclkhdr_304_io_scan_mode)
  );
  rvclkhdr rvclkhdr_305 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_305_io_l1clk),
    .io_clk(rvclkhdr_305_io_clk),
    .io_en(rvclkhdr_305_io_en),
    .io_scan_mode(rvclkhdr_305_io_scan_mode)
  );
  rvclkhdr rvclkhdr_306 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_306_io_l1clk),
    .io_clk(rvclkhdr_306_io_clk),
    .io_en(rvclkhdr_306_io_en),
    .io_scan_mode(rvclkhdr_306_io_scan_mode)
  );
  rvclkhdr rvclkhdr_307 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_307_io_l1clk),
    .io_clk(rvclkhdr_307_io_clk),
    .io_en(rvclkhdr_307_io_en),
    .io_scan_mode(rvclkhdr_307_io_scan_mode)
  );
  rvclkhdr rvclkhdr_308 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_308_io_l1clk),
    .io_clk(rvclkhdr_308_io_clk),
    .io_en(rvclkhdr_308_io_en),
    .io_scan_mode(rvclkhdr_308_io_scan_mode)
  );
  rvclkhdr rvclkhdr_309 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_309_io_l1clk),
    .io_clk(rvclkhdr_309_io_clk),
    .io_en(rvclkhdr_309_io_en),
    .io_scan_mode(rvclkhdr_309_io_scan_mode)
  );
  rvclkhdr rvclkhdr_310 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_310_io_l1clk),
    .io_clk(rvclkhdr_310_io_clk),
    .io_en(rvclkhdr_310_io_en),
    .io_scan_mode(rvclkhdr_310_io_scan_mode)
  );
  rvclkhdr rvclkhdr_311 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_311_io_l1clk),
    .io_clk(rvclkhdr_311_io_clk),
    .io_en(rvclkhdr_311_io_en),
    .io_scan_mode(rvclkhdr_311_io_scan_mode)
  );
  rvclkhdr rvclkhdr_312 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_312_io_l1clk),
    .io_clk(rvclkhdr_312_io_clk),
    .io_en(rvclkhdr_312_io_en),
    .io_scan_mode(rvclkhdr_312_io_scan_mode)
  );
  rvclkhdr rvclkhdr_313 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_313_io_l1clk),
    .io_clk(rvclkhdr_313_io_clk),
    .io_en(rvclkhdr_313_io_en),
    .io_scan_mode(rvclkhdr_313_io_scan_mode)
  );
  rvclkhdr rvclkhdr_314 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_314_io_l1clk),
    .io_clk(rvclkhdr_314_io_clk),
    .io_en(rvclkhdr_314_io_en),
    .io_scan_mode(rvclkhdr_314_io_scan_mode)
  );
  rvclkhdr rvclkhdr_315 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_315_io_l1clk),
    .io_clk(rvclkhdr_315_io_clk),
    .io_en(rvclkhdr_315_io_en),
    .io_scan_mode(rvclkhdr_315_io_scan_mode)
  );
  rvclkhdr rvclkhdr_316 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_316_io_l1clk),
    .io_clk(rvclkhdr_316_io_clk),
    .io_en(rvclkhdr_316_io_en),
    .io_scan_mode(rvclkhdr_316_io_scan_mode)
  );
  rvclkhdr rvclkhdr_317 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_317_io_l1clk),
    .io_clk(rvclkhdr_317_io_clk),
    .io_en(rvclkhdr_317_io_en),
    .io_scan_mode(rvclkhdr_317_io_scan_mode)
  );
  rvclkhdr rvclkhdr_318 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_318_io_l1clk),
    .io_clk(rvclkhdr_318_io_clk),
    .io_en(rvclkhdr_318_io_en),
    .io_scan_mode(rvclkhdr_318_io_scan_mode)
  );
  rvclkhdr rvclkhdr_319 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_319_io_l1clk),
    .io_clk(rvclkhdr_319_io_clk),
    .io_en(rvclkhdr_319_io_en),
    .io_scan_mode(rvclkhdr_319_io_scan_mode)
  );
  rvclkhdr rvclkhdr_320 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_320_io_l1clk),
    .io_clk(rvclkhdr_320_io_clk),
    .io_en(rvclkhdr_320_io_en),
    .io_scan_mode(rvclkhdr_320_io_scan_mode)
  );
  rvclkhdr rvclkhdr_321 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_321_io_l1clk),
    .io_clk(rvclkhdr_321_io_clk),
    .io_en(rvclkhdr_321_io_en),
    .io_scan_mode(rvclkhdr_321_io_scan_mode)
  );
  rvclkhdr rvclkhdr_322 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_322_io_l1clk),
    .io_clk(rvclkhdr_322_io_clk),
    .io_en(rvclkhdr_322_io_en),
    .io_scan_mode(rvclkhdr_322_io_scan_mode)
  );
  rvclkhdr rvclkhdr_323 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_323_io_l1clk),
    .io_clk(rvclkhdr_323_io_clk),
    .io_en(rvclkhdr_323_io_en),
    .io_scan_mode(rvclkhdr_323_io_scan_mode)
  );
  rvclkhdr rvclkhdr_324 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_324_io_l1clk),
    .io_clk(rvclkhdr_324_io_clk),
    .io_en(rvclkhdr_324_io_en),
    .io_scan_mode(rvclkhdr_324_io_scan_mode)
  );
  rvclkhdr rvclkhdr_325 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_325_io_l1clk),
    .io_clk(rvclkhdr_325_io_clk),
    .io_en(rvclkhdr_325_io_en),
    .io_scan_mode(rvclkhdr_325_io_scan_mode)
  );
  rvclkhdr rvclkhdr_326 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_326_io_l1clk),
    .io_clk(rvclkhdr_326_io_clk),
    .io_en(rvclkhdr_326_io_en),
    .io_scan_mode(rvclkhdr_326_io_scan_mode)
  );
  rvclkhdr rvclkhdr_327 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_327_io_l1clk),
    .io_clk(rvclkhdr_327_io_clk),
    .io_en(rvclkhdr_327_io_en),
    .io_scan_mode(rvclkhdr_327_io_scan_mode)
  );
  rvclkhdr rvclkhdr_328 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_328_io_l1clk),
    .io_clk(rvclkhdr_328_io_clk),
    .io_en(rvclkhdr_328_io_en),
    .io_scan_mode(rvclkhdr_328_io_scan_mode)
  );
  rvclkhdr rvclkhdr_329 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_329_io_l1clk),
    .io_clk(rvclkhdr_329_io_clk),
    .io_en(rvclkhdr_329_io_en),
    .io_scan_mode(rvclkhdr_329_io_scan_mode)
  );
  rvclkhdr rvclkhdr_330 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_330_io_l1clk),
    .io_clk(rvclkhdr_330_io_clk),
    .io_en(rvclkhdr_330_io_en),
    .io_scan_mode(rvclkhdr_330_io_scan_mode)
  );
  rvclkhdr rvclkhdr_331 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_331_io_l1clk),
    .io_clk(rvclkhdr_331_io_clk),
    .io_en(rvclkhdr_331_io_en),
    .io_scan_mode(rvclkhdr_331_io_scan_mode)
  );
  rvclkhdr rvclkhdr_332 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_332_io_l1clk),
    .io_clk(rvclkhdr_332_io_clk),
    .io_en(rvclkhdr_332_io_en),
    .io_scan_mode(rvclkhdr_332_io_scan_mode)
  );
  rvclkhdr rvclkhdr_333 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_333_io_l1clk),
    .io_clk(rvclkhdr_333_io_clk),
    .io_en(rvclkhdr_333_io_en),
    .io_scan_mode(rvclkhdr_333_io_scan_mode)
  );
  rvclkhdr rvclkhdr_334 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_334_io_l1clk),
    .io_clk(rvclkhdr_334_io_clk),
    .io_en(rvclkhdr_334_io_en),
    .io_scan_mode(rvclkhdr_334_io_scan_mode)
  );
  rvclkhdr rvclkhdr_335 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_335_io_l1clk),
    .io_clk(rvclkhdr_335_io_clk),
    .io_en(rvclkhdr_335_io_en),
    .io_scan_mode(rvclkhdr_335_io_scan_mode)
  );
  rvclkhdr rvclkhdr_336 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_336_io_l1clk),
    .io_clk(rvclkhdr_336_io_clk),
    .io_en(rvclkhdr_336_io_en),
    .io_scan_mode(rvclkhdr_336_io_scan_mode)
  );
  rvclkhdr rvclkhdr_337 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_337_io_l1clk),
    .io_clk(rvclkhdr_337_io_clk),
    .io_en(rvclkhdr_337_io_en),
    .io_scan_mode(rvclkhdr_337_io_scan_mode)
  );
  rvclkhdr rvclkhdr_338 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_338_io_l1clk),
    .io_clk(rvclkhdr_338_io_clk),
    .io_en(rvclkhdr_338_io_en),
    .io_scan_mode(rvclkhdr_338_io_scan_mode)
  );
  rvclkhdr rvclkhdr_339 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_339_io_l1clk),
    .io_clk(rvclkhdr_339_io_clk),
    .io_en(rvclkhdr_339_io_en),
    .io_scan_mode(rvclkhdr_339_io_scan_mode)
  );
  rvclkhdr rvclkhdr_340 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_340_io_l1clk),
    .io_clk(rvclkhdr_340_io_clk),
    .io_en(rvclkhdr_340_io_en),
    .io_scan_mode(rvclkhdr_340_io_scan_mode)
  );
  rvclkhdr rvclkhdr_341 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_341_io_l1clk),
    .io_clk(rvclkhdr_341_io_clk),
    .io_en(rvclkhdr_341_io_en),
    .io_scan_mode(rvclkhdr_341_io_scan_mode)
  );
  rvclkhdr rvclkhdr_342 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_342_io_l1clk),
    .io_clk(rvclkhdr_342_io_clk),
    .io_en(rvclkhdr_342_io_en),
    .io_scan_mode(rvclkhdr_342_io_scan_mode)
  );
  rvclkhdr rvclkhdr_343 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_343_io_l1clk),
    .io_clk(rvclkhdr_343_io_clk),
    .io_en(rvclkhdr_343_io_en),
    .io_scan_mode(rvclkhdr_343_io_scan_mode)
  );
  rvclkhdr rvclkhdr_344 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_344_io_l1clk),
    .io_clk(rvclkhdr_344_io_clk),
    .io_en(rvclkhdr_344_io_en),
    .io_scan_mode(rvclkhdr_344_io_scan_mode)
  );
  rvclkhdr rvclkhdr_345 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_345_io_l1clk),
    .io_clk(rvclkhdr_345_io_clk),
    .io_en(rvclkhdr_345_io_en),
    .io_scan_mode(rvclkhdr_345_io_scan_mode)
  );
  rvclkhdr rvclkhdr_346 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_346_io_l1clk),
    .io_clk(rvclkhdr_346_io_clk),
    .io_en(rvclkhdr_346_io_en),
    .io_scan_mode(rvclkhdr_346_io_scan_mode)
  );
  rvclkhdr rvclkhdr_347 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_347_io_l1clk),
    .io_clk(rvclkhdr_347_io_clk),
    .io_en(rvclkhdr_347_io_en),
    .io_scan_mode(rvclkhdr_347_io_scan_mode)
  );
  rvclkhdr rvclkhdr_348 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_348_io_l1clk),
    .io_clk(rvclkhdr_348_io_clk),
    .io_en(rvclkhdr_348_io_en),
    .io_scan_mode(rvclkhdr_348_io_scan_mode)
  );
  rvclkhdr rvclkhdr_349 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_349_io_l1clk),
    .io_clk(rvclkhdr_349_io_clk),
    .io_en(rvclkhdr_349_io_en),
    .io_scan_mode(rvclkhdr_349_io_scan_mode)
  );
  rvclkhdr rvclkhdr_350 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_350_io_l1clk),
    .io_clk(rvclkhdr_350_io_clk),
    .io_en(rvclkhdr_350_io_en),
    .io_scan_mode(rvclkhdr_350_io_scan_mode)
  );
  rvclkhdr rvclkhdr_351 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_351_io_l1clk),
    .io_clk(rvclkhdr_351_io_clk),
    .io_en(rvclkhdr_351_io_en),
    .io_scan_mode(rvclkhdr_351_io_scan_mode)
  );
  rvclkhdr rvclkhdr_352 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_352_io_l1clk),
    .io_clk(rvclkhdr_352_io_clk),
    .io_en(rvclkhdr_352_io_en),
    .io_scan_mode(rvclkhdr_352_io_scan_mode)
  );
  rvclkhdr rvclkhdr_353 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_353_io_l1clk),
    .io_clk(rvclkhdr_353_io_clk),
    .io_en(rvclkhdr_353_io_en),
    .io_scan_mode(rvclkhdr_353_io_scan_mode)
  );
  rvclkhdr rvclkhdr_354 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_354_io_l1clk),
    .io_clk(rvclkhdr_354_io_clk),
    .io_en(rvclkhdr_354_io_en),
    .io_scan_mode(rvclkhdr_354_io_scan_mode)
  );
  rvclkhdr rvclkhdr_355 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_355_io_l1clk),
    .io_clk(rvclkhdr_355_io_clk),
    .io_en(rvclkhdr_355_io_en),
    .io_scan_mode(rvclkhdr_355_io_scan_mode)
  );
  rvclkhdr rvclkhdr_356 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_356_io_l1clk),
    .io_clk(rvclkhdr_356_io_clk),
    .io_en(rvclkhdr_356_io_en),
    .io_scan_mode(rvclkhdr_356_io_scan_mode)
  );
  rvclkhdr rvclkhdr_357 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_357_io_l1clk),
    .io_clk(rvclkhdr_357_io_clk),
    .io_en(rvclkhdr_357_io_en),
    .io_scan_mode(rvclkhdr_357_io_scan_mode)
  );
  rvclkhdr rvclkhdr_358 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_358_io_l1clk),
    .io_clk(rvclkhdr_358_io_clk),
    .io_en(rvclkhdr_358_io_en),
    .io_scan_mode(rvclkhdr_358_io_scan_mode)
  );
  rvclkhdr rvclkhdr_359 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_359_io_l1clk),
    .io_clk(rvclkhdr_359_io_clk),
    .io_en(rvclkhdr_359_io_en),
    .io_scan_mode(rvclkhdr_359_io_scan_mode)
  );
  rvclkhdr rvclkhdr_360 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_360_io_l1clk),
    .io_clk(rvclkhdr_360_io_clk),
    .io_en(rvclkhdr_360_io_en),
    .io_scan_mode(rvclkhdr_360_io_scan_mode)
  );
  rvclkhdr rvclkhdr_361 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_361_io_l1clk),
    .io_clk(rvclkhdr_361_io_clk),
    .io_en(rvclkhdr_361_io_en),
    .io_scan_mode(rvclkhdr_361_io_scan_mode)
  );
  rvclkhdr rvclkhdr_362 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_362_io_l1clk),
    .io_clk(rvclkhdr_362_io_clk),
    .io_en(rvclkhdr_362_io_en),
    .io_scan_mode(rvclkhdr_362_io_scan_mode)
  );
  rvclkhdr rvclkhdr_363 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_363_io_l1clk),
    .io_clk(rvclkhdr_363_io_clk),
    .io_en(rvclkhdr_363_io_en),
    .io_scan_mode(rvclkhdr_363_io_scan_mode)
  );
  rvclkhdr rvclkhdr_364 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_364_io_l1clk),
    .io_clk(rvclkhdr_364_io_clk),
    .io_en(rvclkhdr_364_io_en),
    .io_scan_mode(rvclkhdr_364_io_scan_mode)
  );
  rvclkhdr rvclkhdr_365 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_365_io_l1clk),
    .io_clk(rvclkhdr_365_io_clk),
    .io_en(rvclkhdr_365_io_en),
    .io_scan_mode(rvclkhdr_365_io_scan_mode)
  );
  rvclkhdr rvclkhdr_366 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_366_io_l1clk),
    .io_clk(rvclkhdr_366_io_clk),
    .io_en(rvclkhdr_366_io_en),
    .io_scan_mode(rvclkhdr_366_io_scan_mode)
  );
  rvclkhdr rvclkhdr_367 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_367_io_l1clk),
    .io_clk(rvclkhdr_367_io_clk),
    .io_en(rvclkhdr_367_io_en),
    .io_scan_mode(rvclkhdr_367_io_scan_mode)
  );
  rvclkhdr rvclkhdr_368 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_368_io_l1clk),
    .io_clk(rvclkhdr_368_io_clk),
    .io_en(rvclkhdr_368_io_en),
    .io_scan_mode(rvclkhdr_368_io_scan_mode)
  );
  rvclkhdr rvclkhdr_369 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_369_io_l1clk),
    .io_clk(rvclkhdr_369_io_clk),
    .io_en(rvclkhdr_369_io_en),
    .io_scan_mode(rvclkhdr_369_io_scan_mode)
  );
  rvclkhdr rvclkhdr_370 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_370_io_l1clk),
    .io_clk(rvclkhdr_370_io_clk),
    .io_en(rvclkhdr_370_io_en),
    .io_scan_mode(rvclkhdr_370_io_scan_mode)
  );
  rvclkhdr rvclkhdr_371 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_371_io_l1clk),
    .io_clk(rvclkhdr_371_io_clk),
    .io_en(rvclkhdr_371_io_en),
    .io_scan_mode(rvclkhdr_371_io_scan_mode)
  );
  rvclkhdr rvclkhdr_372 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_372_io_l1clk),
    .io_clk(rvclkhdr_372_io_clk),
    .io_en(rvclkhdr_372_io_en),
    .io_scan_mode(rvclkhdr_372_io_scan_mode)
  );
  rvclkhdr rvclkhdr_373 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_373_io_l1clk),
    .io_clk(rvclkhdr_373_io_clk),
    .io_en(rvclkhdr_373_io_en),
    .io_scan_mode(rvclkhdr_373_io_scan_mode)
  );
  rvclkhdr rvclkhdr_374 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_374_io_l1clk),
    .io_clk(rvclkhdr_374_io_clk),
    .io_en(rvclkhdr_374_io_en),
    .io_scan_mode(rvclkhdr_374_io_scan_mode)
  );
  rvclkhdr rvclkhdr_375 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_375_io_l1clk),
    .io_clk(rvclkhdr_375_io_clk),
    .io_en(rvclkhdr_375_io_en),
    .io_scan_mode(rvclkhdr_375_io_scan_mode)
  );
  rvclkhdr rvclkhdr_376 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_376_io_l1clk),
    .io_clk(rvclkhdr_376_io_clk),
    .io_en(rvclkhdr_376_io_en),
    .io_scan_mode(rvclkhdr_376_io_scan_mode)
  );
  rvclkhdr rvclkhdr_377 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_377_io_l1clk),
    .io_clk(rvclkhdr_377_io_clk),
    .io_en(rvclkhdr_377_io_en),
    .io_scan_mode(rvclkhdr_377_io_scan_mode)
  );
  rvclkhdr rvclkhdr_378 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_378_io_l1clk),
    .io_clk(rvclkhdr_378_io_clk),
    .io_en(rvclkhdr_378_io_en),
    .io_scan_mode(rvclkhdr_378_io_scan_mode)
  );
  rvclkhdr rvclkhdr_379 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_379_io_l1clk),
    .io_clk(rvclkhdr_379_io_clk),
    .io_en(rvclkhdr_379_io_en),
    .io_scan_mode(rvclkhdr_379_io_scan_mode)
  );
  rvclkhdr rvclkhdr_380 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_380_io_l1clk),
    .io_clk(rvclkhdr_380_io_clk),
    .io_en(rvclkhdr_380_io_en),
    .io_scan_mode(rvclkhdr_380_io_scan_mode)
  );
  rvclkhdr rvclkhdr_381 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_381_io_l1clk),
    .io_clk(rvclkhdr_381_io_clk),
    .io_en(rvclkhdr_381_io_en),
    .io_scan_mode(rvclkhdr_381_io_scan_mode)
  );
  rvclkhdr rvclkhdr_382 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_382_io_l1clk),
    .io_clk(rvclkhdr_382_io_clk),
    .io_en(rvclkhdr_382_io_en),
    .io_scan_mode(rvclkhdr_382_io_scan_mode)
  );
  rvclkhdr rvclkhdr_383 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_383_io_l1clk),
    .io_clk(rvclkhdr_383_io_clk),
    .io_en(rvclkhdr_383_io_en),
    .io_scan_mode(rvclkhdr_383_io_scan_mode)
  );
  rvclkhdr rvclkhdr_384 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_384_io_l1clk),
    .io_clk(rvclkhdr_384_io_clk),
    .io_en(rvclkhdr_384_io_en),
    .io_scan_mode(rvclkhdr_384_io_scan_mode)
  );
  rvclkhdr rvclkhdr_385 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_385_io_l1clk),
    .io_clk(rvclkhdr_385_io_clk),
    .io_en(rvclkhdr_385_io_en),
    .io_scan_mode(rvclkhdr_385_io_scan_mode)
  );
  rvclkhdr rvclkhdr_386 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_386_io_l1clk),
    .io_clk(rvclkhdr_386_io_clk),
    .io_en(rvclkhdr_386_io_en),
    .io_scan_mode(rvclkhdr_386_io_scan_mode)
  );
  rvclkhdr rvclkhdr_387 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_387_io_l1clk),
    .io_clk(rvclkhdr_387_io_clk),
    .io_en(rvclkhdr_387_io_en),
    .io_scan_mode(rvclkhdr_387_io_scan_mode)
  );
  rvclkhdr rvclkhdr_388 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_388_io_l1clk),
    .io_clk(rvclkhdr_388_io_clk),
    .io_en(rvclkhdr_388_io_en),
    .io_scan_mode(rvclkhdr_388_io_scan_mode)
  );
  rvclkhdr rvclkhdr_389 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_389_io_l1clk),
    .io_clk(rvclkhdr_389_io_clk),
    .io_en(rvclkhdr_389_io_en),
    .io_scan_mode(rvclkhdr_389_io_scan_mode)
  );
  rvclkhdr rvclkhdr_390 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_390_io_l1clk),
    .io_clk(rvclkhdr_390_io_clk),
    .io_en(rvclkhdr_390_io_en),
    .io_scan_mode(rvclkhdr_390_io_scan_mode)
  );
  rvclkhdr rvclkhdr_391 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_391_io_l1clk),
    .io_clk(rvclkhdr_391_io_clk),
    .io_en(rvclkhdr_391_io_en),
    .io_scan_mode(rvclkhdr_391_io_scan_mode)
  );
  rvclkhdr rvclkhdr_392 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_392_io_l1clk),
    .io_clk(rvclkhdr_392_io_clk),
    .io_en(rvclkhdr_392_io_en),
    .io_scan_mode(rvclkhdr_392_io_scan_mode)
  );
  rvclkhdr rvclkhdr_393 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_393_io_l1clk),
    .io_clk(rvclkhdr_393_io_clk),
    .io_en(rvclkhdr_393_io_en),
    .io_scan_mode(rvclkhdr_393_io_scan_mode)
  );
  rvclkhdr rvclkhdr_394 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_394_io_l1clk),
    .io_clk(rvclkhdr_394_io_clk),
    .io_en(rvclkhdr_394_io_en),
    .io_scan_mode(rvclkhdr_394_io_scan_mode)
  );
  rvclkhdr rvclkhdr_395 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_395_io_l1clk),
    .io_clk(rvclkhdr_395_io_clk),
    .io_en(rvclkhdr_395_io_en),
    .io_scan_mode(rvclkhdr_395_io_scan_mode)
  );
  rvclkhdr rvclkhdr_396 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_396_io_l1clk),
    .io_clk(rvclkhdr_396_io_clk),
    .io_en(rvclkhdr_396_io_en),
    .io_scan_mode(rvclkhdr_396_io_scan_mode)
  );
  rvclkhdr rvclkhdr_397 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_397_io_l1clk),
    .io_clk(rvclkhdr_397_io_clk),
    .io_en(rvclkhdr_397_io_en),
    .io_scan_mode(rvclkhdr_397_io_scan_mode)
  );
  rvclkhdr rvclkhdr_398 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_398_io_l1clk),
    .io_clk(rvclkhdr_398_io_clk),
    .io_en(rvclkhdr_398_io_en),
    .io_scan_mode(rvclkhdr_398_io_scan_mode)
  );
  rvclkhdr rvclkhdr_399 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_399_io_l1clk),
    .io_clk(rvclkhdr_399_io_clk),
    .io_en(rvclkhdr_399_io_en),
    .io_scan_mode(rvclkhdr_399_io_scan_mode)
  );
  rvclkhdr rvclkhdr_400 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_400_io_l1clk),
    .io_clk(rvclkhdr_400_io_clk),
    .io_en(rvclkhdr_400_io_en),
    .io_scan_mode(rvclkhdr_400_io_scan_mode)
  );
  rvclkhdr rvclkhdr_401 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_401_io_l1clk),
    .io_clk(rvclkhdr_401_io_clk),
    .io_en(rvclkhdr_401_io_en),
    .io_scan_mode(rvclkhdr_401_io_scan_mode)
  );
  rvclkhdr rvclkhdr_402 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_402_io_l1clk),
    .io_clk(rvclkhdr_402_io_clk),
    .io_en(rvclkhdr_402_io_en),
    .io_scan_mode(rvclkhdr_402_io_scan_mode)
  );
  rvclkhdr rvclkhdr_403 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_403_io_l1clk),
    .io_clk(rvclkhdr_403_io_clk),
    .io_en(rvclkhdr_403_io_en),
    .io_scan_mode(rvclkhdr_403_io_scan_mode)
  );
  rvclkhdr rvclkhdr_404 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_404_io_l1clk),
    .io_clk(rvclkhdr_404_io_clk),
    .io_en(rvclkhdr_404_io_en),
    .io_scan_mode(rvclkhdr_404_io_scan_mode)
  );
  rvclkhdr rvclkhdr_405 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_405_io_l1clk),
    .io_clk(rvclkhdr_405_io_clk),
    .io_en(rvclkhdr_405_io_en),
    .io_scan_mode(rvclkhdr_405_io_scan_mode)
  );
  rvclkhdr rvclkhdr_406 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_406_io_l1clk),
    .io_clk(rvclkhdr_406_io_clk),
    .io_en(rvclkhdr_406_io_en),
    .io_scan_mode(rvclkhdr_406_io_scan_mode)
  );
  rvclkhdr rvclkhdr_407 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_407_io_l1clk),
    .io_clk(rvclkhdr_407_io_clk),
    .io_en(rvclkhdr_407_io_en),
    .io_scan_mode(rvclkhdr_407_io_scan_mode)
  );
  rvclkhdr rvclkhdr_408 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_408_io_l1clk),
    .io_clk(rvclkhdr_408_io_clk),
    .io_en(rvclkhdr_408_io_en),
    .io_scan_mode(rvclkhdr_408_io_scan_mode)
  );
  rvclkhdr rvclkhdr_409 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_409_io_l1clk),
    .io_clk(rvclkhdr_409_io_clk),
    .io_en(rvclkhdr_409_io_en),
    .io_scan_mode(rvclkhdr_409_io_scan_mode)
  );
  rvclkhdr rvclkhdr_410 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_410_io_l1clk),
    .io_clk(rvclkhdr_410_io_clk),
    .io_en(rvclkhdr_410_io_en),
    .io_scan_mode(rvclkhdr_410_io_scan_mode)
  );
  rvclkhdr rvclkhdr_411 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_411_io_l1clk),
    .io_clk(rvclkhdr_411_io_clk),
    .io_en(rvclkhdr_411_io_en),
    .io_scan_mode(rvclkhdr_411_io_scan_mode)
  );
  rvclkhdr rvclkhdr_412 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_412_io_l1clk),
    .io_clk(rvclkhdr_412_io_clk),
    .io_en(rvclkhdr_412_io_en),
    .io_scan_mode(rvclkhdr_412_io_scan_mode)
  );
  rvclkhdr rvclkhdr_413 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_413_io_l1clk),
    .io_clk(rvclkhdr_413_io_clk),
    .io_en(rvclkhdr_413_io_en),
    .io_scan_mode(rvclkhdr_413_io_scan_mode)
  );
  rvclkhdr rvclkhdr_414 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_414_io_l1clk),
    .io_clk(rvclkhdr_414_io_clk),
    .io_en(rvclkhdr_414_io_en),
    .io_scan_mode(rvclkhdr_414_io_scan_mode)
  );
  rvclkhdr rvclkhdr_415 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_415_io_l1clk),
    .io_clk(rvclkhdr_415_io_clk),
    .io_en(rvclkhdr_415_io_en),
    .io_scan_mode(rvclkhdr_415_io_scan_mode)
  );
  rvclkhdr rvclkhdr_416 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_416_io_l1clk),
    .io_clk(rvclkhdr_416_io_clk),
    .io_en(rvclkhdr_416_io_en),
    .io_scan_mode(rvclkhdr_416_io_scan_mode)
  );
  rvclkhdr rvclkhdr_417 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_417_io_l1clk),
    .io_clk(rvclkhdr_417_io_clk),
    .io_en(rvclkhdr_417_io_en),
    .io_scan_mode(rvclkhdr_417_io_scan_mode)
  );
  rvclkhdr rvclkhdr_418 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_418_io_l1clk),
    .io_clk(rvclkhdr_418_io_clk),
    .io_en(rvclkhdr_418_io_en),
    .io_scan_mode(rvclkhdr_418_io_scan_mode)
  );
  rvclkhdr rvclkhdr_419 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_419_io_l1clk),
    .io_clk(rvclkhdr_419_io_clk),
    .io_en(rvclkhdr_419_io_en),
    .io_scan_mode(rvclkhdr_419_io_scan_mode)
  );
  rvclkhdr rvclkhdr_420 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_420_io_l1clk),
    .io_clk(rvclkhdr_420_io_clk),
    .io_en(rvclkhdr_420_io_en),
    .io_scan_mode(rvclkhdr_420_io_scan_mode)
  );
  rvclkhdr rvclkhdr_421 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_421_io_l1clk),
    .io_clk(rvclkhdr_421_io_clk),
    .io_en(rvclkhdr_421_io_en),
    .io_scan_mode(rvclkhdr_421_io_scan_mode)
  );
  rvclkhdr rvclkhdr_422 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_422_io_l1clk),
    .io_clk(rvclkhdr_422_io_clk),
    .io_en(rvclkhdr_422_io_en),
    .io_scan_mode(rvclkhdr_422_io_scan_mode)
  );
  rvclkhdr rvclkhdr_423 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_423_io_l1clk),
    .io_clk(rvclkhdr_423_io_clk),
    .io_en(rvclkhdr_423_io_en),
    .io_scan_mode(rvclkhdr_423_io_scan_mode)
  );
  rvclkhdr rvclkhdr_424 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_424_io_l1clk),
    .io_clk(rvclkhdr_424_io_clk),
    .io_en(rvclkhdr_424_io_en),
    .io_scan_mode(rvclkhdr_424_io_scan_mode)
  );
  rvclkhdr rvclkhdr_425 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_425_io_l1clk),
    .io_clk(rvclkhdr_425_io_clk),
    .io_en(rvclkhdr_425_io_en),
    .io_scan_mode(rvclkhdr_425_io_scan_mode)
  );
  rvclkhdr rvclkhdr_426 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_426_io_l1clk),
    .io_clk(rvclkhdr_426_io_clk),
    .io_en(rvclkhdr_426_io_en),
    .io_scan_mode(rvclkhdr_426_io_scan_mode)
  );
  rvclkhdr rvclkhdr_427 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_427_io_l1clk),
    .io_clk(rvclkhdr_427_io_clk),
    .io_en(rvclkhdr_427_io_en),
    .io_scan_mode(rvclkhdr_427_io_scan_mode)
  );
  rvclkhdr rvclkhdr_428 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_428_io_l1clk),
    .io_clk(rvclkhdr_428_io_clk),
    .io_en(rvclkhdr_428_io_en),
    .io_scan_mode(rvclkhdr_428_io_scan_mode)
  );
  rvclkhdr rvclkhdr_429 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_429_io_l1clk),
    .io_clk(rvclkhdr_429_io_clk),
    .io_en(rvclkhdr_429_io_en),
    .io_scan_mode(rvclkhdr_429_io_scan_mode)
  );
  rvclkhdr rvclkhdr_430 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_430_io_l1clk),
    .io_clk(rvclkhdr_430_io_clk),
    .io_en(rvclkhdr_430_io_en),
    .io_scan_mode(rvclkhdr_430_io_scan_mode)
  );
  rvclkhdr rvclkhdr_431 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_431_io_l1clk),
    .io_clk(rvclkhdr_431_io_clk),
    .io_en(rvclkhdr_431_io_en),
    .io_scan_mode(rvclkhdr_431_io_scan_mode)
  );
  rvclkhdr rvclkhdr_432 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_432_io_l1clk),
    .io_clk(rvclkhdr_432_io_clk),
    .io_en(rvclkhdr_432_io_en),
    .io_scan_mode(rvclkhdr_432_io_scan_mode)
  );
  rvclkhdr rvclkhdr_433 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_433_io_l1clk),
    .io_clk(rvclkhdr_433_io_clk),
    .io_en(rvclkhdr_433_io_en),
    .io_scan_mode(rvclkhdr_433_io_scan_mode)
  );
  rvclkhdr rvclkhdr_434 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_434_io_l1clk),
    .io_clk(rvclkhdr_434_io_clk),
    .io_en(rvclkhdr_434_io_en),
    .io_scan_mode(rvclkhdr_434_io_scan_mode)
  );
  rvclkhdr rvclkhdr_435 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_435_io_l1clk),
    .io_clk(rvclkhdr_435_io_clk),
    .io_en(rvclkhdr_435_io_en),
    .io_scan_mode(rvclkhdr_435_io_scan_mode)
  );
  rvclkhdr rvclkhdr_436 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_436_io_l1clk),
    .io_clk(rvclkhdr_436_io_clk),
    .io_en(rvclkhdr_436_io_en),
    .io_scan_mode(rvclkhdr_436_io_scan_mode)
  );
  rvclkhdr rvclkhdr_437 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_437_io_l1clk),
    .io_clk(rvclkhdr_437_io_clk),
    .io_en(rvclkhdr_437_io_en),
    .io_scan_mode(rvclkhdr_437_io_scan_mode)
  );
  rvclkhdr rvclkhdr_438 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_438_io_l1clk),
    .io_clk(rvclkhdr_438_io_clk),
    .io_en(rvclkhdr_438_io_en),
    .io_scan_mode(rvclkhdr_438_io_scan_mode)
  );
  rvclkhdr rvclkhdr_439 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_439_io_l1clk),
    .io_clk(rvclkhdr_439_io_clk),
    .io_en(rvclkhdr_439_io_en),
    .io_scan_mode(rvclkhdr_439_io_scan_mode)
  );
  rvclkhdr rvclkhdr_440 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_440_io_l1clk),
    .io_clk(rvclkhdr_440_io_clk),
    .io_en(rvclkhdr_440_io_en),
    .io_scan_mode(rvclkhdr_440_io_scan_mode)
  );
  rvclkhdr rvclkhdr_441 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_441_io_l1clk),
    .io_clk(rvclkhdr_441_io_clk),
    .io_en(rvclkhdr_441_io_en),
    .io_scan_mode(rvclkhdr_441_io_scan_mode)
  );
  rvclkhdr rvclkhdr_442 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_442_io_l1clk),
    .io_clk(rvclkhdr_442_io_clk),
    .io_en(rvclkhdr_442_io_en),
    .io_scan_mode(rvclkhdr_442_io_scan_mode)
  );
  rvclkhdr rvclkhdr_443 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_443_io_l1clk),
    .io_clk(rvclkhdr_443_io_clk),
    .io_en(rvclkhdr_443_io_en),
    .io_scan_mode(rvclkhdr_443_io_scan_mode)
  );
  rvclkhdr rvclkhdr_444 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_444_io_l1clk),
    .io_clk(rvclkhdr_444_io_clk),
    .io_en(rvclkhdr_444_io_en),
    .io_scan_mode(rvclkhdr_444_io_scan_mode)
  );
  rvclkhdr rvclkhdr_445 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_445_io_l1clk),
    .io_clk(rvclkhdr_445_io_clk),
    .io_en(rvclkhdr_445_io_en),
    .io_scan_mode(rvclkhdr_445_io_scan_mode)
  );
  rvclkhdr rvclkhdr_446 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_446_io_l1clk),
    .io_clk(rvclkhdr_446_io_clk),
    .io_en(rvclkhdr_446_io_en),
    .io_scan_mode(rvclkhdr_446_io_scan_mode)
  );
  rvclkhdr rvclkhdr_447 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_447_io_l1clk),
    .io_clk(rvclkhdr_447_io_clk),
    .io_en(rvclkhdr_447_io_en),
    .io_scan_mode(rvclkhdr_447_io_scan_mode)
  );
  rvclkhdr rvclkhdr_448 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_448_io_l1clk),
    .io_clk(rvclkhdr_448_io_clk),
    .io_en(rvclkhdr_448_io_en),
    .io_scan_mode(rvclkhdr_448_io_scan_mode)
  );
  rvclkhdr rvclkhdr_449 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_449_io_l1clk),
    .io_clk(rvclkhdr_449_io_clk),
    .io_en(rvclkhdr_449_io_en),
    .io_scan_mode(rvclkhdr_449_io_scan_mode)
  );
  rvclkhdr rvclkhdr_450 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_450_io_l1clk),
    .io_clk(rvclkhdr_450_io_clk),
    .io_en(rvclkhdr_450_io_en),
    .io_scan_mode(rvclkhdr_450_io_scan_mode)
  );
  rvclkhdr rvclkhdr_451 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_451_io_l1clk),
    .io_clk(rvclkhdr_451_io_clk),
    .io_en(rvclkhdr_451_io_en),
    .io_scan_mode(rvclkhdr_451_io_scan_mode)
  );
  rvclkhdr rvclkhdr_452 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_452_io_l1clk),
    .io_clk(rvclkhdr_452_io_clk),
    .io_en(rvclkhdr_452_io_en),
    .io_scan_mode(rvclkhdr_452_io_scan_mode)
  );
  rvclkhdr rvclkhdr_453 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_453_io_l1clk),
    .io_clk(rvclkhdr_453_io_clk),
    .io_en(rvclkhdr_453_io_en),
    .io_scan_mode(rvclkhdr_453_io_scan_mode)
  );
  rvclkhdr rvclkhdr_454 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_454_io_l1clk),
    .io_clk(rvclkhdr_454_io_clk),
    .io_en(rvclkhdr_454_io_en),
    .io_scan_mode(rvclkhdr_454_io_scan_mode)
  );
  rvclkhdr rvclkhdr_455 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_455_io_l1clk),
    .io_clk(rvclkhdr_455_io_clk),
    .io_en(rvclkhdr_455_io_en),
    .io_scan_mode(rvclkhdr_455_io_scan_mode)
  );
  rvclkhdr rvclkhdr_456 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_456_io_l1clk),
    .io_clk(rvclkhdr_456_io_clk),
    .io_en(rvclkhdr_456_io_en),
    .io_scan_mode(rvclkhdr_456_io_scan_mode)
  );
  rvclkhdr rvclkhdr_457 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_457_io_l1clk),
    .io_clk(rvclkhdr_457_io_clk),
    .io_en(rvclkhdr_457_io_en),
    .io_scan_mode(rvclkhdr_457_io_scan_mode)
  );
  rvclkhdr rvclkhdr_458 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_458_io_l1clk),
    .io_clk(rvclkhdr_458_io_clk),
    .io_en(rvclkhdr_458_io_en),
    .io_scan_mode(rvclkhdr_458_io_scan_mode)
  );
  rvclkhdr rvclkhdr_459 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_459_io_l1clk),
    .io_clk(rvclkhdr_459_io_clk),
    .io_en(rvclkhdr_459_io_en),
    .io_scan_mode(rvclkhdr_459_io_scan_mode)
  );
  rvclkhdr rvclkhdr_460 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_460_io_l1clk),
    .io_clk(rvclkhdr_460_io_clk),
    .io_en(rvclkhdr_460_io_en),
    .io_scan_mode(rvclkhdr_460_io_scan_mode)
  );
  rvclkhdr rvclkhdr_461 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_461_io_l1clk),
    .io_clk(rvclkhdr_461_io_clk),
    .io_en(rvclkhdr_461_io_en),
    .io_scan_mode(rvclkhdr_461_io_scan_mode)
  );
  rvclkhdr rvclkhdr_462 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_462_io_l1clk),
    .io_clk(rvclkhdr_462_io_clk),
    .io_en(rvclkhdr_462_io_en),
    .io_scan_mode(rvclkhdr_462_io_scan_mode)
  );
  rvclkhdr rvclkhdr_463 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_463_io_l1clk),
    .io_clk(rvclkhdr_463_io_clk),
    .io_en(rvclkhdr_463_io_en),
    .io_scan_mode(rvclkhdr_463_io_scan_mode)
  );
  rvclkhdr rvclkhdr_464 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_464_io_l1clk),
    .io_clk(rvclkhdr_464_io_clk),
    .io_en(rvclkhdr_464_io_en),
    .io_scan_mode(rvclkhdr_464_io_scan_mode)
  );
  rvclkhdr rvclkhdr_465 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_465_io_l1clk),
    .io_clk(rvclkhdr_465_io_clk),
    .io_en(rvclkhdr_465_io_en),
    .io_scan_mode(rvclkhdr_465_io_scan_mode)
  );
  rvclkhdr rvclkhdr_466 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_466_io_l1clk),
    .io_clk(rvclkhdr_466_io_clk),
    .io_en(rvclkhdr_466_io_en),
    .io_scan_mode(rvclkhdr_466_io_scan_mode)
  );
  rvclkhdr rvclkhdr_467 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_467_io_l1clk),
    .io_clk(rvclkhdr_467_io_clk),
    .io_en(rvclkhdr_467_io_en),
    .io_scan_mode(rvclkhdr_467_io_scan_mode)
  );
  rvclkhdr rvclkhdr_468 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_468_io_l1clk),
    .io_clk(rvclkhdr_468_io_clk),
    .io_en(rvclkhdr_468_io_en),
    .io_scan_mode(rvclkhdr_468_io_scan_mode)
  );
  rvclkhdr rvclkhdr_469 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_469_io_l1clk),
    .io_clk(rvclkhdr_469_io_clk),
    .io_en(rvclkhdr_469_io_en),
    .io_scan_mode(rvclkhdr_469_io_scan_mode)
  );
  rvclkhdr rvclkhdr_470 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_470_io_l1clk),
    .io_clk(rvclkhdr_470_io_clk),
    .io_en(rvclkhdr_470_io_en),
    .io_scan_mode(rvclkhdr_470_io_scan_mode)
  );
  rvclkhdr rvclkhdr_471 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_471_io_l1clk),
    .io_clk(rvclkhdr_471_io_clk),
    .io_en(rvclkhdr_471_io_en),
    .io_scan_mode(rvclkhdr_471_io_scan_mode)
  );
  rvclkhdr rvclkhdr_472 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_472_io_l1clk),
    .io_clk(rvclkhdr_472_io_clk),
    .io_en(rvclkhdr_472_io_en),
    .io_scan_mode(rvclkhdr_472_io_scan_mode)
  );
  rvclkhdr rvclkhdr_473 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_473_io_l1clk),
    .io_clk(rvclkhdr_473_io_clk),
    .io_en(rvclkhdr_473_io_en),
    .io_scan_mode(rvclkhdr_473_io_scan_mode)
  );
  rvclkhdr rvclkhdr_474 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_474_io_l1clk),
    .io_clk(rvclkhdr_474_io_clk),
    .io_en(rvclkhdr_474_io_en),
    .io_scan_mode(rvclkhdr_474_io_scan_mode)
  );
  rvclkhdr rvclkhdr_475 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_475_io_l1clk),
    .io_clk(rvclkhdr_475_io_clk),
    .io_en(rvclkhdr_475_io_en),
    .io_scan_mode(rvclkhdr_475_io_scan_mode)
  );
  rvclkhdr rvclkhdr_476 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_476_io_l1clk),
    .io_clk(rvclkhdr_476_io_clk),
    .io_en(rvclkhdr_476_io_en),
    .io_scan_mode(rvclkhdr_476_io_scan_mode)
  );
  rvclkhdr rvclkhdr_477 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_477_io_l1clk),
    .io_clk(rvclkhdr_477_io_clk),
    .io_en(rvclkhdr_477_io_en),
    .io_scan_mode(rvclkhdr_477_io_scan_mode)
  );
  rvclkhdr rvclkhdr_478 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_478_io_l1clk),
    .io_clk(rvclkhdr_478_io_clk),
    .io_en(rvclkhdr_478_io_en),
    .io_scan_mode(rvclkhdr_478_io_scan_mode)
  );
  rvclkhdr rvclkhdr_479 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_479_io_l1clk),
    .io_clk(rvclkhdr_479_io_clk),
    .io_en(rvclkhdr_479_io_en),
    .io_scan_mode(rvclkhdr_479_io_scan_mode)
  );
  rvclkhdr rvclkhdr_480 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_480_io_l1clk),
    .io_clk(rvclkhdr_480_io_clk),
    .io_en(rvclkhdr_480_io_en),
    .io_scan_mode(rvclkhdr_480_io_scan_mode)
  );
  rvclkhdr rvclkhdr_481 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_481_io_l1clk),
    .io_clk(rvclkhdr_481_io_clk),
    .io_en(rvclkhdr_481_io_en),
    .io_scan_mode(rvclkhdr_481_io_scan_mode)
  );
  rvclkhdr rvclkhdr_482 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_482_io_l1clk),
    .io_clk(rvclkhdr_482_io_clk),
    .io_en(rvclkhdr_482_io_en),
    .io_scan_mode(rvclkhdr_482_io_scan_mode)
  );
  rvclkhdr rvclkhdr_483 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_483_io_l1clk),
    .io_clk(rvclkhdr_483_io_clk),
    .io_en(rvclkhdr_483_io_en),
    .io_scan_mode(rvclkhdr_483_io_scan_mode)
  );
  rvclkhdr rvclkhdr_484 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_484_io_l1clk),
    .io_clk(rvclkhdr_484_io_clk),
    .io_en(rvclkhdr_484_io_en),
    .io_scan_mode(rvclkhdr_484_io_scan_mode)
  );
  rvclkhdr rvclkhdr_485 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_485_io_l1clk),
    .io_clk(rvclkhdr_485_io_clk),
    .io_en(rvclkhdr_485_io_en),
    .io_scan_mode(rvclkhdr_485_io_scan_mode)
  );
  rvclkhdr rvclkhdr_486 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_486_io_l1clk),
    .io_clk(rvclkhdr_486_io_clk),
    .io_en(rvclkhdr_486_io_en),
    .io_scan_mode(rvclkhdr_486_io_scan_mode)
  );
  rvclkhdr rvclkhdr_487 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_487_io_l1clk),
    .io_clk(rvclkhdr_487_io_clk),
    .io_en(rvclkhdr_487_io_en),
    .io_scan_mode(rvclkhdr_487_io_scan_mode)
  );
  rvclkhdr rvclkhdr_488 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_488_io_l1clk),
    .io_clk(rvclkhdr_488_io_clk),
    .io_en(rvclkhdr_488_io_en),
    .io_scan_mode(rvclkhdr_488_io_scan_mode)
  );
  rvclkhdr rvclkhdr_489 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_489_io_l1clk),
    .io_clk(rvclkhdr_489_io_clk),
    .io_en(rvclkhdr_489_io_en),
    .io_scan_mode(rvclkhdr_489_io_scan_mode)
  );
  rvclkhdr rvclkhdr_490 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_490_io_l1clk),
    .io_clk(rvclkhdr_490_io_clk),
    .io_en(rvclkhdr_490_io_en),
    .io_scan_mode(rvclkhdr_490_io_scan_mode)
  );
  rvclkhdr rvclkhdr_491 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_491_io_l1clk),
    .io_clk(rvclkhdr_491_io_clk),
    .io_en(rvclkhdr_491_io_en),
    .io_scan_mode(rvclkhdr_491_io_scan_mode)
  );
  rvclkhdr rvclkhdr_492 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_492_io_l1clk),
    .io_clk(rvclkhdr_492_io_clk),
    .io_en(rvclkhdr_492_io_en),
    .io_scan_mode(rvclkhdr_492_io_scan_mode)
  );
  rvclkhdr rvclkhdr_493 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_493_io_l1clk),
    .io_clk(rvclkhdr_493_io_clk),
    .io_en(rvclkhdr_493_io_en),
    .io_scan_mode(rvclkhdr_493_io_scan_mode)
  );
  rvclkhdr rvclkhdr_494 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_494_io_l1clk),
    .io_clk(rvclkhdr_494_io_clk),
    .io_en(rvclkhdr_494_io_en),
    .io_scan_mode(rvclkhdr_494_io_scan_mode)
  );
  rvclkhdr rvclkhdr_495 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_495_io_l1clk),
    .io_clk(rvclkhdr_495_io_clk),
    .io_en(rvclkhdr_495_io_en),
    .io_scan_mode(rvclkhdr_495_io_scan_mode)
  );
  rvclkhdr rvclkhdr_496 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_496_io_l1clk),
    .io_clk(rvclkhdr_496_io_clk),
    .io_en(rvclkhdr_496_io_en),
    .io_scan_mode(rvclkhdr_496_io_scan_mode)
  );
  rvclkhdr rvclkhdr_497 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_497_io_l1clk),
    .io_clk(rvclkhdr_497_io_clk),
    .io_en(rvclkhdr_497_io_en),
    .io_scan_mode(rvclkhdr_497_io_scan_mode)
  );
  rvclkhdr rvclkhdr_498 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_498_io_l1clk),
    .io_clk(rvclkhdr_498_io_clk),
    .io_en(rvclkhdr_498_io_en),
    .io_scan_mode(rvclkhdr_498_io_scan_mode)
  );
  rvclkhdr rvclkhdr_499 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_499_io_l1clk),
    .io_clk(rvclkhdr_499_io_clk),
    .io_en(rvclkhdr_499_io_en),
    .io_scan_mode(rvclkhdr_499_io_scan_mode)
  );
  rvclkhdr rvclkhdr_500 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_500_io_l1clk),
    .io_clk(rvclkhdr_500_io_clk),
    .io_en(rvclkhdr_500_io_en),
    .io_scan_mode(rvclkhdr_500_io_scan_mode)
  );
  rvclkhdr rvclkhdr_501 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_501_io_l1clk),
    .io_clk(rvclkhdr_501_io_clk),
    .io_en(rvclkhdr_501_io_en),
    .io_scan_mode(rvclkhdr_501_io_scan_mode)
  );
  rvclkhdr rvclkhdr_502 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_502_io_l1clk),
    .io_clk(rvclkhdr_502_io_clk),
    .io_en(rvclkhdr_502_io_en),
    .io_scan_mode(rvclkhdr_502_io_scan_mode)
  );
  rvclkhdr rvclkhdr_503 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_503_io_l1clk),
    .io_clk(rvclkhdr_503_io_clk),
    .io_en(rvclkhdr_503_io_en),
    .io_scan_mode(rvclkhdr_503_io_scan_mode)
  );
  rvclkhdr rvclkhdr_504 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_504_io_l1clk),
    .io_clk(rvclkhdr_504_io_clk),
    .io_en(rvclkhdr_504_io_en),
    .io_scan_mode(rvclkhdr_504_io_scan_mode)
  );
  rvclkhdr rvclkhdr_505 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_505_io_l1clk),
    .io_clk(rvclkhdr_505_io_clk),
    .io_en(rvclkhdr_505_io_en),
    .io_scan_mode(rvclkhdr_505_io_scan_mode)
  );
  rvclkhdr rvclkhdr_506 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_506_io_l1clk),
    .io_clk(rvclkhdr_506_io_clk),
    .io_en(rvclkhdr_506_io_en),
    .io_scan_mode(rvclkhdr_506_io_scan_mode)
  );
  rvclkhdr rvclkhdr_507 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_507_io_l1clk),
    .io_clk(rvclkhdr_507_io_clk),
    .io_en(rvclkhdr_507_io_en),
    .io_scan_mode(rvclkhdr_507_io_scan_mode)
  );
  rvclkhdr rvclkhdr_508 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_508_io_l1clk),
    .io_clk(rvclkhdr_508_io_clk),
    .io_en(rvclkhdr_508_io_en),
    .io_scan_mode(rvclkhdr_508_io_scan_mode)
  );
  rvclkhdr rvclkhdr_509 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_509_io_l1clk),
    .io_clk(rvclkhdr_509_io_clk),
    .io_en(rvclkhdr_509_io_en),
    .io_scan_mode(rvclkhdr_509_io_scan_mode)
  );
  rvclkhdr rvclkhdr_510 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_510_io_l1clk),
    .io_clk(rvclkhdr_510_io_clk),
    .io_en(rvclkhdr_510_io_en),
    .io_scan_mode(rvclkhdr_510_io_scan_mode)
  );
  rvclkhdr rvclkhdr_511 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_511_io_l1clk),
    .io_clk(rvclkhdr_511_io_clk),
    .io_en(rvclkhdr_511_io_en),
    .io_scan_mode(rvclkhdr_511_io_scan_mode)
  );
  rvclkhdr rvclkhdr_512 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_512_io_l1clk),
    .io_clk(rvclkhdr_512_io_clk),
    .io_en(rvclkhdr_512_io_en),
    .io_scan_mode(rvclkhdr_512_io_scan_mode)
  );
  rvclkhdr rvclkhdr_513 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_513_io_l1clk),
    .io_clk(rvclkhdr_513_io_clk),
    .io_en(rvclkhdr_513_io_en),
    .io_scan_mode(rvclkhdr_513_io_scan_mode)
  );
  rvclkhdr rvclkhdr_514 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_514_io_l1clk),
    .io_clk(rvclkhdr_514_io_clk),
    .io_en(rvclkhdr_514_io_en),
    .io_scan_mode(rvclkhdr_514_io_scan_mode)
  );
  rvclkhdr rvclkhdr_515 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_515_io_l1clk),
    .io_clk(rvclkhdr_515_io_clk),
    .io_en(rvclkhdr_515_io_en),
    .io_scan_mode(rvclkhdr_515_io_scan_mode)
  );
  rvclkhdr rvclkhdr_516 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_516_io_l1clk),
    .io_clk(rvclkhdr_516_io_clk),
    .io_en(rvclkhdr_516_io_en),
    .io_scan_mode(rvclkhdr_516_io_scan_mode)
  );
  rvclkhdr rvclkhdr_517 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_517_io_l1clk),
    .io_clk(rvclkhdr_517_io_clk),
    .io_en(rvclkhdr_517_io_en),
    .io_scan_mode(rvclkhdr_517_io_scan_mode)
  );
  rvclkhdr rvclkhdr_518 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_518_io_l1clk),
    .io_clk(rvclkhdr_518_io_clk),
    .io_en(rvclkhdr_518_io_en),
    .io_scan_mode(rvclkhdr_518_io_scan_mode)
  );
  rvclkhdr rvclkhdr_519 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_519_io_l1clk),
    .io_clk(rvclkhdr_519_io_clk),
    .io_en(rvclkhdr_519_io_en),
    .io_scan_mode(rvclkhdr_519_io_scan_mode)
  );
  rvclkhdr rvclkhdr_520 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_520_io_l1clk),
    .io_clk(rvclkhdr_520_io_clk),
    .io_en(rvclkhdr_520_io_en),
    .io_scan_mode(rvclkhdr_520_io_scan_mode)
  );
  rvclkhdr rvclkhdr_521 ( // @[el2_lib.scala 475:23]
    .io_l1clk(rvclkhdr_521_io_l1clk),
    .io_clk(rvclkhdr_521_io_clk),
    .io_en(rvclkhdr_521_io_en),
    .io_scan_mode(rvclkhdr_521_io_scan_mode)
  );
  rvclkhdr rvclkhdr_522 ( // @[el2_lib.scala 461:22]
    .io_l1clk(rvclkhdr_522_io_l1clk),
    .io_clk(rvclkhdr_522_io_clk),
    .io_en(rvclkhdr_522_io_en),
    .io_scan_mode(rvclkhdr_522_io_scan_mode)
  );
  rvclkhdr rvclkhdr_523 ( // @[el2_lib.scala 461:22]
    .io_l1clk(rvclkhdr_523_io_l1clk),
    .io_clk(rvclkhdr_523_io_clk),
    .io_en(rvclkhdr_523_io_en),
    .io_scan_mode(rvclkhdr_523_io_scan_mode)
  );
  rvclkhdr rvclkhdr_524 ( // @[el2_lib.scala 461:22]
    .io_l1clk(rvclkhdr_524_io_l1clk),
    .io_clk(rvclkhdr_524_io_clk),
    .io_en(rvclkhdr_524_io_en),
    .io_scan_mode(rvclkhdr_524_io_scan_mode)
  );
  rvclkhdr rvclkhdr_525 ( // @[el2_lib.scala 461:22]
    .io_l1clk(rvclkhdr_525_io_l1clk),
    .io_clk(rvclkhdr_525_io_clk),
    .io_en(rvclkhdr_525_io_en),
    .io_scan_mode(rvclkhdr_525_io_scan_mode)
  );
  rvclkhdr rvclkhdr_526 ( // @[el2_lib.scala 461:22]
    .io_l1clk(rvclkhdr_526_io_l1clk),
    .io_clk(rvclkhdr_526_io_clk),
    .io_en(rvclkhdr_526_io_en),
    .io_scan_mode(rvclkhdr_526_io_scan_mode)
  );
  rvclkhdr rvclkhdr_527 ( // @[el2_lib.scala 461:22]
    .io_l1clk(rvclkhdr_527_io_l1clk),
    .io_clk(rvclkhdr_527_io_clk),
    .io_en(rvclkhdr_527_io_en),
    .io_scan_mode(rvclkhdr_527_io_scan_mode)
  );
  rvclkhdr rvclkhdr_528 ( // @[el2_lib.scala 461:22]
    .io_l1clk(rvclkhdr_528_io_l1clk),
    .io_clk(rvclkhdr_528_io_clk),
    .io_en(rvclkhdr_528_io_en),
    .io_scan_mode(rvclkhdr_528_io_scan_mode)
  );
  rvclkhdr rvclkhdr_529 ( // @[el2_lib.scala 461:22]
    .io_l1clk(rvclkhdr_529_io_l1clk),
    .io_clk(rvclkhdr_529_io_clk),
    .io_en(rvclkhdr_529_io_en),
    .io_scan_mode(rvclkhdr_529_io_scan_mode)
  );
  rvclkhdr rvclkhdr_530 ( // @[el2_lib.scala 461:22]
    .io_l1clk(rvclkhdr_530_io_l1clk),
    .io_clk(rvclkhdr_530_io_clk),
    .io_en(rvclkhdr_530_io_en),
    .io_scan_mode(rvclkhdr_530_io_scan_mode)
  );
  rvclkhdr rvclkhdr_531 ( // @[el2_lib.scala 461:22]
    .io_l1clk(rvclkhdr_531_io_l1clk),
    .io_clk(rvclkhdr_531_io_clk),
    .io_en(rvclkhdr_531_io_en),
    .io_scan_mode(rvclkhdr_531_io_scan_mode)
  );
  rvclkhdr rvclkhdr_532 ( // @[el2_lib.scala 461:22]
    .io_l1clk(rvclkhdr_532_io_l1clk),
    .io_clk(rvclkhdr_532_io_clk),
    .io_en(rvclkhdr_532_io_en),
    .io_scan_mode(rvclkhdr_532_io_scan_mode)
  );
  rvclkhdr rvclkhdr_533 ( // @[el2_lib.scala 461:22]
    .io_l1clk(rvclkhdr_533_io_l1clk),
    .io_clk(rvclkhdr_533_io_clk),
    .io_en(rvclkhdr_533_io_en),
    .io_scan_mode(rvclkhdr_533_io_scan_mode)
  );
  rvclkhdr rvclkhdr_534 ( // @[el2_lib.scala 461:22]
    .io_l1clk(rvclkhdr_534_io_l1clk),
    .io_clk(rvclkhdr_534_io_clk),
    .io_en(rvclkhdr_534_io_en),
    .io_scan_mode(rvclkhdr_534_io_scan_mode)
  );
  rvclkhdr rvclkhdr_535 ( // @[el2_lib.scala 461:22]
    .io_l1clk(rvclkhdr_535_io_l1clk),
    .io_clk(rvclkhdr_535_io_clk),
    .io_en(rvclkhdr_535_io_en),
    .io_scan_mode(rvclkhdr_535_io_scan_mode)
  );
  rvclkhdr rvclkhdr_536 ( // @[el2_lib.scala 461:22]
    .io_l1clk(rvclkhdr_536_io_l1clk),
    .io_clk(rvclkhdr_536_io_clk),
    .io_en(rvclkhdr_536_io_en),
    .io_scan_mode(rvclkhdr_536_io_scan_mode)
  );
  rvclkhdr rvclkhdr_537 ( // @[el2_lib.scala 461:22]
    .io_l1clk(rvclkhdr_537_io_l1clk),
    .io_clk(rvclkhdr_537_io_clk),
    .io_en(rvclkhdr_537_io_en),
    .io_scan_mode(rvclkhdr_537_io_scan_mode)
  );
  rvclkhdr rvclkhdr_538 ( // @[el2_lib.scala 461:22]
    .io_l1clk(rvclkhdr_538_io_l1clk),
    .io_clk(rvclkhdr_538_io_clk),
    .io_en(rvclkhdr_538_io_en),
    .io_scan_mode(rvclkhdr_538_io_scan_mode)
  );
  rvclkhdr rvclkhdr_539 ( // @[el2_lib.scala 461:22]
    .io_l1clk(rvclkhdr_539_io_l1clk),
    .io_clk(rvclkhdr_539_io_clk),
    .io_en(rvclkhdr_539_io_en),
    .io_scan_mode(rvclkhdr_539_io_scan_mode)
  );
  rvclkhdr rvclkhdr_540 ( // @[el2_lib.scala 461:22]
    .io_l1clk(rvclkhdr_540_io_l1clk),
    .io_clk(rvclkhdr_540_io_clk),
    .io_en(rvclkhdr_540_io_en),
    .io_scan_mode(rvclkhdr_540_io_scan_mode)
  );
  rvclkhdr rvclkhdr_541 ( // @[el2_lib.scala 461:22]
    .io_l1clk(rvclkhdr_541_io_l1clk),
    .io_clk(rvclkhdr_541_io_clk),
    .io_en(rvclkhdr_541_io_en),
    .io_scan_mode(rvclkhdr_541_io_scan_mode)
  );
  rvclkhdr rvclkhdr_542 ( // @[el2_lib.scala 461:22]
    .io_l1clk(rvclkhdr_542_io_l1clk),
    .io_clk(rvclkhdr_542_io_clk),
    .io_en(rvclkhdr_542_io_en),
    .io_scan_mode(rvclkhdr_542_io_scan_mode)
  );
  rvclkhdr rvclkhdr_543 ( // @[el2_lib.scala 461:22]
    .io_l1clk(rvclkhdr_543_io_l1clk),
    .io_clk(rvclkhdr_543_io_clk),
    .io_en(rvclkhdr_543_io_en),
    .io_scan_mode(rvclkhdr_543_io_scan_mode)
  );
  rvclkhdr rvclkhdr_544 ( // @[el2_lib.scala 461:22]
    .io_l1clk(rvclkhdr_544_io_l1clk),
    .io_clk(rvclkhdr_544_io_clk),
    .io_en(rvclkhdr_544_io_en),
    .io_scan_mode(rvclkhdr_544_io_scan_mode)
  );
  rvclkhdr rvclkhdr_545 ( // @[el2_lib.scala 461:22]
    .io_l1clk(rvclkhdr_545_io_l1clk),
    .io_clk(rvclkhdr_545_io_clk),
    .io_en(rvclkhdr_545_io_en),
    .io_scan_mode(rvclkhdr_545_io_scan_mode)
  );
  rvclkhdr rvclkhdr_546 ( // @[el2_lib.scala 461:22]
    .io_l1clk(rvclkhdr_546_io_l1clk),
    .io_clk(rvclkhdr_546_io_clk),
    .io_en(rvclkhdr_546_io_en),
    .io_scan_mode(rvclkhdr_546_io_scan_mode)
  );
  rvclkhdr rvclkhdr_547 ( // @[el2_lib.scala 461:22]
    .io_l1clk(rvclkhdr_547_io_l1clk),
    .io_clk(rvclkhdr_547_io_clk),
    .io_en(rvclkhdr_547_io_en),
    .io_scan_mode(rvclkhdr_547_io_scan_mode)
  );
  rvclkhdr rvclkhdr_548 ( // @[el2_lib.scala 461:22]
    .io_l1clk(rvclkhdr_548_io_l1clk),
    .io_clk(rvclkhdr_548_io_clk),
    .io_en(rvclkhdr_548_io_en),
    .io_scan_mode(rvclkhdr_548_io_scan_mode)
  );
  rvclkhdr rvclkhdr_549 ( // @[el2_lib.scala 461:22]
    .io_l1clk(rvclkhdr_549_io_l1clk),
    .io_clk(rvclkhdr_549_io_clk),
    .io_en(rvclkhdr_549_io_en),
    .io_scan_mode(rvclkhdr_549_io_scan_mode)
  );
  rvclkhdr rvclkhdr_550 ( // @[el2_lib.scala 461:22]
    .io_l1clk(rvclkhdr_550_io_l1clk),
    .io_clk(rvclkhdr_550_io_clk),
    .io_en(rvclkhdr_550_io_en),
    .io_scan_mode(rvclkhdr_550_io_scan_mode)
  );
  rvclkhdr rvclkhdr_551 ( // @[el2_lib.scala 461:22]
    .io_l1clk(rvclkhdr_551_io_l1clk),
    .io_clk(rvclkhdr_551_io_clk),
    .io_en(rvclkhdr_551_io_en),
    .io_scan_mode(rvclkhdr_551_io_scan_mode)
  );
  rvclkhdr rvclkhdr_552 ( // @[el2_lib.scala 461:22]
    .io_l1clk(rvclkhdr_552_io_l1clk),
    .io_clk(rvclkhdr_552_io_clk),
    .io_en(rvclkhdr_552_io_en),
    .io_scan_mode(rvclkhdr_552_io_scan_mode)
  );
  rvclkhdr rvclkhdr_553 ( // @[el2_lib.scala 461:22]
    .io_l1clk(rvclkhdr_553_io_l1clk),
    .io_clk(rvclkhdr_553_io_clk),
    .io_en(rvclkhdr_553_io_en),
    .io_scan_mode(rvclkhdr_553_io_scan_mode)
  );
  assign io_ifu_bp_hit_taken_f = _T_237 & _T_238; // @[el2_ifu_bp_ctl.scala 273:25]
  assign io_ifu_bp_btb_target_f = _T_428 ? rets_out_0[31:1] : bp_btb_target_adder_f[31:1]; // @[el2_ifu_bp_ctl.scala 369:26]
  assign io_ifu_bp_inst_mask_f = _T_274 | _T_275; // @[el2_ifu_bp_ctl.scala 297:25]
  assign io_ifu_bp_fghr_f = fghr; // @[el2_ifu_bp_ctl.scala 337:20]
  assign io_ifu_bp_way_f = tag_match_vway1_expanded_f | _T_212; // @[el2_ifu_bp_ctl.scala 247:19]
  assign io_ifu_bp_ret_f = {_T_294,_T_300}; // @[el2_ifu_bp_ctl.scala 343:19]
  assign io_ifu_bp_hist1_f = bht_force_taken_f | _T_279; // @[el2_ifu_bp_ctl.scala 338:21]
  assign io_ifu_bp_hist0_f = {bht_vbank1_rd_data_f[0],bht_vbank0_rd_data_f[0]}; // @[el2_ifu_bp_ctl.scala 339:21]
  assign io_ifu_bp_pc4_f = {_T_285,_T_288}; // @[el2_ifu_bp_ctl.scala 340:19]
  assign io_ifu_bp_valid_f = vwayhit_f & _T_344; // @[el2_ifu_bp_ctl.scala 342:21]
  assign io_ifu_bp_poffset_f = btb_sel_data_f[15:4]; // @[el2_ifu_bp_ctl.scala 356:23]
  assign io_test = btb_lru_b0_f; // @[el2_ifu_bp_ctl.scala 68:11]
  assign rvclkhdr_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_io_en = io_ifc_fetch_req_f | exu_mp_valid; // @[el2_lib.scala 478:17]
  assign rvclkhdr_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_1_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_1_io_en = _T_375 & io_ic_hit_f; // @[el2_lib.scala 478:17]
  assign rvclkhdr_1_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_2_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_2_io_en = ~rs_hold; // @[el2_lib.scala 478:17]
  assign rvclkhdr_2_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_3_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_3_io_en = rs_push | rs_pop; // @[el2_lib.scala 478:17]
  assign rvclkhdr_3_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_4_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_4_io_en = rs_push | rs_pop; // @[el2_lib.scala 478:17]
  assign rvclkhdr_4_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_5_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_5_io_en = rs_push | rs_pop; // @[el2_lib.scala 478:17]
  assign rvclkhdr_5_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_6_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_6_io_en = rs_push | rs_pop; // @[el2_lib.scala 478:17]
  assign rvclkhdr_6_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_7_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_7_io_en = rs_push | rs_pop; // @[el2_lib.scala 478:17]
  assign rvclkhdr_7_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_8_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_8_io_en = rs_push | rs_pop; // @[el2_lib.scala 478:17]
  assign rvclkhdr_8_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_9_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_9_io_en = _T_472 & io_ifu_bp_hit_taken_f; // @[el2_lib.scala 478:17]
  assign rvclkhdr_9_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_10_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_10_io_en = _T_575 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_10_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_11_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_11_io_en = _T_578 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_11_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_12_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_12_io_en = _T_581 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_12_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_13_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_13_io_en = _T_584 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_13_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_14_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_14_io_en = _T_587 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_14_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_15_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_15_io_en = _T_590 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_15_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_16_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_16_io_en = _T_593 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_16_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_17_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_17_io_en = _T_596 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_17_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_18_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_18_io_en = _T_599 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_18_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_19_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_19_io_en = _T_602 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_19_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_20_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_20_io_en = _T_605 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_20_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_21_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_21_io_en = _T_608 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_21_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_22_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_22_io_en = _T_611 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_22_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_23_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_23_io_en = _T_614 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_23_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_24_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_24_io_en = _T_617 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_24_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_25_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_25_io_en = _T_620 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_25_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_26_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_26_io_en = _T_623 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_26_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_27_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_27_io_en = _T_626 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_27_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_28_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_28_io_en = _T_629 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_28_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_29_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_29_io_en = _T_632 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_29_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_30_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_30_io_en = _T_635 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_30_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_31_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_31_io_en = _T_638 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_31_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_32_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_32_io_en = _T_641 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_32_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_33_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_33_io_en = _T_644 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_33_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_34_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_34_io_en = _T_647 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_34_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_35_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_35_io_en = _T_650 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_35_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_36_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_36_io_en = _T_653 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_36_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_37_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_37_io_en = _T_656 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_37_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_38_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_38_io_en = _T_659 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_38_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_39_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_39_io_en = _T_662 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_39_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_40_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_40_io_en = _T_665 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_40_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_41_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_41_io_en = _T_668 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_41_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_42_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_42_io_en = _T_671 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_42_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_43_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_43_io_en = _T_674 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_43_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_44_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_44_io_en = _T_677 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_44_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_45_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_45_io_en = _T_680 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_45_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_46_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_46_io_en = _T_683 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_46_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_47_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_47_io_en = _T_686 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_47_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_48_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_48_io_en = _T_689 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_48_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_49_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_49_io_en = _T_692 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_49_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_50_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_50_io_en = _T_695 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_50_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_51_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_51_io_en = _T_698 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_51_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_52_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_52_io_en = _T_701 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_52_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_53_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_53_io_en = _T_704 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_53_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_54_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_54_io_en = _T_707 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_54_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_55_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_55_io_en = _T_710 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_55_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_56_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_56_io_en = _T_713 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_56_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_57_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_57_io_en = _T_716 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_57_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_58_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_58_io_en = _T_719 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_58_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_59_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_59_io_en = _T_722 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_59_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_60_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_60_io_en = _T_725 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_60_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_61_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_61_io_en = _T_728 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_61_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_62_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_62_io_en = _T_731 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_62_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_63_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_63_io_en = _T_734 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_63_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_64_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_64_io_en = _T_737 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_64_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_65_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_65_io_en = _T_740 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_65_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_66_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_66_io_en = _T_743 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_66_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_67_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_67_io_en = _T_746 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_67_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_68_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_68_io_en = _T_749 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_68_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_69_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_69_io_en = _T_752 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_69_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_70_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_70_io_en = _T_755 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_70_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_71_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_71_io_en = _T_758 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_71_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_72_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_72_io_en = _T_761 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_72_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_73_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_73_io_en = _T_764 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_73_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_74_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_74_io_en = _T_767 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_74_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_75_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_75_io_en = _T_770 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_75_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_76_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_76_io_en = _T_773 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_76_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_77_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_77_io_en = _T_776 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_77_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_78_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_78_io_en = _T_779 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_78_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_79_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_79_io_en = _T_782 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_79_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_80_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_80_io_en = _T_785 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_80_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_81_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_81_io_en = _T_788 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_81_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_82_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_82_io_en = _T_791 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_82_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_83_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_83_io_en = _T_794 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_83_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_84_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_84_io_en = _T_797 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_84_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_85_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_85_io_en = _T_800 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_85_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_86_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_86_io_en = _T_803 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_86_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_87_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_87_io_en = _T_806 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_87_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_88_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_88_io_en = _T_809 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_88_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_89_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_89_io_en = _T_812 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_89_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_90_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_90_io_en = _T_815 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_90_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_91_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_91_io_en = _T_818 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_91_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_92_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_92_io_en = _T_821 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_92_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_93_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_93_io_en = _T_824 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_93_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_94_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_94_io_en = _T_827 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_94_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_95_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_95_io_en = _T_830 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_95_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_96_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_96_io_en = _T_833 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_96_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_97_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_97_io_en = _T_836 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_97_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_98_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_98_io_en = _T_839 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_98_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_99_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_99_io_en = _T_842 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_99_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_100_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_100_io_en = _T_845 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_100_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_101_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_101_io_en = _T_848 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_101_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_102_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_102_io_en = _T_851 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_102_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_103_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_103_io_en = _T_854 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_103_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_104_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_104_io_en = _T_857 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_104_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_105_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_105_io_en = _T_860 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_105_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_106_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_106_io_en = _T_863 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_106_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_107_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_107_io_en = _T_866 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_107_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_108_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_108_io_en = _T_869 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_108_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_109_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_109_io_en = _T_872 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_109_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_110_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_110_io_en = _T_875 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_110_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_111_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_111_io_en = _T_878 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_111_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_112_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_112_io_en = _T_881 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_112_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_113_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_113_io_en = _T_884 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_113_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_114_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_114_io_en = _T_887 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_114_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_115_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_115_io_en = _T_890 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_115_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_116_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_116_io_en = _T_893 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_116_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_117_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_117_io_en = _T_896 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_117_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_118_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_118_io_en = _T_899 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_118_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_119_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_119_io_en = _T_902 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_119_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_120_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_120_io_en = _T_905 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_120_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_121_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_121_io_en = _T_908 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_121_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_122_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_122_io_en = _T_911 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_122_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_123_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_123_io_en = _T_914 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_123_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_124_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_124_io_en = _T_917 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_124_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_125_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_125_io_en = _T_920 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_125_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_126_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_126_io_en = _T_923 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_126_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_127_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_127_io_en = _T_926 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_127_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_128_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_128_io_en = _T_929 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_128_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_129_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_129_io_en = _T_932 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_129_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_130_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_130_io_en = _T_935 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_130_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_131_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_131_io_en = _T_938 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_131_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_132_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_132_io_en = _T_941 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_132_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_133_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_133_io_en = _T_944 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_133_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_134_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_134_io_en = _T_947 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_134_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_135_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_135_io_en = _T_950 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_135_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_136_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_136_io_en = _T_953 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_136_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_137_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_137_io_en = _T_956 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_137_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_138_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_138_io_en = _T_959 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_138_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_139_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_139_io_en = _T_962 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_139_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_140_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_140_io_en = _T_965 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_140_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_141_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_141_io_en = _T_968 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_141_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_142_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_142_io_en = _T_971 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_142_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_143_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_143_io_en = _T_974 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_143_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_144_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_144_io_en = _T_977 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_144_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_145_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_145_io_en = _T_980 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_145_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_146_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_146_io_en = _T_983 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_146_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_147_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_147_io_en = _T_986 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_147_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_148_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_148_io_en = _T_989 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_148_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_149_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_149_io_en = _T_992 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_149_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_150_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_150_io_en = _T_995 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_150_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_151_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_151_io_en = _T_998 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_151_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_152_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_152_io_en = _T_1001 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_152_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_153_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_153_io_en = _T_1004 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_153_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_154_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_154_io_en = _T_1007 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_154_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_155_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_155_io_en = _T_1010 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_155_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_156_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_156_io_en = _T_1013 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_156_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_157_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_157_io_en = _T_1016 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_157_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_158_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_158_io_en = _T_1019 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_158_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_159_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_159_io_en = _T_1022 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_159_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_160_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_160_io_en = _T_1025 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_160_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_161_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_161_io_en = _T_1028 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_161_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_162_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_162_io_en = _T_1031 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_162_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_163_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_163_io_en = _T_1034 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_163_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_164_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_164_io_en = _T_1037 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_164_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_165_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_165_io_en = _T_1040 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_165_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_166_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_166_io_en = _T_1043 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_166_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_167_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_167_io_en = _T_1046 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_167_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_168_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_168_io_en = _T_1049 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_168_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_169_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_169_io_en = _T_1052 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_169_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_170_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_170_io_en = _T_1055 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_170_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_171_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_171_io_en = _T_1058 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_171_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_172_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_172_io_en = _T_1061 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_172_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_173_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_173_io_en = _T_1064 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_173_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_174_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_174_io_en = _T_1067 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_174_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_175_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_175_io_en = _T_1070 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_175_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_176_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_176_io_en = _T_1073 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_176_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_177_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_177_io_en = _T_1076 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_177_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_178_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_178_io_en = _T_1079 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_178_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_179_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_179_io_en = _T_1082 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_179_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_180_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_180_io_en = _T_1085 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_180_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_181_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_181_io_en = _T_1088 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_181_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_182_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_182_io_en = _T_1091 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_182_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_183_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_183_io_en = _T_1094 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_183_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_184_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_184_io_en = _T_1097 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_184_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_185_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_185_io_en = _T_1100 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_185_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_186_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_186_io_en = _T_1103 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_186_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_187_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_187_io_en = _T_1106 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_187_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_188_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_188_io_en = _T_1109 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_188_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_189_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_189_io_en = _T_1112 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_189_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_190_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_190_io_en = _T_1115 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_190_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_191_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_191_io_en = _T_1118 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_191_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_192_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_192_io_en = _T_1121 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_192_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_193_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_193_io_en = _T_1124 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_193_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_194_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_194_io_en = _T_1127 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_194_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_195_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_195_io_en = _T_1130 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_195_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_196_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_196_io_en = _T_1133 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_196_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_197_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_197_io_en = _T_1136 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_197_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_198_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_198_io_en = _T_1139 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_198_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_199_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_199_io_en = _T_1142 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_199_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_200_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_200_io_en = _T_1145 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_200_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_201_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_201_io_en = _T_1148 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_201_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_202_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_202_io_en = _T_1151 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_202_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_203_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_203_io_en = _T_1154 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_203_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_204_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_204_io_en = _T_1157 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_204_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_205_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_205_io_en = _T_1160 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_205_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_206_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_206_io_en = _T_1163 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_206_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_207_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_207_io_en = _T_1166 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_207_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_208_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_208_io_en = _T_1169 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_208_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_209_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_209_io_en = _T_1172 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_209_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_210_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_210_io_en = _T_1175 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_210_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_211_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_211_io_en = _T_1178 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_211_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_212_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_212_io_en = _T_1181 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_212_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_213_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_213_io_en = _T_1184 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_213_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_214_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_214_io_en = _T_1187 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_214_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_215_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_215_io_en = _T_1190 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_215_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_216_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_216_io_en = _T_1193 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_216_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_217_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_217_io_en = _T_1196 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_217_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_218_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_218_io_en = _T_1199 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_218_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_219_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_219_io_en = _T_1202 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_219_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_220_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_220_io_en = _T_1205 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_220_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_221_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_221_io_en = _T_1208 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_221_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_222_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_222_io_en = _T_1211 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_222_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_223_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_223_io_en = _T_1214 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_223_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_224_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_224_io_en = _T_1217 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_224_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_225_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_225_io_en = _T_1220 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_225_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_226_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_226_io_en = _T_1223 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_226_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_227_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_227_io_en = _T_1226 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_227_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_228_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_228_io_en = _T_1229 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_228_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_229_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_229_io_en = _T_1232 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_229_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_230_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_230_io_en = _T_1235 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_230_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_231_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_231_io_en = _T_1238 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_231_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_232_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_232_io_en = _T_1241 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_232_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_233_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_233_io_en = _T_1244 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_233_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_234_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_234_io_en = _T_1247 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_234_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_235_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_235_io_en = _T_1250 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_235_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_236_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_236_io_en = _T_1253 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_236_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_237_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_237_io_en = _T_1256 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_237_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_238_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_238_io_en = _T_1259 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_238_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_239_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_239_io_en = _T_1262 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_239_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_240_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_240_io_en = _T_1265 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_240_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_241_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_241_io_en = _T_1268 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_241_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_242_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_242_io_en = _T_1271 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_242_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_243_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_243_io_en = _T_1274 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_243_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_244_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_244_io_en = _T_1277 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_244_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_245_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_245_io_en = _T_1280 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_245_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_246_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_246_io_en = _T_1283 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_246_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_247_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_247_io_en = _T_1286 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_247_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_248_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_248_io_en = _T_1289 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_248_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_249_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_249_io_en = _T_1292 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_249_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_250_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_250_io_en = _T_1295 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_250_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_251_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_251_io_en = _T_1298 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_251_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_252_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_252_io_en = _T_1301 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_252_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_253_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_253_io_en = _T_1304 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_253_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_254_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_254_io_en = _T_1307 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_254_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_255_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_255_io_en = _T_1310 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_255_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_256_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_256_io_en = _T_1313 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_256_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_257_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_257_io_en = _T_1316 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_257_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_258_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_258_io_en = _T_1319 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_258_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_259_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_259_io_en = _T_1322 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_259_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_260_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_260_io_en = _T_1325 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_260_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_261_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_261_io_en = _T_1328 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_261_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_262_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_262_io_en = _T_1331 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_262_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_263_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_263_io_en = _T_1334 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_263_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_264_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_264_io_en = _T_1337 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_264_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_265_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_265_io_en = _T_1340 & btb_wr_en_way0; // @[el2_lib.scala 478:17]
  assign rvclkhdr_265_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_266_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_266_io_en = _T_575 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_266_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_267_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_267_io_en = _T_578 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_267_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_268_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_268_io_en = _T_581 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_268_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_269_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_269_io_en = _T_584 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_269_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_270_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_270_io_en = _T_587 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_270_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_271_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_271_io_en = _T_590 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_271_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_272_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_272_io_en = _T_593 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_272_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_273_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_273_io_en = _T_596 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_273_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_274_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_274_io_en = _T_599 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_274_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_275_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_275_io_en = _T_602 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_275_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_276_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_276_io_en = _T_605 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_276_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_277_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_277_io_en = _T_608 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_277_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_278_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_278_io_en = _T_611 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_278_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_279_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_279_io_en = _T_614 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_279_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_280_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_280_io_en = _T_617 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_280_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_281_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_281_io_en = _T_620 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_281_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_282_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_282_io_en = _T_623 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_282_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_283_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_283_io_en = _T_626 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_283_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_284_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_284_io_en = _T_629 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_284_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_285_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_285_io_en = _T_632 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_285_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_286_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_286_io_en = _T_635 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_286_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_287_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_287_io_en = _T_638 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_287_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_288_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_288_io_en = _T_641 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_288_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_289_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_289_io_en = _T_644 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_289_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_290_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_290_io_en = _T_647 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_290_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_291_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_291_io_en = _T_650 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_291_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_292_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_292_io_en = _T_653 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_292_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_293_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_293_io_en = _T_656 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_293_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_294_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_294_io_en = _T_659 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_294_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_295_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_295_io_en = _T_662 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_295_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_296_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_296_io_en = _T_665 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_296_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_297_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_297_io_en = _T_668 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_297_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_298_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_298_io_en = _T_671 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_298_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_299_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_299_io_en = _T_674 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_299_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_300_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_300_io_en = _T_677 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_300_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_301_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_301_io_en = _T_680 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_301_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_302_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_302_io_en = _T_683 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_302_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_303_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_303_io_en = _T_686 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_303_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_304_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_304_io_en = _T_689 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_304_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_305_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_305_io_en = _T_692 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_305_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_306_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_306_io_en = _T_695 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_306_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_307_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_307_io_en = _T_698 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_307_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_308_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_308_io_en = _T_701 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_308_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_309_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_309_io_en = _T_704 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_309_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_310_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_310_io_en = _T_707 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_310_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_311_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_311_io_en = _T_710 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_311_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_312_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_312_io_en = _T_713 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_312_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_313_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_313_io_en = _T_716 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_313_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_314_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_314_io_en = _T_719 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_314_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_315_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_315_io_en = _T_722 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_315_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_316_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_316_io_en = _T_725 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_316_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_317_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_317_io_en = _T_728 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_317_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_318_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_318_io_en = _T_731 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_318_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_319_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_319_io_en = _T_734 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_319_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_320_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_320_io_en = _T_737 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_320_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_321_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_321_io_en = _T_740 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_321_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_322_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_322_io_en = _T_743 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_322_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_323_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_323_io_en = _T_746 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_323_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_324_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_324_io_en = _T_749 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_324_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_325_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_325_io_en = _T_752 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_325_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_326_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_326_io_en = _T_755 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_326_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_327_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_327_io_en = _T_758 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_327_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_328_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_328_io_en = _T_761 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_328_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_329_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_329_io_en = _T_764 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_329_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_330_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_330_io_en = _T_767 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_330_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_331_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_331_io_en = _T_770 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_331_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_332_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_332_io_en = _T_773 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_332_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_333_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_333_io_en = _T_776 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_333_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_334_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_334_io_en = _T_779 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_334_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_335_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_335_io_en = _T_782 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_335_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_336_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_336_io_en = _T_785 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_336_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_337_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_337_io_en = _T_788 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_337_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_338_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_338_io_en = _T_791 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_338_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_339_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_339_io_en = _T_794 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_339_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_340_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_340_io_en = _T_797 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_340_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_341_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_341_io_en = _T_800 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_341_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_342_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_342_io_en = _T_803 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_342_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_343_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_343_io_en = _T_806 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_343_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_344_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_344_io_en = _T_809 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_344_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_345_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_345_io_en = _T_812 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_345_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_346_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_346_io_en = _T_815 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_346_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_347_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_347_io_en = _T_818 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_347_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_348_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_348_io_en = _T_821 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_348_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_349_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_349_io_en = _T_824 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_349_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_350_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_350_io_en = _T_827 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_350_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_351_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_351_io_en = _T_830 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_351_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_352_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_352_io_en = _T_833 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_352_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_353_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_353_io_en = _T_836 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_353_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_354_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_354_io_en = _T_839 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_354_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_355_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_355_io_en = _T_842 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_355_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_356_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_356_io_en = _T_845 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_356_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_357_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_357_io_en = _T_848 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_357_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_358_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_358_io_en = _T_851 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_358_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_359_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_359_io_en = _T_854 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_359_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_360_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_360_io_en = _T_857 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_360_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_361_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_361_io_en = _T_860 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_361_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_362_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_362_io_en = _T_863 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_362_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_363_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_363_io_en = _T_866 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_363_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_364_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_364_io_en = _T_869 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_364_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_365_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_365_io_en = _T_872 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_365_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_366_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_366_io_en = _T_875 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_366_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_367_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_367_io_en = _T_878 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_367_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_368_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_368_io_en = _T_881 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_368_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_369_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_369_io_en = _T_884 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_369_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_370_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_370_io_en = _T_887 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_370_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_371_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_371_io_en = _T_890 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_371_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_372_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_372_io_en = _T_893 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_372_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_373_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_373_io_en = _T_896 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_373_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_374_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_374_io_en = _T_899 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_374_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_375_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_375_io_en = _T_902 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_375_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_376_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_376_io_en = _T_905 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_376_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_377_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_377_io_en = _T_908 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_377_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_378_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_378_io_en = _T_911 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_378_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_379_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_379_io_en = _T_914 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_379_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_380_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_380_io_en = _T_917 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_380_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_381_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_381_io_en = _T_920 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_381_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_382_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_382_io_en = _T_923 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_382_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_383_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_383_io_en = _T_926 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_383_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_384_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_384_io_en = _T_929 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_384_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_385_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_385_io_en = _T_932 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_385_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_386_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_386_io_en = _T_935 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_386_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_387_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_387_io_en = _T_938 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_387_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_388_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_388_io_en = _T_941 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_388_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_389_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_389_io_en = _T_944 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_389_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_390_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_390_io_en = _T_947 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_390_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_391_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_391_io_en = _T_950 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_391_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_392_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_392_io_en = _T_953 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_392_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_393_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_393_io_en = _T_956 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_393_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_394_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_394_io_en = _T_959 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_394_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_395_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_395_io_en = _T_962 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_395_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_396_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_396_io_en = _T_965 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_396_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_397_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_397_io_en = _T_968 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_397_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_398_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_398_io_en = _T_971 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_398_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_399_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_399_io_en = _T_974 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_399_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_400_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_400_io_en = _T_977 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_400_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_401_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_401_io_en = _T_980 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_401_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_402_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_402_io_en = _T_983 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_402_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_403_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_403_io_en = _T_986 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_403_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_404_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_404_io_en = _T_989 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_404_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_405_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_405_io_en = _T_992 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_405_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_406_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_406_io_en = _T_995 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_406_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_407_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_407_io_en = _T_998 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_407_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_408_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_408_io_en = _T_1001 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_408_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_409_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_409_io_en = _T_1004 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_409_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_410_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_410_io_en = _T_1007 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_410_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_411_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_411_io_en = _T_1010 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_411_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_412_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_412_io_en = _T_1013 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_412_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_413_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_413_io_en = _T_1016 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_413_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_414_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_414_io_en = _T_1019 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_414_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_415_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_415_io_en = _T_1022 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_415_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_416_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_416_io_en = _T_1025 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_416_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_417_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_417_io_en = _T_1028 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_417_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_418_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_418_io_en = _T_1031 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_418_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_419_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_419_io_en = _T_1034 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_419_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_420_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_420_io_en = _T_1037 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_420_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_421_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_421_io_en = _T_1040 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_421_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_422_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_422_io_en = _T_1043 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_422_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_423_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_423_io_en = _T_1046 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_423_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_424_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_424_io_en = _T_1049 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_424_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_425_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_425_io_en = _T_1052 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_425_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_426_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_426_io_en = _T_1055 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_426_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_427_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_427_io_en = _T_1058 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_427_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_428_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_428_io_en = _T_1061 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_428_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_429_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_429_io_en = _T_1064 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_429_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_430_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_430_io_en = _T_1067 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_430_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_431_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_431_io_en = _T_1070 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_431_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_432_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_432_io_en = _T_1073 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_432_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_433_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_433_io_en = _T_1076 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_433_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_434_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_434_io_en = _T_1079 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_434_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_435_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_435_io_en = _T_1082 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_435_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_436_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_436_io_en = _T_1085 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_436_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_437_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_437_io_en = _T_1088 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_437_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_438_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_438_io_en = _T_1091 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_438_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_439_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_439_io_en = _T_1094 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_439_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_440_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_440_io_en = _T_1097 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_440_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_441_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_441_io_en = _T_1100 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_441_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_442_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_442_io_en = _T_1103 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_442_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_443_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_443_io_en = _T_1106 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_443_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_444_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_444_io_en = _T_1109 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_444_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_445_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_445_io_en = _T_1112 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_445_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_446_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_446_io_en = _T_1115 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_446_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_447_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_447_io_en = _T_1118 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_447_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_448_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_448_io_en = _T_1121 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_448_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_449_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_449_io_en = _T_1124 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_449_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_450_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_450_io_en = _T_1127 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_450_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_451_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_451_io_en = _T_1130 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_451_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_452_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_452_io_en = _T_1133 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_452_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_453_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_453_io_en = _T_1136 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_453_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_454_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_454_io_en = _T_1139 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_454_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_455_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_455_io_en = _T_1142 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_455_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_456_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_456_io_en = _T_1145 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_456_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_457_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_457_io_en = _T_1148 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_457_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_458_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_458_io_en = _T_1151 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_458_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_459_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_459_io_en = _T_1154 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_459_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_460_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_460_io_en = _T_1157 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_460_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_461_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_461_io_en = _T_1160 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_461_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_462_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_462_io_en = _T_1163 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_462_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_463_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_463_io_en = _T_1166 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_463_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_464_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_464_io_en = _T_1169 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_464_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_465_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_465_io_en = _T_1172 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_465_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_466_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_466_io_en = _T_1175 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_466_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_467_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_467_io_en = _T_1178 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_467_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_468_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_468_io_en = _T_1181 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_468_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_469_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_469_io_en = _T_1184 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_469_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_470_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_470_io_en = _T_1187 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_470_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_471_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_471_io_en = _T_1190 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_471_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_472_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_472_io_en = _T_1193 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_472_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_473_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_473_io_en = _T_1196 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_473_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_474_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_474_io_en = _T_1199 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_474_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_475_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_475_io_en = _T_1202 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_475_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_476_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_476_io_en = _T_1205 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_476_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_477_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_477_io_en = _T_1208 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_477_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_478_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_478_io_en = _T_1211 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_478_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_479_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_479_io_en = _T_1214 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_479_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_480_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_480_io_en = _T_1217 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_480_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_481_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_481_io_en = _T_1220 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_481_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_482_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_482_io_en = _T_1223 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_482_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_483_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_483_io_en = _T_1226 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_483_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_484_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_484_io_en = _T_1229 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_484_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_485_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_485_io_en = _T_1232 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_485_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_486_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_486_io_en = _T_1235 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_486_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_487_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_487_io_en = _T_1238 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_487_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_488_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_488_io_en = _T_1241 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_488_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_489_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_489_io_en = _T_1244 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_489_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_490_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_490_io_en = _T_1247 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_490_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_491_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_491_io_en = _T_1250 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_491_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_492_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_492_io_en = _T_1253 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_492_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_493_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_493_io_en = _T_1256 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_493_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_494_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_494_io_en = _T_1259 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_494_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_495_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_495_io_en = _T_1262 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_495_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_496_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_496_io_en = _T_1265 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_496_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_497_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_497_io_en = _T_1268 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_497_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_498_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_498_io_en = _T_1271 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_498_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_499_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_499_io_en = _T_1274 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_499_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_500_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_500_io_en = _T_1277 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_500_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_501_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_501_io_en = _T_1280 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_501_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_502_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_502_io_en = _T_1283 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_502_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_503_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_503_io_en = _T_1286 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_503_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_504_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_504_io_en = _T_1289 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_504_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_505_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_505_io_en = _T_1292 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_505_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_506_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_506_io_en = _T_1295 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_506_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_507_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_507_io_en = _T_1298 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_507_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_508_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_508_io_en = _T_1301 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_508_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_509_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_509_io_en = _T_1304 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_509_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_510_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_510_io_en = _T_1307 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_510_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_511_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_511_io_en = _T_1310 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_511_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_512_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_512_io_en = _T_1313 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_512_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_513_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_513_io_en = _T_1316 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_513_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_514_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_514_io_en = _T_1319 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_514_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_515_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_515_io_en = _T_1322 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_515_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_516_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_516_io_en = _T_1325 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_516_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_517_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_517_io_en = _T_1328 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_517_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_518_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_518_io_en = _T_1331 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_518_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_519_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_519_io_en = _T_1334 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_519_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_520_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_520_io_en = _T_1337 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_520_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_521_io_clk = clock; // @[el2_lib.scala 477:18]
  assign rvclkhdr_521_io_en = _T_1340 & btb_wr_en_way1; // @[el2_lib.scala 478:17]
  assign rvclkhdr_521_io_scan_mode = io_scan_mode; // @[el2_lib.scala 479:24]
  assign rvclkhdr_522_io_clk = clock; // @[el2_lib.scala 462:17]
  assign rvclkhdr_522_io_en = _T_6211 | _T_6216; // @[el2_lib.scala 463:16]
  assign rvclkhdr_522_io_scan_mode = io_scan_mode; // @[el2_lib.scala 464:23]
  assign rvclkhdr_523_io_clk = clock; // @[el2_lib.scala 462:17]
  assign rvclkhdr_523_io_en = _T_6222 | _T_6227; // @[el2_lib.scala 463:16]
  assign rvclkhdr_523_io_scan_mode = io_scan_mode; // @[el2_lib.scala 464:23]
  assign rvclkhdr_524_io_clk = clock; // @[el2_lib.scala 462:17]
  assign rvclkhdr_524_io_en = _T_6233 | _T_6238; // @[el2_lib.scala 463:16]
  assign rvclkhdr_524_io_scan_mode = io_scan_mode; // @[el2_lib.scala 464:23]
  assign rvclkhdr_525_io_clk = clock; // @[el2_lib.scala 462:17]
  assign rvclkhdr_525_io_en = _T_6244 | _T_6249; // @[el2_lib.scala 463:16]
  assign rvclkhdr_525_io_scan_mode = io_scan_mode; // @[el2_lib.scala 464:23]
  assign rvclkhdr_526_io_clk = clock; // @[el2_lib.scala 462:17]
  assign rvclkhdr_526_io_en = _T_6255 | _T_6260; // @[el2_lib.scala 463:16]
  assign rvclkhdr_526_io_scan_mode = io_scan_mode; // @[el2_lib.scala 464:23]
  assign rvclkhdr_527_io_clk = clock; // @[el2_lib.scala 462:17]
  assign rvclkhdr_527_io_en = _T_6266 | _T_6271; // @[el2_lib.scala 463:16]
  assign rvclkhdr_527_io_scan_mode = io_scan_mode; // @[el2_lib.scala 464:23]
  assign rvclkhdr_528_io_clk = clock; // @[el2_lib.scala 462:17]
  assign rvclkhdr_528_io_en = _T_6277 | _T_6282; // @[el2_lib.scala 463:16]
  assign rvclkhdr_528_io_scan_mode = io_scan_mode; // @[el2_lib.scala 464:23]
  assign rvclkhdr_529_io_clk = clock; // @[el2_lib.scala 462:17]
  assign rvclkhdr_529_io_en = _T_6288 | _T_6293; // @[el2_lib.scala 463:16]
  assign rvclkhdr_529_io_scan_mode = io_scan_mode; // @[el2_lib.scala 464:23]
  assign rvclkhdr_530_io_clk = clock; // @[el2_lib.scala 462:17]
  assign rvclkhdr_530_io_en = _T_6299 | _T_6304; // @[el2_lib.scala 463:16]
  assign rvclkhdr_530_io_scan_mode = io_scan_mode; // @[el2_lib.scala 464:23]
  assign rvclkhdr_531_io_clk = clock; // @[el2_lib.scala 462:17]
  assign rvclkhdr_531_io_en = _T_6310 | _T_6315; // @[el2_lib.scala 463:16]
  assign rvclkhdr_531_io_scan_mode = io_scan_mode; // @[el2_lib.scala 464:23]
  assign rvclkhdr_532_io_clk = clock; // @[el2_lib.scala 462:17]
  assign rvclkhdr_532_io_en = _T_6321 | _T_6326; // @[el2_lib.scala 463:16]
  assign rvclkhdr_532_io_scan_mode = io_scan_mode; // @[el2_lib.scala 464:23]
  assign rvclkhdr_533_io_clk = clock; // @[el2_lib.scala 462:17]
  assign rvclkhdr_533_io_en = _T_6332 | _T_6337; // @[el2_lib.scala 463:16]
  assign rvclkhdr_533_io_scan_mode = io_scan_mode; // @[el2_lib.scala 464:23]
  assign rvclkhdr_534_io_clk = clock; // @[el2_lib.scala 462:17]
  assign rvclkhdr_534_io_en = _T_6343 | _T_6348; // @[el2_lib.scala 463:16]
  assign rvclkhdr_534_io_scan_mode = io_scan_mode; // @[el2_lib.scala 464:23]
  assign rvclkhdr_535_io_clk = clock; // @[el2_lib.scala 462:17]
  assign rvclkhdr_535_io_en = _T_6354 | _T_6359; // @[el2_lib.scala 463:16]
  assign rvclkhdr_535_io_scan_mode = io_scan_mode; // @[el2_lib.scala 464:23]
  assign rvclkhdr_536_io_clk = clock; // @[el2_lib.scala 462:17]
  assign rvclkhdr_536_io_en = _T_6365 | _T_6370; // @[el2_lib.scala 463:16]
  assign rvclkhdr_536_io_scan_mode = io_scan_mode; // @[el2_lib.scala 464:23]
  assign rvclkhdr_537_io_clk = clock; // @[el2_lib.scala 462:17]
  assign rvclkhdr_537_io_en = _T_6376 | _T_6381; // @[el2_lib.scala 463:16]
  assign rvclkhdr_537_io_scan_mode = io_scan_mode; // @[el2_lib.scala 464:23]
  assign rvclkhdr_538_io_clk = clock; // @[el2_lib.scala 462:17]
  assign rvclkhdr_538_io_en = _T_6387 | _T_6392; // @[el2_lib.scala 463:16]
  assign rvclkhdr_538_io_scan_mode = io_scan_mode; // @[el2_lib.scala 464:23]
  assign rvclkhdr_539_io_clk = clock; // @[el2_lib.scala 462:17]
  assign rvclkhdr_539_io_en = _T_6398 | _T_6403; // @[el2_lib.scala 463:16]
  assign rvclkhdr_539_io_scan_mode = io_scan_mode; // @[el2_lib.scala 464:23]
  assign rvclkhdr_540_io_clk = clock; // @[el2_lib.scala 462:17]
  assign rvclkhdr_540_io_en = _T_6409 | _T_6414; // @[el2_lib.scala 463:16]
  assign rvclkhdr_540_io_scan_mode = io_scan_mode; // @[el2_lib.scala 464:23]
  assign rvclkhdr_541_io_clk = clock; // @[el2_lib.scala 462:17]
  assign rvclkhdr_541_io_en = _T_6420 | _T_6425; // @[el2_lib.scala 463:16]
  assign rvclkhdr_541_io_scan_mode = io_scan_mode; // @[el2_lib.scala 464:23]
  assign rvclkhdr_542_io_clk = clock; // @[el2_lib.scala 462:17]
  assign rvclkhdr_542_io_en = _T_6431 | _T_6436; // @[el2_lib.scala 463:16]
  assign rvclkhdr_542_io_scan_mode = io_scan_mode; // @[el2_lib.scala 464:23]
  assign rvclkhdr_543_io_clk = clock; // @[el2_lib.scala 462:17]
  assign rvclkhdr_543_io_en = _T_6442 | _T_6447; // @[el2_lib.scala 463:16]
  assign rvclkhdr_543_io_scan_mode = io_scan_mode; // @[el2_lib.scala 464:23]
  assign rvclkhdr_544_io_clk = clock; // @[el2_lib.scala 462:17]
  assign rvclkhdr_544_io_en = _T_6453 | _T_6458; // @[el2_lib.scala 463:16]
  assign rvclkhdr_544_io_scan_mode = io_scan_mode; // @[el2_lib.scala 464:23]
  assign rvclkhdr_545_io_clk = clock; // @[el2_lib.scala 462:17]
  assign rvclkhdr_545_io_en = _T_6464 | _T_6469; // @[el2_lib.scala 463:16]
  assign rvclkhdr_545_io_scan_mode = io_scan_mode; // @[el2_lib.scala 464:23]
  assign rvclkhdr_546_io_clk = clock; // @[el2_lib.scala 462:17]
  assign rvclkhdr_546_io_en = _T_6475 | _T_6480; // @[el2_lib.scala 463:16]
  assign rvclkhdr_546_io_scan_mode = io_scan_mode; // @[el2_lib.scala 464:23]
  assign rvclkhdr_547_io_clk = clock; // @[el2_lib.scala 462:17]
  assign rvclkhdr_547_io_en = _T_6486 | _T_6491; // @[el2_lib.scala 463:16]
  assign rvclkhdr_547_io_scan_mode = io_scan_mode; // @[el2_lib.scala 464:23]
  assign rvclkhdr_548_io_clk = clock; // @[el2_lib.scala 462:17]
  assign rvclkhdr_548_io_en = _T_6497 | _T_6502; // @[el2_lib.scala 463:16]
  assign rvclkhdr_548_io_scan_mode = io_scan_mode; // @[el2_lib.scala 464:23]
  assign rvclkhdr_549_io_clk = clock; // @[el2_lib.scala 462:17]
  assign rvclkhdr_549_io_en = _T_6508 | _T_6513; // @[el2_lib.scala 463:16]
  assign rvclkhdr_549_io_scan_mode = io_scan_mode; // @[el2_lib.scala 464:23]
  assign rvclkhdr_550_io_clk = clock; // @[el2_lib.scala 462:17]
  assign rvclkhdr_550_io_en = _T_6519 | _T_6524; // @[el2_lib.scala 463:16]
  assign rvclkhdr_550_io_scan_mode = io_scan_mode; // @[el2_lib.scala 464:23]
  assign rvclkhdr_551_io_clk = clock; // @[el2_lib.scala 462:17]
  assign rvclkhdr_551_io_en = _T_6530 | _T_6535; // @[el2_lib.scala 463:16]
  assign rvclkhdr_551_io_scan_mode = io_scan_mode; // @[el2_lib.scala 464:23]
  assign rvclkhdr_552_io_clk = clock; // @[el2_lib.scala 462:17]
  assign rvclkhdr_552_io_en = _T_6541 | _T_6546; // @[el2_lib.scala 463:16]
  assign rvclkhdr_552_io_scan_mode = io_scan_mode; // @[el2_lib.scala 464:23]
  assign rvclkhdr_553_io_clk = clock; // @[el2_lib.scala 462:17]
  assign rvclkhdr_553_io_en = _T_6552 | _T_6557; // @[el2_lib.scala 463:16]
  assign rvclkhdr_553_io_scan_mode = io_scan_mode; // @[el2_lib.scala 464:23]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  leak_one_f_d1 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_0 = _RAND_1[21:0];
  _RAND_2 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_1 = _RAND_2[21:0];
  _RAND_3 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_2 = _RAND_3[21:0];
  _RAND_4 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_3 = _RAND_4[21:0];
  _RAND_5 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_4 = _RAND_5[21:0];
  _RAND_6 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_5 = _RAND_6[21:0];
  _RAND_7 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_6 = _RAND_7[21:0];
  _RAND_8 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_7 = _RAND_8[21:0];
  _RAND_9 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_8 = _RAND_9[21:0];
  _RAND_10 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_9 = _RAND_10[21:0];
  _RAND_11 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_10 = _RAND_11[21:0];
  _RAND_12 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_11 = _RAND_12[21:0];
  _RAND_13 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_12 = _RAND_13[21:0];
  _RAND_14 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_13 = _RAND_14[21:0];
  _RAND_15 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_14 = _RAND_15[21:0];
  _RAND_16 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_15 = _RAND_16[21:0];
  _RAND_17 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_16 = _RAND_17[21:0];
  _RAND_18 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_17 = _RAND_18[21:0];
  _RAND_19 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_18 = _RAND_19[21:0];
  _RAND_20 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_19 = _RAND_20[21:0];
  _RAND_21 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_20 = _RAND_21[21:0];
  _RAND_22 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_21 = _RAND_22[21:0];
  _RAND_23 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_22 = _RAND_23[21:0];
  _RAND_24 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_23 = _RAND_24[21:0];
  _RAND_25 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_24 = _RAND_25[21:0];
  _RAND_26 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_25 = _RAND_26[21:0];
  _RAND_27 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_26 = _RAND_27[21:0];
  _RAND_28 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_27 = _RAND_28[21:0];
  _RAND_29 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_28 = _RAND_29[21:0];
  _RAND_30 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_29 = _RAND_30[21:0];
  _RAND_31 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_30 = _RAND_31[21:0];
  _RAND_32 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_31 = _RAND_32[21:0];
  _RAND_33 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_32 = _RAND_33[21:0];
  _RAND_34 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_33 = _RAND_34[21:0];
  _RAND_35 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_34 = _RAND_35[21:0];
  _RAND_36 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_35 = _RAND_36[21:0];
  _RAND_37 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_36 = _RAND_37[21:0];
  _RAND_38 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_37 = _RAND_38[21:0];
  _RAND_39 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_38 = _RAND_39[21:0];
  _RAND_40 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_39 = _RAND_40[21:0];
  _RAND_41 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_40 = _RAND_41[21:0];
  _RAND_42 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_41 = _RAND_42[21:0];
  _RAND_43 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_42 = _RAND_43[21:0];
  _RAND_44 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_43 = _RAND_44[21:0];
  _RAND_45 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_44 = _RAND_45[21:0];
  _RAND_46 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_45 = _RAND_46[21:0];
  _RAND_47 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_46 = _RAND_47[21:0];
  _RAND_48 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_47 = _RAND_48[21:0];
  _RAND_49 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_48 = _RAND_49[21:0];
  _RAND_50 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_49 = _RAND_50[21:0];
  _RAND_51 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_50 = _RAND_51[21:0];
  _RAND_52 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_51 = _RAND_52[21:0];
  _RAND_53 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_52 = _RAND_53[21:0];
  _RAND_54 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_53 = _RAND_54[21:0];
  _RAND_55 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_54 = _RAND_55[21:0];
  _RAND_56 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_55 = _RAND_56[21:0];
  _RAND_57 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_56 = _RAND_57[21:0];
  _RAND_58 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_57 = _RAND_58[21:0];
  _RAND_59 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_58 = _RAND_59[21:0];
  _RAND_60 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_59 = _RAND_60[21:0];
  _RAND_61 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_60 = _RAND_61[21:0];
  _RAND_62 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_61 = _RAND_62[21:0];
  _RAND_63 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_62 = _RAND_63[21:0];
  _RAND_64 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_63 = _RAND_64[21:0];
  _RAND_65 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_64 = _RAND_65[21:0];
  _RAND_66 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_65 = _RAND_66[21:0];
  _RAND_67 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_66 = _RAND_67[21:0];
  _RAND_68 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_67 = _RAND_68[21:0];
  _RAND_69 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_68 = _RAND_69[21:0];
  _RAND_70 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_69 = _RAND_70[21:0];
  _RAND_71 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_70 = _RAND_71[21:0];
  _RAND_72 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_71 = _RAND_72[21:0];
  _RAND_73 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_72 = _RAND_73[21:0];
  _RAND_74 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_73 = _RAND_74[21:0];
  _RAND_75 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_74 = _RAND_75[21:0];
  _RAND_76 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_75 = _RAND_76[21:0];
  _RAND_77 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_76 = _RAND_77[21:0];
  _RAND_78 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_77 = _RAND_78[21:0];
  _RAND_79 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_78 = _RAND_79[21:0];
  _RAND_80 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_79 = _RAND_80[21:0];
  _RAND_81 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_80 = _RAND_81[21:0];
  _RAND_82 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_81 = _RAND_82[21:0];
  _RAND_83 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_82 = _RAND_83[21:0];
  _RAND_84 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_83 = _RAND_84[21:0];
  _RAND_85 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_84 = _RAND_85[21:0];
  _RAND_86 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_85 = _RAND_86[21:0];
  _RAND_87 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_86 = _RAND_87[21:0];
  _RAND_88 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_87 = _RAND_88[21:0];
  _RAND_89 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_88 = _RAND_89[21:0];
  _RAND_90 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_89 = _RAND_90[21:0];
  _RAND_91 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_90 = _RAND_91[21:0];
  _RAND_92 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_91 = _RAND_92[21:0];
  _RAND_93 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_92 = _RAND_93[21:0];
  _RAND_94 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_93 = _RAND_94[21:0];
  _RAND_95 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_94 = _RAND_95[21:0];
  _RAND_96 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_95 = _RAND_96[21:0];
  _RAND_97 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_96 = _RAND_97[21:0];
  _RAND_98 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_97 = _RAND_98[21:0];
  _RAND_99 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_98 = _RAND_99[21:0];
  _RAND_100 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_99 = _RAND_100[21:0];
  _RAND_101 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_100 = _RAND_101[21:0];
  _RAND_102 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_101 = _RAND_102[21:0];
  _RAND_103 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_102 = _RAND_103[21:0];
  _RAND_104 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_103 = _RAND_104[21:0];
  _RAND_105 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_104 = _RAND_105[21:0];
  _RAND_106 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_105 = _RAND_106[21:0];
  _RAND_107 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_106 = _RAND_107[21:0];
  _RAND_108 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_107 = _RAND_108[21:0];
  _RAND_109 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_108 = _RAND_109[21:0];
  _RAND_110 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_109 = _RAND_110[21:0];
  _RAND_111 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_110 = _RAND_111[21:0];
  _RAND_112 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_111 = _RAND_112[21:0];
  _RAND_113 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_112 = _RAND_113[21:0];
  _RAND_114 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_113 = _RAND_114[21:0];
  _RAND_115 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_114 = _RAND_115[21:0];
  _RAND_116 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_115 = _RAND_116[21:0];
  _RAND_117 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_116 = _RAND_117[21:0];
  _RAND_118 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_117 = _RAND_118[21:0];
  _RAND_119 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_118 = _RAND_119[21:0];
  _RAND_120 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_119 = _RAND_120[21:0];
  _RAND_121 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_120 = _RAND_121[21:0];
  _RAND_122 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_121 = _RAND_122[21:0];
  _RAND_123 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_122 = _RAND_123[21:0];
  _RAND_124 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_123 = _RAND_124[21:0];
  _RAND_125 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_124 = _RAND_125[21:0];
  _RAND_126 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_125 = _RAND_126[21:0];
  _RAND_127 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_126 = _RAND_127[21:0];
  _RAND_128 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_127 = _RAND_128[21:0];
  _RAND_129 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_128 = _RAND_129[21:0];
  _RAND_130 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_129 = _RAND_130[21:0];
  _RAND_131 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_130 = _RAND_131[21:0];
  _RAND_132 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_131 = _RAND_132[21:0];
  _RAND_133 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_132 = _RAND_133[21:0];
  _RAND_134 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_133 = _RAND_134[21:0];
  _RAND_135 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_134 = _RAND_135[21:0];
  _RAND_136 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_135 = _RAND_136[21:0];
  _RAND_137 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_136 = _RAND_137[21:0];
  _RAND_138 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_137 = _RAND_138[21:0];
  _RAND_139 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_138 = _RAND_139[21:0];
  _RAND_140 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_139 = _RAND_140[21:0];
  _RAND_141 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_140 = _RAND_141[21:0];
  _RAND_142 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_141 = _RAND_142[21:0];
  _RAND_143 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_142 = _RAND_143[21:0];
  _RAND_144 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_143 = _RAND_144[21:0];
  _RAND_145 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_144 = _RAND_145[21:0];
  _RAND_146 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_145 = _RAND_146[21:0];
  _RAND_147 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_146 = _RAND_147[21:0];
  _RAND_148 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_147 = _RAND_148[21:0];
  _RAND_149 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_148 = _RAND_149[21:0];
  _RAND_150 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_149 = _RAND_150[21:0];
  _RAND_151 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_150 = _RAND_151[21:0];
  _RAND_152 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_151 = _RAND_152[21:0];
  _RAND_153 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_152 = _RAND_153[21:0];
  _RAND_154 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_153 = _RAND_154[21:0];
  _RAND_155 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_154 = _RAND_155[21:0];
  _RAND_156 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_155 = _RAND_156[21:0];
  _RAND_157 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_156 = _RAND_157[21:0];
  _RAND_158 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_157 = _RAND_158[21:0];
  _RAND_159 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_158 = _RAND_159[21:0];
  _RAND_160 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_159 = _RAND_160[21:0];
  _RAND_161 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_160 = _RAND_161[21:0];
  _RAND_162 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_161 = _RAND_162[21:0];
  _RAND_163 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_162 = _RAND_163[21:0];
  _RAND_164 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_163 = _RAND_164[21:0];
  _RAND_165 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_164 = _RAND_165[21:0];
  _RAND_166 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_165 = _RAND_166[21:0];
  _RAND_167 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_166 = _RAND_167[21:0];
  _RAND_168 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_167 = _RAND_168[21:0];
  _RAND_169 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_168 = _RAND_169[21:0];
  _RAND_170 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_169 = _RAND_170[21:0];
  _RAND_171 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_170 = _RAND_171[21:0];
  _RAND_172 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_171 = _RAND_172[21:0];
  _RAND_173 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_172 = _RAND_173[21:0];
  _RAND_174 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_173 = _RAND_174[21:0];
  _RAND_175 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_174 = _RAND_175[21:0];
  _RAND_176 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_175 = _RAND_176[21:0];
  _RAND_177 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_176 = _RAND_177[21:0];
  _RAND_178 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_177 = _RAND_178[21:0];
  _RAND_179 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_178 = _RAND_179[21:0];
  _RAND_180 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_179 = _RAND_180[21:0];
  _RAND_181 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_180 = _RAND_181[21:0];
  _RAND_182 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_181 = _RAND_182[21:0];
  _RAND_183 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_182 = _RAND_183[21:0];
  _RAND_184 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_183 = _RAND_184[21:0];
  _RAND_185 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_184 = _RAND_185[21:0];
  _RAND_186 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_185 = _RAND_186[21:0];
  _RAND_187 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_186 = _RAND_187[21:0];
  _RAND_188 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_187 = _RAND_188[21:0];
  _RAND_189 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_188 = _RAND_189[21:0];
  _RAND_190 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_189 = _RAND_190[21:0];
  _RAND_191 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_190 = _RAND_191[21:0];
  _RAND_192 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_191 = _RAND_192[21:0];
  _RAND_193 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_192 = _RAND_193[21:0];
  _RAND_194 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_193 = _RAND_194[21:0];
  _RAND_195 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_194 = _RAND_195[21:0];
  _RAND_196 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_195 = _RAND_196[21:0];
  _RAND_197 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_196 = _RAND_197[21:0];
  _RAND_198 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_197 = _RAND_198[21:0];
  _RAND_199 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_198 = _RAND_199[21:0];
  _RAND_200 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_199 = _RAND_200[21:0];
  _RAND_201 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_200 = _RAND_201[21:0];
  _RAND_202 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_201 = _RAND_202[21:0];
  _RAND_203 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_202 = _RAND_203[21:0];
  _RAND_204 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_203 = _RAND_204[21:0];
  _RAND_205 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_204 = _RAND_205[21:0];
  _RAND_206 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_205 = _RAND_206[21:0];
  _RAND_207 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_206 = _RAND_207[21:0];
  _RAND_208 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_207 = _RAND_208[21:0];
  _RAND_209 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_208 = _RAND_209[21:0];
  _RAND_210 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_209 = _RAND_210[21:0];
  _RAND_211 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_210 = _RAND_211[21:0];
  _RAND_212 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_211 = _RAND_212[21:0];
  _RAND_213 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_212 = _RAND_213[21:0];
  _RAND_214 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_213 = _RAND_214[21:0];
  _RAND_215 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_214 = _RAND_215[21:0];
  _RAND_216 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_215 = _RAND_216[21:0];
  _RAND_217 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_216 = _RAND_217[21:0];
  _RAND_218 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_217 = _RAND_218[21:0];
  _RAND_219 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_218 = _RAND_219[21:0];
  _RAND_220 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_219 = _RAND_220[21:0];
  _RAND_221 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_220 = _RAND_221[21:0];
  _RAND_222 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_221 = _RAND_222[21:0];
  _RAND_223 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_222 = _RAND_223[21:0];
  _RAND_224 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_223 = _RAND_224[21:0];
  _RAND_225 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_224 = _RAND_225[21:0];
  _RAND_226 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_225 = _RAND_226[21:0];
  _RAND_227 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_226 = _RAND_227[21:0];
  _RAND_228 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_227 = _RAND_228[21:0];
  _RAND_229 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_228 = _RAND_229[21:0];
  _RAND_230 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_229 = _RAND_230[21:0];
  _RAND_231 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_230 = _RAND_231[21:0];
  _RAND_232 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_231 = _RAND_232[21:0];
  _RAND_233 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_232 = _RAND_233[21:0];
  _RAND_234 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_233 = _RAND_234[21:0];
  _RAND_235 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_234 = _RAND_235[21:0];
  _RAND_236 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_235 = _RAND_236[21:0];
  _RAND_237 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_236 = _RAND_237[21:0];
  _RAND_238 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_237 = _RAND_238[21:0];
  _RAND_239 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_238 = _RAND_239[21:0];
  _RAND_240 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_239 = _RAND_240[21:0];
  _RAND_241 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_240 = _RAND_241[21:0];
  _RAND_242 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_241 = _RAND_242[21:0];
  _RAND_243 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_242 = _RAND_243[21:0];
  _RAND_244 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_243 = _RAND_244[21:0];
  _RAND_245 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_244 = _RAND_245[21:0];
  _RAND_246 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_245 = _RAND_246[21:0];
  _RAND_247 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_246 = _RAND_247[21:0];
  _RAND_248 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_247 = _RAND_248[21:0];
  _RAND_249 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_248 = _RAND_249[21:0];
  _RAND_250 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_249 = _RAND_250[21:0];
  _RAND_251 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_250 = _RAND_251[21:0];
  _RAND_252 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_251 = _RAND_252[21:0];
  _RAND_253 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_252 = _RAND_253[21:0];
  _RAND_254 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_253 = _RAND_254[21:0];
  _RAND_255 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_254 = _RAND_255[21:0];
  _RAND_256 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_255 = _RAND_256[21:0];
  _RAND_257 = {1{`RANDOM}};
  dec_tlu_way_wb_f = _RAND_257[0:0];
  _RAND_258 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_0 = _RAND_258[21:0];
  _RAND_259 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_1 = _RAND_259[21:0];
  _RAND_260 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_2 = _RAND_260[21:0];
  _RAND_261 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_3 = _RAND_261[21:0];
  _RAND_262 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_4 = _RAND_262[21:0];
  _RAND_263 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_5 = _RAND_263[21:0];
  _RAND_264 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_6 = _RAND_264[21:0];
  _RAND_265 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_7 = _RAND_265[21:0];
  _RAND_266 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_8 = _RAND_266[21:0];
  _RAND_267 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_9 = _RAND_267[21:0];
  _RAND_268 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_10 = _RAND_268[21:0];
  _RAND_269 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_11 = _RAND_269[21:0];
  _RAND_270 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_12 = _RAND_270[21:0];
  _RAND_271 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_13 = _RAND_271[21:0];
  _RAND_272 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_14 = _RAND_272[21:0];
  _RAND_273 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_15 = _RAND_273[21:0];
  _RAND_274 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_16 = _RAND_274[21:0];
  _RAND_275 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_17 = _RAND_275[21:0];
  _RAND_276 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_18 = _RAND_276[21:0];
  _RAND_277 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_19 = _RAND_277[21:0];
  _RAND_278 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_20 = _RAND_278[21:0];
  _RAND_279 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_21 = _RAND_279[21:0];
  _RAND_280 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_22 = _RAND_280[21:0];
  _RAND_281 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_23 = _RAND_281[21:0];
  _RAND_282 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_24 = _RAND_282[21:0];
  _RAND_283 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_25 = _RAND_283[21:0];
  _RAND_284 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_26 = _RAND_284[21:0];
  _RAND_285 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_27 = _RAND_285[21:0];
  _RAND_286 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_28 = _RAND_286[21:0];
  _RAND_287 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_29 = _RAND_287[21:0];
  _RAND_288 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_30 = _RAND_288[21:0];
  _RAND_289 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_31 = _RAND_289[21:0];
  _RAND_290 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_32 = _RAND_290[21:0];
  _RAND_291 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_33 = _RAND_291[21:0];
  _RAND_292 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_34 = _RAND_292[21:0];
  _RAND_293 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_35 = _RAND_293[21:0];
  _RAND_294 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_36 = _RAND_294[21:0];
  _RAND_295 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_37 = _RAND_295[21:0];
  _RAND_296 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_38 = _RAND_296[21:0];
  _RAND_297 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_39 = _RAND_297[21:0];
  _RAND_298 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_40 = _RAND_298[21:0];
  _RAND_299 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_41 = _RAND_299[21:0];
  _RAND_300 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_42 = _RAND_300[21:0];
  _RAND_301 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_43 = _RAND_301[21:0];
  _RAND_302 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_44 = _RAND_302[21:0];
  _RAND_303 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_45 = _RAND_303[21:0];
  _RAND_304 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_46 = _RAND_304[21:0];
  _RAND_305 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_47 = _RAND_305[21:0];
  _RAND_306 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_48 = _RAND_306[21:0];
  _RAND_307 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_49 = _RAND_307[21:0];
  _RAND_308 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_50 = _RAND_308[21:0];
  _RAND_309 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_51 = _RAND_309[21:0];
  _RAND_310 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_52 = _RAND_310[21:0];
  _RAND_311 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_53 = _RAND_311[21:0];
  _RAND_312 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_54 = _RAND_312[21:0];
  _RAND_313 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_55 = _RAND_313[21:0];
  _RAND_314 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_56 = _RAND_314[21:0];
  _RAND_315 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_57 = _RAND_315[21:0];
  _RAND_316 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_58 = _RAND_316[21:0];
  _RAND_317 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_59 = _RAND_317[21:0];
  _RAND_318 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_60 = _RAND_318[21:0];
  _RAND_319 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_61 = _RAND_319[21:0];
  _RAND_320 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_62 = _RAND_320[21:0];
  _RAND_321 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_63 = _RAND_321[21:0];
  _RAND_322 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_64 = _RAND_322[21:0];
  _RAND_323 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_65 = _RAND_323[21:0];
  _RAND_324 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_66 = _RAND_324[21:0];
  _RAND_325 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_67 = _RAND_325[21:0];
  _RAND_326 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_68 = _RAND_326[21:0];
  _RAND_327 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_69 = _RAND_327[21:0];
  _RAND_328 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_70 = _RAND_328[21:0];
  _RAND_329 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_71 = _RAND_329[21:0];
  _RAND_330 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_72 = _RAND_330[21:0];
  _RAND_331 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_73 = _RAND_331[21:0];
  _RAND_332 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_74 = _RAND_332[21:0];
  _RAND_333 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_75 = _RAND_333[21:0];
  _RAND_334 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_76 = _RAND_334[21:0];
  _RAND_335 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_77 = _RAND_335[21:0];
  _RAND_336 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_78 = _RAND_336[21:0];
  _RAND_337 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_79 = _RAND_337[21:0];
  _RAND_338 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_80 = _RAND_338[21:0];
  _RAND_339 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_81 = _RAND_339[21:0];
  _RAND_340 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_82 = _RAND_340[21:0];
  _RAND_341 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_83 = _RAND_341[21:0];
  _RAND_342 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_84 = _RAND_342[21:0];
  _RAND_343 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_85 = _RAND_343[21:0];
  _RAND_344 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_86 = _RAND_344[21:0];
  _RAND_345 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_87 = _RAND_345[21:0];
  _RAND_346 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_88 = _RAND_346[21:0];
  _RAND_347 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_89 = _RAND_347[21:0];
  _RAND_348 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_90 = _RAND_348[21:0];
  _RAND_349 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_91 = _RAND_349[21:0];
  _RAND_350 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_92 = _RAND_350[21:0];
  _RAND_351 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_93 = _RAND_351[21:0];
  _RAND_352 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_94 = _RAND_352[21:0];
  _RAND_353 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_95 = _RAND_353[21:0];
  _RAND_354 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_96 = _RAND_354[21:0];
  _RAND_355 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_97 = _RAND_355[21:0];
  _RAND_356 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_98 = _RAND_356[21:0];
  _RAND_357 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_99 = _RAND_357[21:0];
  _RAND_358 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_100 = _RAND_358[21:0];
  _RAND_359 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_101 = _RAND_359[21:0];
  _RAND_360 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_102 = _RAND_360[21:0];
  _RAND_361 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_103 = _RAND_361[21:0];
  _RAND_362 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_104 = _RAND_362[21:0];
  _RAND_363 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_105 = _RAND_363[21:0];
  _RAND_364 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_106 = _RAND_364[21:0];
  _RAND_365 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_107 = _RAND_365[21:0];
  _RAND_366 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_108 = _RAND_366[21:0];
  _RAND_367 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_109 = _RAND_367[21:0];
  _RAND_368 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_110 = _RAND_368[21:0];
  _RAND_369 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_111 = _RAND_369[21:0];
  _RAND_370 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_112 = _RAND_370[21:0];
  _RAND_371 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_113 = _RAND_371[21:0];
  _RAND_372 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_114 = _RAND_372[21:0];
  _RAND_373 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_115 = _RAND_373[21:0];
  _RAND_374 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_116 = _RAND_374[21:0];
  _RAND_375 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_117 = _RAND_375[21:0];
  _RAND_376 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_118 = _RAND_376[21:0];
  _RAND_377 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_119 = _RAND_377[21:0];
  _RAND_378 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_120 = _RAND_378[21:0];
  _RAND_379 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_121 = _RAND_379[21:0];
  _RAND_380 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_122 = _RAND_380[21:0];
  _RAND_381 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_123 = _RAND_381[21:0];
  _RAND_382 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_124 = _RAND_382[21:0];
  _RAND_383 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_125 = _RAND_383[21:0];
  _RAND_384 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_126 = _RAND_384[21:0];
  _RAND_385 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_127 = _RAND_385[21:0];
  _RAND_386 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_128 = _RAND_386[21:0];
  _RAND_387 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_129 = _RAND_387[21:0];
  _RAND_388 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_130 = _RAND_388[21:0];
  _RAND_389 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_131 = _RAND_389[21:0];
  _RAND_390 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_132 = _RAND_390[21:0];
  _RAND_391 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_133 = _RAND_391[21:0];
  _RAND_392 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_134 = _RAND_392[21:0];
  _RAND_393 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_135 = _RAND_393[21:0];
  _RAND_394 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_136 = _RAND_394[21:0];
  _RAND_395 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_137 = _RAND_395[21:0];
  _RAND_396 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_138 = _RAND_396[21:0];
  _RAND_397 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_139 = _RAND_397[21:0];
  _RAND_398 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_140 = _RAND_398[21:0];
  _RAND_399 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_141 = _RAND_399[21:0];
  _RAND_400 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_142 = _RAND_400[21:0];
  _RAND_401 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_143 = _RAND_401[21:0];
  _RAND_402 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_144 = _RAND_402[21:0];
  _RAND_403 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_145 = _RAND_403[21:0];
  _RAND_404 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_146 = _RAND_404[21:0];
  _RAND_405 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_147 = _RAND_405[21:0];
  _RAND_406 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_148 = _RAND_406[21:0];
  _RAND_407 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_149 = _RAND_407[21:0];
  _RAND_408 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_150 = _RAND_408[21:0];
  _RAND_409 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_151 = _RAND_409[21:0];
  _RAND_410 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_152 = _RAND_410[21:0];
  _RAND_411 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_153 = _RAND_411[21:0];
  _RAND_412 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_154 = _RAND_412[21:0];
  _RAND_413 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_155 = _RAND_413[21:0];
  _RAND_414 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_156 = _RAND_414[21:0];
  _RAND_415 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_157 = _RAND_415[21:0];
  _RAND_416 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_158 = _RAND_416[21:0];
  _RAND_417 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_159 = _RAND_417[21:0];
  _RAND_418 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_160 = _RAND_418[21:0];
  _RAND_419 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_161 = _RAND_419[21:0];
  _RAND_420 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_162 = _RAND_420[21:0];
  _RAND_421 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_163 = _RAND_421[21:0];
  _RAND_422 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_164 = _RAND_422[21:0];
  _RAND_423 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_165 = _RAND_423[21:0];
  _RAND_424 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_166 = _RAND_424[21:0];
  _RAND_425 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_167 = _RAND_425[21:0];
  _RAND_426 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_168 = _RAND_426[21:0];
  _RAND_427 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_169 = _RAND_427[21:0];
  _RAND_428 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_170 = _RAND_428[21:0];
  _RAND_429 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_171 = _RAND_429[21:0];
  _RAND_430 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_172 = _RAND_430[21:0];
  _RAND_431 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_173 = _RAND_431[21:0];
  _RAND_432 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_174 = _RAND_432[21:0];
  _RAND_433 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_175 = _RAND_433[21:0];
  _RAND_434 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_176 = _RAND_434[21:0];
  _RAND_435 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_177 = _RAND_435[21:0];
  _RAND_436 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_178 = _RAND_436[21:0];
  _RAND_437 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_179 = _RAND_437[21:0];
  _RAND_438 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_180 = _RAND_438[21:0];
  _RAND_439 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_181 = _RAND_439[21:0];
  _RAND_440 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_182 = _RAND_440[21:0];
  _RAND_441 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_183 = _RAND_441[21:0];
  _RAND_442 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_184 = _RAND_442[21:0];
  _RAND_443 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_185 = _RAND_443[21:0];
  _RAND_444 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_186 = _RAND_444[21:0];
  _RAND_445 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_187 = _RAND_445[21:0];
  _RAND_446 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_188 = _RAND_446[21:0];
  _RAND_447 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_189 = _RAND_447[21:0];
  _RAND_448 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_190 = _RAND_448[21:0];
  _RAND_449 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_191 = _RAND_449[21:0];
  _RAND_450 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_192 = _RAND_450[21:0];
  _RAND_451 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_193 = _RAND_451[21:0];
  _RAND_452 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_194 = _RAND_452[21:0];
  _RAND_453 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_195 = _RAND_453[21:0];
  _RAND_454 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_196 = _RAND_454[21:0];
  _RAND_455 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_197 = _RAND_455[21:0];
  _RAND_456 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_198 = _RAND_456[21:0];
  _RAND_457 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_199 = _RAND_457[21:0];
  _RAND_458 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_200 = _RAND_458[21:0];
  _RAND_459 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_201 = _RAND_459[21:0];
  _RAND_460 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_202 = _RAND_460[21:0];
  _RAND_461 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_203 = _RAND_461[21:0];
  _RAND_462 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_204 = _RAND_462[21:0];
  _RAND_463 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_205 = _RAND_463[21:0];
  _RAND_464 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_206 = _RAND_464[21:0];
  _RAND_465 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_207 = _RAND_465[21:0];
  _RAND_466 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_208 = _RAND_466[21:0];
  _RAND_467 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_209 = _RAND_467[21:0];
  _RAND_468 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_210 = _RAND_468[21:0];
  _RAND_469 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_211 = _RAND_469[21:0];
  _RAND_470 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_212 = _RAND_470[21:0];
  _RAND_471 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_213 = _RAND_471[21:0];
  _RAND_472 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_214 = _RAND_472[21:0];
  _RAND_473 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_215 = _RAND_473[21:0];
  _RAND_474 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_216 = _RAND_474[21:0];
  _RAND_475 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_217 = _RAND_475[21:0];
  _RAND_476 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_218 = _RAND_476[21:0];
  _RAND_477 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_219 = _RAND_477[21:0];
  _RAND_478 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_220 = _RAND_478[21:0];
  _RAND_479 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_221 = _RAND_479[21:0];
  _RAND_480 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_222 = _RAND_480[21:0];
  _RAND_481 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_223 = _RAND_481[21:0];
  _RAND_482 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_224 = _RAND_482[21:0];
  _RAND_483 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_225 = _RAND_483[21:0];
  _RAND_484 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_226 = _RAND_484[21:0];
  _RAND_485 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_227 = _RAND_485[21:0];
  _RAND_486 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_228 = _RAND_486[21:0];
  _RAND_487 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_229 = _RAND_487[21:0];
  _RAND_488 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_230 = _RAND_488[21:0];
  _RAND_489 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_231 = _RAND_489[21:0];
  _RAND_490 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_232 = _RAND_490[21:0];
  _RAND_491 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_233 = _RAND_491[21:0];
  _RAND_492 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_234 = _RAND_492[21:0];
  _RAND_493 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_235 = _RAND_493[21:0];
  _RAND_494 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_236 = _RAND_494[21:0];
  _RAND_495 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_237 = _RAND_495[21:0];
  _RAND_496 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_238 = _RAND_496[21:0];
  _RAND_497 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_239 = _RAND_497[21:0];
  _RAND_498 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_240 = _RAND_498[21:0];
  _RAND_499 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_241 = _RAND_499[21:0];
  _RAND_500 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_242 = _RAND_500[21:0];
  _RAND_501 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_243 = _RAND_501[21:0];
  _RAND_502 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_244 = _RAND_502[21:0];
  _RAND_503 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_245 = _RAND_503[21:0];
  _RAND_504 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_246 = _RAND_504[21:0];
  _RAND_505 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_247 = _RAND_505[21:0];
  _RAND_506 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_248 = _RAND_506[21:0];
  _RAND_507 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_249 = _RAND_507[21:0];
  _RAND_508 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_250 = _RAND_508[21:0];
  _RAND_509 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_251 = _RAND_509[21:0];
  _RAND_510 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_252 = _RAND_510[21:0];
  _RAND_511 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_253 = _RAND_511[21:0];
  _RAND_512 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_254 = _RAND_512[21:0];
  _RAND_513 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_255 = _RAND_513[21:0];
  _RAND_514 = {1{`RANDOM}};
  fghr = _RAND_514[7:0];
  _RAND_515 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_0 = _RAND_515[1:0];
  _RAND_516 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_1 = _RAND_516[1:0];
  _RAND_517 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_2 = _RAND_517[1:0];
  _RAND_518 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_3 = _RAND_518[1:0];
  _RAND_519 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_4 = _RAND_519[1:0];
  _RAND_520 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_5 = _RAND_520[1:0];
  _RAND_521 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_6 = _RAND_521[1:0];
  _RAND_522 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_7 = _RAND_522[1:0];
  _RAND_523 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_8 = _RAND_523[1:0];
  _RAND_524 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_9 = _RAND_524[1:0];
  _RAND_525 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_10 = _RAND_525[1:0];
  _RAND_526 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_11 = _RAND_526[1:0];
  _RAND_527 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_12 = _RAND_527[1:0];
  _RAND_528 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_13 = _RAND_528[1:0];
  _RAND_529 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_14 = _RAND_529[1:0];
  _RAND_530 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_15 = _RAND_530[1:0];
  _RAND_531 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_16 = _RAND_531[1:0];
  _RAND_532 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_17 = _RAND_532[1:0];
  _RAND_533 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_18 = _RAND_533[1:0];
  _RAND_534 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_19 = _RAND_534[1:0];
  _RAND_535 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_20 = _RAND_535[1:0];
  _RAND_536 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_21 = _RAND_536[1:0];
  _RAND_537 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_22 = _RAND_537[1:0];
  _RAND_538 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_23 = _RAND_538[1:0];
  _RAND_539 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_24 = _RAND_539[1:0];
  _RAND_540 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_25 = _RAND_540[1:0];
  _RAND_541 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_26 = _RAND_541[1:0];
  _RAND_542 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_27 = _RAND_542[1:0];
  _RAND_543 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_28 = _RAND_543[1:0];
  _RAND_544 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_29 = _RAND_544[1:0];
  _RAND_545 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_30 = _RAND_545[1:0];
  _RAND_546 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_31 = _RAND_546[1:0];
  _RAND_547 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_32 = _RAND_547[1:0];
  _RAND_548 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_33 = _RAND_548[1:0];
  _RAND_549 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_34 = _RAND_549[1:0];
  _RAND_550 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_35 = _RAND_550[1:0];
  _RAND_551 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_36 = _RAND_551[1:0];
  _RAND_552 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_37 = _RAND_552[1:0];
  _RAND_553 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_38 = _RAND_553[1:0];
  _RAND_554 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_39 = _RAND_554[1:0];
  _RAND_555 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_40 = _RAND_555[1:0];
  _RAND_556 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_41 = _RAND_556[1:0];
  _RAND_557 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_42 = _RAND_557[1:0];
  _RAND_558 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_43 = _RAND_558[1:0];
  _RAND_559 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_44 = _RAND_559[1:0];
  _RAND_560 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_45 = _RAND_560[1:0];
  _RAND_561 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_46 = _RAND_561[1:0];
  _RAND_562 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_47 = _RAND_562[1:0];
  _RAND_563 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_48 = _RAND_563[1:0];
  _RAND_564 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_49 = _RAND_564[1:0];
  _RAND_565 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_50 = _RAND_565[1:0];
  _RAND_566 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_51 = _RAND_566[1:0];
  _RAND_567 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_52 = _RAND_567[1:0];
  _RAND_568 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_53 = _RAND_568[1:0];
  _RAND_569 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_54 = _RAND_569[1:0];
  _RAND_570 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_55 = _RAND_570[1:0];
  _RAND_571 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_56 = _RAND_571[1:0];
  _RAND_572 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_57 = _RAND_572[1:0];
  _RAND_573 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_58 = _RAND_573[1:0];
  _RAND_574 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_59 = _RAND_574[1:0];
  _RAND_575 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_60 = _RAND_575[1:0];
  _RAND_576 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_61 = _RAND_576[1:0];
  _RAND_577 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_62 = _RAND_577[1:0];
  _RAND_578 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_63 = _RAND_578[1:0];
  _RAND_579 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_64 = _RAND_579[1:0];
  _RAND_580 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_65 = _RAND_580[1:0];
  _RAND_581 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_66 = _RAND_581[1:0];
  _RAND_582 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_67 = _RAND_582[1:0];
  _RAND_583 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_68 = _RAND_583[1:0];
  _RAND_584 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_69 = _RAND_584[1:0];
  _RAND_585 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_70 = _RAND_585[1:0];
  _RAND_586 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_71 = _RAND_586[1:0];
  _RAND_587 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_72 = _RAND_587[1:0];
  _RAND_588 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_73 = _RAND_588[1:0];
  _RAND_589 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_74 = _RAND_589[1:0];
  _RAND_590 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_75 = _RAND_590[1:0];
  _RAND_591 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_76 = _RAND_591[1:0];
  _RAND_592 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_77 = _RAND_592[1:0];
  _RAND_593 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_78 = _RAND_593[1:0];
  _RAND_594 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_79 = _RAND_594[1:0];
  _RAND_595 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_80 = _RAND_595[1:0];
  _RAND_596 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_81 = _RAND_596[1:0];
  _RAND_597 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_82 = _RAND_597[1:0];
  _RAND_598 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_83 = _RAND_598[1:0];
  _RAND_599 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_84 = _RAND_599[1:0];
  _RAND_600 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_85 = _RAND_600[1:0];
  _RAND_601 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_86 = _RAND_601[1:0];
  _RAND_602 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_87 = _RAND_602[1:0];
  _RAND_603 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_88 = _RAND_603[1:0];
  _RAND_604 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_89 = _RAND_604[1:0];
  _RAND_605 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_90 = _RAND_605[1:0];
  _RAND_606 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_91 = _RAND_606[1:0];
  _RAND_607 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_92 = _RAND_607[1:0];
  _RAND_608 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_93 = _RAND_608[1:0];
  _RAND_609 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_94 = _RAND_609[1:0];
  _RAND_610 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_95 = _RAND_610[1:0];
  _RAND_611 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_96 = _RAND_611[1:0];
  _RAND_612 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_97 = _RAND_612[1:0];
  _RAND_613 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_98 = _RAND_613[1:0];
  _RAND_614 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_99 = _RAND_614[1:0];
  _RAND_615 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_100 = _RAND_615[1:0];
  _RAND_616 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_101 = _RAND_616[1:0];
  _RAND_617 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_102 = _RAND_617[1:0];
  _RAND_618 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_103 = _RAND_618[1:0];
  _RAND_619 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_104 = _RAND_619[1:0];
  _RAND_620 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_105 = _RAND_620[1:0];
  _RAND_621 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_106 = _RAND_621[1:0];
  _RAND_622 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_107 = _RAND_622[1:0];
  _RAND_623 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_108 = _RAND_623[1:0];
  _RAND_624 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_109 = _RAND_624[1:0];
  _RAND_625 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_110 = _RAND_625[1:0];
  _RAND_626 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_111 = _RAND_626[1:0];
  _RAND_627 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_112 = _RAND_627[1:0];
  _RAND_628 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_113 = _RAND_628[1:0];
  _RAND_629 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_114 = _RAND_629[1:0];
  _RAND_630 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_115 = _RAND_630[1:0];
  _RAND_631 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_116 = _RAND_631[1:0];
  _RAND_632 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_117 = _RAND_632[1:0];
  _RAND_633 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_118 = _RAND_633[1:0];
  _RAND_634 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_119 = _RAND_634[1:0];
  _RAND_635 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_120 = _RAND_635[1:0];
  _RAND_636 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_121 = _RAND_636[1:0];
  _RAND_637 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_122 = _RAND_637[1:0];
  _RAND_638 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_123 = _RAND_638[1:0];
  _RAND_639 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_124 = _RAND_639[1:0];
  _RAND_640 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_125 = _RAND_640[1:0];
  _RAND_641 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_126 = _RAND_641[1:0];
  _RAND_642 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_127 = _RAND_642[1:0];
  _RAND_643 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_128 = _RAND_643[1:0];
  _RAND_644 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_129 = _RAND_644[1:0];
  _RAND_645 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_130 = _RAND_645[1:0];
  _RAND_646 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_131 = _RAND_646[1:0];
  _RAND_647 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_132 = _RAND_647[1:0];
  _RAND_648 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_133 = _RAND_648[1:0];
  _RAND_649 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_134 = _RAND_649[1:0];
  _RAND_650 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_135 = _RAND_650[1:0];
  _RAND_651 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_136 = _RAND_651[1:0];
  _RAND_652 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_137 = _RAND_652[1:0];
  _RAND_653 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_138 = _RAND_653[1:0];
  _RAND_654 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_139 = _RAND_654[1:0];
  _RAND_655 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_140 = _RAND_655[1:0];
  _RAND_656 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_141 = _RAND_656[1:0];
  _RAND_657 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_142 = _RAND_657[1:0];
  _RAND_658 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_143 = _RAND_658[1:0];
  _RAND_659 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_144 = _RAND_659[1:0];
  _RAND_660 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_145 = _RAND_660[1:0];
  _RAND_661 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_146 = _RAND_661[1:0];
  _RAND_662 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_147 = _RAND_662[1:0];
  _RAND_663 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_148 = _RAND_663[1:0];
  _RAND_664 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_149 = _RAND_664[1:0];
  _RAND_665 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_150 = _RAND_665[1:0];
  _RAND_666 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_151 = _RAND_666[1:0];
  _RAND_667 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_152 = _RAND_667[1:0];
  _RAND_668 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_153 = _RAND_668[1:0];
  _RAND_669 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_154 = _RAND_669[1:0];
  _RAND_670 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_155 = _RAND_670[1:0];
  _RAND_671 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_156 = _RAND_671[1:0];
  _RAND_672 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_157 = _RAND_672[1:0];
  _RAND_673 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_158 = _RAND_673[1:0];
  _RAND_674 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_159 = _RAND_674[1:0];
  _RAND_675 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_160 = _RAND_675[1:0];
  _RAND_676 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_161 = _RAND_676[1:0];
  _RAND_677 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_162 = _RAND_677[1:0];
  _RAND_678 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_163 = _RAND_678[1:0];
  _RAND_679 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_164 = _RAND_679[1:0];
  _RAND_680 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_165 = _RAND_680[1:0];
  _RAND_681 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_166 = _RAND_681[1:0];
  _RAND_682 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_167 = _RAND_682[1:0];
  _RAND_683 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_168 = _RAND_683[1:0];
  _RAND_684 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_169 = _RAND_684[1:0];
  _RAND_685 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_170 = _RAND_685[1:0];
  _RAND_686 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_171 = _RAND_686[1:0];
  _RAND_687 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_172 = _RAND_687[1:0];
  _RAND_688 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_173 = _RAND_688[1:0];
  _RAND_689 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_174 = _RAND_689[1:0];
  _RAND_690 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_175 = _RAND_690[1:0];
  _RAND_691 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_176 = _RAND_691[1:0];
  _RAND_692 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_177 = _RAND_692[1:0];
  _RAND_693 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_178 = _RAND_693[1:0];
  _RAND_694 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_179 = _RAND_694[1:0];
  _RAND_695 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_180 = _RAND_695[1:0];
  _RAND_696 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_181 = _RAND_696[1:0];
  _RAND_697 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_182 = _RAND_697[1:0];
  _RAND_698 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_183 = _RAND_698[1:0];
  _RAND_699 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_184 = _RAND_699[1:0];
  _RAND_700 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_185 = _RAND_700[1:0];
  _RAND_701 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_186 = _RAND_701[1:0];
  _RAND_702 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_187 = _RAND_702[1:0];
  _RAND_703 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_188 = _RAND_703[1:0];
  _RAND_704 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_189 = _RAND_704[1:0];
  _RAND_705 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_190 = _RAND_705[1:0];
  _RAND_706 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_191 = _RAND_706[1:0];
  _RAND_707 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_192 = _RAND_707[1:0];
  _RAND_708 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_193 = _RAND_708[1:0];
  _RAND_709 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_194 = _RAND_709[1:0];
  _RAND_710 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_195 = _RAND_710[1:0];
  _RAND_711 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_196 = _RAND_711[1:0];
  _RAND_712 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_197 = _RAND_712[1:0];
  _RAND_713 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_198 = _RAND_713[1:0];
  _RAND_714 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_199 = _RAND_714[1:0];
  _RAND_715 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_200 = _RAND_715[1:0];
  _RAND_716 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_201 = _RAND_716[1:0];
  _RAND_717 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_202 = _RAND_717[1:0];
  _RAND_718 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_203 = _RAND_718[1:0];
  _RAND_719 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_204 = _RAND_719[1:0];
  _RAND_720 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_205 = _RAND_720[1:0];
  _RAND_721 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_206 = _RAND_721[1:0];
  _RAND_722 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_207 = _RAND_722[1:0];
  _RAND_723 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_208 = _RAND_723[1:0];
  _RAND_724 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_209 = _RAND_724[1:0];
  _RAND_725 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_210 = _RAND_725[1:0];
  _RAND_726 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_211 = _RAND_726[1:0];
  _RAND_727 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_212 = _RAND_727[1:0];
  _RAND_728 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_213 = _RAND_728[1:0];
  _RAND_729 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_214 = _RAND_729[1:0];
  _RAND_730 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_215 = _RAND_730[1:0];
  _RAND_731 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_216 = _RAND_731[1:0];
  _RAND_732 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_217 = _RAND_732[1:0];
  _RAND_733 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_218 = _RAND_733[1:0];
  _RAND_734 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_219 = _RAND_734[1:0];
  _RAND_735 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_220 = _RAND_735[1:0];
  _RAND_736 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_221 = _RAND_736[1:0];
  _RAND_737 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_222 = _RAND_737[1:0];
  _RAND_738 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_223 = _RAND_738[1:0];
  _RAND_739 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_224 = _RAND_739[1:0];
  _RAND_740 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_225 = _RAND_740[1:0];
  _RAND_741 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_226 = _RAND_741[1:0];
  _RAND_742 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_227 = _RAND_742[1:0];
  _RAND_743 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_228 = _RAND_743[1:0];
  _RAND_744 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_229 = _RAND_744[1:0];
  _RAND_745 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_230 = _RAND_745[1:0];
  _RAND_746 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_231 = _RAND_746[1:0];
  _RAND_747 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_232 = _RAND_747[1:0];
  _RAND_748 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_233 = _RAND_748[1:0];
  _RAND_749 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_234 = _RAND_749[1:0];
  _RAND_750 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_235 = _RAND_750[1:0];
  _RAND_751 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_236 = _RAND_751[1:0];
  _RAND_752 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_237 = _RAND_752[1:0];
  _RAND_753 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_238 = _RAND_753[1:0];
  _RAND_754 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_239 = _RAND_754[1:0];
  _RAND_755 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_240 = _RAND_755[1:0];
  _RAND_756 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_241 = _RAND_756[1:0];
  _RAND_757 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_242 = _RAND_757[1:0];
  _RAND_758 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_243 = _RAND_758[1:0];
  _RAND_759 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_244 = _RAND_759[1:0];
  _RAND_760 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_245 = _RAND_760[1:0];
  _RAND_761 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_246 = _RAND_761[1:0];
  _RAND_762 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_247 = _RAND_762[1:0];
  _RAND_763 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_248 = _RAND_763[1:0];
  _RAND_764 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_249 = _RAND_764[1:0];
  _RAND_765 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_250 = _RAND_765[1:0];
  _RAND_766 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_251 = _RAND_766[1:0];
  _RAND_767 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_252 = _RAND_767[1:0];
  _RAND_768 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_253 = _RAND_768[1:0];
  _RAND_769 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_254 = _RAND_769[1:0];
  _RAND_770 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_255 = _RAND_770[1:0];
  _RAND_771 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_0 = _RAND_771[1:0];
  _RAND_772 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_1 = _RAND_772[1:0];
  _RAND_773 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_2 = _RAND_773[1:0];
  _RAND_774 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_3 = _RAND_774[1:0];
  _RAND_775 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_4 = _RAND_775[1:0];
  _RAND_776 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_5 = _RAND_776[1:0];
  _RAND_777 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_6 = _RAND_777[1:0];
  _RAND_778 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_7 = _RAND_778[1:0];
  _RAND_779 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_8 = _RAND_779[1:0];
  _RAND_780 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_9 = _RAND_780[1:0];
  _RAND_781 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_10 = _RAND_781[1:0];
  _RAND_782 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_11 = _RAND_782[1:0];
  _RAND_783 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_12 = _RAND_783[1:0];
  _RAND_784 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_13 = _RAND_784[1:0];
  _RAND_785 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_14 = _RAND_785[1:0];
  _RAND_786 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_15 = _RAND_786[1:0];
  _RAND_787 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_16 = _RAND_787[1:0];
  _RAND_788 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_17 = _RAND_788[1:0];
  _RAND_789 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_18 = _RAND_789[1:0];
  _RAND_790 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_19 = _RAND_790[1:0];
  _RAND_791 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_20 = _RAND_791[1:0];
  _RAND_792 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_21 = _RAND_792[1:0];
  _RAND_793 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_22 = _RAND_793[1:0];
  _RAND_794 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_23 = _RAND_794[1:0];
  _RAND_795 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_24 = _RAND_795[1:0];
  _RAND_796 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_25 = _RAND_796[1:0];
  _RAND_797 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_26 = _RAND_797[1:0];
  _RAND_798 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_27 = _RAND_798[1:0];
  _RAND_799 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_28 = _RAND_799[1:0];
  _RAND_800 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_29 = _RAND_800[1:0];
  _RAND_801 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_30 = _RAND_801[1:0];
  _RAND_802 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_31 = _RAND_802[1:0];
  _RAND_803 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_32 = _RAND_803[1:0];
  _RAND_804 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_33 = _RAND_804[1:0];
  _RAND_805 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_34 = _RAND_805[1:0];
  _RAND_806 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_35 = _RAND_806[1:0];
  _RAND_807 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_36 = _RAND_807[1:0];
  _RAND_808 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_37 = _RAND_808[1:0];
  _RAND_809 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_38 = _RAND_809[1:0];
  _RAND_810 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_39 = _RAND_810[1:0];
  _RAND_811 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_40 = _RAND_811[1:0];
  _RAND_812 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_41 = _RAND_812[1:0];
  _RAND_813 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_42 = _RAND_813[1:0];
  _RAND_814 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_43 = _RAND_814[1:0];
  _RAND_815 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_44 = _RAND_815[1:0];
  _RAND_816 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_45 = _RAND_816[1:0];
  _RAND_817 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_46 = _RAND_817[1:0];
  _RAND_818 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_47 = _RAND_818[1:0];
  _RAND_819 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_48 = _RAND_819[1:0];
  _RAND_820 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_49 = _RAND_820[1:0];
  _RAND_821 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_50 = _RAND_821[1:0];
  _RAND_822 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_51 = _RAND_822[1:0];
  _RAND_823 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_52 = _RAND_823[1:0];
  _RAND_824 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_53 = _RAND_824[1:0];
  _RAND_825 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_54 = _RAND_825[1:0];
  _RAND_826 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_55 = _RAND_826[1:0];
  _RAND_827 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_56 = _RAND_827[1:0];
  _RAND_828 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_57 = _RAND_828[1:0];
  _RAND_829 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_58 = _RAND_829[1:0];
  _RAND_830 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_59 = _RAND_830[1:0];
  _RAND_831 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_60 = _RAND_831[1:0];
  _RAND_832 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_61 = _RAND_832[1:0];
  _RAND_833 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_62 = _RAND_833[1:0];
  _RAND_834 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_63 = _RAND_834[1:0];
  _RAND_835 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_64 = _RAND_835[1:0];
  _RAND_836 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_65 = _RAND_836[1:0];
  _RAND_837 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_66 = _RAND_837[1:0];
  _RAND_838 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_67 = _RAND_838[1:0];
  _RAND_839 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_68 = _RAND_839[1:0];
  _RAND_840 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_69 = _RAND_840[1:0];
  _RAND_841 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_70 = _RAND_841[1:0];
  _RAND_842 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_71 = _RAND_842[1:0];
  _RAND_843 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_72 = _RAND_843[1:0];
  _RAND_844 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_73 = _RAND_844[1:0];
  _RAND_845 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_74 = _RAND_845[1:0];
  _RAND_846 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_75 = _RAND_846[1:0];
  _RAND_847 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_76 = _RAND_847[1:0];
  _RAND_848 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_77 = _RAND_848[1:0];
  _RAND_849 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_78 = _RAND_849[1:0];
  _RAND_850 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_79 = _RAND_850[1:0];
  _RAND_851 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_80 = _RAND_851[1:0];
  _RAND_852 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_81 = _RAND_852[1:0];
  _RAND_853 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_82 = _RAND_853[1:0];
  _RAND_854 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_83 = _RAND_854[1:0];
  _RAND_855 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_84 = _RAND_855[1:0];
  _RAND_856 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_85 = _RAND_856[1:0];
  _RAND_857 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_86 = _RAND_857[1:0];
  _RAND_858 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_87 = _RAND_858[1:0];
  _RAND_859 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_88 = _RAND_859[1:0];
  _RAND_860 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_89 = _RAND_860[1:0];
  _RAND_861 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_90 = _RAND_861[1:0];
  _RAND_862 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_91 = _RAND_862[1:0];
  _RAND_863 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_92 = _RAND_863[1:0];
  _RAND_864 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_93 = _RAND_864[1:0];
  _RAND_865 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_94 = _RAND_865[1:0];
  _RAND_866 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_95 = _RAND_866[1:0];
  _RAND_867 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_96 = _RAND_867[1:0];
  _RAND_868 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_97 = _RAND_868[1:0];
  _RAND_869 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_98 = _RAND_869[1:0];
  _RAND_870 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_99 = _RAND_870[1:0];
  _RAND_871 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_100 = _RAND_871[1:0];
  _RAND_872 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_101 = _RAND_872[1:0];
  _RAND_873 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_102 = _RAND_873[1:0];
  _RAND_874 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_103 = _RAND_874[1:0];
  _RAND_875 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_104 = _RAND_875[1:0];
  _RAND_876 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_105 = _RAND_876[1:0];
  _RAND_877 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_106 = _RAND_877[1:0];
  _RAND_878 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_107 = _RAND_878[1:0];
  _RAND_879 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_108 = _RAND_879[1:0];
  _RAND_880 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_109 = _RAND_880[1:0];
  _RAND_881 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_110 = _RAND_881[1:0];
  _RAND_882 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_111 = _RAND_882[1:0];
  _RAND_883 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_112 = _RAND_883[1:0];
  _RAND_884 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_113 = _RAND_884[1:0];
  _RAND_885 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_114 = _RAND_885[1:0];
  _RAND_886 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_115 = _RAND_886[1:0];
  _RAND_887 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_116 = _RAND_887[1:0];
  _RAND_888 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_117 = _RAND_888[1:0];
  _RAND_889 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_118 = _RAND_889[1:0];
  _RAND_890 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_119 = _RAND_890[1:0];
  _RAND_891 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_120 = _RAND_891[1:0];
  _RAND_892 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_121 = _RAND_892[1:0];
  _RAND_893 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_122 = _RAND_893[1:0];
  _RAND_894 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_123 = _RAND_894[1:0];
  _RAND_895 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_124 = _RAND_895[1:0];
  _RAND_896 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_125 = _RAND_896[1:0];
  _RAND_897 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_126 = _RAND_897[1:0];
  _RAND_898 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_127 = _RAND_898[1:0];
  _RAND_899 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_128 = _RAND_899[1:0];
  _RAND_900 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_129 = _RAND_900[1:0];
  _RAND_901 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_130 = _RAND_901[1:0];
  _RAND_902 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_131 = _RAND_902[1:0];
  _RAND_903 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_132 = _RAND_903[1:0];
  _RAND_904 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_133 = _RAND_904[1:0];
  _RAND_905 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_134 = _RAND_905[1:0];
  _RAND_906 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_135 = _RAND_906[1:0];
  _RAND_907 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_136 = _RAND_907[1:0];
  _RAND_908 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_137 = _RAND_908[1:0];
  _RAND_909 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_138 = _RAND_909[1:0];
  _RAND_910 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_139 = _RAND_910[1:0];
  _RAND_911 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_140 = _RAND_911[1:0];
  _RAND_912 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_141 = _RAND_912[1:0];
  _RAND_913 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_142 = _RAND_913[1:0];
  _RAND_914 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_143 = _RAND_914[1:0];
  _RAND_915 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_144 = _RAND_915[1:0];
  _RAND_916 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_145 = _RAND_916[1:0];
  _RAND_917 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_146 = _RAND_917[1:0];
  _RAND_918 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_147 = _RAND_918[1:0];
  _RAND_919 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_148 = _RAND_919[1:0];
  _RAND_920 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_149 = _RAND_920[1:0];
  _RAND_921 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_150 = _RAND_921[1:0];
  _RAND_922 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_151 = _RAND_922[1:0];
  _RAND_923 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_152 = _RAND_923[1:0];
  _RAND_924 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_153 = _RAND_924[1:0];
  _RAND_925 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_154 = _RAND_925[1:0];
  _RAND_926 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_155 = _RAND_926[1:0];
  _RAND_927 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_156 = _RAND_927[1:0];
  _RAND_928 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_157 = _RAND_928[1:0];
  _RAND_929 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_158 = _RAND_929[1:0];
  _RAND_930 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_159 = _RAND_930[1:0];
  _RAND_931 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_160 = _RAND_931[1:0];
  _RAND_932 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_161 = _RAND_932[1:0];
  _RAND_933 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_162 = _RAND_933[1:0];
  _RAND_934 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_163 = _RAND_934[1:0];
  _RAND_935 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_164 = _RAND_935[1:0];
  _RAND_936 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_165 = _RAND_936[1:0];
  _RAND_937 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_166 = _RAND_937[1:0];
  _RAND_938 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_167 = _RAND_938[1:0];
  _RAND_939 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_168 = _RAND_939[1:0];
  _RAND_940 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_169 = _RAND_940[1:0];
  _RAND_941 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_170 = _RAND_941[1:0];
  _RAND_942 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_171 = _RAND_942[1:0];
  _RAND_943 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_172 = _RAND_943[1:0];
  _RAND_944 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_173 = _RAND_944[1:0];
  _RAND_945 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_174 = _RAND_945[1:0];
  _RAND_946 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_175 = _RAND_946[1:0];
  _RAND_947 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_176 = _RAND_947[1:0];
  _RAND_948 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_177 = _RAND_948[1:0];
  _RAND_949 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_178 = _RAND_949[1:0];
  _RAND_950 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_179 = _RAND_950[1:0];
  _RAND_951 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_180 = _RAND_951[1:0];
  _RAND_952 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_181 = _RAND_952[1:0];
  _RAND_953 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_182 = _RAND_953[1:0];
  _RAND_954 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_183 = _RAND_954[1:0];
  _RAND_955 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_184 = _RAND_955[1:0];
  _RAND_956 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_185 = _RAND_956[1:0];
  _RAND_957 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_186 = _RAND_957[1:0];
  _RAND_958 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_187 = _RAND_958[1:0];
  _RAND_959 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_188 = _RAND_959[1:0];
  _RAND_960 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_189 = _RAND_960[1:0];
  _RAND_961 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_190 = _RAND_961[1:0];
  _RAND_962 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_191 = _RAND_962[1:0];
  _RAND_963 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_192 = _RAND_963[1:0];
  _RAND_964 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_193 = _RAND_964[1:0];
  _RAND_965 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_194 = _RAND_965[1:0];
  _RAND_966 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_195 = _RAND_966[1:0];
  _RAND_967 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_196 = _RAND_967[1:0];
  _RAND_968 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_197 = _RAND_968[1:0];
  _RAND_969 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_198 = _RAND_969[1:0];
  _RAND_970 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_199 = _RAND_970[1:0];
  _RAND_971 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_200 = _RAND_971[1:0];
  _RAND_972 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_201 = _RAND_972[1:0];
  _RAND_973 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_202 = _RAND_973[1:0];
  _RAND_974 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_203 = _RAND_974[1:0];
  _RAND_975 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_204 = _RAND_975[1:0];
  _RAND_976 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_205 = _RAND_976[1:0];
  _RAND_977 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_206 = _RAND_977[1:0];
  _RAND_978 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_207 = _RAND_978[1:0];
  _RAND_979 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_208 = _RAND_979[1:0];
  _RAND_980 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_209 = _RAND_980[1:0];
  _RAND_981 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_210 = _RAND_981[1:0];
  _RAND_982 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_211 = _RAND_982[1:0];
  _RAND_983 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_212 = _RAND_983[1:0];
  _RAND_984 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_213 = _RAND_984[1:0];
  _RAND_985 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_214 = _RAND_985[1:0];
  _RAND_986 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_215 = _RAND_986[1:0];
  _RAND_987 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_216 = _RAND_987[1:0];
  _RAND_988 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_217 = _RAND_988[1:0];
  _RAND_989 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_218 = _RAND_989[1:0];
  _RAND_990 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_219 = _RAND_990[1:0];
  _RAND_991 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_220 = _RAND_991[1:0];
  _RAND_992 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_221 = _RAND_992[1:0];
  _RAND_993 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_222 = _RAND_993[1:0];
  _RAND_994 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_223 = _RAND_994[1:0];
  _RAND_995 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_224 = _RAND_995[1:0];
  _RAND_996 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_225 = _RAND_996[1:0];
  _RAND_997 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_226 = _RAND_997[1:0];
  _RAND_998 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_227 = _RAND_998[1:0];
  _RAND_999 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_228 = _RAND_999[1:0];
  _RAND_1000 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_229 = _RAND_1000[1:0];
  _RAND_1001 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_230 = _RAND_1001[1:0];
  _RAND_1002 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_231 = _RAND_1002[1:0];
  _RAND_1003 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_232 = _RAND_1003[1:0];
  _RAND_1004 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_233 = _RAND_1004[1:0];
  _RAND_1005 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_234 = _RAND_1005[1:0];
  _RAND_1006 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_235 = _RAND_1006[1:0];
  _RAND_1007 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_236 = _RAND_1007[1:0];
  _RAND_1008 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_237 = _RAND_1008[1:0];
  _RAND_1009 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_238 = _RAND_1009[1:0];
  _RAND_1010 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_239 = _RAND_1010[1:0];
  _RAND_1011 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_240 = _RAND_1011[1:0];
  _RAND_1012 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_241 = _RAND_1012[1:0];
  _RAND_1013 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_242 = _RAND_1013[1:0];
  _RAND_1014 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_243 = _RAND_1014[1:0];
  _RAND_1015 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_244 = _RAND_1015[1:0];
  _RAND_1016 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_245 = _RAND_1016[1:0];
  _RAND_1017 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_246 = _RAND_1017[1:0];
  _RAND_1018 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_247 = _RAND_1018[1:0];
  _RAND_1019 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_248 = _RAND_1019[1:0];
  _RAND_1020 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_249 = _RAND_1020[1:0];
  _RAND_1021 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_250 = _RAND_1021[1:0];
  _RAND_1022 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_251 = _RAND_1022[1:0];
  _RAND_1023 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_252 = _RAND_1023[1:0];
  _RAND_1024 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_253 = _RAND_1024[1:0];
  _RAND_1025 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_254 = _RAND_1025[1:0];
  _RAND_1026 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_255 = _RAND_1026[1:0];
  _RAND_1027 = {1{`RANDOM}};
  exu_mp_way_f = _RAND_1027[0:0];
  _RAND_1028 = {1{`RANDOM}};
  exu_flush_final_d1 = _RAND_1028[0:0];
  _RAND_1029 = {8{`RANDOM}};
  btb_lru_b0_f = _RAND_1029[255:0];
  _RAND_1030 = {1{`RANDOM}};
  ifc_fetch_adder_prior = _RAND_1030[29:0];
  _RAND_1031 = {1{`RANDOM}};
  rets_out_0 = _RAND_1031[31:0];
  _RAND_1032 = {1{`RANDOM}};
  rets_out_1 = _RAND_1032[31:0];
  _RAND_1033 = {1{`RANDOM}};
  rets_out_2 = _RAND_1033[31:0];
  _RAND_1034 = {1{`RANDOM}};
  rets_out_3 = _RAND_1034[31:0];
  _RAND_1035 = {1{`RANDOM}};
  rets_out_4 = _RAND_1035[31:0];
  _RAND_1036 = {1{`RANDOM}};
  rets_out_5 = _RAND_1036[31:0];
  _RAND_1037 = {1{`RANDOM}};
  rets_out_6 = _RAND_1037[31:0];
  _RAND_1038 = {1{`RANDOM}};
  rets_out_7 = _RAND_1038[31:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    leak_one_f_d1 = 1'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_0 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_1 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_2 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_3 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_4 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_5 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_6 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_7 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_8 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_9 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_10 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_11 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_12 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_13 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_14 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_15 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_16 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_17 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_18 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_19 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_20 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_21 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_22 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_23 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_24 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_25 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_26 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_27 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_28 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_29 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_30 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_31 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_32 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_33 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_34 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_35 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_36 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_37 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_38 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_39 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_40 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_41 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_42 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_43 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_44 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_45 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_46 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_47 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_48 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_49 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_50 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_51 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_52 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_53 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_54 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_55 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_56 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_57 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_58 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_59 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_60 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_61 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_62 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_63 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_64 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_65 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_66 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_67 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_68 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_69 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_70 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_71 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_72 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_73 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_74 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_75 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_76 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_77 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_78 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_79 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_80 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_81 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_82 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_83 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_84 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_85 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_86 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_87 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_88 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_89 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_90 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_91 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_92 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_93 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_94 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_95 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_96 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_97 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_98 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_99 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_100 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_101 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_102 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_103 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_104 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_105 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_106 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_107 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_108 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_109 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_110 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_111 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_112 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_113 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_114 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_115 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_116 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_117 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_118 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_119 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_120 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_121 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_122 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_123 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_124 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_125 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_126 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_127 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_128 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_129 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_130 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_131 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_132 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_133 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_134 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_135 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_136 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_137 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_138 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_139 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_140 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_141 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_142 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_143 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_144 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_145 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_146 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_147 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_148 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_149 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_150 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_151 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_152 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_153 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_154 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_155 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_156 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_157 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_158 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_159 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_160 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_161 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_162 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_163 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_164 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_165 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_166 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_167 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_168 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_169 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_170 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_171 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_172 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_173 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_174 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_175 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_176 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_177 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_178 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_179 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_180 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_181 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_182 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_183 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_184 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_185 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_186 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_187 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_188 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_189 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_190 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_191 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_192 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_193 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_194 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_195 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_196 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_197 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_198 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_199 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_200 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_201 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_202 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_203 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_204 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_205 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_206 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_207 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_208 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_209 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_210 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_211 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_212 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_213 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_214 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_215 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_216 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_217 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_218 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_219 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_220 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_221 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_222 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_223 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_224 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_225 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_226 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_227 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_228 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_229 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_230 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_231 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_232 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_233 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_234 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_235 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_236 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_237 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_238 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_239 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_240 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_241 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_242 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_243 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_244 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_245 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_246 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_247 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_248 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_249 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_250 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_251 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_252 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_253 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_254 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_255 = 22'h0;
  end
  if (reset) begin
    dec_tlu_way_wb_f = 1'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_0 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_1 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_2 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_3 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_4 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_5 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_6 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_7 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_8 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_9 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_10 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_11 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_12 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_13 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_14 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_15 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_16 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_17 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_18 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_19 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_20 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_21 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_22 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_23 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_24 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_25 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_26 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_27 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_28 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_29 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_30 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_31 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_32 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_33 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_34 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_35 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_36 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_37 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_38 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_39 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_40 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_41 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_42 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_43 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_44 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_45 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_46 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_47 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_48 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_49 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_50 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_51 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_52 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_53 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_54 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_55 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_56 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_57 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_58 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_59 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_60 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_61 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_62 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_63 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_64 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_65 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_66 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_67 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_68 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_69 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_70 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_71 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_72 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_73 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_74 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_75 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_76 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_77 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_78 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_79 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_80 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_81 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_82 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_83 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_84 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_85 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_86 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_87 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_88 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_89 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_90 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_91 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_92 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_93 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_94 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_95 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_96 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_97 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_98 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_99 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_100 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_101 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_102 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_103 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_104 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_105 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_106 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_107 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_108 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_109 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_110 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_111 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_112 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_113 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_114 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_115 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_116 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_117 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_118 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_119 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_120 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_121 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_122 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_123 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_124 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_125 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_126 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_127 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_128 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_129 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_130 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_131 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_132 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_133 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_134 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_135 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_136 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_137 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_138 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_139 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_140 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_141 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_142 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_143 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_144 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_145 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_146 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_147 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_148 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_149 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_150 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_151 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_152 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_153 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_154 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_155 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_156 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_157 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_158 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_159 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_160 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_161 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_162 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_163 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_164 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_165 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_166 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_167 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_168 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_169 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_170 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_171 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_172 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_173 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_174 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_175 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_176 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_177 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_178 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_179 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_180 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_181 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_182 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_183 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_184 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_185 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_186 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_187 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_188 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_189 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_190 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_191 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_192 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_193 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_194 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_195 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_196 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_197 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_198 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_199 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_200 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_201 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_202 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_203 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_204 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_205 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_206 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_207 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_208 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_209 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_210 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_211 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_212 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_213 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_214 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_215 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_216 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_217 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_218 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_219 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_220 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_221 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_222 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_223 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_224 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_225 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_226 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_227 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_228 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_229 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_230 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_231 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_232 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_233 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_234 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_235 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_236 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_237 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_238 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_239 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_240 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_241 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_242 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_243 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_244 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_245 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_246 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_247 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_248 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_249 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_250 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_251 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_252 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_253 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_254 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_255 = 22'h0;
  end
  if (reset) begin
    fghr = 8'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_0 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_1 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_2 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_3 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_4 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_5 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_6 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_7 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_8 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_9 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_10 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_11 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_12 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_13 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_14 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_15 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_16 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_17 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_18 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_19 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_20 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_21 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_22 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_23 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_24 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_25 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_26 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_27 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_28 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_29 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_30 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_31 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_32 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_33 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_34 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_35 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_36 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_37 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_38 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_39 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_40 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_41 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_42 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_43 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_44 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_45 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_46 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_47 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_48 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_49 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_50 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_51 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_52 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_53 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_54 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_55 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_56 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_57 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_58 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_59 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_60 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_61 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_62 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_63 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_64 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_65 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_66 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_67 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_68 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_69 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_70 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_71 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_72 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_73 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_74 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_75 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_76 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_77 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_78 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_79 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_80 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_81 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_82 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_83 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_84 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_85 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_86 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_87 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_88 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_89 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_90 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_91 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_92 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_93 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_94 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_95 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_96 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_97 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_98 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_99 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_100 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_101 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_102 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_103 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_104 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_105 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_106 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_107 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_108 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_109 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_110 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_111 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_112 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_113 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_114 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_115 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_116 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_117 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_118 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_119 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_120 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_121 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_122 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_123 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_124 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_125 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_126 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_127 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_128 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_129 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_130 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_131 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_132 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_133 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_134 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_135 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_136 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_137 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_138 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_139 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_140 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_141 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_142 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_143 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_144 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_145 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_146 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_147 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_148 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_149 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_150 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_151 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_152 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_153 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_154 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_155 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_156 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_157 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_158 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_159 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_160 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_161 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_162 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_163 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_164 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_165 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_166 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_167 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_168 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_169 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_170 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_171 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_172 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_173 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_174 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_175 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_176 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_177 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_178 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_179 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_180 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_181 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_182 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_183 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_184 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_185 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_186 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_187 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_188 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_189 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_190 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_191 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_192 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_193 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_194 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_195 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_196 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_197 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_198 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_199 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_200 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_201 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_202 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_203 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_204 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_205 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_206 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_207 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_208 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_209 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_210 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_211 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_212 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_213 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_214 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_215 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_216 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_217 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_218 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_219 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_220 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_221 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_222 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_223 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_224 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_225 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_226 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_227 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_228 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_229 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_230 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_231 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_232 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_233 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_234 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_235 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_236 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_237 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_238 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_239 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_240 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_241 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_242 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_243 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_244 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_245 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_246 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_247 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_248 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_249 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_250 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_251 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_252 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_253 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_254 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_255 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_0 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_1 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_2 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_3 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_4 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_5 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_6 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_7 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_8 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_9 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_10 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_11 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_12 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_13 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_14 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_15 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_16 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_17 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_18 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_19 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_20 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_21 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_22 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_23 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_24 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_25 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_26 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_27 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_28 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_29 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_30 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_31 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_32 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_33 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_34 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_35 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_36 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_37 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_38 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_39 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_40 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_41 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_42 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_43 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_44 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_45 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_46 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_47 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_48 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_49 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_50 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_51 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_52 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_53 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_54 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_55 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_56 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_57 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_58 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_59 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_60 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_61 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_62 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_63 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_64 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_65 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_66 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_67 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_68 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_69 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_70 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_71 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_72 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_73 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_74 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_75 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_76 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_77 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_78 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_79 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_80 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_81 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_82 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_83 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_84 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_85 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_86 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_87 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_88 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_89 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_90 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_91 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_92 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_93 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_94 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_95 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_96 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_97 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_98 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_99 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_100 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_101 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_102 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_103 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_104 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_105 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_106 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_107 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_108 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_109 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_110 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_111 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_112 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_113 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_114 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_115 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_116 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_117 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_118 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_119 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_120 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_121 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_122 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_123 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_124 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_125 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_126 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_127 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_128 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_129 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_130 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_131 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_132 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_133 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_134 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_135 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_136 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_137 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_138 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_139 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_140 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_141 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_142 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_143 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_144 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_145 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_146 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_147 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_148 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_149 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_150 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_151 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_152 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_153 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_154 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_155 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_156 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_157 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_158 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_159 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_160 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_161 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_162 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_163 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_164 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_165 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_166 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_167 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_168 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_169 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_170 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_171 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_172 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_173 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_174 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_175 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_176 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_177 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_178 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_179 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_180 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_181 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_182 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_183 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_184 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_185 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_186 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_187 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_188 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_189 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_190 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_191 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_192 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_193 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_194 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_195 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_196 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_197 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_198 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_199 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_200 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_201 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_202 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_203 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_204 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_205 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_206 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_207 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_208 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_209 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_210 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_211 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_212 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_213 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_214 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_215 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_216 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_217 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_218 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_219 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_220 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_221 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_222 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_223 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_224 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_225 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_226 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_227 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_228 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_229 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_230 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_231 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_232 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_233 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_234 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_235 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_236 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_237 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_238 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_239 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_240 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_241 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_242 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_243 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_244 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_245 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_246 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_247 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_248 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_249 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_250 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_251 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_252 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_253 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_254 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_255 = 2'h0;
  end
  if (reset) begin
    exu_mp_way_f = 1'h0;
  end
  if (reset) begin
    exu_flush_final_d1 = 1'h0;
  end
  if (reset) begin
    btb_lru_b0_f = 256'h0;
  end
  if (reset) begin
    ifc_fetch_adder_prior = 30'h0;
  end
  if (reset) begin
    rets_out_0 = 32'h0;
  end
  if (reset) begin
    rets_out_1 = 32'h0;
  end
  if (reset) begin
    rets_out_2 = 32'h0;
  end
  if (reset) begin
    rets_out_3 = 32'h0;
  end
  if (reset) begin
    rets_out_4 = 32'h0;
  end
  if (reset) begin
    rets_out_5 = 32'h0;
  end
  if (reset) begin
    rets_out_6 = 32'h0;
  end
  if (reset) begin
    rets_out_7 = 32'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      leak_one_f_d1 <= 1'h0;
    end else begin
      leak_one_f_d1 <= _T_40 | _T_41;
    end
  end
  always @(posedge rvclkhdr_10_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_0 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_0 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_11_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_1 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_1 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_12_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_2 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_2 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_13_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_3 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_3 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_14_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_4 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_4 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_15_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_5 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_5 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_16_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_6 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_6 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_17_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_7 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_7 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_18_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_8 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_8 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_19_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_9 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_9 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_20_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_10 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_10 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_21_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_11 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_11 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_22_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_12 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_12 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_23_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_13 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_13 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_24_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_14 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_14 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_25_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_15 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_15 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_26_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_16 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_16 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_27_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_17 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_17 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_28_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_18 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_18 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_29_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_19 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_19 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_30_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_20 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_20 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_31_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_21 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_21 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_32_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_22 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_22 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_33_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_23 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_23 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_34_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_24 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_24 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_35_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_25 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_25 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_36_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_26 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_26 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_37_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_27 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_27 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_38_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_28 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_28 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_39_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_29 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_29 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_40_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_30 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_30 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_41_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_31 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_31 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_42_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_32 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_32 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_43_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_33 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_33 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_44_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_34 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_34 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_45_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_35 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_35 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_46_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_36 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_36 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_47_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_37 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_37 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_48_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_38 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_38 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_49_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_39 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_39 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_50_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_40 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_40 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_51_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_41 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_41 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_52_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_42 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_42 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_53_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_43 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_43 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_54_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_44 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_44 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_55_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_45 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_45 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_56_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_46 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_46 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_57_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_47 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_47 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_58_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_48 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_48 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_59_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_49 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_49 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_60_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_50 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_50 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_61_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_51 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_51 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_62_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_52 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_52 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_63_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_53 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_53 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_64_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_54 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_54 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_65_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_55 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_55 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_66_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_56 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_56 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_67_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_57 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_57 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_68_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_58 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_58 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_69_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_59 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_59 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_70_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_60 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_60 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_71_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_61 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_61 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_72_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_62 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_62 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_73_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_63 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_63 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_74_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_64 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_64 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_75_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_65 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_65 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_76_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_66 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_66 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_77_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_67 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_67 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_78_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_68 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_68 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_79_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_69 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_69 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_80_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_70 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_70 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_81_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_71 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_71 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_82_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_72 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_72 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_83_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_73 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_73 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_84_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_74 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_74 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_85_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_75 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_75 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_76 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_76 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_77 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_77 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_78 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_78 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_79 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_79 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_80 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_80 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_81 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_81 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_82 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_82 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_83 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_83 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_94_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_84 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_84 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_95_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_85 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_85 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_96_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_86 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_86 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_97_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_87 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_87 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_98_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_88 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_88 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_99_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_89 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_89 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_100_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_90 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_90 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_101_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_91 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_91 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_102_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_92 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_92 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_103_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_93 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_93 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_104_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_94 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_94 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_105_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_95 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_95 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_106_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_96 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_96 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_107_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_97 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_97 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_108_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_98 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_98 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_109_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_99 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_99 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_110_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_100 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_100 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_111_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_101 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_101 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_112_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_102 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_102 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_113_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_103 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_103 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_114_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_104 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_104 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_115_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_105 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_105 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_116_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_106 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_106 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_117_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_107 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_107 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_118_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_108 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_108 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_119_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_109 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_109 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_120_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_110 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_110 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_121_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_111 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_111 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_122_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_112 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_112 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_123_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_113 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_113 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_124_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_114 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_114 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_125_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_115 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_115 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_126_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_116 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_116 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_127_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_117 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_117 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_128_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_118 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_118 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_129_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_119 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_119 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_130_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_120 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_120 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_131_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_121 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_121 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_132_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_122 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_122 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_133_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_123 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_123 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_134_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_124 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_124 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_135_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_125 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_125 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_136_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_126 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_126 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_137_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_127 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_127 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_138_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_128 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_128 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_139_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_129 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_129 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_140_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_130 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_130 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_141_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_131 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_131 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_142_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_132 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_132 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_143_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_133 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_133 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_144_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_134 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_134 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_145_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_135 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_135 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_146_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_136 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_136 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_147_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_137 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_137 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_148_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_138 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_138 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_149_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_139 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_139 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_150_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_140 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_140 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_151_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_141 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_141 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_152_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_142 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_142 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_153_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_143 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_143 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_154_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_144 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_144 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_155_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_145 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_145 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_156_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_146 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_146 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_157_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_147 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_147 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_158_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_148 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_148 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_159_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_149 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_149 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_160_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_150 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_150 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_161_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_151 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_151 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_162_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_152 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_152 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_163_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_153 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_153 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_164_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_154 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_154 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_165_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_155 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_155 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_166_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_156 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_156 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_167_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_157 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_157 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_168_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_158 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_158 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_169_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_159 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_159 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_170_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_160 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_160 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_171_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_161 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_161 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_172_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_162 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_162 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_173_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_163 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_163 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_174_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_164 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_164 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_175_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_165 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_165 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_176_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_166 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_166 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_177_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_167 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_167 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_178_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_168 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_168 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_179_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_169 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_169 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_180_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_170 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_170 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_181_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_171 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_171 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_182_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_172 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_172 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_183_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_173 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_173 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_184_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_174 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_174 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_185_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_175 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_175 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_186_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_176 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_176 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_187_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_177 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_177 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_188_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_178 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_178 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_189_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_179 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_179 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_190_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_180 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_180 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_191_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_181 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_181 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_192_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_182 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_182 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_193_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_183 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_183 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_194_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_184 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_184 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_195_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_185 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_185 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_196_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_186 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_186 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_197_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_187 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_187 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_198_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_188 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_188 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_199_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_189 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_189 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_200_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_190 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_190 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_201_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_191 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_191 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_202_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_192 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_192 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_203_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_193 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_193 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_204_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_194 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_194 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_205_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_195 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_195 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_206_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_196 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_196 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_207_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_197 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_197 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_208_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_198 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_198 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_209_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_199 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_199 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_210_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_200 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_200 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_211_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_201 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_201 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_212_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_202 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_202 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_213_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_203 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_203 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_214_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_204 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_204 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_215_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_205 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_205 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_216_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_206 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_206 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_217_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_207 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_207 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_218_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_208 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_208 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_219_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_209 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_209 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_220_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_210 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_210 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_221_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_211 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_211 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_222_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_212 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_212 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_223_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_213 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_213 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_224_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_214 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_214 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_225_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_215 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_215 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_226_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_216 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_216 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_227_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_217 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_217 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_228_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_218 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_218 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_229_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_219 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_219 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_230_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_220 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_220 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_231_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_221 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_221 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_232_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_222 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_222 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_233_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_223 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_223 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_234_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_224 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_224 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_235_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_225 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_225 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_236_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_226 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_226 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_237_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_227 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_227 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_238_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_228 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_228 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_239_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_229 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_229 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_240_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_230 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_230 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_241_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_231 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_231 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_242_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_232 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_232 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_243_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_233 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_233 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_244_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_234 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_234 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_245_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_235 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_235 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_246_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_236 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_236 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_247_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_237 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_237 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_248_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_238 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_238 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_249_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_239 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_239 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_250_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_240 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_240 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_251_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_241 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_241 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_252_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_242 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_242 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_253_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_243 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_243 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_254_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_244 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_244 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_255_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_245 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_245 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_256_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_246 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_246 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_257_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_247 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_247 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_258_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_248 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_248 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_259_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_249 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_249 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_260_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_250 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_250 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_261_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_251 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_251 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_262_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_252 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_252 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_263_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_253 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_253 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_264_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_254 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_254 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_265_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_255 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_255 <= {_T_537,_T_534};
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      dec_tlu_way_wb_f <= 1'h0;
    end else begin
      dec_tlu_way_wb_f <= io_dec_tlu_br0_r_pkt_way;
    end
  end
  always @(posedge rvclkhdr_266_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_0 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_0 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_267_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_1 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_1 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_268_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_2 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_2 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_269_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_3 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_3 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_270_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_4 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_4 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_271_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_5 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_5 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_272_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_6 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_6 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_273_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_7 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_7 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_274_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_8 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_8 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_275_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_9 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_9 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_276_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_10 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_10 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_277_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_11 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_11 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_278_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_12 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_12 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_279_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_13 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_13 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_280_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_14 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_14 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_281_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_15 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_15 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_282_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_16 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_16 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_283_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_17 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_17 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_284_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_18 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_18 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_285_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_19 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_19 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_286_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_20 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_20 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_287_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_21 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_21 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_288_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_22 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_22 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_289_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_23 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_23 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_290_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_24 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_24 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_291_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_25 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_25 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_292_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_26 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_26 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_293_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_27 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_27 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_294_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_28 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_28 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_295_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_29 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_29 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_296_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_30 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_30 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_297_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_31 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_31 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_298_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_32 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_32 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_299_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_33 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_33 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_300_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_34 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_34 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_301_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_35 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_35 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_302_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_36 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_36 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_303_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_37 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_37 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_304_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_38 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_38 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_305_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_39 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_39 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_306_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_40 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_40 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_307_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_41 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_41 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_308_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_42 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_42 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_309_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_43 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_43 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_310_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_44 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_44 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_311_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_45 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_45 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_312_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_46 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_46 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_313_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_47 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_47 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_314_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_48 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_48 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_315_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_49 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_49 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_316_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_50 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_50 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_317_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_51 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_51 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_318_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_52 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_52 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_319_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_53 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_53 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_320_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_54 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_54 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_321_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_55 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_55 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_322_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_56 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_56 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_323_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_57 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_57 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_324_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_58 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_58 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_325_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_59 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_59 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_326_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_60 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_60 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_327_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_61 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_61 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_328_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_62 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_62 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_329_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_63 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_63 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_330_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_64 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_64 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_331_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_65 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_65 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_332_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_66 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_66 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_333_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_67 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_67 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_334_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_68 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_68 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_335_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_69 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_69 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_336_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_70 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_70 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_337_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_71 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_71 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_338_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_72 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_72 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_339_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_73 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_73 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_340_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_74 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_74 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_341_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_75 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_75 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_342_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_76 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_76 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_343_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_77 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_77 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_344_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_78 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_78 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_345_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_79 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_79 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_346_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_80 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_80 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_347_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_81 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_81 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_348_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_82 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_82 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_349_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_83 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_83 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_350_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_84 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_84 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_351_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_85 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_85 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_352_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_86 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_86 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_353_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_87 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_87 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_354_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_88 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_88 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_355_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_89 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_89 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_356_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_90 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_90 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_357_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_91 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_91 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_358_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_92 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_92 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_359_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_93 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_93 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_360_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_94 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_94 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_361_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_95 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_95 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_362_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_96 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_96 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_363_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_97 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_97 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_364_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_98 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_98 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_365_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_99 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_99 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_366_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_100 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_100 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_367_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_101 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_101 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_368_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_102 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_102 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_369_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_103 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_103 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_370_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_104 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_104 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_371_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_105 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_105 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_372_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_106 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_106 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_373_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_107 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_107 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_374_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_108 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_108 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_375_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_109 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_109 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_376_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_110 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_110 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_377_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_111 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_111 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_378_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_112 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_112 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_379_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_113 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_113 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_380_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_114 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_114 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_381_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_115 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_115 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_382_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_116 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_116 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_383_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_117 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_117 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_384_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_118 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_118 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_385_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_119 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_119 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_386_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_120 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_120 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_387_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_121 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_121 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_388_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_122 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_122 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_389_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_123 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_123 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_390_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_124 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_124 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_391_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_125 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_125 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_392_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_126 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_126 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_393_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_127 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_127 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_394_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_128 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_128 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_395_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_129 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_129 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_396_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_130 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_130 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_397_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_131 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_131 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_398_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_132 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_132 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_399_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_133 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_133 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_400_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_134 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_134 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_401_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_135 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_135 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_402_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_136 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_136 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_403_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_137 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_137 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_404_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_138 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_138 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_405_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_139 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_139 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_406_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_140 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_140 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_407_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_141 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_141 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_408_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_142 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_142 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_409_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_143 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_143 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_410_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_144 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_144 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_411_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_145 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_145 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_412_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_146 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_146 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_413_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_147 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_147 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_414_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_148 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_148 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_415_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_149 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_149 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_416_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_150 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_150 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_417_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_151 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_151 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_418_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_152 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_152 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_419_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_153 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_153 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_420_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_154 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_154 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_421_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_155 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_155 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_422_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_156 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_156 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_423_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_157 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_157 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_424_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_158 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_158 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_425_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_159 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_159 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_426_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_160 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_160 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_427_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_161 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_161 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_428_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_162 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_162 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_429_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_163 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_163 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_430_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_164 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_164 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_431_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_165 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_165 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_432_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_166 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_166 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_433_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_167 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_167 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_434_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_168 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_168 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_435_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_169 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_169 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_436_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_170 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_170 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_437_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_171 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_171 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_438_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_172 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_172 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_439_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_173 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_173 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_440_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_174 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_174 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_441_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_175 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_175 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_442_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_176 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_176 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_443_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_177 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_177 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_444_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_178 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_178 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_445_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_179 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_179 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_446_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_180 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_180 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_447_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_181 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_181 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_448_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_182 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_182 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_449_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_183 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_183 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_450_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_184 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_184 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_451_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_185 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_185 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_452_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_186 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_186 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_453_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_187 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_187 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_454_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_188 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_188 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_455_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_189 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_189 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_456_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_190 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_190 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_457_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_191 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_191 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_458_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_192 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_192 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_459_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_193 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_193 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_460_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_194 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_194 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_461_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_195 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_195 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_462_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_196 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_196 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_463_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_197 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_197 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_464_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_198 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_198 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_465_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_199 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_199 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_466_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_200 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_200 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_467_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_201 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_201 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_468_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_202 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_202 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_469_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_203 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_203 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_470_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_204 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_204 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_471_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_205 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_205 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_472_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_206 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_206 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_473_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_207 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_207 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_474_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_208 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_208 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_475_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_209 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_209 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_476_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_210 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_210 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_477_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_211 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_211 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_478_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_212 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_212 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_479_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_213 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_213 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_480_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_214 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_214 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_481_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_215 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_215 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_482_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_216 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_216 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_483_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_217 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_217 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_484_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_218 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_218 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_485_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_219 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_219 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_486_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_220 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_220 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_487_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_221 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_221 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_488_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_222 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_222 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_489_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_223 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_223 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_490_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_224 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_224 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_491_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_225 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_225 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_492_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_226 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_226 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_493_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_227 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_227 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_494_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_228 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_228 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_495_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_229 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_229 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_496_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_230 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_230 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_497_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_231 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_231 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_498_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_232 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_232 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_499_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_233 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_233 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_500_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_234 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_234 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_501_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_235 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_235 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_502_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_236 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_236 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_503_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_237 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_237 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_504_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_238 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_238 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_505_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_239 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_239 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_506_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_240 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_240 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_507_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_241 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_241 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_508_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_242 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_242 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_509_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_243 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_243 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_510_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_244 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_244 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_511_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_245 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_245 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_512_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_246 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_246 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_513_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_247 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_247 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_514_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_248 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_248 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_515_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_249 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_249 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_516_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_250 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_250 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_517_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_251 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_251 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_518_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_252 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_252 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_519_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_253 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_253 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_520_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_254 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_254 <= {_T_537,_T_534};
    end
  end
  always @(posedge rvclkhdr_521_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_255 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_255 <= {_T_537,_T_534};
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      fghr <= 8'h0;
    end else begin
      fghr <= _T_338 | _T_337;
    end
  end
  always @(posedge rvclkhdr_538_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_0 <= 2'h0;
    end else if (bht_bank_sel_1_0_0) begin
      if (_T_8869) begin
        bht_bank_rd_data_out_1_0 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_0 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_538_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_1 <= 2'h0;
    end else if (bht_bank_sel_1_0_1) begin
      if (_T_8878) begin
        bht_bank_rd_data_out_1_1 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_1 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_538_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_2 <= 2'h0;
    end else if (bht_bank_sel_1_0_2) begin
      if (_T_8887) begin
        bht_bank_rd_data_out_1_2 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_2 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_538_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_3 <= 2'h0;
    end else if (bht_bank_sel_1_0_3) begin
      if (_T_8896) begin
        bht_bank_rd_data_out_1_3 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_3 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_538_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_4 <= 2'h0;
    end else if (bht_bank_sel_1_0_4) begin
      if (_T_8905) begin
        bht_bank_rd_data_out_1_4 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_4 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_538_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_5 <= 2'h0;
    end else if (bht_bank_sel_1_0_5) begin
      if (_T_8914) begin
        bht_bank_rd_data_out_1_5 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_5 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_538_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_6 <= 2'h0;
    end else if (bht_bank_sel_1_0_6) begin
      if (_T_8923) begin
        bht_bank_rd_data_out_1_6 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_6 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_538_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_7 <= 2'h0;
    end else if (bht_bank_sel_1_0_7) begin
      if (_T_8932) begin
        bht_bank_rd_data_out_1_7 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_7 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_538_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_8 <= 2'h0;
    end else if (bht_bank_sel_1_0_8) begin
      if (_T_8941) begin
        bht_bank_rd_data_out_1_8 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_8 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_538_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_9 <= 2'h0;
    end else if (bht_bank_sel_1_0_9) begin
      if (_T_8950) begin
        bht_bank_rd_data_out_1_9 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_9 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_538_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_10 <= 2'h0;
    end else if (bht_bank_sel_1_0_10) begin
      if (_T_8959) begin
        bht_bank_rd_data_out_1_10 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_10 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_538_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_11 <= 2'h0;
    end else if (bht_bank_sel_1_0_11) begin
      if (_T_8968) begin
        bht_bank_rd_data_out_1_11 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_11 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_538_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_12 <= 2'h0;
    end else if (bht_bank_sel_1_0_12) begin
      if (_T_8977) begin
        bht_bank_rd_data_out_1_12 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_12 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_538_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_13 <= 2'h0;
    end else if (bht_bank_sel_1_0_13) begin
      if (_T_8986) begin
        bht_bank_rd_data_out_1_13 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_13 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_538_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_14 <= 2'h0;
    end else if (bht_bank_sel_1_0_14) begin
      if (_T_8995) begin
        bht_bank_rd_data_out_1_14 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_14 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_538_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_15 <= 2'h0;
    end else if (bht_bank_sel_1_0_15) begin
      if (_T_9004) begin
        bht_bank_rd_data_out_1_15 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_15 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_539_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_16 <= 2'h0;
    end else if (bht_bank_sel_1_1_0) begin
      if (_T_9013) begin
        bht_bank_rd_data_out_1_16 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_16 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_539_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_17 <= 2'h0;
    end else if (bht_bank_sel_1_1_1) begin
      if (_T_9022) begin
        bht_bank_rd_data_out_1_17 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_17 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_539_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_18 <= 2'h0;
    end else if (bht_bank_sel_1_1_2) begin
      if (_T_9031) begin
        bht_bank_rd_data_out_1_18 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_18 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_539_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_19 <= 2'h0;
    end else if (bht_bank_sel_1_1_3) begin
      if (_T_9040) begin
        bht_bank_rd_data_out_1_19 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_19 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_539_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_20 <= 2'h0;
    end else if (bht_bank_sel_1_1_4) begin
      if (_T_9049) begin
        bht_bank_rd_data_out_1_20 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_20 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_539_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_21 <= 2'h0;
    end else if (bht_bank_sel_1_1_5) begin
      if (_T_9058) begin
        bht_bank_rd_data_out_1_21 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_21 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_539_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_22 <= 2'h0;
    end else if (bht_bank_sel_1_1_6) begin
      if (_T_9067) begin
        bht_bank_rd_data_out_1_22 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_22 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_539_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_23 <= 2'h0;
    end else if (bht_bank_sel_1_1_7) begin
      if (_T_9076) begin
        bht_bank_rd_data_out_1_23 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_23 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_539_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_24 <= 2'h0;
    end else if (bht_bank_sel_1_1_8) begin
      if (_T_9085) begin
        bht_bank_rd_data_out_1_24 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_24 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_539_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_25 <= 2'h0;
    end else if (bht_bank_sel_1_1_9) begin
      if (_T_9094) begin
        bht_bank_rd_data_out_1_25 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_25 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_539_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_26 <= 2'h0;
    end else if (bht_bank_sel_1_1_10) begin
      if (_T_9103) begin
        bht_bank_rd_data_out_1_26 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_26 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_539_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_27 <= 2'h0;
    end else if (bht_bank_sel_1_1_11) begin
      if (_T_9112) begin
        bht_bank_rd_data_out_1_27 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_27 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_539_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_28 <= 2'h0;
    end else if (bht_bank_sel_1_1_12) begin
      if (_T_9121) begin
        bht_bank_rd_data_out_1_28 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_28 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_539_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_29 <= 2'h0;
    end else if (bht_bank_sel_1_1_13) begin
      if (_T_9130) begin
        bht_bank_rd_data_out_1_29 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_29 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_539_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_30 <= 2'h0;
    end else if (bht_bank_sel_1_1_14) begin
      if (_T_9139) begin
        bht_bank_rd_data_out_1_30 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_30 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_539_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_31 <= 2'h0;
    end else if (bht_bank_sel_1_1_15) begin
      if (_T_9148) begin
        bht_bank_rd_data_out_1_31 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_31 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_540_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_32 <= 2'h0;
    end else if (bht_bank_sel_1_2_0) begin
      if (_T_9157) begin
        bht_bank_rd_data_out_1_32 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_32 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_540_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_33 <= 2'h0;
    end else if (bht_bank_sel_1_2_1) begin
      if (_T_9166) begin
        bht_bank_rd_data_out_1_33 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_33 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_540_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_34 <= 2'h0;
    end else if (bht_bank_sel_1_2_2) begin
      if (_T_9175) begin
        bht_bank_rd_data_out_1_34 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_34 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_540_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_35 <= 2'h0;
    end else if (bht_bank_sel_1_2_3) begin
      if (_T_9184) begin
        bht_bank_rd_data_out_1_35 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_35 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_540_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_36 <= 2'h0;
    end else if (bht_bank_sel_1_2_4) begin
      if (_T_9193) begin
        bht_bank_rd_data_out_1_36 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_36 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_540_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_37 <= 2'h0;
    end else if (bht_bank_sel_1_2_5) begin
      if (_T_9202) begin
        bht_bank_rd_data_out_1_37 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_37 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_540_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_38 <= 2'h0;
    end else if (bht_bank_sel_1_2_6) begin
      if (_T_9211) begin
        bht_bank_rd_data_out_1_38 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_38 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_540_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_39 <= 2'h0;
    end else if (bht_bank_sel_1_2_7) begin
      if (_T_9220) begin
        bht_bank_rd_data_out_1_39 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_39 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_540_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_40 <= 2'h0;
    end else if (bht_bank_sel_1_2_8) begin
      if (_T_9229) begin
        bht_bank_rd_data_out_1_40 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_40 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_540_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_41 <= 2'h0;
    end else if (bht_bank_sel_1_2_9) begin
      if (_T_9238) begin
        bht_bank_rd_data_out_1_41 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_41 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_540_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_42 <= 2'h0;
    end else if (bht_bank_sel_1_2_10) begin
      if (_T_9247) begin
        bht_bank_rd_data_out_1_42 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_42 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_540_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_43 <= 2'h0;
    end else if (bht_bank_sel_1_2_11) begin
      if (_T_9256) begin
        bht_bank_rd_data_out_1_43 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_43 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_540_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_44 <= 2'h0;
    end else if (bht_bank_sel_1_2_12) begin
      if (_T_9265) begin
        bht_bank_rd_data_out_1_44 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_44 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_540_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_45 <= 2'h0;
    end else if (bht_bank_sel_1_2_13) begin
      if (_T_9274) begin
        bht_bank_rd_data_out_1_45 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_45 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_540_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_46 <= 2'h0;
    end else if (bht_bank_sel_1_2_14) begin
      if (_T_9283) begin
        bht_bank_rd_data_out_1_46 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_46 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_540_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_47 <= 2'h0;
    end else if (bht_bank_sel_1_2_15) begin
      if (_T_9292) begin
        bht_bank_rd_data_out_1_47 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_47 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_541_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_48 <= 2'h0;
    end else if (bht_bank_sel_1_3_0) begin
      if (_T_9301) begin
        bht_bank_rd_data_out_1_48 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_48 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_541_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_49 <= 2'h0;
    end else if (bht_bank_sel_1_3_1) begin
      if (_T_9310) begin
        bht_bank_rd_data_out_1_49 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_49 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_541_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_50 <= 2'h0;
    end else if (bht_bank_sel_1_3_2) begin
      if (_T_9319) begin
        bht_bank_rd_data_out_1_50 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_50 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_541_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_51 <= 2'h0;
    end else if (bht_bank_sel_1_3_3) begin
      if (_T_9328) begin
        bht_bank_rd_data_out_1_51 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_51 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_541_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_52 <= 2'h0;
    end else if (bht_bank_sel_1_3_4) begin
      if (_T_9337) begin
        bht_bank_rd_data_out_1_52 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_52 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_541_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_53 <= 2'h0;
    end else if (bht_bank_sel_1_3_5) begin
      if (_T_9346) begin
        bht_bank_rd_data_out_1_53 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_53 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_541_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_54 <= 2'h0;
    end else if (bht_bank_sel_1_3_6) begin
      if (_T_9355) begin
        bht_bank_rd_data_out_1_54 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_54 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_541_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_55 <= 2'h0;
    end else if (bht_bank_sel_1_3_7) begin
      if (_T_9364) begin
        bht_bank_rd_data_out_1_55 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_55 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_541_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_56 <= 2'h0;
    end else if (bht_bank_sel_1_3_8) begin
      if (_T_9373) begin
        bht_bank_rd_data_out_1_56 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_56 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_541_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_57 <= 2'h0;
    end else if (bht_bank_sel_1_3_9) begin
      if (_T_9382) begin
        bht_bank_rd_data_out_1_57 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_57 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_541_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_58 <= 2'h0;
    end else if (bht_bank_sel_1_3_10) begin
      if (_T_9391) begin
        bht_bank_rd_data_out_1_58 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_58 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_541_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_59 <= 2'h0;
    end else if (bht_bank_sel_1_3_11) begin
      if (_T_9400) begin
        bht_bank_rd_data_out_1_59 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_59 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_541_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_60 <= 2'h0;
    end else if (bht_bank_sel_1_3_12) begin
      if (_T_9409) begin
        bht_bank_rd_data_out_1_60 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_60 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_541_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_61 <= 2'h0;
    end else if (bht_bank_sel_1_3_13) begin
      if (_T_9418) begin
        bht_bank_rd_data_out_1_61 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_61 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_541_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_62 <= 2'h0;
    end else if (bht_bank_sel_1_3_14) begin
      if (_T_9427) begin
        bht_bank_rd_data_out_1_62 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_62 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_541_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_63 <= 2'h0;
    end else if (bht_bank_sel_1_3_15) begin
      if (_T_9436) begin
        bht_bank_rd_data_out_1_63 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_63 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_542_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_64 <= 2'h0;
    end else if (bht_bank_sel_1_4_0) begin
      if (_T_9445) begin
        bht_bank_rd_data_out_1_64 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_64 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_542_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_65 <= 2'h0;
    end else if (bht_bank_sel_1_4_1) begin
      if (_T_9454) begin
        bht_bank_rd_data_out_1_65 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_65 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_542_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_66 <= 2'h0;
    end else if (bht_bank_sel_1_4_2) begin
      if (_T_9463) begin
        bht_bank_rd_data_out_1_66 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_66 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_542_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_67 <= 2'h0;
    end else if (bht_bank_sel_1_4_3) begin
      if (_T_9472) begin
        bht_bank_rd_data_out_1_67 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_67 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_542_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_68 <= 2'h0;
    end else if (bht_bank_sel_1_4_4) begin
      if (_T_9481) begin
        bht_bank_rd_data_out_1_68 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_68 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_542_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_69 <= 2'h0;
    end else if (bht_bank_sel_1_4_5) begin
      if (_T_9490) begin
        bht_bank_rd_data_out_1_69 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_69 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_542_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_70 <= 2'h0;
    end else if (bht_bank_sel_1_4_6) begin
      if (_T_9499) begin
        bht_bank_rd_data_out_1_70 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_70 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_542_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_71 <= 2'h0;
    end else if (bht_bank_sel_1_4_7) begin
      if (_T_9508) begin
        bht_bank_rd_data_out_1_71 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_71 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_542_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_72 <= 2'h0;
    end else if (bht_bank_sel_1_4_8) begin
      if (_T_9517) begin
        bht_bank_rd_data_out_1_72 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_72 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_542_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_73 <= 2'h0;
    end else if (bht_bank_sel_1_4_9) begin
      if (_T_9526) begin
        bht_bank_rd_data_out_1_73 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_73 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_542_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_74 <= 2'h0;
    end else if (bht_bank_sel_1_4_10) begin
      if (_T_9535) begin
        bht_bank_rd_data_out_1_74 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_74 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_542_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_75 <= 2'h0;
    end else if (bht_bank_sel_1_4_11) begin
      if (_T_9544) begin
        bht_bank_rd_data_out_1_75 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_75 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_542_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_76 <= 2'h0;
    end else if (bht_bank_sel_1_4_12) begin
      if (_T_9553) begin
        bht_bank_rd_data_out_1_76 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_76 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_542_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_77 <= 2'h0;
    end else if (bht_bank_sel_1_4_13) begin
      if (_T_9562) begin
        bht_bank_rd_data_out_1_77 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_77 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_542_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_78 <= 2'h0;
    end else if (bht_bank_sel_1_4_14) begin
      if (_T_9571) begin
        bht_bank_rd_data_out_1_78 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_78 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_542_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_79 <= 2'h0;
    end else if (bht_bank_sel_1_4_15) begin
      if (_T_9580) begin
        bht_bank_rd_data_out_1_79 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_79 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_543_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_80 <= 2'h0;
    end else if (bht_bank_sel_1_5_0) begin
      if (_T_9589) begin
        bht_bank_rd_data_out_1_80 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_80 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_543_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_81 <= 2'h0;
    end else if (bht_bank_sel_1_5_1) begin
      if (_T_9598) begin
        bht_bank_rd_data_out_1_81 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_81 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_543_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_82 <= 2'h0;
    end else if (bht_bank_sel_1_5_2) begin
      if (_T_9607) begin
        bht_bank_rd_data_out_1_82 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_82 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_543_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_83 <= 2'h0;
    end else if (bht_bank_sel_1_5_3) begin
      if (_T_9616) begin
        bht_bank_rd_data_out_1_83 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_83 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_543_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_84 <= 2'h0;
    end else if (bht_bank_sel_1_5_4) begin
      if (_T_9625) begin
        bht_bank_rd_data_out_1_84 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_84 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_543_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_85 <= 2'h0;
    end else if (bht_bank_sel_1_5_5) begin
      if (_T_9634) begin
        bht_bank_rd_data_out_1_85 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_85 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_543_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_86 <= 2'h0;
    end else if (bht_bank_sel_1_5_6) begin
      if (_T_9643) begin
        bht_bank_rd_data_out_1_86 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_86 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_543_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_87 <= 2'h0;
    end else if (bht_bank_sel_1_5_7) begin
      if (_T_9652) begin
        bht_bank_rd_data_out_1_87 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_87 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_543_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_88 <= 2'h0;
    end else if (bht_bank_sel_1_5_8) begin
      if (_T_9661) begin
        bht_bank_rd_data_out_1_88 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_88 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_543_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_89 <= 2'h0;
    end else if (bht_bank_sel_1_5_9) begin
      if (_T_9670) begin
        bht_bank_rd_data_out_1_89 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_89 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_543_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_90 <= 2'h0;
    end else if (bht_bank_sel_1_5_10) begin
      if (_T_9679) begin
        bht_bank_rd_data_out_1_90 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_90 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_543_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_91 <= 2'h0;
    end else if (bht_bank_sel_1_5_11) begin
      if (_T_9688) begin
        bht_bank_rd_data_out_1_91 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_91 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_543_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_92 <= 2'h0;
    end else if (bht_bank_sel_1_5_12) begin
      if (_T_9697) begin
        bht_bank_rd_data_out_1_92 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_92 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_543_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_93 <= 2'h0;
    end else if (bht_bank_sel_1_5_13) begin
      if (_T_9706) begin
        bht_bank_rd_data_out_1_93 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_93 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_543_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_94 <= 2'h0;
    end else if (bht_bank_sel_1_5_14) begin
      if (_T_9715) begin
        bht_bank_rd_data_out_1_94 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_94 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_543_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_95 <= 2'h0;
    end else if (bht_bank_sel_1_5_15) begin
      if (_T_9724) begin
        bht_bank_rd_data_out_1_95 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_95 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_544_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_96 <= 2'h0;
    end else if (bht_bank_sel_1_6_0) begin
      if (_T_9733) begin
        bht_bank_rd_data_out_1_96 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_96 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_544_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_97 <= 2'h0;
    end else if (bht_bank_sel_1_6_1) begin
      if (_T_9742) begin
        bht_bank_rd_data_out_1_97 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_97 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_544_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_98 <= 2'h0;
    end else if (bht_bank_sel_1_6_2) begin
      if (_T_9751) begin
        bht_bank_rd_data_out_1_98 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_98 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_544_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_99 <= 2'h0;
    end else if (bht_bank_sel_1_6_3) begin
      if (_T_9760) begin
        bht_bank_rd_data_out_1_99 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_99 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_544_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_100 <= 2'h0;
    end else if (bht_bank_sel_1_6_4) begin
      if (_T_9769) begin
        bht_bank_rd_data_out_1_100 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_100 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_544_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_101 <= 2'h0;
    end else if (bht_bank_sel_1_6_5) begin
      if (_T_9778) begin
        bht_bank_rd_data_out_1_101 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_101 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_544_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_102 <= 2'h0;
    end else if (bht_bank_sel_1_6_6) begin
      if (_T_9787) begin
        bht_bank_rd_data_out_1_102 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_102 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_544_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_103 <= 2'h0;
    end else if (bht_bank_sel_1_6_7) begin
      if (_T_9796) begin
        bht_bank_rd_data_out_1_103 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_103 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_544_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_104 <= 2'h0;
    end else if (bht_bank_sel_1_6_8) begin
      if (_T_9805) begin
        bht_bank_rd_data_out_1_104 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_104 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_544_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_105 <= 2'h0;
    end else if (bht_bank_sel_1_6_9) begin
      if (_T_9814) begin
        bht_bank_rd_data_out_1_105 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_105 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_544_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_106 <= 2'h0;
    end else if (bht_bank_sel_1_6_10) begin
      if (_T_9823) begin
        bht_bank_rd_data_out_1_106 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_106 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_544_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_107 <= 2'h0;
    end else if (bht_bank_sel_1_6_11) begin
      if (_T_9832) begin
        bht_bank_rd_data_out_1_107 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_107 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_544_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_108 <= 2'h0;
    end else if (bht_bank_sel_1_6_12) begin
      if (_T_9841) begin
        bht_bank_rd_data_out_1_108 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_108 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_544_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_109 <= 2'h0;
    end else if (bht_bank_sel_1_6_13) begin
      if (_T_9850) begin
        bht_bank_rd_data_out_1_109 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_109 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_544_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_110 <= 2'h0;
    end else if (bht_bank_sel_1_6_14) begin
      if (_T_9859) begin
        bht_bank_rd_data_out_1_110 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_110 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_544_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_111 <= 2'h0;
    end else if (bht_bank_sel_1_6_15) begin
      if (_T_9868) begin
        bht_bank_rd_data_out_1_111 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_111 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_545_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_112 <= 2'h0;
    end else if (bht_bank_sel_1_7_0) begin
      if (_T_9877) begin
        bht_bank_rd_data_out_1_112 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_112 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_545_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_113 <= 2'h0;
    end else if (bht_bank_sel_1_7_1) begin
      if (_T_9886) begin
        bht_bank_rd_data_out_1_113 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_113 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_545_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_114 <= 2'h0;
    end else if (bht_bank_sel_1_7_2) begin
      if (_T_9895) begin
        bht_bank_rd_data_out_1_114 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_114 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_545_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_115 <= 2'h0;
    end else if (bht_bank_sel_1_7_3) begin
      if (_T_9904) begin
        bht_bank_rd_data_out_1_115 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_115 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_545_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_116 <= 2'h0;
    end else if (bht_bank_sel_1_7_4) begin
      if (_T_9913) begin
        bht_bank_rd_data_out_1_116 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_116 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_545_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_117 <= 2'h0;
    end else if (bht_bank_sel_1_7_5) begin
      if (_T_9922) begin
        bht_bank_rd_data_out_1_117 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_117 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_545_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_118 <= 2'h0;
    end else if (bht_bank_sel_1_7_6) begin
      if (_T_9931) begin
        bht_bank_rd_data_out_1_118 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_118 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_545_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_119 <= 2'h0;
    end else if (bht_bank_sel_1_7_7) begin
      if (_T_9940) begin
        bht_bank_rd_data_out_1_119 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_119 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_545_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_120 <= 2'h0;
    end else if (bht_bank_sel_1_7_8) begin
      if (_T_9949) begin
        bht_bank_rd_data_out_1_120 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_120 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_545_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_121 <= 2'h0;
    end else if (bht_bank_sel_1_7_9) begin
      if (_T_9958) begin
        bht_bank_rd_data_out_1_121 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_121 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_545_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_122 <= 2'h0;
    end else if (bht_bank_sel_1_7_10) begin
      if (_T_9967) begin
        bht_bank_rd_data_out_1_122 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_122 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_545_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_123 <= 2'h0;
    end else if (bht_bank_sel_1_7_11) begin
      if (_T_9976) begin
        bht_bank_rd_data_out_1_123 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_123 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_545_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_124 <= 2'h0;
    end else if (bht_bank_sel_1_7_12) begin
      if (_T_9985) begin
        bht_bank_rd_data_out_1_124 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_124 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_545_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_125 <= 2'h0;
    end else if (bht_bank_sel_1_7_13) begin
      if (_T_9994) begin
        bht_bank_rd_data_out_1_125 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_125 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_545_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_126 <= 2'h0;
    end else if (bht_bank_sel_1_7_14) begin
      if (_T_10003) begin
        bht_bank_rd_data_out_1_126 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_126 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_545_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_127 <= 2'h0;
    end else if (bht_bank_sel_1_7_15) begin
      if (_T_10012) begin
        bht_bank_rd_data_out_1_127 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_127 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_546_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_128 <= 2'h0;
    end else if (bht_bank_sel_1_8_0) begin
      if (_T_10021) begin
        bht_bank_rd_data_out_1_128 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_128 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_546_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_129 <= 2'h0;
    end else if (bht_bank_sel_1_8_1) begin
      if (_T_10030) begin
        bht_bank_rd_data_out_1_129 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_129 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_546_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_130 <= 2'h0;
    end else if (bht_bank_sel_1_8_2) begin
      if (_T_10039) begin
        bht_bank_rd_data_out_1_130 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_130 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_546_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_131 <= 2'h0;
    end else if (bht_bank_sel_1_8_3) begin
      if (_T_10048) begin
        bht_bank_rd_data_out_1_131 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_131 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_546_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_132 <= 2'h0;
    end else if (bht_bank_sel_1_8_4) begin
      if (_T_10057) begin
        bht_bank_rd_data_out_1_132 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_132 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_546_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_133 <= 2'h0;
    end else if (bht_bank_sel_1_8_5) begin
      if (_T_10066) begin
        bht_bank_rd_data_out_1_133 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_133 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_546_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_134 <= 2'h0;
    end else if (bht_bank_sel_1_8_6) begin
      if (_T_10075) begin
        bht_bank_rd_data_out_1_134 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_134 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_546_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_135 <= 2'h0;
    end else if (bht_bank_sel_1_8_7) begin
      if (_T_10084) begin
        bht_bank_rd_data_out_1_135 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_135 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_546_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_136 <= 2'h0;
    end else if (bht_bank_sel_1_8_8) begin
      if (_T_10093) begin
        bht_bank_rd_data_out_1_136 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_136 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_546_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_137 <= 2'h0;
    end else if (bht_bank_sel_1_8_9) begin
      if (_T_10102) begin
        bht_bank_rd_data_out_1_137 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_137 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_546_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_138 <= 2'h0;
    end else if (bht_bank_sel_1_8_10) begin
      if (_T_10111) begin
        bht_bank_rd_data_out_1_138 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_138 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_546_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_139 <= 2'h0;
    end else if (bht_bank_sel_1_8_11) begin
      if (_T_10120) begin
        bht_bank_rd_data_out_1_139 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_139 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_546_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_140 <= 2'h0;
    end else if (bht_bank_sel_1_8_12) begin
      if (_T_10129) begin
        bht_bank_rd_data_out_1_140 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_140 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_546_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_141 <= 2'h0;
    end else if (bht_bank_sel_1_8_13) begin
      if (_T_10138) begin
        bht_bank_rd_data_out_1_141 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_141 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_546_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_142 <= 2'h0;
    end else if (bht_bank_sel_1_8_14) begin
      if (_T_10147) begin
        bht_bank_rd_data_out_1_142 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_142 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_546_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_143 <= 2'h0;
    end else if (bht_bank_sel_1_8_15) begin
      if (_T_10156) begin
        bht_bank_rd_data_out_1_143 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_143 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_547_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_144 <= 2'h0;
    end else if (bht_bank_sel_1_9_0) begin
      if (_T_10165) begin
        bht_bank_rd_data_out_1_144 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_144 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_547_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_145 <= 2'h0;
    end else if (bht_bank_sel_1_9_1) begin
      if (_T_10174) begin
        bht_bank_rd_data_out_1_145 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_145 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_547_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_146 <= 2'h0;
    end else if (bht_bank_sel_1_9_2) begin
      if (_T_10183) begin
        bht_bank_rd_data_out_1_146 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_146 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_547_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_147 <= 2'h0;
    end else if (bht_bank_sel_1_9_3) begin
      if (_T_10192) begin
        bht_bank_rd_data_out_1_147 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_147 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_547_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_148 <= 2'h0;
    end else if (bht_bank_sel_1_9_4) begin
      if (_T_10201) begin
        bht_bank_rd_data_out_1_148 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_148 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_547_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_149 <= 2'h0;
    end else if (bht_bank_sel_1_9_5) begin
      if (_T_10210) begin
        bht_bank_rd_data_out_1_149 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_149 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_547_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_150 <= 2'h0;
    end else if (bht_bank_sel_1_9_6) begin
      if (_T_10219) begin
        bht_bank_rd_data_out_1_150 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_150 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_547_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_151 <= 2'h0;
    end else if (bht_bank_sel_1_9_7) begin
      if (_T_10228) begin
        bht_bank_rd_data_out_1_151 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_151 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_547_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_152 <= 2'h0;
    end else if (bht_bank_sel_1_9_8) begin
      if (_T_10237) begin
        bht_bank_rd_data_out_1_152 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_152 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_547_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_153 <= 2'h0;
    end else if (bht_bank_sel_1_9_9) begin
      if (_T_10246) begin
        bht_bank_rd_data_out_1_153 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_153 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_547_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_154 <= 2'h0;
    end else if (bht_bank_sel_1_9_10) begin
      if (_T_10255) begin
        bht_bank_rd_data_out_1_154 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_154 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_547_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_155 <= 2'h0;
    end else if (bht_bank_sel_1_9_11) begin
      if (_T_10264) begin
        bht_bank_rd_data_out_1_155 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_155 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_547_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_156 <= 2'h0;
    end else if (bht_bank_sel_1_9_12) begin
      if (_T_10273) begin
        bht_bank_rd_data_out_1_156 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_156 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_547_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_157 <= 2'h0;
    end else if (bht_bank_sel_1_9_13) begin
      if (_T_10282) begin
        bht_bank_rd_data_out_1_157 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_157 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_547_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_158 <= 2'h0;
    end else if (bht_bank_sel_1_9_14) begin
      if (_T_10291) begin
        bht_bank_rd_data_out_1_158 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_158 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_547_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_159 <= 2'h0;
    end else if (bht_bank_sel_1_9_15) begin
      if (_T_10300) begin
        bht_bank_rd_data_out_1_159 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_159 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_548_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_160 <= 2'h0;
    end else if (bht_bank_sel_1_10_0) begin
      if (_T_10309) begin
        bht_bank_rd_data_out_1_160 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_160 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_548_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_161 <= 2'h0;
    end else if (bht_bank_sel_1_10_1) begin
      if (_T_10318) begin
        bht_bank_rd_data_out_1_161 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_161 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_548_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_162 <= 2'h0;
    end else if (bht_bank_sel_1_10_2) begin
      if (_T_10327) begin
        bht_bank_rd_data_out_1_162 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_162 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_548_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_163 <= 2'h0;
    end else if (bht_bank_sel_1_10_3) begin
      if (_T_10336) begin
        bht_bank_rd_data_out_1_163 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_163 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_548_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_164 <= 2'h0;
    end else if (bht_bank_sel_1_10_4) begin
      if (_T_10345) begin
        bht_bank_rd_data_out_1_164 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_164 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_548_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_165 <= 2'h0;
    end else if (bht_bank_sel_1_10_5) begin
      if (_T_10354) begin
        bht_bank_rd_data_out_1_165 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_165 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_548_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_166 <= 2'h0;
    end else if (bht_bank_sel_1_10_6) begin
      if (_T_10363) begin
        bht_bank_rd_data_out_1_166 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_166 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_548_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_167 <= 2'h0;
    end else if (bht_bank_sel_1_10_7) begin
      if (_T_10372) begin
        bht_bank_rd_data_out_1_167 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_167 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_548_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_168 <= 2'h0;
    end else if (bht_bank_sel_1_10_8) begin
      if (_T_10381) begin
        bht_bank_rd_data_out_1_168 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_168 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_548_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_169 <= 2'h0;
    end else if (bht_bank_sel_1_10_9) begin
      if (_T_10390) begin
        bht_bank_rd_data_out_1_169 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_169 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_548_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_170 <= 2'h0;
    end else if (bht_bank_sel_1_10_10) begin
      if (_T_10399) begin
        bht_bank_rd_data_out_1_170 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_170 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_548_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_171 <= 2'h0;
    end else if (bht_bank_sel_1_10_11) begin
      if (_T_10408) begin
        bht_bank_rd_data_out_1_171 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_171 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_548_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_172 <= 2'h0;
    end else if (bht_bank_sel_1_10_12) begin
      if (_T_10417) begin
        bht_bank_rd_data_out_1_172 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_172 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_548_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_173 <= 2'h0;
    end else if (bht_bank_sel_1_10_13) begin
      if (_T_10426) begin
        bht_bank_rd_data_out_1_173 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_173 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_548_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_174 <= 2'h0;
    end else if (bht_bank_sel_1_10_14) begin
      if (_T_10435) begin
        bht_bank_rd_data_out_1_174 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_174 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_548_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_175 <= 2'h0;
    end else if (bht_bank_sel_1_10_15) begin
      if (_T_10444) begin
        bht_bank_rd_data_out_1_175 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_175 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_549_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_176 <= 2'h0;
    end else if (bht_bank_sel_1_11_0) begin
      if (_T_10453) begin
        bht_bank_rd_data_out_1_176 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_176 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_549_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_177 <= 2'h0;
    end else if (bht_bank_sel_1_11_1) begin
      if (_T_10462) begin
        bht_bank_rd_data_out_1_177 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_177 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_549_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_178 <= 2'h0;
    end else if (bht_bank_sel_1_11_2) begin
      if (_T_10471) begin
        bht_bank_rd_data_out_1_178 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_178 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_549_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_179 <= 2'h0;
    end else if (bht_bank_sel_1_11_3) begin
      if (_T_10480) begin
        bht_bank_rd_data_out_1_179 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_179 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_549_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_180 <= 2'h0;
    end else if (bht_bank_sel_1_11_4) begin
      if (_T_10489) begin
        bht_bank_rd_data_out_1_180 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_180 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_549_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_181 <= 2'h0;
    end else if (bht_bank_sel_1_11_5) begin
      if (_T_10498) begin
        bht_bank_rd_data_out_1_181 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_181 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_549_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_182 <= 2'h0;
    end else if (bht_bank_sel_1_11_6) begin
      if (_T_10507) begin
        bht_bank_rd_data_out_1_182 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_182 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_549_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_183 <= 2'h0;
    end else if (bht_bank_sel_1_11_7) begin
      if (_T_10516) begin
        bht_bank_rd_data_out_1_183 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_183 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_549_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_184 <= 2'h0;
    end else if (bht_bank_sel_1_11_8) begin
      if (_T_10525) begin
        bht_bank_rd_data_out_1_184 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_184 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_549_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_185 <= 2'h0;
    end else if (bht_bank_sel_1_11_9) begin
      if (_T_10534) begin
        bht_bank_rd_data_out_1_185 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_185 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_549_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_186 <= 2'h0;
    end else if (bht_bank_sel_1_11_10) begin
      if (_T_10543) begin
        bht_bank_rd_data_out_1_186 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_186 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_549_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_187 <= 2'h0;
    end else if (bht_bank_sel_1_11_11) begin
      if (_T_10552) begin
        bht_bank_rd_data_out_1_187 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_187 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_549_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_188 <= 2'h0;
    end else if (bht_bank_sel_1_11_12) begin
      if (_T_10561) begin
        bht_bank_rd_data_out_1_188 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_188 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_549_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_189 <= 2'h0;
    end else if (bht_bank_sel_1_11_13) begin
      if (_T_10570) begin
        bht_bank_rd_data_out_1_189 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_189 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_549_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_190 <= 2'h0;
    end else if (bht_bank_sel_1_11_14) begin
      if (_T_10579) begin
        bht_bank_rd_data_out_1_190 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_190 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_549_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_191 <= 2'h0;
    end else if (bht_bank_sel_1_11_15) begin
      if (_T_10588) begin
        bht_bank_rd_data_out_1_191 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_191 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_550_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_192 <= 2'h0;
    end else if (bht_bank_sel_1_12_0) begin
      if (_T_10597) begin
        bht_bank_rd_data_out_1_192 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_192 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_550_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_193 <= 2'h0;
    end else if (bht_bank_sel_1_12_1) begin
      if (_T_10606) begin
        bht_bank_rd_data_out_1_193 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_193 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_550_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_194 <= 2'h0;
    end else if (bht_bank_sel_1_12_2) begin
      if (_T_10615) begin
        bht_bank_rd_data_out_1_194 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_194 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_550_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_195 <= 2'h0;
    end else if (bht_bank_sel_1_12_3) begin
      if (_T_10624) begin
        bht_bank_rd_data_out_1_195 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_195 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_550_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_196 <= 2'h0;
    end else if (bht_bank_sel_1_12_4) begin
      if (_T_10633) begin
        bht_bank_rd_data_out_1_196 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_196 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_550_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_197 <= 2'h0;
    end else if (bht_bank_sel_1_12_5) begin
      if (_T_10642) begin
        bht_bank_rd_data_out_1_197 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_197 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_550_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_198 <= 2'h0;
    end else if (bht_bank_sel_1_12_6) begin
      if (_T_10651) begin
        bht_bank_rd_data_out_1_198 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_198 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_550_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_199 <= 2'h0;
    end else if (bht_bank_sel_1_12_7) begin
      if (_T_10660) begin
        bht_bank_rd_data_out_1_199 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_199 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_550_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_200 <= 2'h0;
    end else if (bht_bank_sel_1_12_8) begin
      if (_T_10669) begin
        bht_bank_rd_data_out_1_200 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_200 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_550_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_201 <= 2'h0;
    end else if (bht_bank_sel_1_12_9) begin
      if (_T_10678) begin
        bht_bank_rd_data_out_1_201 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_201 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_550_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_202 <= 2'h0;
    end else if (bht_bank_sel_1_12_10) begin
      if (_T_10687) begin
        bht_bank_rd_data_out_1_202 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_202 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_550_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_203 <= 2'h0;
    end else if (bht_bank_sel_1_12_11) begin
      if (_T_10696) begin
        bht_bank_rd_data_out_1_203 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_203 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_550_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_204 <= 2'h0;
    end else if (bht_bank_sel_1_12_12) begin
      if (_T_10705) begin
        bht_bank_rd_data_out_1_204 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_204 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_550_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_205 <= 2'h0;
    end else if (bht_bank_sel_1_12_13) begin
      if (_T_10714) begin
        bht_bank_rd_data_out_1_205 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_205 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_550_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_206 <= 2'h0;
    end else if (bht_bank_sel_1_12_14) begin
      if (_T_10723) begin
        bht_bank_rd_data_out_1_206 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_206 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_550_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_207 <= 2'h0;
    end else if (bht_bank_sel_1_12_15) begin
      if (_T_10732) begin
        bht_bank_rd_data_out_1_207 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_207 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_551_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_208 <= 2'h0;
    end else if (bht_bank_sel_1_13_0) begin
      if (_T_10741) begin
        bht_bank_rd_data_out_1_208 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_208 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_551_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_209 <= 2'h0;
    end else if (bht_bank_sel_1_13_1) begin
      if (_T_10750) begin
        bht_bank_rd_data_out_1_209 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_209 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_551_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_210 <= 2'h0;
    end else if (bht_bank_sel_1_13_2) begin
      if (_T_10759) begin
        bht_bank_rd_data_out_1_210 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_210 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_551_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_211 <= 2'h0;
    end else if (bht_bank_sel_1_13_3) begin
      if (_T_10768) begin
        bht_bank_rd_data_out_1_211 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_211 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_551_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_212 <= 2'h0;
    end else if (bht_bank_sel_1_13_4) begin
      if (_T_10777) begin
        bht_bank_rd_data_out_1_212 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_212 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_551_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_213 <= 2'h0;
    end else if (bht_bank_sel_1_13_5) begin
      if (_T_10786) begin
        bht_bank_rd_data_out_1_213 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_213 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_551_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_214 <= 2'h0;
    end else if (bht_bank_sel_1_13_6) begin
      if (_T_10795) begin
        bht_bank_rd_data_out_1_214 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_214 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_551_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_215 <= 2'h0;
    end else if (bht_bank_sel_1_13_7) begin
      if (_T_10804) begin
        bht_bank_rd_data_out_1_215 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_215 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_551_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_216 <= 2'h0;
    end else if (bht_bank_sel_1_13_8) begin
      if (_T_10813) begin
        bht_bank_rd_data_out_1_216 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_216 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_551_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_217 <= 2'h0;
    end else if (bht_bank_sel_1_13_9) begin
      if (_T_10822) begin
        bht_bank_rd_data_out_1_217 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_217 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_551_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_218 <= 2'h0;
    end else if (bht_bank_sel_1_13_10) begin
      if (_T_10831) begin
        bht_bank_rd_data_out_1_218 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_218 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_551_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_219 <= 2'h0;
    end else if (bht_bank_sel_1_13_11) begin
      if (_T_10840) begin
        bht_bank_rd_data_out_1_219 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_219 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_551_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_220 <= 2'h0;
    end else if (bht_bank_sel_1_13_12) begin
      if (_T_10849) begin
        bht_bank_rd_data_out_1_220 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_220 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_551_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_221 <= 2'h0;
    end else if (bht_bank_sel_1_13_13) begin
      if (_T_10858) begin
        bht_bank_rd_data_out_1_221 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_221 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_551_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_222 <= 2'h0;
    end else if (bht_bank_sel_1_13_14) begin
      if (_T_10867) begin
        bht_bank_rd_data_out_1_222 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_222 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_551_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_223 <= 2'h0;
    end else if (bht_bank_sel_1_13_15) begin
      if (_T_10876) begin
        bht_bank_rd_data_out_1_223 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_223 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_552_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_224 <= 2'h0;
    end else if (bht_bank_sel_1_14_0) begin
      if (_T_10885) begin
        bht_bank_rd_data_out_1_224 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_224 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_552_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_225 <= 2'h0;
    end else if (bht_bank_sel_1_14_1) begin
      if (_T_10894) begin
        bht_bank_rd_data_out_1_225 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_225 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_552_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_226 <= 2'h0;
    end else if (bht_bank_sel_1_14_2) begin
      if (_T_10903) begin
        bht_bank_rd_data_out_1_226 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_226 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_552_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_227 <= 2'h0;
    end else if (bht_bank_sel_1_14_3) begin
      if (_T_10912) begin
        bht_bank_rd_data_out_1_227 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_227 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_552_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_228 <= 2'h0;
    end else if (bht_bank_sel_1_14_4) begin
      if (_T_10921) begin
        bht_bank_rd_data_out_1_228 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_228 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_552_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_229 <= 2'h0;
    end else if (bht_bank_sel_1_14_5) begin
      if (_T_10930) begin
        bht_bank_rd_data_out_1_229 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_229 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_552_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_230 <= 2'h0;
    end else if (bht_bank_sel_1_14_6) begin
      if (_T_10939) begin
        bht_bank_rd_data_out_1_230 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_230 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_552_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_231 <= 2'h0;
    end else if (bht_bank_sel_1_14_7) begin
      if (_T_10948) begin
        bht_bank_rd_data_out_1_231 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_231 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_552_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_232 <= 2'h0;
    end else if (bht_bank_sel_1_14_8) begin
      if (_T_10957) begin
        bht_bank_rd_data_out_1_232 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_232 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_552_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_233 <= 2'h0;
    end else if (bht_bank_sel_1_14_9) begin
      if (_T_10966) begin
        bht_bank_rd_data_out_1_233 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_233 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_552_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_234 <= 2'h0;
    end else if (bht_bank_sel_1_14_10) begin
      if (_T_10975) begin
        bht_bank_rd_data_out_1_234 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_234 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_552_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_235 <= 2'h0;
    end else if (bht_bank_sel_1_14_11) begin
      if (_T_10984) begin
        bht_bank_rd_data_out_1_235 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_235 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_552_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_236 <= 2'h0;
    end else if (bht_bank_sel_1_14_12) begin
      if (_T_10993) begin
        bht_bank_rd_data_out_1_236 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_236 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_552_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_237 <= 2'h0;
    end else if (bht_bank_sel_1_14_13) begin
      if (_T_11002) begin
        bht_bank_rd_data_out_1_237 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_237 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_552_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_238 <= 2'h0;
    end else if (bht_bank_sel_1_14_14) begin
      if (_T_11011) begin
        bht_bank_rd_data_out_1_238 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_238 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_552_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_239 <= 2'h0;
    end else if (bht_bank_sel_1_14_15) begin
      if (_T_11020) begin
        bht_bank_rd_data_out_1_239 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_239 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_553_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_240 <= 2'h0;
    end else if (bht_bank_sel_1_15_0) begin
      if (_T_11029) begin
        bht_bank_rd_data_out_1_240 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_240 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_553_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_241 <= 2'h0;
    end else if (bht_bank_sel_1_15_1) begin
      if (_T_11038) begin
        bht_bank_rd_data_out_1_241 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_241 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_553_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_242 <= 2'h0;
    end else if (bht_bank_sel_1_15_2) begin
      if (_T_11047) begin
        bht_bank_rd_data_out_1_242 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_242 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_553_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_243 <= 2'h0;
    end else if (bht_bank_sel_1_15_3) begin
      if (_T_11056) begin
        bht_bank_rd_data_out_1_243 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_243 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_553_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_244 <= 2'h0;
    end else if (bht_bank_sel_1_15_4) begin
      if (_T_11065) begin
        bht_bank_rd_data_out_1_244 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_244 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_553_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_245 <= 2'h0;
    end else if (bht_bank_sel_1_15_5) begin
      if (_T_11074) begin
        bht_bank_rd_data_out_1_245 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_245 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_553_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_246 <= 2'h0;
    end else if (bht_bank_sel_1_15_6) begin
      if (_T_11083) begin
        bht_bank_rd_data_out_1_246 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_246 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_553_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_247 <= 2'h0;
    end else if (bht_bank_sel_1_15_7) begin
      if (_T_11092) begin
        bht_bank_rd_data_out_1_247 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_247 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_553_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_248 <= 2'h0;
    end else if (bht_bank_sel_1_15_8) begin
      if (_T_11101) begin
        bht_bank_rd_data_out_1_248 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_248 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_553_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_249 <= 2'h0;
    end else if (bht_bank_sel_1_15_9) begin
      if (_T_11110) begin
        bht_bank_rd_data_out_1_249 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_249 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_553_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_250 <= 2'h0;
    end else if (bht_bank_sel_1_15_10) begin
      if (_T_11119) begin
        bht_bank_rd_data_out_1_250 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_250 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_553_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_251 <= 2'h0;
    end else if (bht_bank_sel_1_15_11) begin
      if (_T_11128) begin
        bht_bank_rd_data_out_1_251 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_251 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_553_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_252 <= 2'h0;
    end else if (bht_bank_sel_1_15_12) begin
      if (_T_11137) begin
        bht_bank_rd_data_out_1_252 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_252 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_553_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_253 <= 2'h0;
    end else if (bht_bank_sel_1_15_13) begin
      if (_T_11146) begin
        bht_bank_rd_data_out_1_253 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_253 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_553_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_254 <= 2'h0;
    end else if (bht_bank_sel_1_15_14) begin
      if (_T_11155) begin
        bht_bank_rd_data_out_1_254 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_254 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_553_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_255 <= 2'h0;
    end else if (bht_bank_sel_1_15_15) begin
      if (_T_11164) begin
        bht_bank_rd_data_out_1_255 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_255 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_522_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_0 <= 2'h0;
    end else if (bht_bank_sel_0_0_0) begin
      if (_T_6565) begin
        bht_bank_rd_data_out_0_0 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_0 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_522_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_1 <= 2'h0;
    end else if (bht_bank_sel_0_0_1) begin
      if (_T_6574) begin
        bht_bank_rd_data_out_0_1 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_1 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_522_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_2 <= 2'h0;
    end else if (bht_bank_sel_0_0_2) begin
      if (_T_6583) begin
        bht_bank_rd_data_out_0_2 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_2 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_522_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_3 <= 2'h0;
    end else if (bht_bank_sel_0_0_3) begin
      if (_T_6592) begin
        bht_bank_rd_data_out_0_3 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_3 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_522_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_4 <= 2'h0;
    end else if (bht_bank_sel_0_0_4) begin
      if (_T_6601) begin
        bht_bank_rd_data_out_0_4 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_4 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_522_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_5 <= 2'h0;
    end else if (bht_bank_sel_0_0_5) begin
      if (_T_6610) begin
        bht_bank_rd_data_out_0_5 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_5 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_522_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_6 <= 2'h0;
    end else if (bht_bank_sel_0_0_6) begin
      if (_T_6619) begin
        bht_bank_rd_data_out_0_6 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_6 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_522_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_7 <= 2'h0;
    end else if (bht_bank_sel_0_0_7) begin
      if (_T_6628) begin
        bht_bank_rd_data_out_0_7 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_7 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_522_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_8 <= 2'h0;
    end else if (bht_bank_sel_0_0_8) begin
      if (_T_6637) begin
        bht_bank_rd_data_out_0_8 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_8 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_522_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_9 <= 2'h0;
    end else if (bht_bank_sel_0_0_9) begin
      if (_T_6646) begin
        bht_bank_rd_data_out_0_9 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_9 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_522_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_10 <= 2'h0;
    end else if (bht_bank_sel_0_0_10) begin
      if (_T_6655) begin
        bht_bank_rd_data_out_0_10 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_10 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_522_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_11 <= 2'h0;
    end else if (bht_bank_sel_0_0_11) begin
      if (_T_6664) begin
        bht_bank_rd_data_out_0_11 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_11 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_522_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_12 <= 2'h0;
    end else if (bht_bank_sel_0_0_12) begin
      if (_T_6673) begin
        bht_bank_rd_data_out_0_12 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_12 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_522_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_13 <= 2'h0;
    end else if (bht_bank_sel_0_0_13) begin
      if (_T_6682) begin
        bht_bank_rd_data_out_0_13 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_13 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_522_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_14 <= 2'h0;
    end else if (bht_bank_sel_0_0_14) begin
      if (_T_6691) begin
        bht_bank_rd_data_out_0_14 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_14 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_522_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_15 <= 2'h0;
    end else if (bht_bank_sel_0_0_15) begin
      if (_T_6700) begin
        bht_bank_rd_data_out_0_15 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_15 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_523_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_16 <= 2'h0;
    end else if (bht_bank_sel_0_1_0) begin
      if (_T_6709) begin
        bht_bank_rd_data_out_0_16 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_16 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_523_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_17 <= 2'h0;
    end else if (bht_bank_sel_0_1_1) begin
      if (_T_6718) begin
        bht_bank_rd_data_out_0_17 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_17 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_523_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_18 <= 2'h0;
    end else if (bht_bank_sel_0_1_2) begin
      if (_T_6727) begin
        bht_bank_rd_data_out_0_18 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_18 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_523_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_19 <= 2'h0;
    end else if (bht_bank_sel_0_1_3) begin
      if (_T_6736) begin
        bht_bank_rd_data_out_0_19 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_19 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_523_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_20 <= 2'h0;
    end else if (bht_bank_sel_0_1_4) begin
      if (_T_6745) begin
        bht_bank_rd_data_out_0_20 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_20 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_523_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_21 <= 2'h0;
    end else if (bht_bank_sel_0_1_5) begin
      if (_T_6754) begin
        bht_bank_rd_data_out_0_21 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_21 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_523_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_22 <= 2'h0;
    end else if (bht_bank_sel_0_1_6) begin
      if (_T_6763) begin
        bht_bank_rd_data_out_0_22 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_22 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_523_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_23 <= 2'h0;
    end else if (bht_bank_sel_0_1_7) begin
      if (_T_6772) begin
        bht_bank_rd_data_out_0_23 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_23 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_523_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_24 <= 2'h0;
    end else if (bht_bank_sel_0_1_8) begin
      if (_T_6781) begin
        bht_bank_rd_data_out_0_24 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_24 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_523_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_25 <= 2'h0;
    end else if (bht_bank_sel_0_1_9) begin
      if (_T_6790) begin
        bht_bank_rd_data_out_0_25 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_25 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_523_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_26 <= 2'h0;
    end else if (bht_bank_sel_0_1_10) begin
      if (_T_6799) begin
        bht_bank_rd_data_out_0_26 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_26 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_523_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_27 <= 2'h0;
    end else if (bht_bank_sel_0_1_11) begin
      if (_T_6808) begin
        bht_bank_rd_data_out_0_27 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_27 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_523_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_28 <= 2'h0;
    end else if (bht_bank_sel_0_1_12) begin
      if (_T_6817) begin
        bht_bank_rd_data_out_0_28 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_28 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_523_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_29 <= 2'h0;
    end else if (bht_bank_sel_0_1_13) begin
      if (_T_6826) begin
        bht_bank_rd_data_out_0_29 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_29 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_523_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_30 <= 2'h0;
    end else if (bht_bank_sel_0_1_14) begin
      if (_T_6835) begin
        bht_bank_rd_data_out_0_30 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_30 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_523_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_31 <= 2'h0;
    end else if (bht_bank_sel_0_1_15) begin
      if (_T_6844) begin
        bht_bank_rd_data_out_0_31 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_31 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_524_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_32 <= 2'h0;
    end else if (bht_bank_sel_0_2_0) begin
      if (_T_6853) begin
        bht_bank_rd_data_out_0_32 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_32 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_524_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_33 <= 2'h0;
    end else if (bht_bank_sel_0_2_1) begin
      if (_T_6862) begin
        bht_bank_rd_data_out_0_33 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_33 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_524_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_34 <= 2'h0;
    end else if (bht_bank_sel_0_2_2) begin
      if (_T_6871) begin
        bht_bank_rd_data_out_0_34 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_34 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_524_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_35 <= 2'h0;
    end else if (bht_bank_sel_0_2_3) begin
      if (_T_6880) begin
        bht_bank_rd_data_out_0_35 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_35 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_524_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_36 <= 2'h0;
    end else if (bht_bank_sel_0_2_4) begin
      if (_T_6889) begin
        bht_bank_rd_data_out_0_36 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_36 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_524_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_37 <= 2'h0;
    end else if (bht_bank_sel_0_2_5) begin
      if (_T_6898) begin
        bht_bank_rd_data_out_0_37 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_37 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_524_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_38 <= 2'h0;
    end else if (bht_bank_sel_0_2_6) begin
      if (_T_6907) begin
        bht_bank_rd_data_out_0_38 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_38 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_524_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_39 <= 2'h0;
    end else if (bht_bank_sel_0_2_7) begin
      if (_T_6916) begin
        bht_bank_rd_data_out_0_39 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_39 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_524_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_40 <= 2'h0;
    end else if (bht_bank_sel_0_2_8) begin
      if (_T_6925) begin
        bht_bank_rd_data_out_0_40 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_40 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_524_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_41 <= 2'h0;
    end else if (bht_bank_sel_0_2_9) begin
      if (_T_6934) begin
        bht_bank_rd_data_out_0_41 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_41 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_524_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_42 <= 2'h0;
    end else if (bht_bank_sel_0_2_10) begin
      if (_T_6943) begin
        bht_bank_rd_data_out_0_42 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_42 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_524_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_43 <= 2'h0;
    end else if (bht_bank_sel_0_2_11) begin
      if (_T_6952) begin
        bht_bank_rd_data_out_0_43 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_43 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_524_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_44 <= 2'h0;
    end else if (bht_bank_sel_0_2_12) begin
      if (_T_6961) begin
        bht_bank_rd_data_out_0_44 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_44 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_524_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_45 <= 2'h0;
    end else if (bht_bank_sel_0_2_13) begin
      if (_T_6970) begin
        bht_bank_rd_data_out_0_45 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_45 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_524_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_46 <= 2'h0;
    end else if (bht_bank_sel_0_2_14) begin
      if (_T_6979) begin
        bht_bank_rd_data_out_0_46 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_46 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_524_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_47 <= 2'h0;
    end else if (bht_bank_sel_0_2_15) begin
      if (_T_6988) begin
        bht_bank_rd_data_out_0_47 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_47 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_525_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_48 <= 2'h0;
    end else if (bht_bank_sel_0_3_0) begin
      if (_T_6997) begin
        bht_bank_rd_data_out_0_48 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_48 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_525_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_49 <= 2'h0;
    end else if (bht_bank_sel_0_3_1) begin
      if (_T_7006) begin
        bht_bank_rd_data_out_0_49 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_49 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_525_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_50 <= 2'h0;
    end else if (bht_bank_sel_0_3_2) begin
      if (_T_7015) begin
        bht_bank_rd_data_out_0_50 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_50 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_525_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_51 <= 2'h0;
    end else if (bht_bank_sel_0_3_3) begin
      if (_T_7024) begin
        bht_bank_rd_data_out_0_51 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_51 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_525_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_52 <= 2'h0;
    end else if (bht_bank_sel_0_3_4) begin
      if (_T_7033) begin
        bht_bank_rd_data_out_0_52 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_52 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_525_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_53 <= 2'h0;
    end else if (bht_bank_sel_0_3_5) begin
      if (_T_7042) begin
        bht_bank_rd_data_out_0_53 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_53 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_525_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_54 <= 2'h0;
    end else if (bht_bank_sel_0_3_6) begin
      if (_T_7051) begin
        bht_bank_rd_data_out_0_54 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_54 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_525_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_55 <= 2'h0;
    end else if (bht_bank_sel_0_3_7) begin
      if (_T_7060) begin
        bht_bank_rd_data_out_0_55 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_55 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_525_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_56 <= 2'h0;
    end else if (bht_bank_sel_0_3_8) begin
      if (_T_7069) begin
        bht_bank_rd_data_out_0_56 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_56 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_525_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_57 <= 2'h0;
    end else if (bht_bank_sel_0_3_9) begin
      if (_T_7078) begin
        bht_bank_rd_data_out_0_57 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_57 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_525_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_58 <= 2'h0;
    end else if (bht_bank_sel_0_3_10) begin
      if (_T_7087) begin
        bht_bank_rd_data_out_0_58 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_58 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_525_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_59 <= 2'h0;
    end else if (bht_bank_sel_0_3_11) begin
      if (_T_7096) begin
        bht_bank_rd_data_out_0_59 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_59 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_525_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_60 <= 2'h0;
    end else if (bht_bank_sel_0_3_12) begin
      if (_T_7105) begin
        bht_bank_rd_data_out_0_60 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_60 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_525_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_61 <= 2'h0;
    end else if (bht_bank_sel_0_3_13) begin
      if (_T_7114) begin
        bht_bank_rd_data_out_0_61 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_61 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_525_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_62 <= 2'h0;
    end else if (bht_bank_sel_0_3_14) begin
      if (_T_7123) begin
        bht_bank_rd_data_out_0_62 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_62 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_525_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_63 <= 2'h0;
    end else if (bht_bank_sel_0_3_15) begin
      if (_T_7132) begin
        bht_bank_rd_data_out_0_63 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_63 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_526_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_64 <= 2'h0;
    end else if (bht_bank_sel_0_4_0) begin
      if (_T_7141) begin
        bht_bank_rd_data_out_0_64 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_64 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_526_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_65 <= 2'h0;
    end else if (bht_bank_sel_0_4_1) begin
      if (_T_7150) begin
        bht_bank_rd_data_out_0_65 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_65 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_526_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_66 <= 2'h0;
    end else if (bht_bank_sel_0_4_2) begin
      if (_T_7159) begin
        bht_bank_rd_data_out_0_66 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_66 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_526_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_67 <= 2'h0;
    end else if (bht_bank_sel_0_4_3) begin
      if (_T_7168) begin
        bht_bank_rd_data_out_0_67 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_67 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_526_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_68 <= 2'h0;
    end else if (bht_bank_sel_0_4_4) begin
      if (_T_7177) begin
        bht_bank_rd_data_out_0_68 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_68 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_526_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_69 <= 2'h0;
    end else if (bht_bank_sel_0_4_5) begin
      if (_T_7186) begin
        bht_bank_rd_data_out_0_69 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_69 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_526_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_70 <= 2'h0;
    end else if (bht_bank_sel_0_4_6) begin
      if (_T_7195) begin
        bht_bank_rd_data_out_0_70 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_70 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_526_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_71 <= 2'h0;
    end else if (bht_bank_sel_0_4_7) begin
      if (_T_7204) begin
        bht_bank_rd_data_out_0_71 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_71 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_526_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_72 <= 2'h0;
    end else if (bht_bank_sel_0_4_8) begin
      if (_T_7213) begin
        bht_bank_rd_data_out_0_72 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_72 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_526_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_73 <= 2'h0;
    end else if (bht_bank_sel_0_4_9) begin
      if (_T_7222) begin
        bht_bank_rd_data_out_0_73 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_73 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_526_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_74 <= 2'h0;
    end else if (bht_bank_sel_0_4_10) begin
      if (_T_7231) begin
        bht_bank_rd_data_out_0_74 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_74 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_526_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_75 <= 2'h0;
    end else if (bht_bank_sel_0_4_11) begin
      if (_T_7240) begin
        bht_bank_rd_data_out_0_75 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_75 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_526_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_76 <= 2'h0;
    end else if (bht_bank_sel_0_4_12) begin
      if (_T_7249) begin
        bht_bank_rd_data_out_0_76 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_76 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_526_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_77 <= 2'h0;
    end else if (bht_bank_sel_0_4_13) begin
      if (_T_7258) begin
        bht_bank_rd_data_out_0_77 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_77 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_526_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_78 <= 2'h0;
    end else if (bht_bank_sel_0_4_14) begin
      if (_T_7267) begin
        bht_bank_rd_data_out_0_78 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_78 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_526_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_79 <= 2'h0;
    end else if (bht_bank_sel_0_4_15) begin
      if (_T_7276) begin
        bht_bank_rd_data_out_0_79 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_79 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_527_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_80 <= 2'h0;
    end else if (bht_bank_sel_0_5_0) begin
      if (_T_7285) begin
        bht_bank_rd_data_out_0_80 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_80 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_527_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_81 <= 2'h0;
    end else if (bht_bank_sel_0_5_1) begin
      if (_T_7294) begin
        bht_bank_rd_data_out_0_81 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_81 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_527_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_82 <= 2'h0;
    end else if (bht_bank_sel_0_5_2) begin
      if (_T_7303) begin
        bht_bank_rd_data_out_0_82 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_82 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_527_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_83 <= 2'h0;
    end else if (bht_bank_sel_0_5_3) begin
      if (_T_7312) begin
        bht_bank_rd_data_out_0_83 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_83 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_527_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_84 <= 2'h0;
    end else if (bht_bank_sel_0_5_4) begin
      if (_T_7321) begin
        bht_bank_rd_data_out_0_84 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_84 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_527_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_85 <= 2'h0;
    end else if (bht_bank_sel_0_5_5) begin
      if (_T_7330) begin
        bht_bank_rd_data_out_0_85 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_85 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_527_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_86 <= 2'h0;
    end else if (bht_bank_sel_0_5_6) begin
      if (_T_7339) begin
        bht_bank_rd_data_out_0_86 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_86 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_527_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_87 <= 2'h0;
    end else if (bht_bank_sel_0_5_7) begin
      if (_T_7348) begin
        bht_bank_rd_data_out_0_87 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_87 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_527_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_88 <= 2'h0;
    end else if (bht_bank_sel_0_5_8) begin
      if (_T_7357) begin
        bht_bank_rd_data_out_0_88 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_88 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_527_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_89 <= 2'h0;
    end else if (bht_bank_sel_0_5_9) begin
      if (_T_7366) begin
        bht_bank_rd_data_out_0_89 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_89 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_527_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_90 <= 2'h0;
    end else if (bht_bank_sel_0_5_10) begin
      if (_T_7375) begin
        bht_bank_rd_data_out_0_90 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_90 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_527_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_91 <= 2'h0;
    end else if (bht_bank_sel_0_5_11) begin
      if (_T_7384) begin
        bht_bank_rd_data_out_0_91 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_91 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_527_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_92 <= 2'h0;
    end else if (bht_bank_sel_0_5_12) begin
      if (_T_7393) begin
        bht_bank_rd_data_out_0_92 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_92 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_527_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_93 <= 2'h0;
    end else if (bht_bank_sel_0_5_13) begin
      if (_T_7402) begin
        bht_bank_rd_data_out_0_93 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_93 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_527_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_94 <= 2'h0;
    end else if (bht_bank_sel_0_5_14) begin
      if (_T_7411) begin
        bht_bank_rd_data_out_0_94 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_94 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_527_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_95 <= 2'h0;
    end else if (bht_bank_sel_0_5_15) begin
      if (_T_7420) begin
        bht_bank_rd_data_out_0_95 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_95 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_528_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_96 <= 2'h0;
    end else if (bht_bank_sel_0_6_0) begin
      if (_T_7429) begin
        bht_bank_rd_data_out_0_96 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_96 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_528_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_97 <= 2'h0;
    end else if (bht_bank_sel_0_6_1) begin
      if (_T_7438) begin
        bht_bank_rd_data_out_0_97 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_97 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_528_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_98 <= 2'h0;
    end else if (bht_bank_sel_0_6_2) begin
      if (_T_7447) begin
        bht_bank_rd_data_out_0_98 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_98 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_528_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_99 <= 2'h0;
    end else if (bht_bank_sel_0_6_3) begin
      if (_T_7456) begin
        bht_bank_rd_data_out_0_99 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_99 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_528_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_100 <= 2'h0;
    end else if (bht_bank_sel_0_6_4) begin
      if (_T_7465) begin
        bht_bank_rd_data_out_0_100 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_100 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_528_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_101 <= 2'h0;
    end else if (bht_bank_sel_0_6_5) begin
      if (_T_7474) begin
        bht_bank_rd_data_out_0_101 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_101 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_528_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_102 <= 2'h0;
    end else if (bht_bank_sel_0_6_6) begin
      if (_T_7483) begin
        bht_bank_rd_data_out_0_102 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_102 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_528_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_103 <= 2'h0;
    end else if (bht_bank_sel_0_6_7) begin
      if (_T_7492) begin
        bht_bank_rd_data_out_0_103 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_103 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_528_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_104 <= 2'h0;
    end else if (bht_bank_sel_0_6_8) begin
      if (_T_7501) begin
        bht_bank_rd_data_out_0_104 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_104 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_528_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_105 <= 2'h0;
    end else if (bht_bank_sel_0_6_9) begin
      if (_T_7510) begin
        bht_bank_rd_data_out_0_105 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_105 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_528_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_106 <= 2'h0;
    end else if (bht_bank_sel_0_6_10) begin
      if (_T_7519) begin
        bht_bank_rd_data_out_0_106 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_106 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_528_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_107 <= 2'h0;
    end else if (bht_bank_sel_0_6_11) begin
      if (_T_7528) begin
        bht_bank_rd_data_out_0_107 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_107 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_528_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_108 <= 2'h0;
    end else if (bht_bank_sel_0_6_12) begin
      if (_T_7537) begin
        bht_bank_rd_data_out_0_108 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_108 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_528_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_109 <= 2'h0;
    end else if (bht_bank_sel_0_6_13) begin
      if (_T_7546) begin
        bht_bank_rd_data_out_0_109 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_109 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_528_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_110 <= 2'h0;
    end else if (bht_bank_sel_0_6_14) begin
      if (_T_7555) begin
        bht_bank_rd_data_out_0_110 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_110 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_528_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_111 <= 2'h0;
    end else if (bht_bank_sel_0_6_15) begin
      if (_T_7564) begin
        bht_bank_rd_data_out_0_111 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_111 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_529_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_112 <= 2'h0;
    end else if (bht_bank_sel_0_7_0) begin
      if (_T_7573) begin
        bht_bank_rd_data_out_0_112 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_112 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_529_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_113 <= 2'h0;
    end else if (bht_bank_sel_0_7_1) begin
      if (_T_7582) begin
        bht_bank_rd_data_out_0_113 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_113 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_529_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_114 <= 2'h0;
    end else if (bht_bank_sel_0_7_2) begin
      if (_T_7591) begin
        bht_bank_rd_data_out_0_114 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_114 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_529_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_115 <= 2'h0;
    end else if (bht_bank_sel_0_7_3) begin
      if (_T_7600) begin
        bht_bank_rd_data_out_0_115 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_115 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_529_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_116 <= 2'h0;
    end else if (bht_bank_sel_0_7_4) begin
      if (_T_7609) begin
        bht_bank_rd_data_out_0_116 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_116 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_529_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_117 <= 2'h0;
    end else if (bht_bank_sel_0_7_5) begin
      if (_T_7618) begin
        bht_bank_rd_data_out_0_117 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_117 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_529_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_118 <= 2'h0;
    end else if (bht_bank_sel_0_7_6) begin
      if (_T_7627) begin
        bht_bank_rd_data_out_0_118 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_118 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_529_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_119 <= 2'h0;
    end else if (bht_bank_sel_0_7_7) begin
      if (_T_7636) begin
        bht_bank_rd_data_out_0_119 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_119 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_529_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_120 <= 2'h0;
    end else if (bht_bank_sel_0_7_8) begin
      if (_T_7645) begin
        bht_bank_rd_data_out_0_120 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_120 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_529_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_121 <= 2'h0;
    end else if (bht_bank_sel_0_7_9) begin
      if (_T_7654) begin
        bht_bank_rd_data_out_0_121 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_121 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_529_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_122 <= 2'h0;
    end else if (bht_bank_sel_0_7_10) begin
      if (_T_7663) begin
        bht_bank_rd_data_out_0_122 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_122 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_529_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_123 <= 2'h0;
    end else if (bht_bank_sel_0_7_11) begin
      if (_T_7672) begin
        bht_bank_rd_data_out_0_123 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_123 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_529_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_124 <= 2'h0;
    end else if (bht_bank_sel_0_7_12) begin
      if (_T_7681) begin
        bht_bank_rd_data_out_0_124 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_124 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_529_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_125 <= 2'h0;
    end else if (bht_bank_sel_0_7_13) begin
      if (_T_7690) begin
        bht_bank_rd_data_out_0_125 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_125 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_529_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_126 <= 2'h0;
    end else if (bht_bank_sel_0_7_14) begin
      if (_T_7699) begin
        bht_bank_rd_data_out_0_126 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_126 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_529_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_127 <= 2'h0;
    end else if (bht_bank_sel_0_7_15) begin
      if (_T_7708) begin
        bht_bank_rd_data_out_0_127 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_127 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_530_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_128 <= 2'h0;
    end else if (bht_bank_sel_0_8_0) begin
      if (_T_7717) begin
        bht_bank_rd_data_out_0_128 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_128 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_530_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_129 <= 2'h0;
    end else if (bht_bank_sel_0_8_1) begin
      if (_T_7726) begin
        bht_bank_rd_data_out_0_129 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_129 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_530_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_130 <= 2'h0;
    end else if (bht_bank_sel_0_8_2) begin
      if (_T_7735) begin
        bht_bank_rd_data_out_0_130 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_130 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_530_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_131 <= 2'h0;
    end else if (bht_bank_sel_0_8_3) begin
      if (_T_7744) begin
        bht_bank_rd_data_out_0_131 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_131 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_530_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_132 <= 2'h0;
    end else if (bht_bank_sel_0_8_4) begin
      if (_T_7753) begin
        bht_bank_rd_data_out_0_132 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_132 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_530_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_133 <= 2'h0;
    end else if (bht_bank_sel_0_8_5) begin
      if (_T_7762) begin
        bht_bank_rd_data_out_0_133 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_133 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_530_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_134 <= 2'h0;
    end else if (bht_bank_sel_0_8_6) begin
      if (_T_7771) begin
        bht_bank_rd_data_out_0_134 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_134 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_530_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_135 <= 2'h0;
    end else if (bht_bank_sel_0_8_7) begin
      if (_T_7780) begin
        bht_bank_rd_data_out_0_135 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_135 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_530_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_136 <= 2'h0;
    end else if (bht_bank_sel_0_8_8) begin
      if (_T_7789) begin
        bht_bank_rd_data_out_0_136 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_136 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_530_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_137 <= 2'h0;
    end else if (bht_bank_sel_0_8_9) begin
      if (_T_7798) begin
        bht_bank_rd_data_out_0_137 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_137 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_530_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_138 <= 2'h0;
    end else if (bht_bank_sel_0_8_10) begin
      if (_T_7807) begin
        bht_bank_rd_data_out_0_138 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_138 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_530_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_139 <= 2'h0;
    end else if (bht_bank_sel_0_8_11) begin
      if (_T_7816) begin
        bht_bank_rd_data_out_0_139 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_139 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_530_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_140 <= 2'h0;
    end else if (bht_bank_sel_0_8_12) begin
      if (_T_7825) begin
        bht_bank_rd_data_out_0_140 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_140 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_530_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_141 <= 2'h0;
    end else if (bht_bank_sel_0_8_13) begin
      if (_T_7834) begin
        bht_bank_rd_data_out_0_141 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_141 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_530_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_142 <= 2'h0;
    end else if (bht_bank_sel_0_8_14) begin
      if (_T_7843) begin
        bht_bank_rd_data_out_0_142 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_142 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_530_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_143 <= 2'h0;
    end else if (bht_bank_sel_0_8_15) begin
      if (_T_7852) begin
        bht_bank_rd_data_out_0_143 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_143 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_531_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_144 <= 2'h0;
    end else if (bht_bank_sel_0_9_0) begin
      if (_T_7861) begin
        bht_bank_rd_data_out_0_144 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_144 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_531_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_145 <= 2'h0;
    end else if (bht_bank_sel_0_9_1) begin
      if (_T_7870) begin
        bht_bank_rd_data_out_0_145 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_145 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_531_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_146 <= 2'h0;
    end else if (bht_bank_sel_0_9_2) begin
      if (_T_7879) begin
        bht_bank_rd_data_out_0_146 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_146 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_531_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_147 <= 2'h0;
    end else if (bht_bank_sel_0_9_3) begin
      if (_T_7888) begin
        bht_bank_rd_data_out_0_147 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_147 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_531_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_148 <= 2'h0;
    end else if (bht_bank_sel_0_9_4) begin
      if (_T_7897) begin
        bht_bank_rd_data_out_0_148 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_148 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_531_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_149 <= 2'h0;
    end else if (bht_bank_sel_0_9_5) begin
      if (_T_7906) begin
        bht_bank_rd_data_out_0_149 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_149 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_531_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_150 <= 2'h0;
    end else if (bht_bank_sel_0_9_6) begin
      if (_T_7915) begin
        bht_bank_rd_data_out_0_150 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_150 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_531_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_151 <= 2'h0;
    end else if (bht_bank_sel_0_9_7) begin
      if (_T_7924) begin
        bht_bank_rd_data_out_0_151 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_151 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_531_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_152 <= 2'h0;
    end else if (bht_bank_sel_0_9_8) begin
      if (_T_7933) begin
        bht_bank_rd_data_out_0_152 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_152 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_531_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_153 <= 2'h0;
    end else if (bht_bank_sel_0_9_9) begin
      if (_T_7942) begin
        bht_bank_rd_data_out_0_153 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_153 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_531_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_154 <= 2'h0;
    end else if (bht_bank_sel_0_9_10) begin
      if (_T_7951) begin
        bht_bank_rd_data_out_0_154 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_154 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_531_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_155 <= 2'h0;
    end else if (bht_bank_sel_0_9_11) begin
      if (_T_7960) begin
        bht_bank_rd_data_out_0_155 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_155 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_531_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_156 <= 2'h0;
    end else if (bht_bank_sel_0_9_12) begin
      if (_T_7969) begin
        bht_bank_rd_data_out_0_156 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_156 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_531_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_157 <= 2'h0;
    end else if (bht_bank_sel_0_9_13) begin
      if (_T_7978) begin
        bht_bank_rd_data_out_0_157 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_157 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_531_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_158 <= 2'h0;
    end else if (bht_bank_sel_0_9_14) begin
      if (_T_7987) begin
        bht_bank_rd_data_out_0_158 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_158 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_531_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_159 <= 2'h0;
    end else if (bht_bank_sel_0_9_15) begin
      if (_T_7996) begin
        bht_bank_rd_data_out_0_159 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_159 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_532_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_160 <= 2'h0;
    end else if (bht_bank_sel_0_10_0) begin
      if (_T_8005) begin
        bht_bank_rd_data_out_0_160 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_160 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_532_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_161 <= 2'h0;
    end else if (bht_bank_sel_0_10_1) begin
      if (_T_8014) begin
        bht_bank_rd_data_out_0_161 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_161 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_532_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_162 <= 2'h0;
    end else if (bht_bank_sel_0_10_2) begin
      if (_T_8023) begin
        bht_bank_rd_data_out_0_162 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_162 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_532_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_163 <= 2'h0;
    end else if (bht_bank_sel_0_10_3) begin
      if (_T_8032) begin
        bht_bank_rd_data_out_0_163 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_163 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_532_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_164 <= 2'h0;
    end else if (bht_bank_sel_0_10_4) begin
      if (_T_8041) begin
        bht_bank_rd_data_out_0_164 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_164 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_532_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_165 <= 2'h0;
    end else if (bht_bank_sel_0_10_5) begin
      if (_T_8050) begin
        bht_bank_rd_data_out_0_165 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_165 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_532_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_166 <= 2'h0;
    end else if (bht_bank_sel_0_10_6) begin
      if (_T_8059) begin
        bht_bank_rd_data_out_0_166 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_166 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_532_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_167 <= 2'h0;
    end else if (bht_bank_sel_0_10_7) begin
      if (_T_8068) begin
        bht_bank_rd_data_out_0_167 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_167 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_532_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_168 <= 2'h0;
    end else if (bht_bank_sel_0_10_8) begin
      if (_T_8077) begin
        bht_bank_rd_data_out_0_168 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_168 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_532_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_169 <= 2'h0;
    end else if (bht_bank_sel_0_10_9) begin
      if (_T_8086) begin
        bht_bank_rd_data_out_0_169 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_169 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_532_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_170 <= 2'h0;
    end else if (bht_bank_sel_0_10_10) begin
      if (_T_8095) begin
        bht_bank_rd_data_out_0_170 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_170 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_532_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_171 <= 2'h0;
    end else if (bht_bank_sel_0_10_11) begin
      if (_T_8104) begin
        bht_bank_rd_data_out_0_171 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_171 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_532_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_172 <= 2'h0;
    end else if (bht_bank_sel_0_10_12) begin
      if (_T_8113) begin
        bht_bank_rd_data_out_0_172 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_172 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_532_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_173 <= 2'h0;
    end else if (bht_bank_sel_0_10_13) begin
      if (_T_8122) begin
        bht_bank_rd_data_out_0_173 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_173 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_532_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_174 <= 2'h0;
    end else if (bht_bank_sel_0_10_14) begin
      if (_T_8131) begin
        bht_bank_rd_data_out_0_174 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_174 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_532_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_175 <= 2'h0;
    end else if (bht_bank_sel_0_10_15) begin
      if (_T_8140) begin
        bht_bank_rd_data_out_0_175 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_175 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_533_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_176 <= 2'h0;
    end else if (bht_bank_sel_0_11_0) begin
      if (_T_8149) begin
        bht_bank_rd_data_out_0_176 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_176 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_533_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_177 <= 2'h0;
    end else if (bht_bank_sel_0_11_1) begin
      if (_T_8158) begin
        bht_bank_rd_data_out_0_177 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_177 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_533_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_178 <= 2'h0;
    end else if (bht_bank_sel_0_11_2) begin
      if (_T_8167) begin
        bht_bank_rd_data_out_0_178 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_178 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_533_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_179 <= 2'h0;
    end else if (bht_bank_sel_0_11_3) begin
      if (_T_8176) begin
        bht_bank_rd_data_out_0_179 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_179 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_533_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_180 <= 2'h0;
    end else if (bht_bank_sel_0_11_4) begin
      if (_T_8185) begin
        bht_bank_rd_data_out_0_180 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_180 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_533_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_181 <= 2'h0;
    end else if (bht_bank_sel_0_11_5) begin
      if (_T_8194) begin
        bht_bank_rd_data_out_0_181 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_181 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_533_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_182 <= 2'h0;
    end else if (bht_bank_sel_0_11_6) begin
      if (_T_8203) begin
        bht_bank_rd_data_out_0_182 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_182 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_533_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_183 <= 2'h0;
    end else if (bht_bank_sel_0_11_7) begin
      if (_T_8212) begin
        bht_bank_rd_data_out_0_183 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_183 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_533_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_184 <= 2'h0;
    end else if (bht_bank_sel_0_11_8) begin
      if (_T_8221) begin
        bht_bank_rd_data_out_0_184 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_184 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_533_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_185 <= 2'h0;
    end else if (bht_bank_sel_0_11_9) begin
      if (_T_8230) begin
        bht_bank_rd_data_out_0_185 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_185 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_533_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_186 <= 2'h0;
    end else if (bht_bank_sel_0_11_10) begin
      if (_T_8239) begin
        bht_bank_rd_data_out_0_186 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_186 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_533_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_187 <= 2'h0;
    end else if (bht_bank_sel_0_11_11) begin
      if (_T_8248) begin
        bht_bank_rd_data_out_0_187 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_187 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_533_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_188 <= 2'h0;
    end else if (bht_bank_sel_0_11_12) begin
      if (_T_8257) begin
        bht_bank_rd_data_out_0_188 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_188 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_533_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_189 <= 2'h0;
    end else if (bht_bank_sel_0_11_13) begin
      if (_T_8266) begin
        bht_bank_rd_data_out_0_189 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_189 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_533_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_190 <= 2'h0;
    end else if (bht_bank_sel_0_11_14) begin
      if (_T_8275) begin
        bht_bank_rd_data_out_0_190 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_190 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_533_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_191 <= 2'h0;
    end else if (bht_bank_sel_0_11_15) begin
      if (_T_8284) begin
        bht_bank_rd_data_out_0_191 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_191 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_534_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_192 <= 2'h0;
    end else if (bht_bank_sel_0_12_0) begin
      if (_T_8293) begin
        bht_bank_rd_data_out_0_192 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_192 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_534_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_193 <= 2'h0;
    end else if (bht_bank_sel_0_12_1) begin
      if (_T_8302) begin
        bht_bank_rd_data_out_0_193 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_193 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_534_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_194 <= 2'h0;
    end else if (bht_bank_sel_0_12_2) begin
      if (_T_8311) begin
        bht_bank_rd_data_out_0_194 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_194 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_534_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_195 <= 2'h0;
    end else if (bht_bank_sel_0_12_3) begin
      if (_T_8320) begin
        bht_bank_rd_data_out_0_195 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_195 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_534_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_196 <= 2'h0;
    end else if (bht_bank_sel_0_12_4) begin
      if (_T_8329) begin
        bht_bank_rd_data_out_0_196 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_196 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_534_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_197 <= 2'h0;
    end else if (bht_bank_sel_0_12_5) begin
      if (_T_8338) begin
        bht_bank_rd_data_out_0_197 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_197 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_534_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_198 <= 2'h0;
    end else if (bht_bank_sel_0_12_6) begin
      if (_T_8347) begin
        bht_bank_rd_data_out_0_198 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_198 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_534_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_199 <= 2'h0;
    end else if (bht_bank_sel_0_12_7) begin
      if (_T_8356) begin
        bht_bank_rd_data_out_0_199 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_199 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_534_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_200 <= 2'h0;
    end else if (bht_bank_sel_0_12_8) begin
      if (_T_8365) begin
        bht_bank_rd_data_out_0_200 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_200 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_534_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_201 <= 2'h0;
    end else if (bht_bank_sel_0_12_9) begin
      if (_T_8374) begin
        bht_bank_rd_data_out_0_201 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_201 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_534_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_202 <= 2'h0;
    end else if (bht_bank_sel_0_12_10) begin
      if (_T_8383) begin
        bht_bank_rd_data_out_0_202 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_202 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_534_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_203 <= 2'h0;
    end else if (bht_bank_sel_0_12_11) begin
      if (_T_8392) begin
        bht_bank_rd_data_out_0_203 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_203 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_534_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_204 <= 2'h0;
    end else if (bht_bank_sel_0_12_12) begin
      if (_T_8401) begin
        bht_bank_rd_data_out_0_204 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_204 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_534_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_205 <= 2'h0;
    end else if (bht_bank_sel_0_12_13) begin
      if (_T_8410) begin
        bht_bank_rd_data_out_0_205 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_205 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_534_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_206 <= 2'h0;
    end else if (bht_bank_sel_0_12_14) begin
      if (_T_8419) begin
        bht_bank_rd_data_out_0_206 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_206 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_534_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_207 <= 2'h0;
    end else if (bht_bank_sel_0_12_15) begin
      if (_T_8428) begin
        bht_bank_rd_data_out_0_207 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_207 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_535_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_208 <= 2'h0;
    end else if (bht_bank_sel_0_13_0) begin
      if (_T_8437) begin
        bht_bank_rd_data_out_0_208 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_208 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_535_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_209 <= 2'h0;
    end else if (bht_bank_sel_0_13_1) begin
      if (_T_8446) begin
        bht_bank_rd_data_out_0_209 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_209 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_535_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_210 <= 2'h0;
    end else if (bht_bank_sel_0_13_2) begin
      if (_T_8455) begin
        bht_bank_rd_data_out_0_210 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_210 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_535_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_211 <= 2'h0;
    end else if (bht_bank_sel_0_13_3) begin
      if (_T_8464) begin
        bht_bank_rd_data_out_0_211 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_211 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_535_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_212 <= 2'h0;
    end else if (bht_bank_sel_0_13_4) begin
      if (_T_8473) begin
        bht_bank_rd_data_out_0_212 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_212 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_535_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_213 <= 2'h0;
    end else if (bht_bank_sel_0_13_5) begin
      if (_T_8482) begin
        bht_bank_rd_data_out_0_213 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_213 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_535_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_214 <= 2'h0;
    end else if (bht_bank_sel_0_13_6) begin
      if (_T_8491) begin
        bht_bank_rd_data_out_0_214 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_214 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_535_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_215 <= 2'h0;
    end else if (bht_bank_sel_0_13_7) begin
      if (_T_8500) begin
        bht_bank_rd_data_out_0_215 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_215 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_535_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_216 <= 2'h0;
    end else if (bht_bank_sel_0_13_8) begin
      if (_T_8509) begin
        bht_bank_rd_data_out_0_216 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_216 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_535_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_217 <= 2'h0;
    end else if (bht_bank_sel_0_13_9) begin
      if (_T_8518) begin
        bht_bank_rd_data_out_0_217 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_217 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_535_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_218 <= 2'h0;
    end else if (bht_bank_sel_0_13_10) begin
      if (_T_8527) begin
        bht_bank_rd_data_out_0_218 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_218 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_535_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_219 <= 2'h0;
    end else if (bht_bank_sel_0_13_11) begin
      if (_T_8536) begin
        bht_bank_rd_data_out_0_219 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_219 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_535_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_220 <= 2'h0;
    end else if (bht_bank_sel_0_13_12) begin
      if (_T_8545) begin
        bht_bank_rd_data_out_0_220 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_220 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_535_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_221 <= 2'h0;
    end else if (bht_bank_sel_0_13_13) begin
      if (_T_8554) begin
        bht_bank_rd_data_out_0_221 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_221 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_535_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_222 <= 2'h0;
    end else if (bht_bank_sel_0_13_14) begin
      if (_T_8563) begin
        bht_bank_rd_data_out_0_222 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_222 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_535_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_223 <= 2'h0;
    end else if (bht_bank_sel_0_13_15) begin
      if (_T_8572) begin
        bht_bank_rd_data_out_0_223 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_223 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_536_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_224 <= 2'h0;
    end else if (bht_bank_sel_0_14_0) begin
      if (_T_8581) begin
        bht_bank_rd_data_out_0_224 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_224 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_536_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_225 <= 2'h0;
    end else if (bht_bank_sel_0_14_1) begin
      if (_T_8590) begin
        bht_bank_rd_data_out_0_225 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_225 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_536_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_226 <= 2'h0;
    end else if (bht_bank_sel_0_14_2) begin
      if (_T_8599) begin
        bht_bank_rd_data_out_0_226 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_226 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_536_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_227 <= 2'h0;
    end else if (bht_bank_sel_0_14_3) begin
      if (_T_8608) begin
        bht_bank_rd_data_out_0_227 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_227 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_536_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_228 <= 2'h0;
    end else if (bht_bank_sel_0_14_4) begin
      if (_T_8617) begin
        bht_bank_rd_data_out_0_228 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_228 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_536_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_229 <= 2'h0;
    end else if (bht_bank_sel_0_14_5) begin
      if (_T_8626) begin
        bht_bank_rd_data_out_0_229 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_229 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_536_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_230 <= 2'h0;
    end else if (bht_bank_sel_0_14_6) begin
      if (_T_8635) begin
        bht_bank_rd_data_out_0_230 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_230 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_536_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_231 <= 2'h0;
    end else if (bht_bank_sel_0_14_7) begin
      if (_T_8644) begin
        bht_bank_rd_data_out_0_231 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_231 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_536_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_232 <= 2'h0;
    end else if (bht_bank_sel_0_14_8) begin
      if (_T_8653) begin
        bht_bank_rd_data_out_0_232 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_232 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_536_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_233 <= 2'h0;
    end else if (bht_bank_sel_0_14_9) begin
      if (_T_8662) begin
        bht_bank_rd_data_out_0_233 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_233 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_536_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_234 <= 2'h0;
    end else if (bht_bank_sel_0_14_10) begin
      if (_T_8671) begin
        bht_bank_rd_data_out_0_234 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_234 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_536_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_235 <= 2'h0;
    end else if (bht_bank_sel_0_14_11) begin
      if (_T_8680) begin
        bht_bank_rd_data_out_0_235 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_235 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_536_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_236 <= 2'h0;
    end else if (bht_bank_sel_0_14_12) begin
      if (_T_8689) begin
        bht_bank_rd_data_out_0_236 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_236 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_536_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_237 <= 2'h0;
    end else if (bht_bank_sel_0_14_13) begin
      if (_T_8698) begin
        bht_bank_rd_data_out_0_237 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_237 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_536_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_238 <= 2'h0;
    end else if (bht_bank_sel_0_14_14) begin
      if (_T_8707) begin
        bht_bank_rd_data_out_0_238 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_238 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_536_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_239 <= 2'h0;
    end else if (bht_bank_sel_0_14_15) begin
      if (_T_8716) begin
        bht_bank_rd_data_out_0_239 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_239 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_537_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_240 <= 2'h0;
    end else if (bht_bank_sel_0_15_0) begin
      if (_T_8725) begin
        bht_bank_rd_data_out_0_240 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_240 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_537_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_241 <= 2'h0;
    end else if (bht_bank_sel_0_15_1) begin
      if (_T_8734) begin
        bht_bank_rd_data_out_0_241 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_241 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_537_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_242 <= 2'h0;
    end else if (bht_bank_sel_0_15_2) begin
      if (_T_8743) begin
        bht_bank_rd_data_out_0_242 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_242 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_537_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_243 <= 2'h0;
    end else if (bht_bank_sel_0_15_3) begin
      if (_T_8752) begin
        bht_bank_rd_data_out_0_243 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_243 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_537_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_244 <= 2'h0;
    end else if (bht_bank_sel_0_15_4) begin
      if (_T_8761) begin
        bht_bank_rd_data_out_0_244 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_244 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_537_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_245 <= 2'h0;
    end else if (bht_bank_sel_0_15_5) begin
      if (_T_8770) begin
        bht_bank_rd_data_out_0_245 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_245 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_537_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_246 <= 2'h0;
    end else if (bht_bank_sel_0_15_6) begin
      if (_T_8779) begin
        bht_bank_rd_data_out_0_246 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_246 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_537_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_247 <= 2'h0;
    end else if (bht_bank_sel_0_15_7) begin
      if (_T_8788) begin
        bht_bank_rd_data_out_0_247 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_247 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_537_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_248 <= 2'h0;
    end else if (bht_bank_sel_0_15_8) begin
      if (_T_8797) begin
        bht_bank_rd_data_out_0_248 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_248 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_537_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_249 <= 2'h0;
    end else if (bht_bank_sel_0_15_9) begin
      if (_T_8806) begin
        bht_bank_rd_data_out_0_249 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_249 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_537_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_250 <= 2'h0;
    end else if (bht_bank_sel_0_15_10) begin
      if (_T_8815) begin
        bht_bank_rd_data_out_0_250 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_250 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_537_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_251 <= 2'h0;
    end else if (bht_bank_sel_0_15_11) begin
      if (_T_8824) begin
        bht_bank_rd_data_out_0_251 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_251 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_537_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_252 <= 2'h0;
    end else if (bht_bank_sel_0_15_12) begin
      if (_T_8833) begin
        bht_bank_rd_data_out_0_252 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_252 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_537_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_253 <= 2'h0;
    end else if (bht_bank_sel_0_15_13) begin
      if (_T_8842) begin
        bht_bank_rd_data_out_0_253 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_253 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_537_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_254 <= 2'h0;
    end else if (bht_bank_sel_0_15_14) begin
      if (_T_8851) begin
        bht_bank_rd_data_out_0_254 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_254 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge rvclkhdr_537_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_255 <= 2'h0;
    end else if (bht_bank_sel_0_15_15) begin
      if (_T_8860) begin
        bht_bank_rd_data_out_0_255 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_255 <= io_exu_mp_pkt_hist;
      end
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      exu_mp_way_f <= 1'h0;
    end else begin
      exu_mp_way_f <= io_exu_mp_pkt_way;
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      exu_flush_final_d1 <= 1'h0;
    end else begin
      exu_flush_final_d1 <= io_exu_flush_final;
    end
  end
  always @(posedge rvclkhdr_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_lru_b0_f <= 256'h0;
    end else begin
      btb_lru_b0_f <= _T_182 | _T_184;
    end
  end
  always @(posedge rvclkhdr_1_io_l1clk or posedge reset) begin
    if (reset) begin
      ifc_fetch_adder_prior <= 30'h0;
    end else begin
      ifc_fetch_adder_prior <= io_ifc_fetch_addr_f[30:1];
    end
  end
  always @(posedge rvclkhdr_2_io_l1clk or posedge reset) begin
    if (reset) begin
      rets_out_0 <= 32'h0;
    end else begin
      rets_out_0 <= _T_481 | _T_482;
    end
  end
  always @(posedge rvclkhdr_3_io_l1clk or posedge reset) begin
    if (reset) begin
      rets_out_1 <= 32'h0;
    end else begin
      rets_out_1 <= _T_486 | _T_487;
    end
  end
  always @(posedge rvclkhdr_4_io_l1clk or posedge reset) begin
    if (reset) begin
      rets_out_2 <= 32'h0;
    end else begin
      rets_out_2 <= _T_491 | _T_492;
    end
  end
  always @(posedge rvclkhdr_5_io_l1clk or posedge reset) begin
    if (reset) begin
      rets_out_3 <= 32'h0;
    end else begin
      rets_out_3 <= _T_496 | _T_497;
    end
  end
  always @(posedge rvclkhdr_6_io_l1clk or posedge reset) begin
    if (reset) begin
      rets_out_4 <= 32'h0;
    end else begin
      rets_out_4 <= _T_501 | _T_502;
    end
  end
  always @(posedge rvclkhdr_7_io_l1clk or posedge reset) begin
    if (reset) begin
      rets_out_5 <= 32'h0;
    end else begin
      rets_out_5 <= _T_506 | _T_507;
    end
  end
  always @(posedge rvclkhdr_8_io_l1clk or posedge reset) begin
    if (reset) begin
      rets_out_6 <= 32'h0;
    end else begin
      rets_out_6 <= _T_511 | _T_512;
    end
  end
  always @(posedge rvclkhdr_9_io_l1clk or posedge reset) begin
    if (reset) begin
      rets_out_7 <= 32'h0;
    end else begin
      rets_out_7 <= rets_out_6;
    end
  end
endmodule
