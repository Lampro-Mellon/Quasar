module pic_ctrl(
  input         clock,
  input         reset,
  input         io_scan_mode,
  input         io_free_clk,
  input         io_clk_override,
  input         io_io_clk_override,
  input  [31:0] io_extintsrc_req,
  input         io_lsu_pic_picm_wren,
  input         io_lsu_pic_picm_rden,
  input         io_lsu_pic_picm_mken,
  input  [31:0] io_lsu_pic_picm_rdaddr,
  input  [31:0] io_lsu_pic_picm_wraddr,
  input  [31:0] io_lsu_pic_picm_wr_data,
  output [31:0] io_lsu_pic_picm_rd_data,
  output [7:0]  io_dec_pic_pic_claimid,
  output [3:0]  io_dec_pic_pic_pl,
  output        io_dec_pic_mhwakeup,
  input  [3:0]  io_dec_pic_dec_tlu_meicurpl,
  input  [3:0]  io_dec_pic_dec_tlu_meipt,
  output        io_dec_pic_mexintpend
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] picm_raddr_ff; // @[pic_ctrl.scala 101:56]
  reg [31:0] picm_waddr_ff; // @[pic_ctrl.scala 102:57]
  reg  picm_wren_ff; // @[pic_ctrl.scala 103:53]
  reg  picm_rden_ff; // @[pic_ctrl.scala 104:53]
  reg  picm_mken_ff; // @[pic_ctrl.scala 105:53]
  reg [31:0] picm_wr_data_ff; // @[pic_ctrl.scala 106:58]
  reg [1:0] gw_config_reg_31; // @[Reg.scala 27:20]
  wire  waddr_intenable_base_match = picm_waddr_ff[31:7] == 25'h1e01840; // @[pic_ctrl.scala 133:71]
  wire  _T_465 = picm_waddr_ff[6:2] == 5'h1f; // @[pic_ctrl.scala 158:139]
  wire  _T_466 = waddr_intenable_base_match & _T_465; // @[pic_ctrl.scala 158:106]
  wire  intenable_reg_we_31 = _T_466 & picm_wren_ff; // @[pic_ctrl.scala 158:153]
  wire  _T_1239 = gw_config_reg_31[1] | intenable_reg_we_31; // @[pic_ctrl.scala 170:95]
  reg  intenable_reg_31; // @[Reg.scala 27:20]
  wire  _T_1240 = _T_1239 | intenable_reg_31; // @[pic_ctrl.scala 170:117]
  wire  addr_clear_gw_base_match = picm_waddr_ff[31:7] == 25'h1e018a0; // @[pic_ctrl.scala 131:71]
  wire  _T_838 = addr_clear_gw_base_match & _T_465; // @[pic_ctrl.scala 162:106]
  wire  gw_clear_reg_we_31 = _T_838 & picm_wren_ff; // @[pic_ctrl.scala 162:153]
  wire  _T_1241 = _T_1240 | gw_clear_reg_we_31; // @[pic_ctrl.scala 170:136]
  reg [1:0] gw_config_reg_30; // @[Reg.scala 27:20]
  wire  _T_462 = picm_waddr_ff[6:2] == 5'h1e; // @[pic_ctrl.scala 158:139]
  wire  _T_463 = waddr_intenable_base_match & _T_462; // @[pic_ctrl.scala 158:106]
  wire  intenable_reg_we_30 = _T_463 & picm_wren_ff; // @[pic_ctrl.scala 158:153]
  wire  _T_1235 = gw_config_reg_30[1] | intenable_reg_we_30; // @[pic_ctrl.scala 170:95]
  reg  intenable_reg_30; // @[Reg.scala 27:20]
  wire  _T_1236 = _T_1235 | intenable_reg_30; // @[pic_ctrl.scala 170:117]
  wire  _T_835 = addr_clear_gw_base_match & _T_462; // @[pic_ctrl.scala 162:106]
  wire  gw_clear_reg_we_30 = _T_835 & picm_wren_ff; // @[pic_ctrl.scala 162:153]
  wire  _T_1237 = _T_1236 | gw_clear_reg_we_30; // @[pic_ctrl.scala 170:136]
  reg [1:0] gw_config_reg_29; // @[Reg.scala 27:20]
  wire  _T_459 = picm_waddr_ff[6:2] == 5'h1d; // @[pic_ctrl.scala 158:139]
  wire  _T_460 = waddr_intenable_base_match & _T_459; // @[pic_ctrl.scala 158:106]
  wire  intenable_reg_we_29 = _T_460 & picm_wren_ff; // @[pic_ctrl.scala 158:153]
  wire  _T_1231 = gw_config_reg_29[1] | intenable_reg_we_29; // @[pic_ctrl.scala 170:95]
  reg  intenable_reg_29; // @[Reg.scala 27:20]
  wire  _T_1232 = _T_1231 | intenable_reg_29; // @[pic_ctrl.scala 170:117]
  wire  _T_832 = addr_clear_gw_base_match & _T_459; // @[pic_ctrl.scala 162:106]
  wire  gw_clear_reg_we_29 = _T_832 & picm_wren_ff; // @[pic_ctrl.scala 162:153]
  wire  _T_1233 = _T_1232 | gw_clear_reg_we_29; // @[pic_ctrl.scala 170:136]
  reg [1:0] gw_config_reg_28; // @[Reg.scala 27:20]
  wire  _T_456 = picm_waddr_ff[6:2] == 5'h1c; // @[pic_ctrl.scala 158:139]
  wire  _T_457 = waddr_intenable_base_match & _T_456; // @[pic_ctrl.scala 158:106]
  wire  intenable_reg_we_28 = _T_457 & picm_wren_ff; // @[pic_ctrl.scala 158:153]
  wire  _T_1227 = gw_config_reg_28[1] | intenable_reg_we_28; // @[pic_ctrl.scala 170:95]
  reg  intenable_reg_28; // @[Reg.scala 27:20]
  wire  _T_1228 = _T_1227 | intenable_reg_28; // @[pic_ctrl.scala 170:117]
  wire  _T_829 = addr_clear_gw_base_match & _T_456; // @[pic_ctrl.scala 162:106]
  wire  gw_clear_reg_we_28 = _T_829 & picm_wren_ff; // @[pic_ctrl.scala 162:153]
  wire  _T_1229 = _T_1228 | gw_clear_reg_we_28; // @[pic_ctrl.scala 170:136]
  reg [1:0] gw_config_reg_27; // @[Reg.scala 27:20]
  wire  _T_453 = picm_waddr_ff[6:2] == 5'h1b; // @[pic_ctrl.scala 158:139]
  wire  _T_454 = waddr_intenable_base_match & _T_453; // @[pic_ctrl.scala 158:106]
  wire  intenable_reg_we_27 = _T_454 & picm_wren_ff; // @[pic_ctrl.scala 158:153]
  wire  _T_1223 = gw_config_reg_27[1] | intenable_reg_we_27; // @[pic_ctrl.scala 170:95]
  reg  intenable_reg_27; // @[Reg.scala 27:20]
  wire  _T_1224 = _T_1223 | intenable_reg_27; // @[pic_ctrl.scala 170:117]
  wire  _T_826 = addr_clear_gw_base_match & _T_453; // @[pic_ctrl.scala 162:106]
  wire  gw_clear_reg_we_27 = _T_826 & picm_wren_ff; // @[pic_ctrl.scala 162:153]
  wire  _T_1225 = _T_1224 | gw_clear_reg_we_27; // @[pic_ctrl.scala 170:136]
  reg [1:0] gw_config_reg_26; // @[Reg.scala 27:20]
  wire  _T_450 = picm_waddr_ff[6:2] == 5'h1a; // @[pic_ctrl.scala 158:139]
  wire  _T_451 = waddr_intenable_base_match & _T_450; // @[pic_ctrl.scala 158:106]
  wire  intenable_reg_we_26 = _T_451 & picm_wren_ff; // @[pic_ctrl.scala 158:153]
  wire  _T_1219 = gw_config_reg_26[1] | intenable_reg_we_26; // @[pic_ctrl.scala 170:95]
  reg  intenable_reg_26; // @[Reg.scala 27:20]
  wire  _T_1220 = _T_1219 | intenable_reg_26; // @[pic_ctrl.scala 170:117]
  wire  _T_823 = addr_clear_gw_base_match & _T_450; // @[pic_ctrl.scala 162:106]
  wire  gw_clear_reg_we_26 = _T_823 & picm_wren_ff; // @[pic_ctrl.scala 162:153]
  wire  _T_1221 = _T_1220 | gw_clear_reg_we_26; // @[pic_ctrl.scala 170:136]
  reg [1:0] gw_config_reg_25; // @[Reg.scala 27:20]
  wire  _T_447 = picm_waddr_ff[6:2] == 5'h19; // @[pic_ctrl.scala 158:139]
  wire  _T_448 = waddr_intenable_base_match & _T_447; // @[pic_ctrl.scala 158:106]
  wire  intenable_reg_we_25 = _T_448 & picm_wren_ff; // @[pic_ctrl.scala 158:153]
  wire  _T_1215 = gw_config_reg_25[1] | intenable_reg_we_25; // @[pic_ctrl.scala 170:95]
  reg  intenable_reg_25; // @[Reg.scala 27:20]
  wire  _T_1216 = _T_1215 | intenable_reg_25; // @[pic_ctrl.scala 170:117]
  wire  _T_820 = addr_clear_gw_base_match & _T_447; // @[pic_ctrl.scala 162:106]
  wire  gw_clear_reg_we_25 = _T_820 & picm_wren_ff; // @[pic_ctrl.scala 162:153]
  wire  _T_1217 = _T_1216 | gw_clear_reg_we_25; // @[pic_ctrl.scala 170:136]
  reg [1:0] gw_config_reg_24; // @[Reg.scala 27:20]
  wire  _T_444 = picm_waddr_ff[6:2] == 5'h18; // @[pic_ctrl.scala 158:139]
  wire  _T_445 = waddr_intenable_base_match & _T_444; // @[pic_ctrl.scala 158:106]
  wire  intenable_reg_we_24 = _T_445 & picm_wren_ff; // @[pic_ctrl.scala 158:153]
  wire  _T_1211 = gw_config_reg_24[1] | intenable_reg_we_24; // @[pic_ctrl.scala 170:95]
  reg  intenable_reg_24; // @[Reg.scala 27:20]
  wire  _T_1212 = _T_1211 | intenable_reg_24; // @[pic_ctrl.scala 170:117]
  wire  _T_817 = addr_clear_gw_base_match & _T_444; // @[pic_ctrl.scala 162:106]
  wire  gw_clear_reg_we_24 = _T_817 & picm_wren_ff; // @[pic_ctrl.scala 162:153]
  wire  _T_1213 = _T_1212 | gw_clear_reg_we_24; // @[pic_ctrl.scala 170:136]
  reg [1:0] gw_config_reg_23; // @[Reg.scala 27:20]
  wire  _T_441 = picm_waddr_ff[6:2] == 5'h17; // @[pic_ctrl.scala 158:139]
  wire  _T_442 = waddr_intenable_base_match & _T_441; // @[pic_ctrl.scala 158:106]
  wire  intenable_reg_we_23 = _T_442 & picm_wren_ff; // @[pic_ctrl.scala 158:153]
  wire  _T_1207 = gw_config_reg_23[1] | intenable_reg_we_23; // @[pic_ctrl.scala 170:95]
  reg  intenable_reg_23; // @[Reg.scala 27:20]
  wire  _T_1208 = _T_1207 | intenable_reg_23; // @[pic_ctrl.scala 170:117]
  wire  _T_814 = addr_clear_gw_base_match & _T_441; // @[pic_ctrl.scala 162:106]
  wire  gw_clear_reg_we_23 = _T_814 & picm_wren_ff; // @[pic_ctrl.scala 162:153]
  wire  _T_1209 = _T_1208 | gw_clear_reg_we_23; // @[pic_ctrl.scala 170:136]
  reg [1:0] gw_config_reg_22; // @[Reg.scala 27:20]
  wire  _T_438 = picm_waddr_ff[6:2] == 5'h16; // @[pic_ctrl.scala 158:139]
  wire  _T_439 = waddr_intenable_base_match & _T_438; // @[pic_ctrl.scala 158:106]
  wire  intenable_reg_we_22 = _T_439 & picm_wren_ff; // @[pic_ctrl.scala 158:153]
  wire  _T_1203 = gw_config_reg_22[1] | intenable_reg_we_22; // @[pic_ctrl.scala 170:95]
  reg  intenable_reg_22; // @[Reg.scala 27:20]
  wire  _T_1204 = _T_1203 | intenable_reg_22; // @[pic_ctrl.scala 170:117]
  wire  _T_811 = addr_clear_gw_base_match & _T_438; // @[pic_ctrl.scala 162:106]
  wire  gw_clear_reg_we_22 = _T_811 & picm_wren_ff; // @[pic_ctrl.scala 162:153]
  wire  _T_1205 = _T_1204 | gw_clear_reg_we_22; // @[pic_ctrl.scala 170:136]
  wire [9:0] _T_1250 = {_T_1241,_T_1237,_T_1233,_T_1229,_T_1225,_T_1221,_T_1217,_T_1213,_T_1209,_T_1205}; // @[Cat.scala 29:58]
  reg [1:0] gw_config_reg_21; // @[Reg.scala 27:20]
  wire  _T_435 = picm_waddr_ff[6:2] == 5'h15; // @[pic_ctrl.scala 158:139]
  wire  _T_436 = waddr_intenable_base_match & _T_435; // @[pic_ctrl.scala 158:106]
  wire  intenable_reg_we_21 = _T_436 & picm_wren_ff; // @[pic_ctrl.scala 158:153]
  wire  _T_1199 = gw_config_reg_21[1] | intenable_reg_we_21; // @[pic_ctrl.scala 170:95]
  reg  intenable_reg_21; // @[Reg.scala 27:20]
  wire  _T_1200 = _T_1199 | intenable_reg_21; // @[pic_ctrl.scala 170:117]
  wire  _T_808 = addr_clear_gw_base_match & _T_435; // @[pic_ctrl.scala 162:106]
  wire  gw_clear_reg_we_21 = _T_808 & picm_wren_ff; // @[pic_ctrl.scala 162:153]
  wire  _T_1201 = _T_1200 | gw_clear_reg_we_21; // @[pic_ctrl.scala 170:136]
  reg [1:0] gw_config_reg_20; // @[Reg.scala 27:20]
  wire  _T_432 = picm_waddr_ff[6:2] == 5'h14; // @[pic_ctrl.scala 158:139]
  wire  _T_433 = waddr_intenable_base_match & _T_432; // @[pic_ctrl.scala 158:106]
  wire  intenable_reg_we_20 = _T_433 & picm_wren_ff; // @[pic_ctrl.scala 158:153]
  wire  _T_1195 = gw_config_reg_20[1] | intenable_reg_we_20; // @[pic_ctrl.scala 170:95]
  reg  intenable_reg_20; // @[Reg.scala 27:20]
  wire  _T_1196 = _T_1195 | intenable_reg_20; // @[pic_ctrl.scala 170:117]
  wire  _T_805 = addr_clear_gw_base_match & _T_432; // @[pic_ctrl.scala 162:106]
  wire  gw_clear_reg_we_20 = _T_805 & picm_wren_ff; // @[pic_ctrl.scala 162:153]
  wire  _T_1197 = _T_1196 | gw_clear_reg_we_20; // @[pic_ctrl.scala 170:136]
  reg [1:0] gw_config_reg_19; // @[Reg.scala 27:20]
  wire  _T_429 = picm_waddr_ff[6:2] == 5'h13; // @[pic_ctrl.scala 158:139]
  wire  _T_430 = waddr_intenable_base_match & _T_429; // @[pic_ctrl.scala 158:106]
  wire  intenable_reg_we_19 = _T_430 & picm_wren_ff; // @[pic_ctrl.scala 158:153]
  wire  _T_1191 = gw_config_reg_19[1] | intenable_reg_we_19; // @[pic_ctrl.scala 170:95]
  reg  intenable_reg_19; // @[Reg.scala 27:20]
  wire  _T_1192 = _T_1191 | intenable_reg_19; // @[pic_ctrl.scala 170:117]
  wire  _T_802 = addr_clear_gw_base_match & _T_429; // @[pic_ctrl.scala 162:106]
  wire  gw_clear_reg_we_19 = _T_802 & picm_wren_ff; // @[pic_ctrl.scala 162:153]
  wire  _T_1193 = _T_1192 | gw_clear_reg_we_19; // @[pic_ctrl.scala 170:136]
  reg [1:0] gw_config_reg_18; // @[Reg.scala 27:20]
  wire  _T_426 = picm_waddr_ff[6:2] == 5'h12; // @[pic_ctrl.scala 158:139]
  wire  _T_427 = waddr_intenable_base_match & _T_426; // @[pic_ctrl.scala 158:106]
  wire  intenable_reg_we_18 = _T_427 & picm_wren_ff; // @[pic_ctrl.scala 158:153]
  wire  _T_1187 = gw_config_reg_18[1] | intenable_reg_we_18; // @[pic_ctrl.scala 170:95]
  reg  intenable_reg_18; // @[Reg.scala 27:20]
  wire  _T_1188 = _T_1187 | intenable_reg_18; // @[pic_ctrl.scala 170:117]
  wire  _T_799 = addr_clear_gw_base_match & _T_426; // @[pic_ctrl.scala 162:106]
  wire  gw_clear_reg_we_18 = _T_799 & picm_wren_ff; // @[pic_ctrl.scala 162:153]
  wire  _T_1189 = _T_1188 | gw_clear_reg_we_18; // @[pic_ctrl.scala 170:136]
  reg [1:0] gw_config_reg_17; // @[Reg.scala 27:20]
  wire  _T_423 = picm_waddr_ff[6:2] == 5'h11; // @[pic_ctrl.scala 158:139]
  wire  _T_424 = waddr_intenable_base_match & _T_423; // @[pic_ctrl.scala 158:106]
  wire  intenable_reg_we_17 = _T_424 & picm_wren_ff; // @[pic_ctrl.scala 158:153]
  wire  _T_1183 = gw_config_reg_17[1] | intenable_reg_we_17; // @[pic_ctrl.scala 170:95]
  reg  intenable_reg_17; // @[Reg.scala 27:20]
  wire  _T_1184 = _T_1183 | intenable_reg_17; // @[pic_ctrl.scala 170:117]
  wire  _T_796 = addr_clear_gw_base_match & _T_423; // @[pic_ctrl.scala 162:106]
  wire  gw_clear_reg_we_17 = _T_796 & picm_wren_ff; // @[pic_ctrl.scala 162:153]
  wire  _T_1185 = _T_1184 | gw_clear_reg_we_17; // @[pic_ctrl.scala 170:136]
  reg [1:0] gw_config_reg_16; // @[Reg.scala 27:20]
  wire  _T_420 = picm_waddr_ff[6:2] == 5'h10; // @[pic_ctrl.scala 158:139]
  wire  _T_421 = waddr_intenable_base_match & _T_420; // @[pic_ctrl.scala 158:106]
  wire  intenable_reg_we_16 = _T_421 & picm_wren_ff; // @[pic_ctrl.scala 158:153]
  wire  _T_1179 = gw_config_reg_16[1] | intenable_reg_we_16; // @[pic_ctrl.scala 170:95]
  reg  intenable_reg_16; // @[Reg.scala 27:20]
  wire  _T_1180 = _T_1179 | intenable_reg_16; // @[pic_ctrl.scala 170:117]
  wire  _T_793 = addr_clear_gw_base_match & _T_420; // @[pic_ctrl.scala 162:106]
  wire  gw_clear_reg_we_16 = _T_793 & picm_wren_ff; // @[pic_ctrl.scala 162:153]
  wire  _T_1181 = _T_1180 | gw_clear_reg_we_16; // @[pic_ctrl.scala 170:136]
  reg [1:0] gw_config_reg_15; // @[Reg.scala 27:20]
  wire  _T_417 = picm_waddr_ff[6:2] == 5'hf; // @[pic_ctrl.scala 158:139]
  wire  _T_418 = waddr_intenable_base_match & _T_417; // @[pic_ctrl.scala 158:106]
  wire  intenable_reg_we_15 = _T_418 & picm_wren_ff; // @[pic_ctrl.scala 158:153]
  wire  _T_1175 = gw_config_reg_15[1] | intenable_reg_we_15; // @[pic_ctrl.scala 170:95]
  reg  intenable_reg_15; // @[Reg.scala 27:20]
  wire  _T_1176 = _T_1175 | intenable_reg_15; // @[pic_ctrl.scala 170:117]
  wire  _T_790 = addr_clear_gw_base_match & _T_417; // @[pic_ctrl.scala 162:106]
  wire  gw_clear_reg_we_15 = _T_790 & picm_wren_ff; // @[pic_ctrl.scala 162:153]
  wire  _T_1177 = _T_1176 | gw_clear_reg_we_15; // @[pic_ctrl.scala 170:136]
  reg [1:0] gw_config_reg_14; // @[Reg.scala 27:20]
  wire  _T_414 = picm_waddr_ff[6:2] == 5'he; // @[pic_ctrl.scala 158:139]
  wire  _T_415 = waddr_intenable_base_match & _T_414; // @[pic_ctrl.scala 158:106]
  wire  intenable_reg_we_14 = _T_415 & picm_wren_ff; // @[pic_ctrl.scala 158:153]
  wire  _T_1171 = gw_config_reg_14[1] | intenable_reg_we_14; // @[pic_ctrl.scala 170:95]
  reg  intenable_reg_14; // @[Reg.scala 27:20]
  wire  _T_1172 = _T_1171 | intenable_reg_14; // @[pic_ctrl.scala 170:117]
  wire  _T_787 = addr_clear_gw_base_match & _T_414; // @[pic_ctrl.scala 162:106]
  wire  gw_clear_reg_we_14 = _T_787 & picm_wren_ff; // @[pic_ctrl.scala 162:153]
  wire  _T_1173 = _T_1172 | gw_clear_reg_we_14; // @[pic_ctrl.scala 170:136]
  reg [1:0] gw_config_reg_13; // @[Reg.scala 27:20]
  wire  _T_411 = picm_waddr_ff[6:2] == 5'hd; // @[pic_ctrl.scala 158:139]
  wire  _T_412 = waddr_intenable_base_match & _T_411; // @[pic_ctrl.scala 158:106]
  wire  intenable_reg_we_13 = _T_412 & picm_wren_ff; // @[pic_ctrl.scala 158:153]
  wire  _T_1167 = gw_config_reg_13[1] | intenable_reg_we_13; // @[pic_ctrl.scala 170:95]
  reg  intenable_reg_13; // @[Reg.scala 27:20]
  wire  _T_1168 = _T_1167 | intenable_reg_13; // @[pic_ctrl.scala 170:117]
  wire  _T_784 = addr_clear_gw_base_match & _T_411; // @[pic_ctrl.scala 162:106]
  wire  gw_clear_reg_we_13 = _T_784 & picm_wren_ff; // @[pic_ctrl.scala 162:153]
  wire  _T_1169 = _T_1168 | gw_clear_reg_we_13; // @[pic_ctrl.scala 170:136]
  wire [18:0] _T_1259 = {_T_1250,_T_1201,_T_1197,_T_1193,_T_1189,_T_1185,_T_1181,_T_1177,_T_1173,_T_1169}; // @[Cat.scala 29:58]
  reg [1:0] gw_config_reg_12; // @[Reg.scala 27:20]
  wire  _T_408 = picm_waddr_ff[6:2] == 5'hc; // @[pic_ctrl.scala 158:139]
  wire  _T_409 = waddr_intenable_base_match & _T_408; // @[pic_ctrl.scala 158:106]
  wire  intenable_reg_we_12 = _T_409 & picm_wren_ff; // @[pic_ctrl.scala 158:153]
  wire  _T_1163 = gw_config_reg_12[1] | intenable_reg_we_12; // @[pic_ctrl.scala 170:95]
  reg  intenable_reg_12; // @[Reg.scala 27:20]
  wire  _T_1164 = _T_1163 | intenable_reg_12; // @[pic_ctrl.scala 170:117]
  wire  _T_781 = addr_clear_gw_base_match & _T_408; // @[pic_ctrl.scala 162:106]
  wire  gw_clear_reg_we_12 = _T_781 & picm_wren_ff; // @[pic_ctrl.scala 162:153]
  wire  _T_1165 = _T_1164 | gw_clear_reg_we_12; // @[pic_ctrl.scala 170:136]
  reg [1:0] gw_config_reg_11; // @[Reg.scala 27:20]
  wire  _T_405 = picm_waddr_ff[6:2] == 5'hb; // @[pic_ctrl.scala 158:139]
  wire  _T_406 = waddr_intenable_base_match & _T_405; // @[pic_ctrl.scala 158:106]
  wire  intenable_reg_we_11 = _T_406 & picm_wren_ff; // @[pic_ctrl.scala 158:153]
  wire  _T_1159 = gw_config_reg_11[1] | intenable_reg_we_11; // @[pic_ctrl.scala 170:95]
  reg  intenable_reg_11; // @[Reg.scala 27:20]
  wire  _T_1160 = _T_1159 | intenable_reg_11; // @[pic_ctrl.scala 170:117]
  wire  _T_778 = addr_clear_gw_base_match & _T_405; // @[pic_ctrl.scala 162:106]
  wire  gw_clear_reg_we_11 = _T_778 & picm_wren_ff; // @[pic_ctrl.scala 162:153]
  wire  _T_1161 = _T_1160 | gw_clear_reg_we_11; // @[pic_ctrl.scala 170:136]
  reg [1:0] gw_config_reg_10; // @[Reg.scala 27:20]
  wire  _T_402 = picm_waddr_ff[6:2] == 5'ha; // @[pic_ctrl.scala 158:139]
  wire  _T_403 = waddr_intenable_base_match & _T_402; // @[pic_ctrl.scala 158:106]
  wire  intenable_reg_we_10 = _T_403 & picm_wren_ff; // @[pic_ctrl.scala 158:153]
  wire  _T_1155 = gw_config_reg_10[1] | intenable_reg_we_10; // @[pic_ctrl.scala 170:95]
  reg  intenable_reg_10; // @[Reg.scala 27:20]
  wire  _T_1156 = _T_1155 | intenable_reg_10; // @[pic_ctrl.scala 170:117]
  wire  _T_775 = addr_clear_gw_base_match & _T_402; // @[pic_ctrl.scala 162:106]
  wire  gw_clear_reg_we_10 = _T_775 & picm_wren_ff; // @[pic_ctrl.scala 162:153]
  wire  _T_1157 = _T_1156 | gw_clear_reg_we_10; // @[pic_ctrl.scala 170:136]
  reg [1:0] gw_config_reg_9; // @[Reg.scala 27:20]
  wire  _T_399 = picm_waddr_ff[6:2] == 5'h9; // @[pic_ctrl.scala 158:139]
  wire  _T_400 = waddr_intenable_base_match & _T_399; // @[pic_ctrl.scala 158:106]
  wire  intenable_reg_we_9 = _T_400 & picm_wren_ff; // @[pic_ctrl.scala 158:153]
  wire  _T_1151 = gw_config_reg_9[1] | intenable_reg_we_9; // @[pic_ctrl.scala 170:95]
  reg  intenable_reg_9; // @[Reg.scala 27:20]
  wire  _T_1152 = _T_1151 | intenable_reg_9; // @[pic_ctrl.scala 170:117]
  wire  _T_772 = addr_clear_gw_base_match & _T_399; // @[pic_ctrl.scala 162:106]
  wire  gw_clear_reg_we_9 = _T_772 & picm_wren_ff; // @[pic_ctrl.scala 162:153]
  wire  _T_1153 = _T_1152 | gw_clear_reg_we_9; // @[pic_ctrl.scala 170:136]
  reg [1:0] gw_config_reg_8; // @[Reg.scala 27:20]
  wire  _T_396 = picm_waddr_ff[6:2] == 5'h8; // @[pic_ctrl.scala 158:139]
  wire  _T_397 = waddr_intenable_base_match & _T_396; // @[pic_ctrl.scala 158:106]
  wire  intenable_reg_we_8 = _T_397 & picm_wren_ff; // @[pic_ctrl.scala 158:153]
  wire  _T_1147 = gw_config_reg_8[1] | intenable_reg_we_8; // @[pic_ctrl.scala 170:95]
  reg  intenable_reg_8; // @[Reg.scala 27:20]
  wire  _T_1148 = _T_1147 | intenable_reg_8; // @[pic_ctrl.scala 170:117]
  wire  _T_769 = addr_clear_gw_base_match & _T_396; // @[pic_ctrl.scala 162:106]
  wire  gw_clear_reg_we_8 = _T_769 & picm_wren_ff; // @[pic_ctrl.scala 162:153]
  wire  _T_1149 = _T_1148 | gw_clear_reg_we_8; // @[pic_ctrl.scala 170:136]
  reg [1:0] gw_config_reg_7; // @[Reg.scala 27:20]
  wire  _T_393 = picm_waddr_ff[6:2] == 5'h7; // @[pic_ctrl.scala 158:139]
  wire  _T_394 = waddr_intenable_base_match & _T_393; // @[pic_ctrl.scala 158:106]
  wire  intenable_reg_we_7 = _T_394 & picm_wren_ff; // @[pic_ctrl.scala 158:153]
  wire  _T_1143 = gw_config_reg_7[1] | intenable_reg_we_7; // @[pic_ctrl.scala 170:95]
  reg  intenable_reg_7; // @[Reg.scala 27:20]
  wire  _T_1144 = _T_1143 | intenable_reg_7; // @[pic_ctrl.scala 170:117]
  wire  _T_766 = addr_clear_gw_base_match & _T_393; // @[pic_ctrl.scala 162:106]
  wire  gw_clear_reg_we_7 = _T_766 & picm_wren_ff; // @[pic_ctrl.scala 162:153]
  wire  _T_1145 = _T_1144 | gw_clear_reg_we_7; // @[pic_ctrl.scala 170:136]
  reg [1:0] gw_config_reg_6; // @[Reg.scala 27:20]
  wire  _T_390 = picm_waddr_ff[6:2] == 5'h6; // @[pic_ctrl.scala 158:139]
  wire  _T_391 = waddr_intenable_base_match & _T_390; // @[pic_ctrl.scala 158:106]
  wire  intenable_reg_we_6 = _T_391 & picm_wren_ff; // @[pic_ctrl.scala 158:153]
  wire  _T_1139 = gw_config_reg_6[1] | intenable_reg_we_6; // @[pic_ctrl.scala 170:95]
  reg  intenable_reg_6; // @[Reg.scala 27:20]
  wire  _T_1140 = _T_1139 | intenable_reg_6; // @[pic_ctrl.scala 170:117]
  wire  _T_763 = addr_clear_gw_base_match & _T_390; // @[pic_ctrl.scala 162:106]
  wire  gw_clear_reg_we_6 = _T_763 & picm_wren_ff; // @[pic_ctrl.scala 162:153]
  wire  _T_1141 = _T_1140 | gw_clear_reg_we_6; // @[pic_ctrl.scala 170:136]
  reg [1:0] gw_config_reg_5; // @[Reg.scala 27:20]
  wire  _T_387 = picm_waddr_ff[6:2] == 5'h5; // @[pic_ctrl.scala 158:139]
  wire  _T_388 = waddr_intenable_base_match & _T_387; // @[pic_ctrl.scala 158:106]
  wire  intenable_reg_we_5 = _T_388 & picm_wren_ff; // @[pic_ctrl.scala 158:153]
  wire  _T_1135 = gw_config_reg_5[1] | intenable_reg_we_5; // @[pic_ctrl.scala 170:95]
  reg  intenable_reg_5; // @[Reg.scala 27:20]
  wire  _T_1136 = _T_1135 | intenable_reg_5; // @[pic_ctrl.scala 170:117]
  wire  _T_760 = addr_clear_gw_base_match & _T_387; // @[pic_ctrl.scala 162:106]
  wire  gw_clear_reg_we_5 = _T_760 & picm_wren_ff; // @[pic_ctrl.scala 162:153]
  wire  _T_1137 = _T_1136 | gw_clear_reg_we_5; // @[pic_ctrl.scala 170:136]
  reg [1:0] gw_config_reg_4; // @[Reg.scala 27:20]
  wire  _T_384 = picm_waddr_ff[6:2] == 5'h4; // @[pic_ctrl.scala 158:139]
  wire  _T_385 = waddr_intenable_base_match & _T_384; // @[pic_ctrl.scala 158:106]
  wire  intenable_reg_we_4 = _T_385 & picm_wren_ff; // @[pic_ctrl.scala 158:153]
  wire  _T_1131 = gw_config_reg_4[1] | intenable_reg_we_4; // @[pic_ctrl.scala 170:95]
  reg  intenable_reg_4; // @[Reg.scala 27:20]
  wire  _T_1132 = _T_1131 | intenable_reg_4; // @[pic_ctrl.scala 170:117]
  wire  _T_757 = addr_clear_gw_base_match & _T_384; // @[pic_ctrl.scala 162:106]
  wire  gw_clear_reg_we_4 = _T_757 & picm_wren_ff; // @[pic_ctrl.scala 162:153]
  wire  _T_1133 = _T_1132 | gw_clear_reg_we_4; // @[pic_ctrl.scala 170:136]
  wire [27:0] _T_1268 = {_T_1259,_T_1165,_T_1161,_T_1157,_T_1153,_T_1149,_T_1145,_T_1141,_T_1137,_T_1133}; // @[Cat.scala 29:58]
  reg [1:0] gw_config_reg_3; // @[Reg.scala 27:20]
  wire  _T_381 = picm_waddr_ff[6:2] == 5'h3; // @[pic_ctrl.scala 158:139]
  wire  _T_382 = waddr_intenable_base_match & _T_381; // @[pic_ctrl.scala 158:106]
  wire  intenable_reg_we_3 = _T_382 & picm_wren_ff; // @[pic_ctrl.scala 158:153]
  wire  _T_1127 = gw_config_reg_3[1] | intenable_reg_we_3; // @[pic_ctrl.scala 170:95]
  reg  intenable_reg_3; // @[Reg.scala 27:20]
  wire  _T_1128 = _T_1127 | intenable_reg_3; // @[pic_ctrl.scala 170:117]
  wire  _T_754 = addr_clear_gw_base_match & _T_381; // @[pic_ctrl.scala 162:106]
  wire  gw_clear_reg_we_3 = _T_754 & picm_wren_ff; // @[pic_ctrl.scala 162:153]
  wire  _T_1129 = _T_1128 | gw_clear_reg_we_3; // @[pic_ctrl.scala 170:136]
  reg [1:0] gw_config_reg_2; // @[Reg.scala 27:20]
  wire  _T_378 = picm_waddr_ff[6:2] == 5'h2; // @[pic_ctrl.scala 158:139]
  wire  _T_379 = waddr_intenable_base_match & _T_378; // @[pic_ctrl.scala 158:106]
  wire  intenable_reg_we_2 = _T_379 & picm_wren_ff; // @[pic_ctrl.scala 158:153]
  wire  _T_1123 = gw_config_reg_2[1] | intenable_reg_we_2; // @[pic_ctrl.scala 170:95]
  reg  intenable_reg_2; // @[Reg.scala 27:20]
  wire  _T_1124 = _T_1123 | intenable_reg_2; // @[pic_ctrl.scala 170:117]
  wire  _T_751 = addr_clear_gw_base_match & _T_378; // @[pic_ctrl.scala 162:106]
  wire  gw_clear_reg_we_2 = _T_751 & picm_wren_ff; // @[pic_ctrl.scala 162:153]
  wire  _T_1125 = _T_1124 | gw_clear_reg_we_2; // @[pic_ctrl.scala 170:136]
  reg [1:0] gw_config_reg_1; // @[Reg.scala 27:20]
  wire  _T_375 = picm_waddr_ff[6:2] == 5'h1; // @[pic_ctrl.scala 158:139]
  wire  _T_376 = waddr_intenable_base_match & _T_375; // @[pic_ctrl.scala 158:106]
  wire  intenable_reg_we_1 = _T_376 & picm_wren_ff; // @[pic_ctrl.scala 158:153]
  wire  _T_1119 = gw_config_reg_1[1] | intenable_reg_we_1; // @[pic_ctrl.scala 170:95]
  reg  intenable_reg_1; // @[Reg.scala 27:20]
  wire  _T_1120 = _T_1119 | intenable_reg_1; // @[pic_ctrl.scala 170:117]
  wire  _T_748 = addr_clear_gw_base_match & _T_375; // @[pic_ctrl.scala 162:106]
  wire  gw_clear_reg_we_1 = _T_748 & picm_wren_ff; // @[pic_ctrl.scala 162:153]
  wire  _T_1121 = _T_1120 | gw_clear_reg_we_1; // @[pic_ctrl.scala 170:136]
  wire [31:0] intenable_clk_enable = {_T_1268,_T_1129,_T_1125,_T_1121,1'h0}; // @[Cat.scala 29:58]
  wire  _T_7 = |intenable_clk_enable[3:0]; // @[pic_ctrl.scala 116:72]
  wire  intenable_clk_enable_grp_0 = _T_7 | io_io_clk_override; // @[pic_ctrl.scala 116:76]
  wire  _T_11 = |intenable_clk_enable[7:4]; // @[pic_ctrl.scala 116:72]
  wire  intenable_clk_enable_grp_1 = _T_11 | io_io_clk_override; // @[pic_ctrl.scala 116:76]
  wire  _T_15 = |intenable_clk_enable[11:8]; // @[pic_ctrl.scala 116:72]
  wire  intenable_clk_enable_grp_2 = _T_15 | io_io_clk_override; // @[pic_ctrl.scala 116:76]
  wire  _T_19 = |intenable_clk_enable[15:12]; // @[pic_ctrl.scala 116:72]
  wire  intenable_clk_enable_grp_3 = _T_19 | io_io_clk_override; // @[pic_ctrl.scala 116:76]
  wire  _T_23 = |intenable_clk_enable[19:16]; // @[pic_ctrl.scala 116:72]
  wire  intenable_clk_enable_grp_4 = _T_23 | io_io_clk_override; // @[pic_ctrl.scala 116:76]
  wire  _T_27 = |intenable_clk_enable[23:20]; // @[pic_ctrl.scala 116:72]
  wire  intenable_clk_enable_grp_5 = _T_27 | io_io_clk_override; // @[pic_ctrl.scala 116:76]
  wire  _T_31 = |intenable_clk_enable[27:24]; // @[pic_ctrl.scala 116:72]
  wire  intenable_clk_enable_grp_6 = _T_31 | io_io_clk_override; // @[pic_ctrl.scala 116:76]
  wire  _T_35 = |intenable_clk_enable[31:28]; // @[pic_ctrl.scala 113:87]
  wire  intenable_clk_enable_grp_7 = _T_35 | io_io_clk_override; // @[pic_ctrl.scala 113:91]
  wire [31:0] _T_38 = picm_raddr_ff ^ 32'hf00c2000; // @[pic_ctrl.scala 122:59]
  wire [31:0] temp_raddr_intenable_base_match = ~_T_38; // @[pic_ctrl.scala 122:43]
  wire  raddr_intenable_base_match = &temp_raddr_intenable_base_match[31:7]; // @[pic_ctrl.scala 123:89]
  wire  raddr_intpriority_base_match = picm_raddr_ff[31:7] == 25'h1e01800; // @[pic_ctrl.scala 125:71]
  wire  raddr_config_gw_base_match = picm_raddr_ff[31:7] == 25'h1e01880; // @[pic_ctrl.scala 126:71]
  wire  raddr_config_pic_match = picm_raddr_ff == 32'hf00c3000; // @[pic_ctrl.scala 127:71]
  wire  addr_intpend_base_match = picm_raddr_ff[31:6] == 26'h3c03040; // @[pic_ctrl.scala 128:71]
  wire  waddr_config_pic_match = picm_waddr_ff == 32'hf00c3000; // @[pic_ctrl.scala 130:71]
  wire  waddr_intpriority_base_match = picm_waddr_ff[31:7] == 25'h1e01800; // @[pic_ctrl.scala 132:71]
  wire  waddr_config_gw_base_match = picm_waddr_ff[31:7] == 25'h1e01880; // @[pic_ctrl.scala 134:71]
  wire  _T_49 = picm_rden_ff & picm_wren_ff; // @[pic_ctrl.scala 135:53]
  wire  _T_50 = picm_raddr_ff == picm_waddr_ff; // @[pic_ctrl.scala 135:86]
  wire  picm_bypass_ff = _T_49 & _T_50; // @[pic_ctrl.scala 135:68]
  wire  _T_53 = raddr_intpriority_base_match & picm_rden_ff; // @[pic_ctrl.scala 141:108]
  wire  _T_56 = raddr_intenable_base_match & picm_rden_ff; // @[pic_ctrl.scala 142:104]
  wire  _T_59 = raddr_config_gw_base_match & picm_rden_ff; // @[pic_ctrl.scala 143:108]
  reg  _T_66; // @[Reg.scala 27:20]
  reg  extintsrc_req_sync_1; // @[Reg.scala 27:20]
  reg  _T_70; // @[Reg.scala 27:20]
  reg  extintsrc_req_sync_2; // @[Reg.scala 27:20]
  reg  _T_74; // @[Reg.scala 27:20]
  reg  extintsrc_req_sync_3; // @[Reg.scala 27:20]
  reg  _T_78; // @[Reg.scala 27:20]
  reg  extintsrc_req_sync_4; // @[Reg.scala 27:20]
  reg  _T_82; // @[Reg.scala 27:20]
  reg  extintsrc_req_sync_5; // @[Reg.scala 27:20]
  reg  _T_86; // @[Reg.scala 27:20]
  reg  extintsrc_req_sync_6; // @[Reg.scala 27:20]
  reg  _T_90; // @[Reg.scala 27:20]
  reg  extintsrc_req_sync_7; // @[Reg.scala 27:20]
  reg  _T_94; // @[Reg.scala 27:20]
  reg  extintsrc_req_sync_8; // @[Reg.scala 27:20]
  reg  _T_98; // @[Reg.scala 27:20]
  reg  extintsrc_req_sync_9; // @[Reg.scala 27:20]
  reg  _T_102; // @[Reg.scala 27:20]
  reg  extintsrc_req_sync_10; // @[Reg.scala 27:20]
  reg  _T_106; // @[Reg.scala 27:20]
  reg  extintsrc_req_sync_11; // @[Reg.scala 27:20]
  reg  _T_110; // @[Reg.scala 27:20]
  reg  extintsrc_req_sync_12; // @[Reg.scala 27:20]
  reg  _T_114; // @[Reg.scala 27:20]
  reg  extintsrc_req_sync_13; // @[Reg.scala 27:20]
  reg  _T_118; // @[Reg.scala 27:20]
  reg  extintsrc_req_sync_14; // @[Reg.scala 27:20]
  reg  _T_122; // @[Reg.scala 27:20]
  reg  extintsrc_req_sync_15; // @[Reg.scala 27:20]
  reg  _T_126; // @[Reg.scala 27:20]
  reg  extintsrc_req_sync_16; // @[Reg.scala 27:20]
  reg  _T_130; // @[Reg.scala 27:20]
  reg  extintsrc_req_sync_17; // @[Reg.scala 27:20]
  reg  _T_134; // @[Reg.scala 27:20]
  reg  extintsrc_req_sync_18; // @[Reg.scala 27:20]
  reg  _T_138; // @[Reg.scala 27:20]
  reg  extintsrc_req_sync_19; // @[Reg.scala 27:20]
  reg  _T_142; // @[Reg.scala 27:20]
  reg  extintsrc_req_sync_20; // @[Reg.scala 27:20]
  reg  _T_146; // @[Reg.scala 27:20]
  reg  extintsrc_req_sync_21; // @[Reg.scala 27:20]
  reg  _T_150; // @[Reg.scala 27:20]
  reg  extintsrc_req_sync_22; // @[Reg.scala 27:20]
  reg  _T_154; // @[Reg.scala 27:20]
  reg  extintsrc_req_sync_23; // @[Reg.scala 27:20]
  reg  _T_158; // @[Reg.scala 27:20]
  reg  extintsrc_req_sync_24; // @[Reg.scala 27:20]
  reg  _T_162; // @[Reg.scala 27:20]
  reg  extintsrc_req_sync_25; // @[Reg.scala 27:20]
  reg  _T_166; // @[Reg.scala 27:20]
  reg  extintsrc_req_sync_26; // @[Reg.scala 27:20]
  reg  _T_170; // @[Reg.scala 27:20]
  reg  extintsrc_req_sync_27; // @[Reg.scala 27:20]
  reg  _T_174; // @[Reg.scala 27:20]
  reg  extintsrc_req_sync_28; // @[Reg.scala 27:20]
  reg  _T_178; // @[Reg.scala 27:20]
  reg  extintsrc_req_sync_29; // @[Reg.scala 27:20]
  reg  _T_182; // @[Reg.scala 27:20]
  reg  extintsrc_req_sync_30; // @[Reg.scala 27:20]
  reg  _T_186; // @[Reg.scala 27:20]
  reg  extintsrc_req_sync_31; // @[Reg.scala 27:20]
  wire  _T_190 = waddr_intpriority_base_match & _T_375; // @[pic_ctrl.scala 156:106]
  wire  intpriority_reg_we_1 = _T_190 & picm_wren_ff; // @[pic_ctrl.scala 156:153]
  wire  _T_193 = waddr_intpriority_base_match & _T_378; // @[pic_ctrl.scala 156:106]
  wire  intpriority_reg_we_2 = _T_193 & picm_wren_ff; // @[pic_ctrl.scala 156:153]
  wire  _T_196 = waddr_intpriority_base_match & _T_381; // @[pic_ctrl.scala 156:106]
  wire  intpriority_reg_we_3 = _T_196 & picm_wren_ff; // @[pic_ctrl.scala 156:153]
  wire  _T_199 = waddr_intpriority_base_match & _T_384; // @[pic_ctrl.scala 156:106]
  wire  intpriority_reg_we_4 = _T_199 & picm_wren_ff; // @[pic_ctrl.scala 156:153]
  wire  _T_202 = waddr_intpriority_base_match & _T_387; // @[pic_ctrl.scala 156:106]
  wire  intpriority_reg_we_5 = _T_202 & picm_wren_ff; // @[pic_ctrl.scala 156:153]
  wire  _T_205 = waddr_intpriority_base_match & _T_390; // @[pic_ctrl.scala 156:106]
  wire  intpriority_reg_we_6 = _T_205 & picm_wren_ff; // @[pic_ctrl.scala 156:153]
  wire  _T_208 = waddr_intpriority_base_match & _T_393; // @[pic_ctrl.scala 156:106]
  wire  intpriority_reg_we_7 = _T_208 & picm_wren_ff; // @[pic_ctrl.scala 156:153]
  wire  _T_211 = waddr_intpriority_base_match & _T_396; // @[pic_ctrl.scala 156:106]
  wire  intpriority_reg_we_8 = _T_211 & picm_wren_ff; // @[pic_ctrl.scala 156:153]
  wire  _T_214 = waddr_intpriority_base_match & _T_399; // @[pic_ctrl.scala 156:106]
  wire  intpriority_reg_we_9 = _T_214 & picm_wren_ff; // @[pic_ctrl.scala 156:153]
  wire  _T_217 = waddr_intpriority_base_match & _T_402; // @[pic_ctrl.scala 156:106]
  wire  intpriority_reg_we_10 = _T_217 & picm_wren_ff; // @[pic_ctrl.scala 156:153]
  wire  _T_220 = waddr_intpriority_base_match & _T_405; // @[pic_ctrl.scala 156:106]
  wire  intpriority_reg_we_11 = _T_220 & picm_wren_ff; // @[pic_ctrl.scala 156:153]
  wire  _T_223 = waddr_intpriority_base_match & _T_408; // @[pic_ctrl.scala 156:106]
  wire  intpriority_reg_we_12 = _T_223 & picm_wren_ff; // @[pic_ctrl.scala 156:153]
  wire  _T_226 = waddr_intpriority_base_match & _T_411; // @[pic_ctrl.scala 156:106]
  wire  intpriority_reg_we_13 = _T_226 & picm_wren_ff; // @[pic_ctrl.scala 156:153]
  wire  _T_229 = waddr_intpriority_base_match & _T_414; // @[pic_ctrl.scala 156:106]
  wire  intpriority_reg_we_14 = _T_229 & picm_wren_ff; // @[pic_ctrl.scala 156:153]
  wire  _T_232 = waddr_intpriority_base_match & _T_417; // @[pic_ctrl.scala 156:106]
  wire  intpriority_reg_we_15 = _T_232 & picm_wren_ff; // @[pic_ctrl.scala 156:153]
  wire  _T_235 = waddr_intpriority_base_match & _T_420; // @[pic_ctrl.scala 156:106]
  wire  intpriority_reg_we_16 = _T_235 & picm_wren_ff; // @[pic_ctrl.scala 156:153]
  wire  _T_238 = waddr_intpriority_base_match & _T_423; // @[pic_ctrl.scala 156:106]
  wire  intpriority_reg_we_17 = _T_238 & picm_wren_ff; // @[pic_ctrl.scala 156:153]
  wire  _T_241 = waddr_intpriority_base_match & _T_426; // @[pic_ctrl.scala 156:106]
  wire  intpriority_reg_we_18 = _T_241 & picm_wren_ff; // @[pic_ctrl.scala 156:153]
  wire  _T_244 = waddr_intpriority_base_match & _T_429; // @[pic_ctrl.scala 156:106]
  wire  intpriority_reg_we_19 = _T_244 & picm_wren_ff; // @[pic_ctrl.scala 156:153]
  wire  _T_247 = waddr_intpriority_base_match & _T_432; // @[pic_ctrl.scala 156:106]
  wire  intpriority_reg_we_20 = _T_247 & picm_wren_ff; // @[pic_ctrl.scala 156:153]
  wire  _T_250 = waddr_intpriority_base_match & _T_435; // @[pic_ctrl.scala 156:106]
  wire  intpriority_reg_we_21 = _T_250 & picm_wren_ff; // @[pic_ctrl.scala 156:153]
  wire  _T_253 = waddr_intpriority_base_match & _T_438; // @[pic_ctrl.scala 156:106]
  wire  intpriority_reg_we_22 = _T_253 & picm_wren_ff; // @[pic_ctrl.scala 156:153]
  wire  _T_256 = waddr_intpriority_base_match & _T_441; // @[pic_ctrl.scala 156:106]
  wire  intpriority_reg_we_23 = _T_256 & picm_wren_ff; // @[pic_ctrl.scala 156:153]
  wire  _T_259 = waddr_intpriority_base_match & _T_444; // @[pic_ctrl.scala 156:106]
  wire  intpriority_reg_we_24 = _T_259 & picm_wren_ff; // @[pic_ctrl.scala 156:153]
  wire  _T_262 = waddr_intpriority_base_match & _T_447; // @[pic_ctrl.scala 156:106]
  wire  intpriority_reg_we_25 = _T_262 & picm_wren_ff; // @[pic_ctrl.scala 156:153]
  wire  _T_265 = waddr_intpriority_base_match & _T_450; // @[pic_ctrl.scala 156:106]
  wire  intpriority_reg_we_26 = _T_265 & picm_wren_ff; // @[pic_ctrl.scala 156:153]
  wire  _T_268 = waddr_intpriority_base_match & _T_453; // @[pic_ctrl.scala 156:106]
  wire  intpriority_reg_we_27 = _T_268 & picm_wren_ff; // @[pic_ctrl.scala 156:153]
  wire  _T_271 = waddr_intpriority_base_match & _T_456; // @[pic_ctrl.scala 156:106]
  wire  intpriority_reg_we_28 = _T_271 & picm_wren_ff; // @[pic_ctrl.scala 156:153]
  wire  _T_274 = waddr_intpriority_base_match & _T_459; // @[pic_ctrl.scala 156:106]
  wire  intpriority_reg_we_29 = _T_274 & picm_wren_ff; // @[pic_ctrl.scala 156:153]
  wire  _T_277 = waddr_intpriority_base_match & _T_462; // @[pic_ctrl.scala 156:106]
  wire  intpriority_reg_we_30 = _T_277 & picm_wren_ff; // @[pic_ctrl.scala 156:153]
  wire  _T_280 = waddr_intpriority_base_match & _T_465; // @[pic_ctrl.scala 156:106]
  wire  intpriority_reg_we_31 = _T_280 & picm_wren_ff; // @[pic_ctrl.scala 156:153]
  wire  _T_282 = picm_raddr_ff[6:2] == 5'h1; // @[pic_ctrl.scala 157:139]
  wire  _T_283 = raddr_intpriority_base_match & _T_282; // @[pic_ctrl.scala 157:106]
  wire  intpriority_reg_re_1 = _T_283 & picm_rden_ff; // @[pic_ctrl.scala 157:153]
  wire  _T_285 = picm_raddr_ff[6:2] == 5'h2; // @[pic_ctrl.scala 157:139]
  wire  _T_286 = raddr_intpriority_base_match & _T_285; // @[pic_ctrl.scala 157:106]
  wire  intpriority_reg_re_2 = _T_286 & picm_rden_ff; // @[pic_ctrl.scala 157:153]
  wire  _T_288 = picm_raddr_ff[6:2] == 5'h3; // @[pic_ctrl.scala 157:139]
  wire  _T_289 = raddr_intpriority_base_match & _T_288; // @[pic_ctrl.scala 157:106]
  wire  intpriority_reg_re_3 = _T_289 & picm_rden_ff; // @[pic_ctrl.scala 157:153]
  wire  _T_291 = picm_raddr_ff[6:2] == 5'h4; // @[pic_ctrl.scala 157:139]
  wire  _T_292 = raddr_intpriority_base_match & _T_291; // @[pic_ctrl.scala 157:106]
  wire  intpriority_reg_re_4 = _T_292 & picm_rden_ff; // @[pic_ctrl.scala 157:153]
  wire  _T_294 = picm_raddr_ff[6:2] == 5'h5; // @[pic_ctrl.scala 157:139]
  wire  _T_295 = raddr_intpriority_base_match & _T_294; // @[pic_ctrl.scala 157:106]
  wire  intpriority_reg_re_5 = _T_295 & picm_rden_ff; // @[pic_ctrl.scala 157:153]
  wire  _T_297 = picm_raddr_ff[6:2] == 5'h6; // @[pic_ctrl.scala 157:139]
  wire  _T_298 = raddr_intpriority_base_match & _T_297; // @[pic_ctrl.scala 157:106]
  wire  intpriority_reg_re_6 = _T_298 & picm_rden_ff; // @[pic_ctrl.scala 157:153]
  wire  _T_300 = picm_raddr_ff[6:2] == 5'h7; // @[pic_ctrl.scala 157:139]
  wire  _T_301 = raddr_intpriority_base_match & _T_300; // @[pic_ctrl.scala 157:106]
  wire  intpriority_reg_re_7 = _T_301 & picm_rden_ff; // @[pic_ctrl.scala 157:153]
  wire  _T_303 = picm_raddr_ff[6:2] == 5'h8; // @[pic_ctrl.scala 157:139]
  wire  _T_304 = raddr_intpriority_base_match & _T_303; // @[pic_ctrl.scala 157:106]
  wire  intpriority_reg_re_8 = _T_304 & picm_rden_ff; // @[pic_ctrl.scala 157:153]
  wire  _T_306 = picm_raddr_ff[6:2] == 5'h9; // @[pic_ctrl.scala 157:139]
  wire  _T_307 = raddr_intpriority_base_match & _T_306; // @[pic_ctrl.scala 157:106]
  wire  intpriority_reg_re_9 = _T_307 & picm_rden_ff; // @[pic_ctrl.scala 157:153]
  wire  _T_309 = picm_raddr_ff[6:2] == 5'ha; // @[pic_ctrl.scala 157:139]
  wire  _T_310 = raddr_intpriority_base_match & _T_309; // @[pic_ctrl.scala 157:106]
  wire  intpriority_reg_re_10 = _T_310 & picm_rden_ff; // @[pic_ctrl.scala 157:153]
  wire  _T_312 = picm_raddr_ff[6:2] == 5'hb; // @[pic_ctrl.scala 157:139]
  wire  _T_313 = raddr_intpriority_base_match & _T_312; // @[pic_ctrl.scala 157:106]
  wire  intpriority_reg_re_11 = _T_313 & picm_rden_ff; // @[pic_ctrl.scala 157:153]
  wire  _T_315 = picm_raddr_ff[6:2] == 5'hc; // @[pic_ctrl.scala 157:139]
  wire  _T_316 = raddr_intpriority_base_match & _T_315; // @[pic_ctrl.scala 157:106]
  wire  intpriority_reg_re_12 = _T_316 & picm_rden_ff; // @[pic_ctrl.scala 157:153]
  wire  _T_318 = picm_raddr_ff[6:2] == 5'hd; // @[pic_ctrl.scala 157:139]
  wire  _T_319 = raddr_intpriority_base_match & _T_318; // @[pic_ctrl.scala 157:106]
  wire  intpriority_reg_re_13 = _T_319 & picm_rden_ff; // @[pic_ctrl.scala 157:153]
  wire  _T_321 = picm_raddr_ff[6:2] == 5'he; // @[pic_ctrl.scala 157:139]
  wire  _T_322 = raddr_intpriority_base_match & _T_321; // @[pic_ctrl.scala 157:106]
  wire  intpriority_reg_re_14 = _T_322 & picm_rden_ff; // @[pic_ctrl.scala 157:153]
  wire  _T_324 = picm_raddr_ff[6:2] == 5'hf; // @[pic_ctrl.scala 157:139]
  wire  _T_325 = raddr_intpriority_base_match & _T_324; // @[pic_ctrl.scala 157:106]
  wire  intpriority_reg_re_15 = _T_325 & picm_rden_ff; // @[pic_ctrl.scala 157:153]
  wire  _T_327 = picm_raddr_ff[6:2] == 5'h10; // @[pic_ctrl.scala 157:139]
  wire  _T_328 = raddr_intpriority_base_match & _T_327; // @[pic_ctrl.scala 157:106]
  wire  intpriority_reg_re_16 = _T_328 & picm_rden_ff; // @[pic_ctrl.scala 157:153]
  wire  _T_330 = picm_raddr_ff[6:2] == 5'h11; // @[pic_ctrl.scala 157:139]
  wire  _T_331 = raddr_intpriority_base_match & _T_330; // @[pic_ctrl.scala 157:106]
  wire  intpriority_reg_re_17 = _T_331 & picm_rden_ff; // @[pic_ctrl.scala 157:153]
  wire  _T_333 = picm_raddr_ff[6:2] == 5'h12; // @[pic_ctrl.scala 157:139]
  wire  _T_334 = raddr_intpriority_base_match & _T_333; // @[pic_ctrl.scala 157:106]
  wire  intpriority_reg_re_18 = _T_334 & picm_rden_ff; // @[pic_ctrl.scala 157:153]
  wire  _T_336 = picm_raddr_ff[6:2] == 5'h13; // @[pic_ctrl.scala 157:139]
  wire  _T_337 = raddr_intpriority_base_match & _T_336; // @[pic_ctrl.scala 157:106]
  wire  intpriority_reg_re_19 = _T_337 & picm_rden_ff; // @[pic_ctrl.scala 157:153]
  wire  _T_339 = picm_raddr_ff[6:2] == 5'h14; // @[pic_ctrl.scala 157:139]
  wire  _T_340 = raddr_intpriority_base_match & _T_339; // @[pic_ctrl.scala 157:106]
  wire  intpriority_reg_re_20 = _T_340 & picm_rden_ff; // @[pic_ctrl.scala 157:153]
  wire  _T_342 = picm_raddr_ff[6:2] == 5'h15; // @[pic_ctrl.scala 157:139]
  wire  _T_343 = raddr_intpriority_base_match & _T_342; // @[pic_ctrl.scala 157:106]
  wire  intpriority_reg_re_21 = _T_343 & picm_rden_ff; // @[pic_ctrl.scala 157:153]
  wire  _T_345 = picm_raddr_ff[6:2] == 5'h16; // @[pic_ctrl.scala 157:139]
  wire  _T_346 = raddr_intpriority_base_match & _T_345; // @[pic_ctrl.scala 157:106]
  wire  intpriority_reg_re_22 = _T_346 & picm_rden_ff; // @[pic_ctrl.scala 157:153]
  wire  _T_348 = picm_raddr_ff[6:2] == 5'h17; // @[pic_ctrl.scala 157:139]
  wire  _T_349 = raddr_intpriority_base_match & _T_348; // @[pic_ctrl.scala 157:106]
  wire  intpriority_reg_re_23 = _T_349 & picm_rden_ff; // @[pic_ctrl.scala 157:153]
  wire  _T_351 = picm_raddr_ff[6:2] == 5'h18; // @[pic_ctrl.scala 157:139]
  wire  _T_352 = raddr_intpriority_base_match & _T_351; // @[pic_ctrl.scala 157:106]
  wire  intpriority_reg_re_24 = _T_352 & picm_rden_ff; // @[pic_ctrl.scala 157:153]
  wire  _T_354 = picm_raddr_ff[6:2] == 5'h19; // @[pic_ctrl.scala 157:139]
  wire  _T_355 = raddr_intpriority_base_match & _T_354; // @[pic_ctrl.scala 157:106]
  wire  intpriority_reg_re_25 = _T_355 & picm_rden_ff; // @[pic_ctrl.scala 157:153]
  wire  _T_357 = picm_raddr_ff[6:2] == 5'h1a; // @[pic_ctrl.scala 157:139]
  wire  _T_358 = raddr_intpriority_base_match & _T_357; // @[pic_ctrl.scala 157:106]
  wire  intpriority_reg_re_26 = _T_358 & picm_rden_ff; // @[pic_ctrl.scala 157:153]
  wire  _T_360 = picm_raddr_ff[6:2] == 5'h1b; // @[pic_ctrl.scala 157:139]
  wire  _T_361 = raddr_intpriority_base_match & _T_360; // @[pic_ctrl.scala 157:106]
  wire  intpriority_reg_re_27 = _T_361 & picm_rden_ff; // @[pic_ctrl.scala 157:153]
  wire  _T_363 = picm_raddr_ff[6:2] == 5'h1c; // @[pic_ctrl.scala 157:139]
  wire  _T_364 = raddr_intpriority_base_match & _T_363; // @[pic_ctrl.scala 157:106]
  wire  intpriority_reg_re_28 = _T_364 & picm_rden_ff; // @[pic_ctrl.scala 157:153]
  wire  _T_366 = picm_raddr_ff[6:2] == 5'h1d; // @[pic_ctrl.scala 157:139]
  wire  _T_367 = raddr_intpriority_base_match & _T_366; // @[pic_ctrl.scala 157:106]
  wire  intpriority_reg_re_29 = _T_367 & picm_rden_ff; // @[pic_ctrl.scala 157:153]
  wire  _T_369 = picm_raddr_ff[6:2] == 5'h1e; // @[pic_ctrl.scala 157:139]
  wire  _T_370 = raddr_intpriority_base_match & _T_369; // @[pic_ctrl.scala 157:106]
  wire  intpriority_reg_re_30 = _T_370 & picm_rden_ff; // @[pic_ctrl.scala 157:153]
  wire  _T_372 = picm_raddr_ff[6:2] == 5'h1f; // @[pic_ctrl.scala 157:139]
  wire  _T_373 = raddr_intpriority_base_match & _T_372; // @[pic_ctrl.scala 157:106]
  wire  intpriority_reg_re_31 = _T_373 & picm_rden_ff; // @[pic_ctrl.scala 157:153]
  wire  _T_469 = raddr_intenable_base_match & _T_282; // @[pic_ctrl.scala 159:106]
  wire  intenable_reg_re_1 = _T_469 & picm_rden_ff; // @[pic_ctrl.scala 159:153]
  wire  _T_472 = raddr_intenable_base_match & _T_285; // @[pic_ctrl.scala 159:106]
  wire  intenable_reg_re_2 = _T_472 & picm_rden_ff; // @[pic_ctrl.scala 159:153]
  wire  _T_475 = raddr_intenable_base_match & _T_288; // @[pic_ctrl.scala 159:106]
  wire  intenable_reg_re_3 = _T_475 & picm_rden_ff; // @[pic_ctrl.scala 159:153]
  wire  _T_478 = raddr_intenable_base_match & _T_291; // @[pic_ctrl.scala 159:106]
  wire  intenable_reg_re_4 = _T_478 & picm_rden_ff; // @[pic_ctrl.scala 159:153]
  wire  _T_481 = raddr_intenable_base_match & _T_294; // @[pic_ctrl.scala 159:106]
  wire  intenable_reg_re_5 = _T_481 & picm_rden_ff; // @[pic_ctrl.scala 159:153]
  wire  _T_484 = raddr_intenable_base_match & _T_297; // @[pic_ctrl.scala 159:106]
  wire  intenable_reg_re_6 = _T_484 & picm_rden_ff; // @[pic_ctrl.scala 159:153]
  wire  _T_487 = raddr_intenable_base_match & _T_300; // @[pic_ctrl.scala 159:106]
  wire  intenable_reg_re_7 = _T_487 & picm_rden_ff; // @[pic_ctrl.scala 159:153]
  wire  _T_490 = raddr_intenable_base_match & _T_303; // @[pic_ctrl.scala 159:106]
  wire  intenable_reg_re_8 = _T_490 & picm_rden_ff; // @[pic_ctrl.scala 159:153]
  wire  _T_493 = raddr_intenable_base_match & _T_306; // @[pic_ctrl.scala 159:106]
  wire  intenable_reg_re_9 = _T_493 & picm_rden_ff; // @[pic_ctrl.scala 159:153]
  wire  _T_496 = raddr_intenable_base_match & _T_309; // @[pic_ctrl.scala 159:106]
  wire  intenable_reg_re_10 = _T_496 & picm_rden_ff; // @[pic_ctrl.scala 159:153]
  wire  _T_499 = raddr_intenable_base_match & _T_312; // @[pic_ctrl.scala 159:106]
  wire  intenable_reg_re_11 = _T_499 & picm_rden_ff; // @[pic_ctrl.scala 159:153]
  wire  _T_502 = raddr_intenable_base_match & _T_315; // @[pic_ctrl.scala 159:106]
  wire  intenable_reg_re_12 = _T_502 & picm_rden_ff; // @[pic_ctrl.scala 159:153]
  wire  _T_505 = raddr_intenable_base_match & _T_318; // @[pic_ctrl.scala 159:106]
  wire  intenable_reg_re_13 = _T_505 & picm_rden_ff; // @[pic_ctrl.scala 159:153]
  wire  _T_508 = raddr_intenable_base_match & _T_321; // @[pic_ctrl.scala 159:106]
  wire  intenable_reg_re_14 = _T_508 & picm_rden_ff; // @[pic_ctrl.scala 159:153]
  wire  _T_511 = raddr_intenable_base_match & _T_324; // @[pic_ctrl.scala 159:106]
  wire  intenable_reg_re_15 = _T_511 & picm_rden_ff; // @[pic_ctrl.scala 159:153]
  wire  _T_514 = raddr_intenable_base_match & _T_327; // @[pic_ctrl.scala 159:106]
  wire  intenable_reg_re_16 = _T_514 & picm_rden_ff; // @[pic_ctrl.scala 159:153]
  wire  _T_517 = raddr_intenable_base_match & _T_330; // @[pic_ctrl.scala 159:106]
  wire  intenable_reg_re_17 = _T_517 & picm_rden_ff; // @[pic_ctrl.scala 159:153]
  wire  _T_520 = raddr_intenable_base_match & _T_333; // @[pic_ctrl.scala 159:106]
  wire  intenable_reg_re_18 = _T_520 & picm_rden_ff; // @[pic_ctrl.scala 159:153]
  wire  _T_523 = raddr_intenable_base_match & _T_336; // @[pic_ctrl.scala 159:106]
  wire  intenable_reg_re_19 = _T_523 & picm_rden_ff; // @[pic_ctrl.scala 159:153]
  wire  _T_526 = raddr_intenable_base_match & _T_339; // @[pic_ctrl.scala 159:106]
  wire  intenable_reg_re_20 = _T_526 & picm_rden_ff; // @[pic_ctrl.scala 159:153]
  wire  _T_529 = raddr_intenable_base_match & _T_342; // @[pic_ctrl.scala 159:106]
  wire  intenable_reg_re_21 = _T_529 & picm_rden_ff; // @[pic_ctrl.scala 159:153]
  wire  _T_532 = raddr_intenable_base_match & _T_345; // @[pic_ctrl.scala 159:106]
  wire  intenable_reg_re_22 = _T_532 & picm_rden_ff; // @[pic_ctrl.scala 159:153]
  wire  _T_535 = raddr_intenable_base_match & _T_348; // @[pic_ctrl.scala 159:106]
  wire  intenable_reg_re_23 = _T_535 & picm_rden_ff; // @[pic_ctrl.scala 159:153]
  wire  _T_538 = raddr_intenable_base_match & _T_351; // @[pic_ctrl.scala 159:106]
  wire  intenable_reg_re_24 = _T_538 & picm_rden_ff; // @[pic_ctrl.scala 159:153]
  wire  _T_541 = raddr_intenable_base_match & _T_354; // @[pic_ctrl.scala 159:106]
  wire  intenable_reg_re_25 = _T_541 & picm_rden_ff; // @[pic_ctrl.scala 159:153]
  wire  _T_544 = raddr_intenable_base_match & _T_357; // @[pic_ctrl.scala 159:106]
  wire  intenable_reg_re_26 = _T_544 & picm_rden_ff; // @[pic_ctrl.scala 159:153]
  wire  _T_547 = raddr_intenable_base_match & _T_360; // @[pic_ctrl.scala 159:106]
  wire  intenable_reg_re_27 = _T_547 & picm_rden_ff; // @[pic_ctrl.scala 159:153]
  wire  _T_550 = raddr_intenable_base_match & _T_363; // @[pic_ctrl.scala 159:106]
  wire  intenable_reg_re_28 = _T_550 & picm_rden_ff; // @[pic_ctrl.scala 159:153]
  wire  _T_553 = raddr_intenable_base_match & _T_366; // @[pic_ctrl.scala 159:106]
  wire  intenable_reg_re_29 = _T_553 & picm_rden_ff; // @[pic_ctrl.scala 159:153]
  wire  _T_556 = raddr_intenable_base_match & _T_369; // @[pic_ctrl.scala 159:106]
  wire  intenable_reg_re_30 = _T_556 & picm_rden_ff; // @[pic_ctrl.scala 159:153]
  wire  _T_559 = raddr_intenable_base_match & _T_372; // @[pic_ctrl.scala 159:106]
  wire  intenable_reg_re_31 = _T_559 & picm_rden_ff; // @[pic_ctrl.scala 159:153]
  wire  _T_562 = waddr_config_gw_base_match & _T_375; // @[pic_ctrl.scala 160:106]
  wire  gw_config_reg_we_1 = _T_562 & picm_wren_ff; // @[pic_ctrl.scala 160:153]
  wire  _T_565 = waddr_config_gw_base_match & _T_378; // @[pic_ctrl.scala 160:106]
  wire  gw_config_reg_we_2 = _T_565 & picm_wren_ff; // @[pic_ctrl.scala 160:153]
  wire  _T_568 = waddr_config_gw_base_match & _T_381; // @[pic_ctrl.scala 160:106]
  wire  gw_config_reg_we_3 = _T_568 & picm_wren_ff; // @[pic_ctrl.scala 160:153]
  wire  _T_571 = waddr_config_gw_base_match & _T_384; // @[pic_ctrl.scala 160:106]
  wire  gw_config_reg_we_4 = _T_571 & picm_wren_ff; // @[pic_ctrl.scala 160:153]
  wire  _T_574 = waddr_config_gw_base_match & _T_387; // @[pic_ctrl.scala 160:106]
  wire  gw_config_reg_we_5 = _T_574 & picm_wren_ff; // @[pic_ctrl.scala 160:153]
  wire  _T_577 = waddr_config_gw_base_match & _T_390; // @[pic_ctrl.scala 160:106]
  wire  gw_config_reg_we_6 = _T_577 & picm_wren_ff; // @[pic_ctrl.scala 160:153]
  wire  _T_580 = waddr_config_gw_base_match & _T_393; // @[pic_ctrl.scala 160:106]
  wire  gw_config_reg_we_7 = _T_580 & picm_wren_ff; // @[pic_ctrl.scala 160:153]
  wire  _T_583 = waddr_config_gw_base_match & _T_396; // @[pic_ctrl.scala 160:106]
  wire  gw_config_reg_we_8 = _T_583 & picm_wren_ff; // @[pic_ctrl.scala 160:153]
  wire  _T_586 = waddr_config_gw_base_match & _T_399; // @[pic_ctrl.scala 160:106]
  wire  gw_config_reg_we_9 = _T_586 & picm_wren_ff; // @[pic_ctrl.scala 160:153]
  wire  _T_589 = waddr_config_gw_base_match & _T_402; // @[pic_ctrl.scala 160:106]
  wire  gw_config_reg_we_10 = _T_589 & picm_wren_ff; // @[pic_ctrl.scala 160:153]
  wire  _T_592 = waddr_config_gw_base_match & _T_405; // @[pic_ctrl.scala 160:106]
  wire  gw_config_reg_we_11 = _T_592 & picm_wren_ff; // @[pic_ctrl.scala 160:153]
  wire  _T_595 = waddr_config_gw_base_match & _T_408; // @[pic_ctrl.scala 160:106]
  wire  gw_config_reg_we_12 = _T_595 & picm_wren_ff; // @[pic_ctrl.scala 160:153]
  wire  _T_598 = waddr_config_gw_base_match & _T_411; // @[pic_ctrl.scala 160:106]
  wire  gw_config_reg_we_13 = _T_598 & picm_wren_ff; // @[pic_ctrl.scala 160:153]
  wire  _T_601 = waddr_config_gw_base_match & _T_414; // @[pic_ctrl.scala 160:106]
  wire  gw_config_reg_we_14 = _T_601 & picm_wren_ff; // @[pic_ctrl.scala 160:153]
  wire  _T_604 = waddr_config_gw_base_match & _T_417; // @[pic_ctrl.scala 160:106]
  wire  gw_config_reg_we_15 = _T_604 & picm_wren_ff; // @[pic_ctrl.scala 160:153]
  wire  _T_607 = waddr_config_gw_base_match & _T_420; // @[pic_ctrl.scala 160:106]
  wire  gw_config_reg_we_16 = _T_607 & picm_wren_ff; // @[pic_ctrl.scala 160:153]
  wire  _T_610 = waddr_config_gw_base_match & _T_423; // @[pic_ctrl.scala 160:106]
  wire  gw_config_reg_we_17 = _T_610 & picm_wren_ff; // @[pic_ctrl.scala 160:153]
  wire  _T_613 = waddr_config_gw_base_match & _T_426; // @[pic_ctrl.scala 160:106]
  wire  gw_config_reg_we_18 = _T_613 & picm_wren_ff; // @[pic_ctrl.scala 160:153]
  wire  _T_616 = waddr_config_gw_base_match & _T_429; // @[pic_ctrl.scala 160:106]
  wire  gw_config_reg_we_19 = _T_616 & picm_wren_ff; // @[pic_ctrl.scala 160:153]
  wire  _T_619 = waddr_config_gw_base_match & _T_432; // @[pic_ctrl.scala 160:106]
  wire  gw_config_reg_we_20 = _T_619 & picm_wren_ff; // @[pic_ctrl.scala 160:153]
  wire  _T_622 = waddr_config_gw_base_match & _T_435; // @[pic_ctrl.scala 160:106]
  wire  gw_config_reg_we_21 = _T_622 & picm_wren_ff; // @[pic_ctrl.scala 160:153]
  wire  _T_625 = waddr_config_gw_base_match & _T_438; // @[pic_ctrl.scala 160:106]
  wire  gw_config_reg_we_22 = _T_625 & picm_wren_ff; // @[pic_ctrl.scala 160:153]
  wire  _T_628 = waddr_config_gw_base_match & _T_441; // @[pic_ctrl.scala 160:106]
  wire  gw_config_reg_we_23 = _T_628 & picm_wren_ff; // @[pic_ctrl.scala 160:153]
  wire  _T_631 = waddr_config_gw_base_match & _T_444; // @[pic_ctrl.scala 160:106]
  wire  gw_config_reg_we_24 = _T_631 & picm_wren_ff; // @[pic_ctrl.scala 160:153]
  wire  _T_634 = waddr_config_gw_base_match & _T_447; // @[pic_ctrl.scala 160:106]
  wire  gw_config_reg_we_25 = _T_634 & picm_wren_ff; // @[pic_ctrl.scala 160:153]
  wire  _T_637 = waddr_config_gw_base_match & _T_450; // @[pic_ctrl.scala 160:106]
  wire  gw_config_reg_we_26 = _T_637 & picm_wren_ff; // @[pic_ctrl.scala 160:153]
  wire  _T_640 = waddr_config_gw_base_match & _T_453; // @[pic_ctrl.scala 160:106]
  wire  gw_config_reg_we_27 = _T_640 & picm_wren_ff; // @[pic_ctrl.scala 160:153]
  wire  _T_643 = waddr_config_gw_base_match & _T_456; // @[pic_ctrl.scala 160:106]
  wire  gw_config_reg_we_28 = _T_643 & picm_wren_ff; // @[pic_ctrl.scala 160:153]
  wire  _T_646 = waddr_config_gw_base_match & _T_459; // @[pic_ctrl.scala 160:106]
  wire  gw_config_reg_we_29 = _T_646 & picm_wren_ff; // @[pic_ctrl.scala 160:153]
  wire  _T_649 = waddr_config_gw_base_match & _T_462; // @[pic_ctrl.scala 160:106]
  wire  gw_config_reg_we_30 = _T_649 & picm_wren_ff; // @[pic_ctrl.scala 160:153]
  wire  _T_652 = waddr_config_gw_base_match & _T_465; // @[pic_ctrl.scala 160:106]
  wire  gw_config_reg_we_31 = _T_652 & picm_wren_ff; // @[pic_ctrl.scala 160:153]
  wire  _T_655 = raddr_config_gw_base_match & _T_282; // @[pic_ctrl.scala 161:106]
  wire  gw_config_reg_re_1 = _T_655 & picm_rden_ff; // @[pic_ctrl.scala 161:153]
  wire  _T_658 = raddr_config_gw_base_match & _T_285; // @[pic_ctrl.scala 161:106]
  wire  gw_config_reg_re_2 = _T_658 & picm_rden_ff; // @[pic_ctrl.scala 161:153]
  wire  _T_661 = raddr_config_gw_base_match & _T_288; // @[pic_ctrl.scala 161:106]
  wire  gw_config_reg_re_3 = _T_661 & picm_rden_ff; // @[pic_ctrl.scala 161:153]
  wire  _T_664 = raddr_config_gw_base_match & _T_291; // @[pic_ctrl.scala 161:106]
  wire  gw_config_reg_re_4 = _T_664 & picm_rden_ff; // @[pic_ctrl.scala 161:153]
  wire  _T_667 = raddr_config_gw_base_match & _T_294; // @[pic_ctrl.scala 161:106]
  wire  gw_config_reg_re_5 = _T_667 & picm_rden_ff; // @[pic_ctrl.scala 161:153]
  wire  _T_670 = raddr_config_gw_base_match & _T_297; // @[pic_ctrl.scala 161:106]
  wire  gw_config_reg_re_6 = _T_670 & picm_rden_ff; // @[pic_ctrl.scala 161:153]
  wire  _T_673 = raddr_config_gw_base_match & _T_300; // @[pic_ctrl.scala 161:106]
  wire  gw_config_reg_re_7 = _T_673 & picm_rden_ff; // @[pic_ctrl.scala 161:153]
  wire  _T_676 = raddr_config_gw_base_match & _T_303; // @[pic_ctrl.scala 161:106]
  wire  gw_config_reg_re_8 = _T_676 & picm_rden_ff; // @[pic_ctrl.scala 161:153]
  wire  _T_679 = raddr_config_gw_base_match & _T_306; // @[pic_ctrl.scala 161:106]
  wire  gw_config_reg_re_9 = _T_679 & picm_rden_ff; // @[pic_ctrl.scala 161:153]
  wire  _T_682 = raddr_config_gw_base_match & _T_309; // @[pic_ctrl.scala 161:106]
  wire  gw_config_reg_re_10 = _T_682 & picm_rden_ff; // @[pic_ctrl.scala 161:153]
  wire  _T_685 = raddr_config_gw_base_match & _T_312; // @[pic_ctrl.scala 161:106]
  wire  gw_config_reg_re_11 = _T_685 & picm_rden_ff; // @[pic_ctrl.scala 161:153]
  wire  _T_688 = raddr_config_gw_base_match & _T_315; // @[pic_ctrl.scala 161:106]
  wire  gw_config_reg_re_12 = _T_688 & picm_rden_ff; // @[pic_ctrl.scala 161:153]
  wire  _T_691 = raddr_config_gw_base_match & _T_318; // @[pic_ctrl.scala 161:106]
  wire  gw_config_reg_re_13 = _T_691 & picm_rden_ff; // @[pic_ctrl.scala 161:153]
  wire  _T_694 = raddr_config_gw_base_match & _T_321; // @[pic_ctrl.scala 161:106]
  wire  gw_config_reg_re_14 = _T_694 & picm_rden_ff; // @[pic_ctrl.scala 161:153]
  wire  _T_697 = raddr_config_gw_base_match & _T_324; // @[pic_ctrl.scala 161:106]
  wire  gw_config_reg_re_15 = _T_697 & picm_rden_ff; // @[pic_ctrl.scala 161:153]
  wire  _T_700 = raddr_config_gw_base_match & _T_327; // @[pic_ctrl.scala 161:106]
  wire  gw_config_reg_re_16 = _T_700 & picm_rden_ff; // @[pic_ctrl.scala 161:153]
  wire  _T_703 = raddr_config_gw_base_match & _T_330; // @[pic_ctrl.scala 161:106]
  wire  gw_config_reg_re_17 = _T_703 & picm_rden_ff; // @[pic_ctrl.scala 161:153]
  wire  _T_706 = raddr_config_gw_base_match & _T_333; // @[pic_ctrl.scala 161:106]
  wire  gw_config_reg_re_18 = _T_706 & picm_rden_ff; // @[pic_ctrl.scala 161:153]
  wire  _T_709 = raddr_config_gw_base_match & _T_336; // @[pic_ctrl.scala 161:106]
  wire  gw_config_reg_re_19 = _T_709 & picm_rden_ff; // @[pic_ctrl.scala 161:153]
  wire  _T_712 = raddr_config_gw_base_match & _T_339; // @[pic_ctrl.scala 161:106]
  wire  gw_config_reg_re_20 = _T_712 & picm_rden_ff; // @[pic_ctrl.scala 161:153]
  wire  _T_715 = raddr_config_gw_base_match & _T_342; // @[pic_ctrl.scala 161:106]
  wire  gw_config_reg_re_21 = _T_715 & picm_rden_ff; // @[pic_ctrl.scala 161:153]
  wire  _T_718 = raddr_config_gw_base_match & _T_345; // @[pic_ctrl.scala 161:106]
  wire  gw_config_reg_re_22 = _T_718 & picm_rden_ff; // @[pic_ctrl.scala 161:153]
  wire  _T_721 = raddr_config_gw_base_match & _T_348; // @[pic_ctrl.scala 161:106]
  wire  gw_config_reg_re_23 = _T_721 & picm_rden_ff; // @[pic_ctrl.scala 161:153]
  wire  _T_724 = raddr_config_gw_base_match & _T_351; // @[pic_ctrl.scala 161:106]
  wire  gw_config_reg_re_24 = _T_724 & picm_rden_ff; // @[pic_ctrl.scala 161:153]
  wire  _T_727 = raddr_config_gw_base_match & _T_354; // @[pic_ctrl.scala 161:106]
  wire  gw_config_reg_re_25 = _T_727 & picm_rden_ff; // @[pic_ctrl.scala 161:153]
  wire  _T_730 = raddr_config_gw_base_match & _T_357; // @[pic_ctrl.scala 161:106]
  wire  gw_config_reg_re_26 = _T_730 & picm_rden_ff; // @[pic_ctrl.scala 161:153]
  wire  _T_733 = raddr_config_gw_base_match & _T_360; // @[pic_ctrl.scala 161:106]
  wire  gw_config_reg_re_27 = _T_733 & picm_rden_ff; // @[pic_ctrl.scala 161:153]
  wire  _T_736 = raddr_config_gw_base_match & _T_363; // @[pic_ctrl.scala 161:106]
  wire  gw_config_reg_re_28 = _T_736 & picm_rden_ff; // @[pic_ctrl.scala 161:153]
  wire  _T_739 = raddr_config_gw_base_match & _T_366; // @[pic_ctrl.scala 161:106]
  wire  gw_config_reg_re_29 = _T_739 & picm_rden_ff; // @[pic_ctrl.scala 161:153]
  wire  _T_742 = raddr_config_gw_base_match & _T_369; // @[pic_ctrl.scala 161:106]
  wire  gw_config_reg_re_30 = _T_742 & picm_rden_ff; // @[pic_ctrl.scala 161:153]
  wire  _T_745 = raddr_config_gw_base_match & _T_372; // @[pic_ctrl.scala 161:106]
  wire  gw_config_reg_re_31 = _T_745 & picm_rden_ff; // @[pic_ctrl.scala 161:153]
  reg [3:0] intpriority_reg_1; // @[Reg.scala 27:20]
  reg [3:0] intpriority_reg_2; // @[Reg.scala 27:20]
  reg [3:0] intpriority_reg_3; // @[Reg.scala 27:20]
  reg [3:0] intpriority_reg_4; // @[Reg.scala 27:20]
  reg [3:0] intpriority_reg_5; // @[Reg.scala 27:20]
  reg [3:0] intpriority_reg_6; // @[Reg.scala 27:20]
  reg [3:0] intpriority_reg_7; // @[Reg.scala 27:20]
  reg [3:0] intpriority_reg_8; // @[Reg.scala 27:20]
  reg [3:0] intpriority_reg_9; // @[Reg.scala 27:20]
  reg [3:0] intpriority_reg_10; // @[Reg.scala 27:20]
  reg [3:0] intpriority_reg_11; // @[Reg.scala 27:20]
  reg [3:0] intpriority_reg_12; // @[Reg.scala 27:20]
  reg [3:0] intpriority_reg_13; // @[Reg.scala 27:20]
  reg [3:0] intpriority_reg_14; // @[Reg.scala 27:20]
  reg [3:0] intpriority_reg_15; // @[Reg.scala 27:20]
  reg [3:0] intpriority_reg_16; // @[Reg.scala 27:20]
  reg [3:0] intpriority_reg_17; // @[Reg.scala 27:20]
  reg [3:0] intpriority_reg_18; // @[Reg.scala 27:20]
  reg [3:0] intpriority_reg_19; // @[Reg.scala 27:20]
  reg [3:0] intpriority_reg_20; // @[Reg.scala 27:20]
  reg [3:0] intpriority_reg_21; // @[Reg.scala 27:20]
  reg [3:0] intpriority_reg_22; // @[Reg.scala 27:20]
  reg [3:0] intpriority_reg_23; // @[Reg.scala 27:20]
  reg [3:0] intpriority_reg_24; // @[Reg.scala 27:20]
  reg [3:0] intpriority_reg_25; // @[Reg.scala 27:20]
  reg [3:0] intpriority_reg_26; // @[Reg.scala 27:20]
  reg [3:0] intpriority_reg_27; // @[Reg.scala 27:20]
  reg [3:0] intpriority_reg_28; // @[Reg.scala 27:20]
  reg [3:0] intpriority_reg_29; // @[Reg.scala 27:20]
  reg [3:0] intpriority_reg_30; // @[Reg.scala 27:20]
  reg [3:0] intpriority_reg_31; // @[Reg.scala 27:20]
  wire  _T_1279 = extintsrc_req_sync_1 ^ gw_config_reg_1[0]; // @[lib.scala 117:50]
  wire  _T_1280 = ~gw_clear_reg_we_1; // @[lib.scala 117:92]
  reg  _T_1283; // @[Reg.scala 27:20]
  wire  _T_1281 = _T_1283 & _T_1280; // @[lib.scala 117:90]
  wire  _T_1282 = _T_1279 | _T_1281; // @[lib.scala 117:72]
  wire  _T_1286 = _T_1279 | _T_1283; // @[lib.scala 119:78]
  wire  extintsrc_req_gw_1 = gw_config_reg_1[1] ? _T_1286 : _T_1279; // @[lib.scala 119:8]
  wire  _T_1294 = extintsrc_req_sync_2 ^ gw_config_reg_2[0]; // @[lib.scala 117:50]
  wire  _T_1295 = ~gw_clear_reg_we_2; // @[lib.scala 117:92]
  reg  _T_1298; // @[Reg.scala 27:20]
  wire  _T_1296 = _T_1298 & _T_1295; // @[lib.scala 117:90]
  wire  _T_1297 = _T_1294 | _T_1296; // @[lib.scala 117:72]
  wire  _T_1301 = _T_1294 | _T_1298; // @[lib.scala 119:78]
  wire  extintsrc_req_gw_2 = gw_config_reg_2[1] ? _T_1301 : _T_1294; // @[lib.scala 119:8]
  wire  _T_1309 = extintsrc_req_sync_3 ^ gw_config_reg_3[0]; // @[lib.scala 117:50]
  wire  _T_1310 = ~gw_clear_reg_we_3; // @[lib.scala 117:92]
  reg  _T_1313; // @[Reg.scala 27:20]
  wire  _T_1311 = _T_1313 & _T_1310; // @[lib.scala 117:90]
  wire  _T_1312 = _T_1309 | _T_1311; // @[lib.scala 117:72]
  wire  _T_1316 = _T_1309 | _T_1313; // @[lib.scala 119:78]
  wire  extintsrc_req_gw_3 = gw_config_reg_3[1] ? _T_1316 : _T_1309; // @[lib.scala 119:8]
  wire  _T_1324 = extintsrc_req_sync_4 ^ gw_config_reg_4[0]; // @[lib.scala 117:50]
  wire  _T_1325 = ~gw_clear_reg_we_4; // @[lib.scala 117:92]
  reg  _T_1328; // @[Reg.scala 27:20]
  wire  _T_1326 = _T_1328 & _T_1325; // @[lib.scala 117:90]
  wire  _T_1327 = _T_1324 | _T_1326; // @[lib.scala 117:72]
  wire  _T_1331 = _T_1324 | _T_1328; // @[lib.scala 119:78]
  wire  extintsrc_req_gw_4 = gw_config_reg_4[1] ? _T_1331 : _T_1324; // @[lib.scala 119:8]
  wire  _T_1339 = extintsrc_req_sync_5 ^ gw_config_reg_5[0]; // @[lib.scala 117:50]
  wire  _T_1340 = ~gw_clear_reg_we_5; // @[lib.scala 117:92]
  reg  _T_1343; // @[Reg.scala 27:20]
  wire  _T_1341 = _T_1343 & _T_1340; // @[lib.scala 117:90]
  wire  _T_1342 = _T_1339 | _T_1341; // @[lib.scala 117:72]
  wire  _T_1346 = _T_1339 | _T_1343; // @[lib.scala 119:78]
  wire  extintsrc_req_gw_5 = gw_config_reg_5[1] ? _T_1346 : _T_1339; // @[lib.scala 119:8]
  wire  _T_1354 = extintsrc_req_sync_6 ^ gw_config_reg_6[0]; // @[lib.scala 117:50]
  wire  _T_1355 = ~gw_clear_reg_we_6; // @[lib.scala 117:92]
  reg  _T_1358; // @[Reg.scala 27:20]
  wire  _T_1356 = _T_1358 & _T_1355; // @[lib.scala 117:90]
  wire  _T_1357 = _T_1354 | _T_1356; // @[lib.scala 117:72]
  wire  _T_1361 = _T_1354 | _T_1358; // @[lib.scala 119:78]
  wire  extintsrc_req_gw_6 = gw_config_reg_6[1] ? _T_1361 : _T_1354; // @[lib.scala 119:8]
  wire  _T_1369 = extintsrc_req_sync_7 ^ gw_config_reg_7[0]; // @[lib.scala 117:50]
  wire  _T_1370 = ~gw_clear_reg_we_7; // @[lib.scala 117:92]
  reg  _T_1373; // @[Reg.scala 27:20]
  wire  _T_1371 = _T_1373 & _T_1370; // @[lib.scala 117:90]
  wire  _T_1372 = _T_1369 | _T_1371; // @[lib.scala 117:72]
  wire  _T_1376 = _T_1369 | _T_1373; // @[lib.scala 119:78]
  wire  extintsrc_req_gw_7 = gw_config_reg_7[1] ? _T_1376 : _T_1369; // @[lib.scala 119:8]
  wire  _T_1384 = extintsrc_req_sync_8 ^ gw_config_reg_8[0]; // @[lib.scala 117:50]
  wire  _T_1385 = ~gw_clear_reg_we_8; // @[lib.scala 117:92]
  reg  _T_1388; // @[Reg.scala 27:20]
  wire  _T_1386 = _T_1388 & _T_1385; // @[lib.scala 117:90]
  wire  _T_1387 = _T_1384 | _T_1386; // @[lib.scala 117:72]
  wire  _T_1391 = _T_1384 | _T_1388; // @[lib.scala 119:78]
  wire  extintsrc_req_gw_8 = gw_config_reg_8[1] ? _T_1391 : _T_1384; // @[lib.scala 119:8]
  wire  _T_1399 = extintsrc_req_sync_9 ^ gw_config_reg_9[0]; // @[lib.scala 117:50]
  wire  _T_1400 = ~gw_clear_reg_we_9; // @[lib.scala 117:92]
  reg  _T_1403; // @[Reg.scala 27:20]
  wire  _T_1401 = _T_1403 & _T_1400; // @[lib.scala 117:90]
  wire  _T_1402 = _T_1399 | _T_1401; // @[lib.scala 117:72]
  wire  _T_1406 = _T_1399 | _T_1403; // @[lib.scala 119:78]
  wire  extintsrc_req_gw_9 = gw_config_reg_9[1] ? _T_1406 : _T_1399; // @[lib.scala 119:8]
  wire  _T_1414 = extintsrc_req_sync_10 ^ gw_config_reg_10[0]; // @[lib.scala 117:50]
  wire  _T_1415 = ~gw_clear_reg_we_10; // @[lib.scala 117:92]
  reg  _T_1418; // @[Reg.scala 27:20]
  wire  _T_1416 = _T_1418 & _T_1415; // @[lib.scala 117:90]
  wire  _T_1417 = _T_1414 | _T_1416; // @[lib.scala 117:72]
  wire  _T_1421 = _T_1414 | _T_1418; // @[lib.scala 119:78]
  wire  extintsrc_req_gw_10 = gw_config_reg_10[1] ? _T_1421 : _T_1414; // @[lib.scala 119:8]
  wire  _T_1429 = extintsrc_req_sync_11 ^ gw_config_reg_11[0]; // @[lib.scala 117:50]
  wire  _T_1430 = ~gw_clear_reg_we_11; // @[lib.scala 117:92]
  reg  _T_1433; // @[Reg.scala 27:20]
  wire  _T_1431 = _T_1433 & _T_1430; // @[lib.scala 117:90]
  wire  _T_1432 = _T_1429 | _T_1431; // @[lib.scala 117:72]
  wire  _T_1436 = _T_1429 | _T_1433; // @[lib.scala 119:78]
  wire  extintsrc_req_gw_11 = gw_config_reg_11[1] ? _T_1436 : _T_1429; // @[lib.scala 119:8]
  wire  _T_1444 = extintsrc_req_sync_12 ^ gw_config_reg_12[0]; // @[lib.scala 117:50]
  wire  _T_1445 = ~gw_clear_reg_we_12; // @[lib.scala 117:92]
  reg  _T_1448; // @[Reg.scala 27:20]
  wire  _T_1446 = _T_1448 & _T_1445; // @[lib.scala 117:90]
  wire  _T_1447 = _T_1444 | _T_1446; // @[lib.scala 117:72]
  wire  _T_1451 = _T_1444 | _T_1448; // @[lib.scala 119:78]
  wire  extintsrc_req_gw_12 = gw_config_reg_12[1] ? _T_1451 : _T_1444; // @[lib.scala 119:8]
  wire  _T_1459 = extintsrc_req_sync_13 ^ gw_config_reg_13[0]; // @[lib.scala 117:50]
  wire  _T_1460 = ~gw_clear_reg_we_13; // @[lib.scala 117:92]
  reg  _T_1463; // @[Reg.scala 27:20]
  wire  _T_1461 = _T_1463 & _T_1460; // @[lib.scala 117:90]
  wire  _T_1462 = _T_1459 | _T_1461; // @[lib.scala 117:72]
  wire  _T_1466 = _T_1459 | _T_1463; // @[lib.scala 119:78]
  wire  extintsrc_req_gw_13 = gw_config_reg_13[1] ? _T_1466 : _T_1459; // @[lib.scala 119:8]
  wire  _T_1474 = extintsrc_req_sync_14 ^ gw_config_reg_14[0]; // @[lib.scala 117:50]
  wire  _T_1475 = ~gw_clear_reg_we_14; // @[lib.scala 117:92]
  reg  _T_1478; // @[Reg.scala 27:20]
  wire  _T_1476 = _T_1478 & _T_1475; // @[lib.scala 117:90]
  wire  _T_1477 = _T_1474 | _T_1476; // @[lib.scala 117:72]
  wire  _T_1481 = _T_1474 | _T_1478; // @[lib.scala 119:78]
  wire  extintsrc_req_gw_14 = gw_config_reg_14[1] ? _T_1481 : _T_1474; // @[lib.scala 119:8]
  wire  _T_1489 = extintsrc_req_sync_15 ^ gw_config_reg_15[0]; // @[lib.scala 117:50]
  wire  _T_1490 = ~gw_clear_reg_we_15; // @[lib.scala 117:92]
  reg  _T_1493; // @[Reg.scala 27:20]
  wire  _T_1491 = _T_1493 & _T_1490; // @[lib.scala 117:90]
  wire  _T_1492 = _T_1489 | _T_1491; // @[lib.scala 117:72]
  wire  _T_1496 = _T_1489 | _T_1493; // @[lib.scala 119:78]
  wire  extintsrc_req_gw_15 = gw_config_reg_15[1] ? _T_1496 : _T_1489; // @[lib.scala 119:8]
  wire  _T_1504 = extintsrc_req_sync_16 ^ gw_config_reg_16[0]; // @[lib.scala 117:50]
  wire  _T_1505 = ~gw_clear_reg_we_16; // @[lib.scala 117:92]
  reg  _T_1508; // @[Reg.scala 27:20]
  wire  _T_1506 = _T_1508 & _T_1505; // @[lib.scala 117:90]
  wire  _T_1507 = _T_1504 | _T_1506; // @[lib.scala 117:72]
  wire  _T_1511 = _T_1504 | _T_1508; // @[lib.scala 119:78]
  wire  extintsrc_req_gw_16 = gw_config_reg_16[1] ? _T_1511 : _T_1504; // @[lib.scala 119:8]
  wire  _T_1519 = extintsrc_req_sync_17 ^ gw_config_reg_17[0]; // @[lib.scala 117:50]
  wire  _T_1520 = ~gw_clear_reg_we_17; // @[lib.scala 117:92]
  reg  _T_1523; // @[Reg.scala 27:20]
  wire  _T_1521 = _T_1523 & _T_1520; // @[lib.scala 117:90]
  wire  _T_1522 = _T_1519 | _T_1521; // @[lib.scala 117:72]
  wire  _T_1526 = _T_1519 | _T_1523; // @[lib.scala 119:78]
  wire  extintsrc_req_gw_17 = gw_config_reg_17[1] ? _T_1526 : _T_1519; // @[lib.scala 119:8]
  wire  _T_1534 = extintsrc_req_sync_18 ^ gw_config_reg_18[0]; // @[lib.scala 117:50]
  wire  _T_1535 = ~gw_clear_reg_we_18; // @[lib.scala 117:92]
  reg  _T_1538; // @[Reg.scala 27:20]
  wire  _T_1536 = _T_1538 & _T_1535; // @[lib.scala 117:90]
  wire  _T_1537 = _T_1534 | _T_1536; // @[lib.scala 117:72]
  wire  _T_1541 = _T_1534 | _T_1538; // @[lib.scala 119:78]
  wire  extintsrc_req_gw_18 = gw_config_reg_18[1] ? _T_1541 : _T_1534; // @[lib.scala 119:8]
  wire  _T_1549 = extintsrc_req_sync_19 ^ gw_config_reg_19[0]; // @[lib.scala 117:50]
  wire  _T_1550 = ~gw_clear_reg_we_19; // @[lib.scala 117:92]
  reg  _T_1553; // @[Reg.scala 27:20]
  wire  _T_1551 = _T_1553 & _T_1550; // @[lib.scala 117:90]
  wire  _T_1552 = _T_1549 | _T_1551; // @[lib.scala 117:72]
  wire  _T_1556 = _T_1549 | _T_1553; // @[lib.scala 119:78]
  wire  extintsrc_req_gw_19 = gw_config_reg_19[1] ? _T_1556 : _T_1549; // @[lib.scala 119:8]
  wire  _T_1564 = extintsrc_req_sync_20 ^ gw_config_reg_20[0]; // @[lib.scala 117:50]
  wire  _T_1565 = ~gw_clear_reg_we_20; // @[lib.scala 117:92]
  reg  _T_1568; // @[Reg.scala 27:20]
  wire  _T_1566 = _T_1568 & _T_1565; // @[lib.scala 117:90]
  wire  _T_1567 = _T_1564 | _T_1566; // @[lib.scala 117:72]
  wire  _T_1571 = _T_1564 | _T_1568; // @[lib.scala 119:78]
  wire  extintsrc_req_gw_20 = gw_config_reg_20[1] ? _T_1571 : _T_1564; // @[lib.scala 119:8]
  wire  _T_1579 = extintsrc_req_sync_21 ^ gw_config_reg_21[0]; // @[lib.scala 117:50]
  wire  _T_1580 = ~gw_clear_reg_we_21; // @[lib.scala 117:92]
  reg  _T_1583; // @[Reg.scala 27:20]
  wire  _T_1581 = _T_1583 & _T_1580; // @[lib.scala 117:90]
  wire  _T_1582 = _T_1579 | _T_1581; // @[lib.scala 117:72]
  wire  _T_1586 = _T_1579 | _T_1583; // @[lib.scala 119:78]
  wire  extintsrc_req_gw_21 = gw_config_reg_21[1] ? _T_1586 : _T_1579; // @[lib.scala 119:8]
  wire  _T_1594 = extintsrc_req_sync_22 ^ gw_config_reg_22[0]; // @[lib.scala 117:50]
  wire  _T_1595 = ~gw_clear_reg_we_22; // @[lib.scala 117:92]
  reg  _T_1598; // @[Reg.scala 27:20]
  wire  _T_1596 = _T_1598 & _T_1595; // @[lib.scala 117:90]
  wire  _T_1597 = _T_1594 | _T_1596; // @[lib.scala 117:72]
  wire  _T_1601 = _T_1594 | _T_1598; // @[lib.scala 119:78]
  wire  extintsrc_req_gw_22 = gw_config_reg_22[1] ? _T_1601 : _T_1594; // @[lib.scala 119:8]
  wire  _T_1609 = extintsrc_req_sync_23 ^ gw_config_reg_23[0]; // @[lib.scala 117:50]
  wire  _T_1610 = ~gw_clear_reg_we_23; // @[lib.scala 117:92]
  reg  _T_1613; // @[Reg.scala 27:20]
  wire  _T_1611 = _T_1613 & _T_1610; // @[lib.scala 117:90]
  wire  _T_1612 = _T_1609 | _T_1611; // @[lib.scala 117:72]
  wire  _T_1616 = _T_1609 | _T_1613; // @[lib.scala 119:78]
  wire  extintsrc_req_gw_23 = gw_config_reg_23[1] ? _T_1616 : _T_1609; // @[lib.scala 119:8]
  wire  _T_1624 = extintsrc_req_sync_24 ^ gw_config_reg_24[0]; // @[lib.scala 117:50]
  wire  _T_1625 = ~gw_clear_reg_we_24; // @[lib.scala 117:92]
  reg  _T_1628; // @[Reg.scala 27:20]
  wire  _T_1626 = _T_1628 & _T_1625; // @[lib.scala 117:90]
  wire  _T_1627 = _T_1624 | _T_1626; // @[lib.scala 117:72]
  wire  _T_1631 = _T_1624 | _T_1628; // @[lib.scala 119:78]
  wire  extintsrc_req_gw_24 = gw_config_reg_24[1] ? _T_1631 : _T_1624; // @[lib.scala 119:8]
  wire  _T_1639 = extintsrc_req_sync_25 ^ gw_config_reg_25[0]; // @[lib.scala 117:50]
  wire  _T_1640 = ~gw_clear_reg_we_25; // @[lib.scala 117:92]
  reg  _T_1643; // @[Reg.scala 27:20]
  wire  _T_1641 = _T_1643 & _T_1640; // @[lib.scala 117:90]
  wire  _T_1642 = _T_1639 | _T_1641; // @[lib.scala 117:72]
  wire  _T_1646 = _T_1639 | _T_1643; // @[lib.scala 119:78]
  wire  extintsrc_req_gw_25 = gw_config_reg_25[1] ? _T_1646 : _T_1639; // @[lib.scala 119:8]
  wire  _T_1654 = extintsrc_req_sync_26 ^ gw_config_reg_26[0]; // @[lib.scala 117:50]
  wire  _T_1655 = ~gw_clear_reg_we_26; // @[lib.scala 117:92]
  reg  _T_1658; // @[Reg.scala 27:20]
  wire  _T_1656 = _T_1658 & _T_1655; // @[lib.scala 117:90]
  wire  _T_1657 = _T_1654 | _T_1656; // @[lib.scala 117:72]
  wire  _T_1661 = _T_1654 | _T_1658; // @[lib.scala 119:78]
  wire  extintsrc_req_gw_26 = gw_config_reg_26[1] ? _T_1661 : _T_1654; // @[lib.scala 119:8]
  wire  _T_1669 = extintsrc_req_sync_27 ^ gw_config_reg_27[0]; // @[lib.scala 117:50]
  wire  _T_1670 = ~gw_clear_reg_we_27; // @[lib.scala 117:92]
  reg  _T_1673; // @[Reg.scala 27:20]
  wire  _T_1671 = _T_1673 & _T_1670; // @[lib.scala 117:90]
  wire  _T_1672 = _T_1669 | _T_1671; // @[lib.scala 117:72]
  wire  _T_1676 = _T_1669 | _T_1673; // @[lib.scala 119:78]
  wire  extintsrc_req_gw_27 = gw_config_reg_27[1] ? _T_1676 : _T_1669; // @[lib.scala 119:8]
  wire  _T_1684 = extintsrc_req_sync_28 ^ gw_config_reg_28[0]; // @[lib.scala 117:50]
  wire  _T_1685 = ~gw_clear_reg_we_28; // @[lib.scala 117:92]
  reg  _T_1688; // @[Reg.scala 27:20]
  wire  _T_1686 = _T_1688 & _T_1685; // @[lib.scala 117:90]
  wire  _T_1687 = _T_1684 | _T_1686; // @[lib.scala 117:72]
  wire  _T_1691 = _T_1684 | _T_1688; // @[lib.scala 119:78]
  wire  extintsrc_req_gw_28 = gw_config_reg_28[1] ? _T_1691 : _T_1684; // @[lib.scala 119:8]
  wire  _T_1699 = extintsrc_req_sync_29 ^ gw_config_reg_29[0]; // @[lib.scala 117:50]
  wire  _T_1700 = ~gw_clear_reg_we_29; // @[lib.scala 117:92]
  reg  _T_1703; // @[Reg.scala 27:20]
  wire  _T_1701 = _T_1703 & _T_1700; // @[lib.scala 117:90]
  wire  _T_1702 = _T_1699 | _T_1701; // @[lib.scala 117:72]
  wire  _T_1706 = _T_1699 | _T_1703; // @[lib.scala 119:78]
  wire  extintsrc_req_gw_29 = gw_config_reg_29[1] ? _T_1706 : _T_1699; // @[lib.scala 119:8]
  wire  _T_1714 = extintsrc_req_sync_30 ^ gw_config_reg_30[0]; // @[lib.scala 117:50]
  wire  _T_1715 = ~gw_clear_reg_we_30; // @[lib.scala 117:92]
  reg  _T_1718; // @[Reg.scala 27:20]
  wire  _T_1716 = _T_1718 & _T_1715; // @[lib.scala 117:90]
  wire  _T_1717 = _T_1714 | _T_1716; // @[lib.scala 117:72]
  wire  _T_1721 = _T_1714 | _T_1718; // @[lib.scala 119:78]
  wire  extintsrc_req_gw_30 = gw_config_reg_30[1] ? _T_1721 : _T_1714; // @[lib.scala 119:8]
  wire  _T_1729 = extintsrc_req_sync_31 ^ gw_config_reg_31[0]; // @[lib.scala 117:50]
  wire  _T_1730 = ~gw_clear_reg_we_31; // @[lib.scala 117:92]
  reg  _T_1733; // @[Reg.scala 27:20]
  wire  _T_1731 = _T_1733 & _T_1730; // @[lib.scala 117:90]
  wire  _T_1732 = _T_1729 | _T_1731; // @[lib.scala 117:72]
  wire  _T_1736 = _T_1729 | _T_1733; // @[lib.scala 119:78]
  wire  extintsrc_req_gw_31 = gw_config_reg_31[1] ? _T_1736 : _T_1729; // @[lib.scala 119:8]
  reg  config_reg; // @[Reg.scala 27:20]
  wire [3:0] intpriority_reg_0 = 4'h0; // @[pic_ctrl.scala 163:32 pic_ctrl.scala 164:208]
  wire [3:0] _T_1742 = ~intpriority_reg_1; // @[pic_ctrl.scala 176:89]
  wire [3:0] intpriority_reg_inv_1 = config_reg ? _T_1742 : intpriority_reg_1; // @[pic_ctrl.scala 176:70]
  wire [3:0] _T_1745 = ~intpriority_reg_2; // @[pic_ctrl.scala 176:89]
  wire [3:0] intpriority_reg_inv_2 = config_reg ? _T_1745 : intpriority_reg_2; // @[pic_ctrl.scala 176:70]
  wire [3:0] _T_1748 = ~intpriority_reg_3; // @[pic_ctrl.scala 176:89]
  wire [3:0] intpriority_reg_inv_3 = config_reg ? _T_1748 : intpriority_reg_3; // @[pic_ctrl.scala 176:70]
  wire [3:0] _T_1751 = ~intpriority_reg_4; // @[pic_ctrl.scala 176:89]
  wire [3:0] intpriority_reg_inv_4 = config_reg ? _T_1751 : intpriority_reg_4; // @[pic_ctrl.scala 176:70]
  wire [3:0] _T_1754 = ~intpriority_reg_5; // @[pic_ctrl.scala 176:89]
  wire [3:0] intpriority_reg_inv_5 = config_reg ? _T_1754 : intpriority_reg_5; // @[pic_ctrl.scala 176:70]
  wire [3:0] _T_1757 = ~intpriority_reg_6; // @[pic_ctrl.scala 176:89]
  wire [3:0] intpriority_reg_inv_6 = config_reg ? _T_1757 : intpriority_reg_6; // @[pic_ctrl.scala 176:70]
  wire [3:0] _T_1760 = ~intpriority_reg_7; // @[pic_ctrl.scala 176:89]
  wire [3:0] intpriority_reg_inv_7 = config_reg ? _T_1760 : intpriority_reg_7; // @[pic_ctrl.scala 176:70]
  wire [3:0] _T_1763 = ~intpriority_reg_8; // @[pic_ctrl.scala 176:89]
  wire [3:0] intpriority_reg_inv_8 = config_reg ? _T_1763 : intpriority_reg_8; // @[pic_ctrl.scala 176:70]
  wire [3:0] _T_1766 = ~intpriority_reg_9; // @[pic_ctrl.scala 176:89]
  wire [3:0] intpriority_reg_inv_9 = config_reg ? _T_1766 : intpriority_reg_9; // @[pic_ctrl.scala 176:70]
  wire [3:0] _T_1769 = ~intpriority_reg_10; // @[pic_ctrl.scala 176:89]
  wire [3:0] intpriority_reg_inv_10 = config_reg ? _T_1769 : intpriority_reg_10; // @[pic_ctrl.scala 176:70]
  wire [3:0] _T_1772 = ~intpriority_reg_11; // @[pic_ctrl.scala 176:89]
  wire [3:0] intpriority_reg_inv_11 = config_reg ? _T_1772 : intpriority_reg_11; // @[pic_ctrl.scala 176:70]
  wire [3:0] _T_1775 = ~intpriority_reg_12; // @[pic_ctrl.scala 176:89]
  wire [3:0] intpriority_reg_inv_12 = config_reg ? _T_1775 : intpriority_reg_12; // @[pic_ctrl.scala 176:70]
  wire [3:0] _T_1778 = ~intpriority_reg_13; // @[pic_ctrl.scala 176:89]
  wire [3:0] intpriority_reg_inv_13 = config_reg ? _T_1778 : intpriority_reg_13; // @[pic_ctrl.scala 176:70]
  wire [3:0] _T_1781 = ~intpriority_reg_14; // @[pic_ctrl.scala 176:89]
  wire [3:0] intpriority_reg_inv_14 = config_reg ? _T_1781 : intpriority_reg_14; // @[pic_ctrl.scala 176:70]
  wire [3:0] _T_1784 = ~intpriority_reg_15; // @[pic_ctrl.scala 176:89]
  wire [3:0] intpriority_reg_inv_15 = config_reg ? _T_1784 : intpriority_reg_15; // @[pic_ctrl.scala 176:70]
  wire [3:0] _T_1787 = ~intpriority_reg_16; // @[pic_ctrl.scala 176:89]
  wire [3:0] intpriority_reg_inv_16 = config_reg ? _T_1787 : intpriority_reg_16; // @[pic_ctrl.scala 176:70]
  wire [3:0] _T_1790 = ~intpriority_reg_17; // @[pic_ctrl.scala 176:89]
  wire [3:0] intpriority_reg_inv_17 = config_reg ? _T_1790 : intpriority_reg_17; // @[pic_ctrl.scala 176:70]
  wire [3:0] _T_1793 = ~intpriority_reg_18; // @[pic_ctrl.scala 176:89]
  wire [3:0] intpriority_reg_inv_18 = config_reg ? _T_1793 : intpriority_reg_18; // @[pic_ctrl.scala 176:70]
  wire [3:0] _T_1796 = ~intpriority_reg_19; // @[pic_ctrl.scala 176:89]
  wire [3:0] intpriority_reg_inv_19 = config_reg ? _T_1796 : intpriority_reg_19; // @[pic_ctrl.scala 176:70]
  wire [3:0] _T_1799 = ~intpriority_reg_20; // @[pic_ctrl.scala 176:89]
  wire [3:0] intpriority_reg_inv_20 = config_reg ? _T_1799 : intpriority_reg_20; // @[pic_ctrl.scala 176:70]
  wire [3:0] _T_1802 = ~intpriority_reg_21; // @[pic_ctrl.scala 176:89]
  wire [3:0] intpriority_reg_inv_21 = config_reg ? _T_1802 : intpriority_reg_21; // @[pic_ctrl.scala 176:70]
  wire [3:0] _T_1805 = ~intpriority_reg_22; // @[pic_ctrl.scala 176:89]
  wire [3:0] intpriority_reg_inv_22 = config_reg ? _T_1805 : intpriority_reg_22; // @[pic_ctrl.scala 176:70]
  wire [3:0] _T_1808 = ~intpriority_reg_23; // @[pic_ctrl.scala 176:89]
  wire [3:0] intpriority_reg_inv_23 = config_reg ? _T_1808 : intpriority_reg_23; // @[pic_ctrl.scala 176:70]
  wire [3:0] _T_1811 = ~intpriority_reg_24; // @[pic_ctrl.scala 176:89]
  wire [3:0] intpriority_reg_inv_24 = config_reg ? _T_1811 : intpriority_reg_24; // @[pic_ctrl.scala 176:70]
  wire [3:0] _T_1814 = ~intpriority_reg_25; // @[pic_ctrl.scala 176:89]
  wire [3:0] intpriority_reg_inv_25 = config_reg ? _T_1814 : intpriority_reg_25; // @[pic_ctrl.scala 176:70]
  wire [3:0] _T_1817 = ~intpriority_reg_26; // @[pic_ctrl.scala 176:89]
  wire [3:0] intpriority_reg_inv_26 = config_reg ? _T_1817 : intpriority_reg_26; // @[pic_ctrl.scala 176:70]
  wire [3:0] _T_1820 = ~intpriority_reg_27; // @[pic_ctrl.scala 176:89]
  wire [3:0] intpriority_reg_inv_27 = config_reg ? _T_1820 : intpriority_reg_27; // @[pic_ctrl.scala 176:70]
  wire [3:0] _T_1823 = ~intpriority_reg_28; // @[pic_ctrl.scala 176:89]
  wire [3:0] intpriority_reg_inv_28 = config_reg ? _T_1823 : intpriority_reg_28; // @[pic_ctrl.scala 176:70]
  wire [3:0] _T_1826 = ~intpriority_reg_29; // @[pic_ctrl.scala 176:89]
  wire [3:0] intpriority_reg_inv_29 = config_reg ? _T_1826 : intpriority_reg_29; // @[pic_ctrl.scala 176:70]
  wire [3:0] _T_1829 = ~intpriority_reg_30; // @[pic_ctrl.scala 176:89]
  wire [3:0] intpriority_reg_inv_30 = config_reg ? _T_1829 : intpriority_reg_30; // @[pic_ctrl.scala 176:70]
  wire [3:0] _T_1832 = ~intpriority_reg_31; // @[pic_ctrl.scala 176:89]
  wire [3:0] intpriority_reg_inv_31 = config_reg ? _T_1832 : intpriority_reg_31; // @[pic_ctrl.scala 176:70]
  wire  _T_1838 = extintsrc_req_gw_1 & intenable_reg_1; // @[pic_ctrl.scala 177:109]
  wire [3:0] _T_1840 = _T_1838 ? 4'hf : 4'h0; // @[Bitwise.scala 72:12]
  wire [3:0] intpend_w_prior_en_1 = _T_1840 & intpriority_reg_inv_1; // @[pic_ctrl.scala 177:129]
  wire  _T_1842 = extintsrc_req_gw_2 & intenable_reg_2; // @[pic_ctrl.scala 177:109]
  wire [3:0] _T_1844 = _T_1842 ? 4'hf : 4'h0; // @[Bitwise.scala 72:12]
  wire [3:0] intpend_w_prior_en_2 = _T_1844 & intpriority_reg_inv_2; // @[pic_ctrl.scala 177:129]
  wire  _T_1846 = extintsrc_req_gw_3 & intenable_reg_3; // @[pic_ctrl.scala 177:109]
  wire [3:0] _T_1848 = _T_1846 ? 4'hf : 4'h0; // @[Bitwise.scala 72:12]
  wire [3:0] intpend_w_prior_en_3 = _T_1848 & intpriority_reg_inv_3; // @[pic_ctrl.scala 177:129]
  wire  _T_1850 = extintsrc_req_gw_4 & intenable_reg_4; // @[pic_ctrl.scala 177:109]
  wire [3:0] _T_1852 = _T_1850 ? 4'hf : 4'h0; // @[Bitwise.scala 72:12]
  wire [3:0] intpend_w_prior_en_4 = _T_1852 & intpriority_reg_inv_4; // @[pic_ctrl.scala 177:129]
  wire  _T_1854 = extintsrc_req_gw_5 & intenable_reg_5; // @[pic_ctrl.scala 177:109]
  wire [3:0] _T_1856 = _T_1854 ? 4'hf : 4'h0; // @[Bitwise.scala 72:12]
  wire [3:0] intpend_w_prior_en_5 = _T_1856 & intpriority_reg_inv_5; // @[pic_ctrl.scala 177:129]
  wire  _T_1858 = extintsrc_req_gw_6 & intenable_reg_6; // @[pic_ctrl.scala 177:109]
  wire [3:0] _T_1860 = _T_1858 ? 4'hf : 4'h0; // @[Bitwise.scala 72:12]
  wire [3:0] intpend_w_prior_en_6 = _T_1860 & intpriority_reg_inv_6; // @[pic_ctrl.scala 177:129]
  wire  _T_1862 = extintsrc_req_gw_7 & intenable_reg_7; // @[pic_ctrl.scala 177:109]
  wire [3:0] _T_1864 = _T_1862 ? 4'hf : 4'h0; // @[Bitwise.scala 72:12]
  wire [3:0] intpend_w_prior_en_7 = _T_1864 & intpriority_reg_inv_7; // @[pic_ctrl.scala 177:129]
  wire  _T_1866 = extintsrc_req_gw_8 & intenable_reg_8; // @[pic_ctrl.scala 177:109]
  wire [3:0] _T_1868 = _T_1866 ? 4'hf : 4'h0; // @[Bitwise.scala 72:12]
  wire [3:0] intpend_w_prior_en_8 = _T_1868 & intpriority_reg_inv_8; // @[pic_ctrl.scala 177:129]
  wire  _T_1870 = extintsrc_req_gw_9 & intenable_reg_9; // @[pic_ctrl.scala 177:109]
  wire [3:0] _T_1872 = _T_1870 ? 4'hf : 4'h0; // @[Bitwise.scala 72:12]
  wire [3:0] intpend_w_prior_en_9 = _T_1872 & intpriority_reg_inv_9; // @[pic_ctrl.scala 177:129]
  wire  _T_1874 = extintsrc_req_gw_10 & intenable_reg_10; // @[pic_ctrl.scala 177:109]
  wire [3:0] _T_1876 = _T_1874 ? 4'hf : 4'h0; // @[Bitwise.scala 72:12]
  wire [3:0] intpend_w_prior_en_10 = _T_1876 & intpriority_reg_inv_10; // @[pic_ctrl.scala 177:129]
  wire  _T_1878 = extintsrc_req_gw_11 & intenable_reg_11; // @[pic_ctrl.scala 177:109]
  wire [3:0] _T_1880 = _T_1878 ? 4'hf : 4'h0; // @[Bitwise.scala 72:12]
  wire [3:0] intpend_w_prior_en_11 = _T_1880 & intpriority_reg_inv_11; // @[pic_ctrl.scala 177:129]
  wire  _T_1882 = extintsrc_req_gw_12 & intenable_reg_12; // @[pic_ctrl.scala 177:109]
  wire [3:0] _T_1884 = _T_1882 ? 4'hf : 4'h0; // @[Bitwise.scala 72:12]
  wire [3:0] intpend_w_prior_en_12 = _T_1884 & intpriority_reg_inv_12; // @[pic_ctrl.scala 177:129]
  wire  _T_1886 = extintsrc_req_gw_13 & intenable_reg_13; // @[pic_ctrl.scala 177:109]
  wire [3:0] _T_1888 = _T_1886 ? 4'hf : 4'h0; // @[Bitwise.scala 72:12]
  wire [3:0] intpend_w_prior_en_13 = _T_1888 & intpriority_reg_inv_13; // @[pic_ctrl.scala 177:129]
  wire  _T_1890 = extintsrc_req_gw_14 & intenable_reg_14; // @[pic_ctrl.scala 177:109]
  wire [3:0] _T_1892 = _T_1890 ? 4'hf : 4'h0; // @[Bitwise.scala 72:12]
  wire [3:0] intpend_w_prior_en_14 = _T_1892 & intpriority_reg_inv_14; // @[pic_ctrl.scala 177:129]
  wire  _T_1894 = extintsrc_req_gw_15 & intenable_reg_15; // @[pic_ctrl.scala 177:109]
  wire [3:0] _T_1896 = _T_1894 ? 4'hf : 4'h0; // @[Bitwise.scala 72:12]
  wire [3:0] intpend_w_prior_en_15 = _T_1896 & intpriority_reg_inv_15; // @[pic_ctrl.scala 177:129]
  wire  _T_1898 = extintsrc_req_gw_16 & intenable_reg_16; // @[pic_ctrl.scala 177:109]
  wire [3:0] _T_1900 = _T_1898 ? 4'hf : 4'h0; // @[Bitwise.scala 72:12]
  wire [3:0] intpend_w_prior_en_16 = _T_1900 & intpriority_reg_inv_16; // @[pic_ctrl.scala 177:129]
  wire  _T_1902 = extintsrc_req_gw_17 & intenable_reg_17; // @[pic_ctrl.scala 177:109]
  wire [3:0] _T_1904 = _T_1902 ? 4'hf : 4'h0; // @[Bitwise.scala 72:12]
  wire [3:0] intpend_w_prior_en_17 = _T_1904 & intpriority_reg_inv_17; // @[pic_ctrl.scala 177:129]
  wire  _T_1906 = extintsrc_req_gw_18 & intenable_reg_18; // @[pic_ctrl.scala 177:109]
  wire [3:0] _T_1908 = _T_1906 ? 4'hf : 4'h0; // @[Bitwise.scala 72:12]
  wire [3:0] intpend_w_prior_en_18 = _T_1908 & intpriority_reg_inv_18; // @[pic_ctrl.scala 177:129]
  wire  _T_1910 = extintsrc_req_gw_19 & intenable_reg_19; // @[pic_ctrl.scala 177:109]
  wire [3:0] _T_1912 = _T_1910 ? 4'hf : 4'h0; // @[Bitwise.scala 72:12]
  wire [3:0] intpend_w_prior_en_19 = _T_1912 & intpriority_reg_inv_19; // @[pic_ctrl.scala 177:129]
  wire  _T_1914 = extintsrc_req_gw_20 & intenable_reg_20; // @[pic_ctrl.scala 177:109]
  wire [3:0] _T_1916 = _T_1914 ? 4'hf : 4'h0; // @[Bitwise.scala 72:12]
  wire [3:0] intpend_w_prior_en_20 = _T_1916 & intpriority_reg_inv_20; // @[pic_ctrl.scala 177:129]
  wire  _T_1918 = extintsrc_req_gw_21 & intenable_reg_21; // @[pic_ctrl.scala 177:109]
  wire [3:0] _T_1920 = _T_1918 ? 4'hf : 4'h0; // @[Bitwise.scala 72:12]
  wire [3:0] intpend_w_prior_en_21 = _T_1920 & intpriority_reg_inv_21; // @[pic_ctrl.scala 177:129]
  wire  _T_1922 = extintsrc_req_gw_22 & intenable_reg_22; // @[pic_ctrl.scala 177:109]
  wire [3:0] _T_1924 = _T_1922 ? 4'hf : 4'h0; // @[Bitwise.scala 72:12]
  wire [3:0] intpend_w_prior_en_22 = _T_1924 & intpriority_reg_inv_22; // @[pic_ctrl.scala 177:129]
  wire  _T_1926 = extintsrc_req_gw_23 & intenable_reg_23; // @[pic_ctrl.scala 177:109]
  wire [3:0] _T_1928 = _T_1926 ? 4'hf : 4'h0; // @[Bitwise.scala 72:12]
  wire [3:0] intpend_w_prior_en_23 = _T_1928 & intpriority_reg_inv_23; // @[pic_ctrl.scala 177:129]
  wire  _T_1930 = extintsrc_req_gw_24 & intenable_reg_24; // @[pic_ctrl.scala 177:109]
  wire [3:0] _T_1932 = _T_1930 ? 4'hf : 4'h0; // @[Bitwise.scala 72:12]
  wire [3:0] intpend_w_prior_en_24 = _T_1932 & intpriority_reg_inv_24; // @[pic_ctrl.scala 177:129]
  wire  _T_1934 = extintsrc_req_gw_25 & intenable_reg_25; // @[pic_ctrl.scala 177:109]
  wire [3:0] _T_1936 = _T_1934 ? 4'hf : 4'h0; // @[Bitwise.scala 72:12]
  wire [3:0] intpend_w_prior_en_25 = _T_1936 & intpriority_reg_inv_25; // @[pic_ctrl.scala 177:129]
  wire  _T_1938 = extintsrc_req_gw_26 & intenable_reg_26; // @[pic_ctrl.scala 177:109]
  wire [3:0] _T_1940 = _T_1938 ? 4'hf : 4'h0; // @[Bitwise.scala 72:12]
  wire [3:0] intpend_w_prior_en_26 = _T_1940 & intpriority_reg_inv_26; // @[pic_ctrl.scala 177:129]
  wire  _T_1942 = extintsrc_req_gw_27 & intenable_reg_27; // @[pic_ctrl.scala 177:109]
  wire [3:0] _T_1944 = _T_1942 ? 4'hf : 4'h0; // @[Bitwise.scala 72:12]
  wire [3:0] intpend_w_prior_en_27 = _T_1944 & intpriority_reg_inv_27; // @[pic_ctrl.scala 177:129]
  wire  _T_1946 = extintsrc_req_gw_28 & intenable_reg_28; // @[pic_ctrl.scala 177:109]
  wire [3:0] _T_1948 = _T_1946 ? 4'hf : 4'h0; // @[Bitwise.scala 72:12]
  wire [3:0] intpend_w_prior_en_28 = _T_1948 & intpriority_reg_inv_28; // @[pic_ctrl.scala 177:129]
  wire  _T_1950 = extintsrc_req_gw_29 & intenable_reg_29; // @[pic_ctrl.scala 177:109]
  wire [3:0] _T_1952 = _T_1950 ? 4'hf : 4'h0; // @[Bitwise.scala 72:12]
  wire [3:0] intpend_w_prior_en_29 = _T_1952 & intpriority_reg_inv_29; // @[pic_ctrl.scala 177:129]
  wire  _T_1954 = extintsrc_req_gw_30 & intenable_reg_30; // @[pic_ctrl.scala 177:109]
  wire [3:0] _T_1956 = _T_1954 ? 4'hf : 4'h0; // @[Bitwise.scala 72:12]
  wire [3:0] intpend_w_prior_en_30 = _T_1956 & intpriority_reg_inv_30; // @[pic_ctrl.scala 177:129]
  wire  _T_1958 = extintsrc_req_gw_31 & intenable_reg_31; // @[pic_ctrl.scala 177:109]
  wire [3:0] _T_1960 = _T_1958 ? 4'hf : 4'h0; // @[Bitwise.scala 72:12]
  wire [3:0] intpend_w_prior_en_31 = _T_1960 & intpriority_reg_inv_31; // @[pic_ctrl.scala 177:129]
  wire [7:0] _T_1964 = 8'hff; // @[Bitwise.scala 72:12]
  wire [3:0] level_intpend_w_prior_en_0_0 = 4'h0; // @[pic_ctrl.scala 229:40 pic_ctrl.scala 233:38 pic_ctrl.scala 236:33]
  wire [3:0] _T_1841 = intpend_w_prior_en_1; // @[pic_ctrl.scala 70:42 pic_ctrl.scala 177:63]
  wire [3:0] level_intpend_w_prior_en_0_1 = intpend_w_prior_en_1; // @[pic_ctrl.scala 229:40 pic_ctrl.scala 233:38 pic_ctrl.scala 236:33]
  wire  _T_1966 = intpriority_reg_0 < _T_1841; // @[pic_ctrl.scala 27:20]
  wire [7:0] intpend_id_1 = 8'h1; // @[pic_ctrl.scala 71:42 pic_ctrl.scala 178:55]
  wire [7:0] level_intpend_id_0_1 = 8'h1; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30 pic_ctrl.scala 237:33]
  wire [7:0] intpend_id_0 = 8'h0; // @[pic_ctrl.scala 71:42 pic_ctrl.scala 178:55]
  wire [7:0] level_intpend_id_0_0 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30 pic_ctrl.scala 237:33]
  wire [7:0] out_id = _T_1966 ? intpend_id_1 : intpend_id_0; // @[pic_ctrl.scala 27:9]
  wire [3:0] out_priority = _T_1966 ? _T_1841 : intpriority_reg_0; // @[pic_ctrl.scala 27:49]
  wire [3:0] _T_1845 = intpend_w_prior_en_2; // @[pic_ctrl.scala 70:42 pic_ctrl.scala 177:63]
  wire [3:0] level_intpend_w_prior_en_0_2 = intpend_w_prior_en_2; // @[pic_ctrl.scala 229:40 pic_ctrl.scala 233:38 pic_ctrl.scala 236:33]
  wire [3:0] _T_1849 = intpend_w_prior_en_3; // @[pic_ctrl.scala 70:42 pic_ctrl.scala 177:63]
  wire [3:0] level_intpend_w_prior_en_0_3 = intpend_w_prior_en_3; // @[pic_ctrl.scala 229:40 pic_ctrl.scala 233:38 pic_ctrl.scala 236:33]
  wire  _T_1968 = _T_1845 < _T_1849; // @[pic_ctrl.scala 27:20]
  wire [7:0] intpend_id_3 = 8'h3; // @[pic_ctrl.scala 71:42 pic_ctrl.scala 178:55]
  wire [7:0] level_intpend_id_0_3 = 8'h3; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30 pic_ctrl.scala 237:33]
  wire [7:0] intpend_id_2 = 8'h2; // @[pic_ctrl.scala 71:42 pic_ctrl.scala 178:55]
  wire [7:0] level_intpend_id_0_2 = 8'h2; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30 pic_ctrl.scala 237:33]
  wire [7:0] out_id_1 = _T_1968 ? intpend_id_3 : intpend_id_2; // @[pic_ctrl.scala 27:9]
  wire [3:0] out_priority_1 = _T_1968 ? _T_1849 : _T_1845; // @[pic_ctrl.scala 27:49]
  wire [3:0] _T_1853 = intpend_w_prior_en_4; // @[pic_ctrl.scala 70:42 pic_ctrl.scala 177:63]
  wire [3:0] level_intpend_w_prior_en_0_4 = intpend_w_prior_en_4; // @[pic_ctrl.scala 229:40 pic_ctrl.scala 233:38 pic_ctrl.scala 236:33]
  wire [3:0] _T_1857 = intpend_w_prior_en_5; // @[pic_ctrl.scala 70:42 pic_ctrl.scala 177:63]
  wire [3:0] level_intpend_w_prior_en_0_5 = intpend_w_prior_en_5; // @[pic_ctrl.scala 229:40 pic_ctrl.scala 233:38 pic_ctrl.scala 236:33]
  wire  _T_1970 = _T_1853 < _T_1857; // @[pic_ctrl.scala 27:20]
  wire [7:0] intpend_id_5 = 8'h5; // @[pic_ctrl.scala 71:42 pic_ctrl.scala 178:55]
  wire [7:0] level_intpend_id_0_5 = 8'h5; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30 pic_ctrl.scala 237:33]
  wire [7:0] intpend_id_4 = 8'h4; // @[pic_ctrl.scala 71:42 pic_ctrl.scala 178:55]
  wire [7:0] level_intpend_id_0_4 = 8'h4; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30 pic_ctrl.scala 237:33]
  wire [7:0] out_id_2 = _T_1970 ? intpend_id_5 : intpend_id_4; // @[pic_ctrl.scala 27:9]
  wire [3:0] out_priority_2 = _T_1970 ? _T_1857 : _T_1853; // @[pic_ctrl.scala 27:49]
  wire [3:0] _T_1861 = intpend_w_prior_en_6; // @[pic_ctrl.scala 70:42 pic_ctrl.scala 177:63]
  wire [3:0] level_intpend_w_prior_en_0_6 = intpend_w_prior_en_6; // @[pic_ctrl.scala 229:40 pic_ctrl.scala 233:38 pic_ctrl.scala 236:33]
  wire [3:0] _T_1865 = intpend_w_prior_en_7; // @[pic_ctrl.scala 70:42 pic_ctrl.scala 177:63]
  wire [3:0] level_intpend_w_prior_en_0_7 = intpend_w_prior_en_7; // @[pic_ctrl.scala 229:40 pic_ctrl.scala 233:38 pic_ctrl.scala 236:33]
  wire  _T_1972 = _T_1861 < _T_1865; // @[pic_ctrl.scala 27:20]
  wire [7:0] intpend_id_7 = 8'h7; // @[pic_ctrl.scala 71:42 pic_ctrl.scala 178:55]
  wire [7:0] level_intpend_id_0_7 = 8'h7; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30 pic_ctrl.scala 237:33]
  wire [7:0] intpend_id_6 = 8'h6; // @[pic_ctrl.scala 71:42 pic_ctrl.scala 178:55]
  wire [7:0] level_intpend_id_0_6 = 8'h6; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30 pic_ctrl.scala 237:33]
  wire [7:0] out_id_3 = _T_1972 ? intpend_id_7 : intpend_id_6; // @[pic_ctrl.scala 27:9]
  wire [3:0] out_priority_3 = _T_1972 ? _T_1865 : _T_1861; // @[pic_ctrl.scala 27:49]
  wire [3:0] _T_1869 = intpend_w_prior_en_8; // @[pic_ctrl.scala 70:42 pic_ctrl.scala 177:63]
  wire [3:0] level_intpend_w_prior_en_0_8 = intpend_w_prior_en_8; // @[pic_ctrl.scala 229:40 pic_ctrl.scala 233:38 pic_ctrl.scala 236:33]
  wire [3:0] _T_1873 = intpend_w_prior_en_9; // @[pic_ctrl.scala 70:42 pic_ctrl.scala 177:63]
  wire [3:0] level_intpend_w_prior_en_0_9 = intpend_w_prior_en_9; // @[pic_ctrl.scala 229:40 pic_ctrl.scala 233:38 pic_ctrl.scala 236:33]
  wire  _T_1974 = _T_1869 < _T_1873; // @[pic_ctrl.scala 27:20]
  wire [7:0] intpend_id_9 = 8'h9; // @[pic_ctrl.scala 71:42 pic_ctrl.scala 178:55]
  wire [7:0] level_intpend_id_0_9 = 8'h9; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30 pic_ctrl.scala 237:33]
  wire [7:0] intpend_id_8 = 8'h8; // @[pic_ctrl.scala 71:42 pic_ctrl.scala 178:55]
  wire [7:0] level_intpend_id_0_8 = 8'h8; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30 pic_ctrl.scala 237:33]
  wire [7:0] out_id_4 = _T_1974 ? intpend_id_9 : intpend_id_8; // @[pic_ctrl.scala 27:9]
  wire [3:0] out_priority_4 = _T_1974 ? _T_1873 : _T_1869; // @[pic_ctrl.scala 27:49]
  wire [3:0] _T_1877 = intpend_w_prior_en_10; // @[pic_ctrl.scala 70:42 pic_ctrl.scala 177:63]
  wire [3:0] level_intpend_w_prior_en_0_10 = intpend_w_prior_en_10; // @[pic_ctrl.scala 229:40 pic_ctrl.scala 233:38 pic_ctrl.scala 236:33]
  wire [3:0] _T_1881 = intpend_w_prior_en_11; // @[pic_ctrl.scala 70:42 pic_ctrl.scala 177:63]
  wire [3:0] level_intpend_w_prior_en_0_11 = intpend_w_prior_en_11; // @[pic_ctrl.scala 229:40 pic_ctrl.scala 233:38 pic_ctrl.scala 236:33]
  wire  _T_1976 = _T_1877 < _T_1881; // @[pic_ctrl.scala 27:20]
  wire [7:0] intpend_id_11 = 8'hb; // @[pic_ctrl.scala 71:42 pic_ctrl.scala 178:55]
  wire [7:0] level_intpend_id_0_11 = 8'hb; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30 pic_ctrl.scala 237:33]
  wire [7:0] intpend_id_10 = 8'ha; // @[pic_ctrl.scala 71:42 pic_ctrl.scala 178:55]
  wire [7:0] level_intpend_id_0_10 = 8'ha; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30 pic_ctrl.scala 237:33]
  wire [7:0] out_id_5 = _T_1976 ? intpend_id_11 : intpend_id_10; // @[pic_ctrl.scala 27:9]
  wire [3:0] out_priority_5 = _T_1976 ? _T_1881 : _T_1877; // @[pic_ctrl.scala 27:49]
  wire [3:0] _T_1885 = intpend_w_prior_en_12; // @[pic_ctrl.scala 70:42 pic_ctrl.scala 177:63]
  wire [3:0] level_intpend_w_prior_en_0_12 = intpend_w_prior_en_12; // @[pic_ctrl.scala 229:40 pic_ctrl.scala 233:38 pic_ctrl.scala 236:33]
  wire [3:0] _T_1889 = intpend_w_prior_en_13; // @[pic_ctrl.scala 70:42 pic_ctrl.scala 177:63]
  wire [3:0] level_intpend_w_prior_en_0_13 = intpend_w_prior_en_13; // @[pic_ctrl.scala 229:40 pic_ctrl.scala 233:38 pic_ctrl.scala 236:33]
  wire  _T_1978 = _T_1885 < _T_1889; // @[pic_ctrl.scala 27:20]
  wire [7:0] intpend_id_13 = 8'hd; // @[pic_ctrl.scala 71:42 pic_ctrl.scala 178:55]
  wire [7:0] level_intpend_id_0_13 = 8'hd; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30 pic_ctrl.scala 237:33]
  wire [7:0] intpend_id_12 = 8'hc; // @[pic_ctrl.scala 71:42 pic_ctrl.scala 178:55]
  wire [7:0] level_intpend_id_0_12 = 8'hc; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30 pic_ctrl.scala 237:33]
  wire [7:0] out_id_6 = _T_1978 ? intpend_id_13 : intpend_id_12; // @[pic_ctrl.scala 27:9]
  wire [3:0] out_priority_6 = _T_1978 ? _T_1889 : _T_1885; // @[pic_ctrl.scala 27:49]
  wire [3:0] _T_1893 = intpend_w_prior_en_14; // @[pic_ctrl.scala 70:42 pic_ctrl.scala 177:63]
  wire [3:0] level_intpend_w_prior_en_0_14 = intpend_w_prior_en_14; // @[pic_ctrl.scala 229:40 pic_ctrl.scala 233:38 pic_ctrl.scala 236:33]
  wire [3:0] _T_1897 = intpend_w_prior_en_15; // @[pic_ctrl.scala 70:42 pic_ctrl.scala 177:63]
  wire [3:0] level_intpend_w_prior_en_0_15 = intpend_w_prior_en_15; // @[pic_ctrl.scala 229:40 pic_ctrl.scala 233:38 pic_ctrl.scala 236:33]
  wire  _T_1980 = _T_1893 < _T_1897; // @[pic_ctrl.scala 27:20]
  wire [7:0] intpend_id_15 = 8'hf; // @[pic_ctrl.scala 71:42 pic_ctrl.scala 178:55]
  wire [7:0] level_intpend_id_0_15 = 8'hf; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30 pic_ctrl.scala 237:33]
  wire [7:0] intpend_id_14 = 8'he; // @[pic_ctrl.scala 71:42 pic_ctrl.scala 178:55]
  wire [7:0] level_intpend_id_0_14 = 8'he; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30 pic_ctrl.scala 237:33]
  wire [7:0] out_id_7 = _T_1980 ? intpend_id_15 : intpend_id_14; // @[pic_ctrl.scala 27:9]
  wire [3:0] out_priority_7 = _T_1980 ? _T_1897 : _T_1893; // @[pic_ctrl.scala 27:49]
  wire [3:0] _T_1901 = intpend_w_prior_en_16; // @[pic_ctrl.scala 70:42 pic_ctrl.scala 177:63]
  wire [3:0] level_intpend_w_prior_en_0_16 = intpend_w_prior_en_16; // @[pic_ctrl.scala 229:40 pic_ctrl.scala 233:38 pic_ctrl.scala 236:33]
  wire [3:0] _T_1905 = intpend_w_prior_en_17; // @[pic_ctrl.scala 70:42 pic_ctrl.scala 177:63]
  wire [3:0] level_intpend_w_prior_en_0_17 = intpend_w_prior_en_17; // @[pic_ctrl.scala 229:40 pic_ctrl.scala 233:38 pic_ctrl.scala 236:33]
  wire  _T_1982 = _T_1901 < _T_1905; // @[pic_ctrl.scala 27:20]
  wire [7:0] intpend_id_17 = 8'h11; // @[pic_ctrl.scala 71:42 pic_ctrl.scala 178:55]
  wire [7:0] level_intpend_id_0_17 = 8'h11; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30 pic_ctrl.scala 237:33]
  wire [7:0] intpend_id_16 = 8'h10; // @[pic_ctrl.scala 71:42 pic_ctrl.scala 178:55]
  wire [7:0] level_intpend_id_0_16 = 8'h10; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30 pic_ctrl.scala 237:33]
  wire [7:0] out_id_8 = _T_1982 ? intpend_id_17 : intpend_id_16; // @[pic_ctrl.scala 27:9]
  wire [3:0] out_priority_8 = _T_1982 ? _T_1905 : _T_1901; // @[pic_ctrl.scala 27:49]
  wire [3:0] _T_1909 = intpend_w_prior_en_18; // @[pic_ctrl.scala 70:42 pic_ctrl.scala 177:63]
  wire [3:0] level_intpend_w_prior_en_0_18 = intpend_w_prior_en_18; // @[pic_ctrl.scala 229:40 pic_ctrl.scala 233:38 pic_ctrl.scala 236:33]
  wire [3:0] _T_1913 = intpend_w_prior_en_19; // @[pic_ctrl.scala 70:42 pic_ctrl.scala 177:63]
  wire [3:0] level_intpend_w_prior_en_0_19 = intpend_w_prior_en_19; // @[pic_ctrl.scala 229:40 pic_ctrl.scala 233:38 pic_ctrl.scala 236:33]
  wire  _T_1984 = _T_1909 < _T_1913; // @[pic_ctrl.scala 27:20]
  wire [7:0] intpend_id_19 = 8'h13; // @[pic_ctrl.scala 71:42 pic_ctrl.scala 178:55]
  wire [7:0] level_intpend_id_0_19 = 8'h13; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30 pic_ctrl.scala 237:33]
  wire [7:0] intpend_id_18 = 8'h12; // @[pic_ctrl.scala 71:42 pic_ctrl.scala 178:55]
  wire [7:0] level_intpend_id_0_18 = 8'h12; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30 pic_ctrl.scala 237:33]
  wire [7:0] out_id_9 = _T_1984 ? intpend_id_19 : intpend_id_18; // @[pic_ctrl.scala 27:9]
  wire [3:0] out_priority_9 = _T_1984 ? _T_1913 : _T_1909; // @[pic_ctrl.scala 27:49]
  wire [3:0] _T_1917 = intpend_w_prior_en_20; // @[pic_ctrl.scala 70:42 pic_ctrl.scala 177:63]
  wire [3:0] level_intpend_w_prior_en_0_20 = intpend_w_prior_en_20; // @[pic_ctrl.scala 229:40 pic_ctrl.scala 233:38 pic_ctrl.scala 236:33]
  wire [3:0] _T_1921 = intpend_w_prior_en_21; // @[pic_ctrl.scala 70:42 pic_ctrl.scala 177:63]
  wire [3:0] level_intpend_w_prior_en_0_21 = intpend_w_prior_en_21; // @[pic_ctrl.scala 229:40 pic_ctrl.scala 233:38 pic_ctrl.scala 236:33]
  wire  _T_1986 = _T_1917 < _T_1921; // @[pic_ctrl.scala 27:20]
  wire [7:0] intpend_id_21 = 8'h15; // @[pic_ctrl.scala 71:42 pic_ctrl.scala 178:55]
  wire [7:0] level_intpend_id_0_21 = 8'h15; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30 pic_ctrl.scala 237:33]
  wire [7:0] intpend_id_20 = 8'h14; // @[pic_ctrl.scala 71:42 pic_ctrl.scala 178:55]
  wire [7:0] level_intpend_id_0_20 = 8'h14; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30 pic_ctrl.scala 237:33]
  wire [7:0] out_id_10 = _T_1986 ? intpend_id_21 : intpend_id_20; // @[pic_ctrl.scala 27:9]
  wire [3:0] out_priority_10 = _T_1986 ? _T_1921 : _T_1917; // @[pic_ctrl.scala 27:49]
  wire [3:0] _T_1925 = intpend_w_prior_en_22; // @[pic_ctrl.scala 70:42 pic_ctrl.scala 177:63]
  wire [3:0] level_intpend_w_prior_en_0_22 = intpend_w_prior_en_22; // @[pic_ctrl.scala 229:40 pic_ctrl.scala 233:38 pic_ctrl.scala 236:33]
  wire [3:0] _T_1929 = intpend_w_prior_en_23; // @[pic_ctrl.scala 70:42 pic_ctrl.scala 177:63]
  wire [3:0] level_intpend_w_prior_en_0_23 = intpend_w_prior_en_23; // @[pic_ctrl.scala 229:40 pic_ctrl.scala 233:38 pic_ctrl.scala 236:33]
  wire  _T_1988 = _T_1925 < _T_1929; // @[pic_ctrl.scala 27:20]
  wire [7:0] intpend_id_23 = 8'h17; // @[pic_ctrl.scala 71:42 pic_ctrl.scala 178:55]
  wire [7:0] level_intpend_id_0_23 = 8'h17; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30 pic_ctrl.scala 237:33]
  wire [7:0] intpend_id_22 = 8'h16; // @[pic_ctrl.scala 71:42 pic_ctrl.scala 178:55]
  wire [7:0] level_intpend_id_0_22 = 8'h16; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30 pic_ctrl.scala 237:33]
  wire [7:0] out_id_11 = _T_1988 ? intpend_id_23 : intpend_id_22; // @[pic_ctrl.scala 27:9]
  wire [3:0] out_priority_11 = _T_1988 ? _T_1929 : _T_1925; // @[pic_ctrl.scala 27:49]
  wire [3:0] _T_1933 = intpend_w_prior_en_24; // @[pic_ctrl.scala 70:42 pic_ctrl.scala 177:63]
  wire [3:0] level_intpend_w_prior_en_0_24 = intpend_w_prior_en_24; // @[pic_ctrl.scala 229:40 pic_ctrl.scala 233:38 pic_ctrl.scala 236:33]
  wire [3:0] _T_1937 = intpend_w_prior_en_25; // @[pic_ctrl.scala 70:42 pic_ctrl.scala 177:63]
  wire [3:0] level_intpend_w_prior_en_0_25 = intpend_w_prior_en_25; // @[pic_ctrl.scala 229:40 pic_ctrl.scala 233:38 pic_ctrl.scala 236:33]
  wire  _T_1990 = _T_1933 < _T_1937; // @[pic_ctrl.scala 27:20]
  wire [7:0] intpend_id_25 = 8'h19; // @[pic_ctrl.scala 71:42 pic_ctrl.scala 178:55]
  wire [7:0] level_intpend_id_0_25 = 8'h19; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30 pic_ctrl.scala 237:33]
  wire [7:0] intpend_id_24 = 8'h18; // @[pic_ctrl.scala 71:42 pic_ctrl.scala 178:55]
  wire [7:0] level_intpend_id_0_24 = 8'h18; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30 pic_ctrl.scala 237:33]
  wire [7:0] out_id_12 = _T_1990 ? intpend_id_25 : intpend_id_24; // @[pic_ctrl.scala 27:9]
  wire [3:0] out_priority_12 = _T_1990 ? _T_1937 : _T_1933; // @[pic_ctrl.scala 27:49]
  wire [3:0] _T_1941 = intpend_w_prior_en_26; // @[pic_ctrl.scala 70:42 pic_ctrl.scala 177:63]
  wire [3:0] level_intpend_w_prior_en_0_26 = intpend_w_prior_en_26; // @[pic_ctrl.scala 229:40 pic_ctrl.scala 233:38 pic_ctrl.scala 236:33]
  wire [3:0] _T_1945 = intpend_w_prior_en_27; // @[pic_ctrl.scala 70:42 pic_ctrl.scala 177:63]
  wire [3:0] level_intpend_w_prior_en_0_27 = intpend_w_prior_en_27; // @[pic_ctrl.scala 229:40 pic_ctrl.scala 233:38 pic_ctrl.scala 236:33]
  wire  _T_1992 = _T_1941 < _T_1945; // @[pic_ctrl.scala 27:20]
  wire [7:0] intpend_id_27 = 8'h1b; // @[pic_ctrl.scala 71:42 pic_ctrl.scala 178:55]
  wire [7:0] level_intpend_id_0_27 = 8'h1b; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30 pic_ctrl.scala 237:33]
  wire [7:0] intpend_id_26 = 8'h1a; // @[pic_ctrl.scala 71:42 pic_ctrl.scala 178:55]
  wire [7:0] level_intpend_id_0_26 = 8'h1a; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30 pic_ctrl.scala 237:33]
  wire [7:0] out_id_13 = _T_1992 ? intpend_id_27 : intpend_id_26; // @[pic_ctrl.scala 27:9]
  wire [3:0] out_priority_13 = _T_1992 ? _T_1945 : _T_1941; // @[pic_ctrl.scala 27:49]
  wire [3:0] _T_1949 = intpend_w_prior_en_28; // @[pic_ctrl.scala 70:42 pic_ctrl.scala 177:63]
  wire [3:0] level_intpend_w_prior_en_0_28 = intpend_w_prior_en_28; // @[pic_ctrl.scala 229:40 pic_ctrl.scala 233:38 pic_ctrl.scala 236:33]
  wire [3:0] _T_1953 = intpend_w_prior_en_29; // @[pic_ctrl.scala 70:42 pic_ctrl.scala 177:63]
  wire [3:0] level_intpend_w_prior_en_0_29 = intpend_w_prior_en_29; // @[pic_ctrl.scala 229:40 pic_ctrl.scala 233:38 pic_ctrl.scala 236:33]
  wire  _T_1994 = _T_1949 < _T_1953; // @[pic_ctrl.scala 27:20]
  wire [7:0] intpend_id_29 = 8'h1d; // @[pic_ctrl.scala 71:42 pic_ctrl.scala 178:55]
  wire [7:0] level_intpend_id_0_29 = 8'h1d; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30 pic_ctrl.scala 237:33]
  wire [7:0] intpend_id_28 = 8'h1c; // @[pic_ctrl.scala 71:42 pic_ctrl.scala 178:55]
  wire [7:0] level_intpend_id_0_28 = 8'h1c; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30 pic_ctrl.scala 237:33]
  wire [7:0] out_id_14 = _T_1994 ? intpend_id_29 : intpend_id_28; // @[pic_ctrl.scala 27:9]
  wire [3:0] out_priority_14 = _T_1994 ? _T_1953 : _T_1949; // @[pic_ctrl.scala 27:49]
  wire [3:0] _T_1957 = intpend_w_prior_en_30; // @[pic_ctrl.scala 70:42 pic_ctrl.scala 177:63]
  wire [3:0] level_intpend_w_prior_en_0_30 = intpend_w_prior_en_30; // @[pic_ctrl.scala 229:40 pic_ctrl.scala 233:38 pic_ctrl.scala 236:33]
  wire [3:0] _T_1961 = intpend_w_prior_en_31; // @[pic_ctrl.scala 70:42 pic_ctrl.scala 177:63]
  wire [3:0] level_intpend_w_prior_en_0_31 = intpend_w_prior_en_31; // @[pic_ctrl.scala 229:40 pic_ctrl.scala 233:38 pic_ctrl.scala 236:33]
  wire  _T_1996 = _T_1957 < _T_1961; // @[pic_ctrl.scala 27:20]
  wire [7:0] intpend_id_31 = 8'h1f; // @[pic_ctrl.scala 71:42 pic_ctrl.scala 178:55]
  wire [7:0] level_intpend_id_0_31 = 8'h1f; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30 pic_ctrl.scala 237:33]
  wire [7:0] intpend_id_30 = 8'h1e; // @[pic_ctrl.scala 71:42 pic_ctrl.scala 178:55]
  wire [7:0] level_intpend_id_0_30 = 8'h1e; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30 pic_ctrl.scala 237:33]
  wire [7:0] out_id_15 = _T_1996 ? intpend_id_31 : intpend_id_30; // @[pic_ctrl.scala 27:9]
  wire [3:0] out_priority_15 = _T_1996 ? _T_1961 : _T_1957; // @[pic_ctrl.scala 27:49]
  wire [3:0] level_intpend_w_prior_en_0_32 = 4'h0; // @[pic_ctrl.scala 229:40 pic_ctrl.scala 233:38 pic_ctrl.scala 236:33]
  wire [3:0] level_intpend_w_prior_en_0_33 = 4'h0; // @[pic_ctrl.scala 229:40 pic_ctrl.scala 233:38 pic_ctrl.scala 236:33]
  wire  _T_1998 = intpriority_reg_0 < intpriority_reg_0; // @[pic_ctrl.scala 27:20]
  wire [7:0] level_intpend_id_0_33 = 8'hff; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30 pic_ctrl.scala 237:33]
  wire [7:0] level_intpend_id_0_32 = 8'hff; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30 pic_ctrl.scala 237:33]
  wire [7:0] out_id_16 = _T_1998 ? _T_1964 : _T_1964; // @[pic_ctrl.scala 27:9]
  wire  _T_2000 = out_priority < out_priority_1; // @[pic_ctrl.scala 27:20]
  wire [7:0] level_intpend_id_1_1 = out_id_1; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30 pic_ctrl.scala 248:43]
  wire [7:0] level_intpend_id_1_0 = out_id; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30 pic_ctrl.scala 248:43]
  wire [7:0] out_id_17 = _T_2000 ? level_intpend_id_1_1 : level_intpend_id_1_0; // @[pic_ctrl.scala 27:9]
  wire [3:0] out_priority_17 = _T_2000 ? out_priority_1 : out_priority; // @[pic_ctrl.scala 27:49]
  wire  _T_2002 = out_priority_2 < out_priority_3; // @[pic_ctrl.scala 27:20]
  wire [7:0] level_intpend_id_1_3 = out_id_3; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30 pic_ctrl.scala 248:43]
  wire [7:0] level_intpend_id_1_2 = out_id_2; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30 pic_ctrl.scala 248:43]
  wire [7:0] out_id_18 = _T_2002 ? level_intpend_id_1_3 : level_intpend_id_1_2; // @[pic_ctrl.scala 27:9]
  wire [3:0] out_priority_18 = _T_2002 ? out_priority_3 : out_priority_2; // @[pic_ctrl.scala 27:49]
  wire  _T_2004 = out_priority_4 < out_priority_5; // @[pic_ctrl.scala 27:20]
  wire [7:0] level_intpend_id_1_5 = out_id_5; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30 pic_ctrl.scala 248:43]
  wire [7:0] level_intpend_id_1_4 = out_id_4; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30 pic_ctrl.scala 248:43]
  wire [7:0] out_id_19 = _T_2004 ? level_intpend_id_1_5 : level_intpend_id_1_4; // @[pic_ctrl.scala 27:9]
  wire [3:0] out_priority_19 = _T_2004 ? out_priority_5 : out_priority_4; // @[pic_ctrl.scala 27:49]
  wire  _T_2006 = out_priority_6 < out_priority_7; // @[pic_ctrl.scala 27:20]
  wire [7:0] level_intpend_id_1_7 = out_id_7; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30 pic_ctrl.scala 248:43]
  wire [7:0] level_intpend_id_1_6 = out_id_6; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30 pic_ctrl.scala 248:43]
  wire [7:0] out_id_20 = _T_2006 ? level_intpend_id_1_7 : level_intpend_id_1_6; // @[pic_ctrl.scala 27:9]
  wire [3:0] out_priority_20 = _T_2006 ? out_priority_7 : out_priority_6; // @[pic_ctrl.scala 27:49]
  wire  _T_2008 = out_priority_8 < out_priority_9; // @[pic_ctrl.scala 27:20]
  wire [7:0] level_intpend_id_1_9 = out_id_9; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30 pic_ctrl.scala 248:43]
  wire [7:0] level_intpend_id_1_8 = out_id_8; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30 pic_ctrl.scala 248:43]
  wire [7:0] out_id_21 = _T_2008 ? level_intpend_id_1_9 : level_intpend_id_1_8; // @[pic_ctrl.scala 27:9]
  wire [3:0] out_priority_21 = _T_2008 ? out_priority_9 : out_priority_8; // @[pic_ctrl.scala 27:49]
  wire  _T_2010 = out_priority_10 < out_priority_11; // @[pic_ctrl.scala 27:20]
  wire [7:0] level_intpend_id_1_11 = out_id_11; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30 pic_ctrl.scala 248:43]
  wire [7:0] level_intpend_id_1_10 = out_id_10; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30 pic_ctrl.scala 248:43]
  wire [7:0] out_id_22 = _T_2010 ? level_intpend_id_1_11 : level_intpend_id_1_10; // @[pic_ctrl.scala 27:9]
  wire [3:0] out_priority_22 = _T_2010 ? out_priority_11 : out_priority_10; // @[pic_ctrl.scala 27:49]
  wire  _T_2012 = out_priority_12 < out_priority_13; // @[pic_ctrl.scala 27:20]
  wire [7:0] level_intpend_id_1_13 = out_id_13; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30 pic_ctrl.scala 248:43]
  wire [7:0] level_intpend_id_1_12 = out_id_12; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30 pic_ctrl.scala 248:43]
  wire [7:0] out_id_23 = _T_2012 ? level_intpend_id_1_13 : level_intpend_id_1_12; // @[pic_ctrl.scala 27:9]
  wire [3:0] out_priority_23 = _T_2012 ? out_priority_13 : out_priority_12; // @[pic_ctrl.scala 27:49]
  wire  _T_2014 = out_priority_14 < out_priority_15; // @[pic_ctrl.scala 27:20]
  wire [7:0] level_intpend_id_1_15 = out_id_15; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30 pic_ctrl.scala 248:43]
  wire [7:0] level_intpend_id_1_14 = out_id_14; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30 pic_ctrl.scala 248:43]
  wire [7:0] out_id_24 = _T_2014 ? level_intpend_id_1_15 : level_intpend_id_1_14; // @[pic_ctrl.scala 27:9]
  wire [3:0] out_priority_24 = _T_2014 ? out_priority_15 : out_priority_14; // @[pic_ctrl.scala 27:49]
  wire [7:0] level_intpend_id_1_17 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30 pic_ctrl.scala 245:46]
  wire [7:0] level_intpend_id_1_16 = out_id_16; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30 pic_ctrl.scala 248:43]
  wire [7:0] out_id_25 = level_intpend_id_1_16; // @[pic_ctrl.scala 27:9]
  wire  _T_2018 = out_priority_17 < out_priority_18; // @[pic_ctrl.scala 27:20]
  wire [7:0] level_intpend_id_2_1 = out_id_18; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30 pic_ctrl.scala 248:43]
  wire [7:0] level_intpend_id_2_0 = out_id_17; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30 pic_ctrl.scala 248:43]
  wire [7:0] out_id_26 = _T_2018 ? level_intpend_id_2_1 : level_intpend_id_2_0; // @[pic_ctrl.scala 27:9]
  wire [3:0] out_priority_26 = _T_2018 ? out_priority_18 : out_priority_17; // @[pic_ctrl.scala 27:49]
  wire  _T_2020 = out_priority_19 < out_priority_20; // @[pic_ctrl.scala 27:20]
  wire [7:0] level_intpend_id_2_3 = out_id_20; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30 pic_ctrl.scala 248:43]
  wire [7:0] level_intpend_id_2_2 = out_id_19; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30 pic_ctrl.scala 248:43]
  wire [7:0] out_id_27 = _T_2020 ? level_intpend_id_2_3 : level_intpend_id_2_2; // @[pic_ctrl.scala 27:9]
  wire [3:0] out_priority_27 = _T_2020 ? out_priority_20 : out_priority_19; // @[pic_ctrl.scala 27:49]
  wire  _T_2022 = out_priority_21 < out_priority_22; // @[pic_ctrl.scala 27:20]
  wire [7:0] level_intpend_id_2_5 = out_id_22; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30 pic_ctrl.scala 248:43]
  wire [7:0] level_intpend_id_2_4 = out_id_21; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30 pic_ctrl.scala 248:43]
  wire [7:0] out_id_28 = _T_2022 ? level_intpend_id_2_5 : level_intpend_id_2_4; // @[pic_ctrl.scala 27:9]
  wire [3:0] out_priority_28 = _T_2022 ? out_priority_22 : out_priority_21; // @[pic_ctrl.scala 27:49]
  wire  _T_2024 = out_priority_23 < out_priority_24; // @[pic_ctrl.scala 27:20]
  wire [7:0] level_intpend_id_2_7 = out_id_24; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30 pic_ctrl.scala 248:43]
  wire [7:0] level_intpend_id_2_6 = out_id_23; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30 pic_ctrl.scala 248:43]
  wire [7:0] out_id_29 = _T_2024 ? level_intpend_id_2_7 : level_intpend_id_2_6; // @[pic_ctrl.scala 27:9]
  wire [3:0] out_priority_29 = _T_2024 ? out_priority_24 : out_priority_23; // @[pic_ctrl.scala 27:49]
  wire [7:0] level_intpend_id_2_9 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30 pic_ctrl.scala 245:46]
  wire [7:0] level_intpend_id_2_8 = level_intpend_id_1_16; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30 pic_ctrl.scala 248:43]
  wire [7:0] out_id_30 = out_id_25; // @[pic_ctrl.scala 27:9]
  wire  _T_2028 = out_priority_26 < out_priority_27; // @[pic_ctrl.scala 27:20]
  wire [7:0] level_intpend_id_3_1 = out_id_27; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30 pic_ctrl.scala 248:43]
  wire [7:0] level_intpend_id_3_0 = out_id_26; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30 pic_ctrl.scala 248:43]
  wire [7:0] out_id_31 = _T_2028 ? level_intpend_id_3_1 : level_intpend_id_3_0; // @[pic_ctrl.scala 27:9]
  wire [3:0] out_priority_31 = _T_2028 ? out_priority_27 : out_priority_26; // @[pic_ctrl.scala 27:49]
  wire  _T_2030 = out_priority_28 < out_priority_29; // @[pic_ctrl.scala 27:20]
  wire [7:0] level_intpend_id_3_3 = out_id_29; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30 pic_ctrl.scala 248:43]
  wire [7:0] level_intpend_id_3_2 = out_id_28; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30 pic_ctrl.scala 248:43]
  wire [7:0] out_id_32 = _T_2030 ? level_intpend_id_3_3 : level_intpend_id_3_2; // @[pic_ctrl.scala 27:9]
  wire [3:0] out_priority_32 = _T_2030 ? out_priority_29 : out_priority_28; // @[pic_ctrl.scala 27:49]
  wire [7:0] level_intpend_id_3_5 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30 pic_ctrl.scala 245:46]
  wire [7:0] level_intpend_id_3_4 = out_id_25; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30 pic_ctrl.scala 248:43]
  wire [7:0] out_id_33 = out_id_30; // @[pic_ctrl.scala 27:9]
  wire  _T_2034 = out_priority_31 < out_priority_32; // @[pic_ctrl.scala 27:20]
  wire [7:0] level_intpend_id_4_1 = out_id_32; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30 pic_ctrl.scala 248:43]
  wire [7:0] level_intpend_id_4_0 = out_id_31; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30 pic_ctrl.scala 248:43]
  wire [7:0] out_id_34 = _T_2034 ? level_intpend_id_4_1 : level_intpend_id_4_0; // @[pic_ctrl.scala 27:9]
  wire [3:0] out_priority_34 = _T_2034 ? out_priority_32 : out_priority_31; // @[pic_ctrl.scala 27:49]
  wire [7:0] level_intpend_id_4_3 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30 pic_ctrl.scala 245:46]
  wire [7:0] level_intpend_id_4_2 = out_id_30; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30 pic_ctrl.scala 248:43]
  wire  config_reg_we = waddr_config_pic_match & picm_wren_ff; // @[pic_ctrl.scala 265:47]
  wire  config_reg_re = raddr_config_pic_match & picm_rden_ff; // @[pic_ctrl.scala 266:47]
  wire [3:0] level_intpend_w_prior_en_5_0 = out_priority_34; // @[pic_ctrl.scala 229:40 pic_ctrl.scala 233:38 pic_ctrl.scala 249:43]
  wire [3:0] selected_int_priority = out_priority_34; // @[pic_ctrl.scala 253:29]
  wire [3:0] _T_2041 = ~level_intpend_w_prior_en_5_0; // @[pic_ctrl.scala 277:38]
  wire [3:0] pl_in_q = config_reg ? _T_2041 : level_intpend_w_prior_en_5_0; // @[pic_ctrl.scala 277:20]
  reg [7:0] _T_2042; // @[pic_ctrl.scala 278:59]
  reg [3:0] _T_2043; // @[pic_ctrl.scala 279:54]
  wire [3:0] _T_2045 = ~io_dec_pic_dec_tlu_meipt; // @[pic_ctrl.scala 280:40]
  wire [3:0] meipt_inv = config_reg ? _T_2045 : io_dec_pic_dec_tlu_meipt; // @[pic_ctrl.scala 280:22]
  wire [3:0] _T_2047 = ~io_dec_pic_dec_tlu_meicurpl; // @[pic_ctrl.scala 281:43]
  wire [3:0] meicurpl_inv = config_reg ? _T_2047 : io_dec_pic_dec_tlu_meicurpl; // @[pic_ctrl.scala 281:25]
  wire  _T_2048 = level_intpend_w_prior_en_5_0 > meipt_inv; // @[pic_ctrl.scala 282:47]
  wire  _T_2049 = level_intpend_w_prior_en_5_0 > meicurpl_inv; // @[pic_ctrl.scala 282:86]
  reg  _T_2050; // @[pic_ctrl.scala 283:58]
  wire [3:0] maxint = config_reg ? 4'h0 : 4'hf; // @[pic_ctrl.scala 284:19]
  reg  _T_2052; // @[pic_ctrl.scala 286:56]
  wire  intpend_reg_read = addr_intpend_base_match & picm_rden_ff; // @[pic_ctrl.scala 292:60]
  wire [9:0] _T_2062 = {extintsrc_req_gw_31,extintsrc_req_gw_30,extintsrc_req_gw_29,extintsrc_req_gw_28,extintsrc_req_gw_27,extintsrc_req_gw_26,extintsrc_req_gw_25,extintsrc_req_gw_24,extintsrc_req_gw_23,extintsrc_req_gw_22}; // @[Cat.scala 29:58]
  wire [18:0] _T_2071 = {_T_2062,extintsrc_req_gw_21,extintsrc_req_gw_20,extintsrc_req_gw_19,extintsrc_req_gw_18,extintsrc_req_gw_17,extintsrc_req_gw_16,extintsrc_req_gw_15,extintsrc_req_gw_14,extintsrc_req_gw_13}; // @[Cat.scala 29:58]
  wire [27:0] _T_2080 = {_T_2071,extintsrc_req_gw_12,extintsrc_req_gw_11,extintsrc_req_gw_10,extintsrc_req_gw_9,extintsrc_req_gw_8,extintsrc_req_gw_7,extintsrc_req_gw_6,extintsrc_req_gw_5,extintsrc_req_gw_4}; // @[Cat.scala 29:58]
  wire [63:0] intpend_reg_extended = {32'h0,_T_2080,extintsrc_req_gw_3,extintsrc_req_gw_2,extintsrc_req_gw_1,1'h0}; // @[Cat.scala 29:58]
  wire  _T_2087 = picm_raddr_ff[5:2] == 4'h0; // @[pic_ctrl.scala 300:105]
  wire  _T_2088 = intpend_reg_read & _T_2087; // @[pic_ctrl.scala 300:83]
  wire [31:0] _T_2090 = _T_2088 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] intpend_rd_part_out_0 = _T_2090 & intpend_reg_extended[31:0]; // @[pic_ctrl.scala 300:121]
  wire  _T_2094 = picm_raddr_ff[5:2] == 4'h1; // @[pic_ctrl.scala 300:105]
  wire  _T_2095 = intpend_reg_read & _T_2094; // @[pic_ctrl.scala 300:83]
  wire [31:0] _T_2097 = _T_2095 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] intpend_rd_part_out_1 = _T_2097 & intpend_reg_extended[63:32]; // @[pic_ctrl.scala 300:121]
  wire [31:0] intpend_rd_out = intpend_rd_part_out_0 | intpend_rd_part_out_1; // @[pic_ctrl.scala 301:58]
  wire  _T_2132 = intenable_reg_re_31 & intenable_reg_31; // @[Mux.scala 98:16]
  wire  _T_2133 = intenable_reg_re_30 ? intenable_reg_30 : _T_2132; // @[Mux.scala 98:16]
  wire  _T_2134 = intenable_reg_re_29 ? intenable_reg_29 : _T_2133; // @[Mux.scala 98:16]
  wire  _T_2135 = intenable_reg_re_28 ? intenable_reg_28 : _T_2134; // @[Mux.scala 98:16]
  wire  _T_2136 = intenable_reg_re_27 ? intenable_reg_27 : _T_2135; // @[Mux.scala 98:16]
  wire  _T_2137 = intenable_reg_re_26 ? intenable_reg_26 : _T_2136; // @[Mux.scala 98:16]
  wire  _T_2138 = intenable_reg_re_25 ? intenable_reg_25 : _T_2137; // @[Mux.scala 98:16]
  wire  _T_2139 = intenable_reg_re_24 ? intenable_reg_24 : _T_2138; // @[Mux.scala 98:16]
  wire  _T_2140 = intenable_reg_re_23 ? intenable_reg_23 : _T_2139; // @[Mux.scala 98:16]
  wire  _T_2141 = intenable_reg_re_22 ? intenable_reg_22 : _T_2140; // @[Mux.scala 98:16]
  wire  _T_2142 = intenable_reg_re_21 ? intenable_reg_21 : _T_2141; // @[Mux.scala 98:16]
  wire  _T_2143 = intenable_reg_re_20 ? intenable_reg_20 : _T_2142; // @[Mux.scala 98:16]
  wire  _T_2144 = intenable_reg_re_19 ? intenable_reg_19 : _T_2143; // @[Mux.scala 98:16]
  wire  _T_2145 = intenable_reg_re_18 ? intenable_reg_18 : _T_2144; // @[Mux.scala 98:16]
  wire  _T_2146 = intenable_reg_re_17 ? intenable_reg_17 : _T_2145; // @[Mux.scala 98:16]
  wire  _T_2147 = intenable_reg_re_16 ? intenable_reg_16 : _T_2146; // @[Mux.scala 98:16]
  wire  _T_2148 = intenable_reg_re_15 ? intenable_reg_15 : _T_2147; // @[Mux.scala 98:16]
  wire  _T_2149 = intenable_reg_re_14 ? intenable_reg_14 : _T_2148; // @[Mux.scala 98:16]
  wire  _T_2150 = intenable_reg_re_13 ? intenable_reg_13 : _T_2149; // @[Mux.scala 98:16]
  wire  _T_2151 = intenable_reg_re_12 ? intenable_reg_12 : _T_2150; // @[Mux.scala 98:16]
  wire  _T_2152 = intenable_reg_re_11 ? intenable_reg_11 : _T_2151; // @[Mux.scala 98:16]
  wire  _T_2153 = intenable_reg_re_10 ? intenable_reg_10 : _T_2152; // @[Mux.scala 98:16]
  wire  _T_2154 = intenable_reg_re_9 ? intenable_reg_9 : _T_2153; // @[Mux.scala 98:16]
  wire  _T_2155 = intenable_reg_re_8 ? intenable_reg_8 : _T_2154; // @[Mux.scala 98:16]
  wire  _T_2156 = intenable_reg_re_7 ? intenable_reg_7 : _T_2155; // @[Mux.scala 98:16]
  wire  _T_2157 = intenable_reg_re_6 ? intenable_reg_6 : _T_2156; // @[Mux.scala 98:16]
  wire  _T_2158 = intenable_reg_re_5 ? intenable_reg_5 : _T_2157; // @[Mux.scala 98:16]
  wire  _T_2159 = intenable_reg_re_4 ? intenable_reg_4 : _T_2158; // @[Mux.scala 98:16]
  wire  _T_2160 = intenable_reg_re_3 ? intenable_reg_3 : _T_2159; // @[Mux.scala 98:16]
  wire  _T_2161 = intenable_reg_re_2 ? intenable_reg_2 : _T_2160; // @[Mux.scala 98:16]
  wire  intenable_rd_out = intenable_reg_re_1 ? intenable_reg_1 : _T_2161; // @[Mux.scala 98:16]
  wire [3:0] _T_2194 = intpriority_reg_re_31 ? intpriority_reg_31 : 4'h0; // @[Mux.scala 98:16]
  wire [3:0] _T_2195 = intpriority_reg_re_30 ? intpriority_reg_30 : _T_2194; // @[Mux.scala 98:16]
  wire [3:0] _T_2196 = intpriority_reg_re_29 ? intpriority_reg_29 : _T_2195; // @[Mux.scala 98:16]
  wire [3:0] _T_2197 = intpriority_reg_re_28 ? intpriority_reg_28 : _T_2196; // @[Mux.scala 98:16]
  wire [3:0] _T_2198 = intpriority_reg_re_27 ? intpriority_reg_27 : _T_2197; // @[Mux.scala 98:16]
  wire [3:0] _T_2199 = intpriority_reg_re_26 ? intpriority_reg_26 : _T_2198; // @[Mux.scala 98:16]
  wire [3:0] _T_2200 = intpriority_reg_re_25 ? intpriority_reg_25 : _T_2199; // @[Mux.scala 98:16]
  wire [3:0] _T_2201 = intpriority_reg_re_24 ? intpriority_reg_24 : _T_2200; // @[Mux.scala 98:16]
  wire [3:0] _T_2202 = intpriority_reg_re_23 ? intpriority_reg_23 : _T_2201; // @[Mux.scala 98:16]
  wire [3:0] _T_2203 = intpriority_reg_re_22 ? intpriority_reg_22 : _T_2202; // @[Mux.scala 98:16]
  wire [3:0] _T_2204 = intpriority_reg_re_21 ? intpriority_reg_21 : _T_2203; // @[Mux.scala 98:16]
  wire [3:0] _T_2205 = intpriority_reg_re_20 ? intpriority_reg_20 : _T_2204; // @[Mux.scala 98:16]
  wire [3:0] _T_2206 = intpriority_reg_re_19 ? intpriority_reg_19 : _T_2205; // @[Mux.scala 98:16]
  wire [3:0] _T_2207 = intpriority_reg_re_18 ? intpriority_reg_18 : _T_2206; // @[Mux.scala 98:16]
  wire [3:0] _T_2208 = intpriority_reg_re_17 ? intpriority_reg_17 : _T_2207; // @[Mux.scala 98:16]
  wire [3:0] _T_2209 = intpriority_reg_re_16 ? intpriority_reg_16 : _T_2208; // @[Mux.scala 98:16]
  wire [3:0] _T_2210 = intpriority_reg_re_15 ? intpriority_reg_15 : _T_2209; // @[Mux.scala 98:16]
  wire [3:0] _T_2211 = intpriority_reg_re_14 ? intpriority_reg_14 : _T_2210; // @[Mux.scala 98:16]
  wire [3:0] _T_2212 = intpriority_reg_re_13 ? intpriority_reg_13 : _T_2211; // @[Mux.scala 98:16]
  wire [3:0] _T_2213 = intpriority_reg_re_12 ? intpriority_reg_12 : _T_2212; // @[Mux.scala 98:16]
  wire [3:0] _T_2214 = intpriority_reg_re_11 ? intpriority_reg_11 : _T_2213; // @[Mux.scala 98:16]
  wire [3:0] _T_2215 = intpriority_reg_re_10 ? intpriority_reg_10 : _T_2214; // @[Mux.scala 98:16]
  wire [3:0] _T_2216 = intpriority_reg_re_9 ? intpriority_reg_9 : _T_2215; // @[Mux.scala 98:16]
  wire [3:0] _T_2217 = intpriority_reg_re_8 ? intpriority_reg_8 : _T_2216; // @[Mux.scala 98:16]
  wire [3:0] _T_2218 = intpriority_reg_re_7 ? intpriority_reg_7 : _T_2217; // @[Mux.scala 98:16]
  wire [3:0] _T_2219 = intpriority_reg_re_6 ? intpriority_reg_6 : _T_2218; // @[Mux.scala 98:16]
  wire [3:0] _T_2220 = intpriority_reg_re_5 ? intpriority_reg_5 : _T_2219; // @[Mux.scala 98:16]
  wire [3:0] _T_2221 = intpriority_reg_re_4 ? intpriority_reg_4 : _T_2220; // @[Mux.scala 98:16]
  wire [3:0] _T_2222 = intpriority_reg_re_3 ? intpriority_reg_3 : _T_2221; // @[Mux.scala 98:16]
  wire [3:0] _T_2223 = intpriority_reg_re_2 ? intpriority_reg_2 : _T_2222; // @[Mux.scala 98:16]
  wire [3:0] intpriority_rd_out = intpriority_reg_re_1 ? intpriority_reg_1 : _T_2223; // @[Mux.scala 98:16]
  wire [1:0] _T_2256 = gw_config_reg_re_31 ? gw_config_reg_31 : 2'h0; // @[Mux.scala 98:16]
  wire [1:0] _T_2257 = gw_config_reg_re_30 ? gw_config_reg_30 : _T_2256; // @[Mux.scala 98:16]
  wire [1:0] _T_2258 = gw_config_reg_re_29 ? gw_config_reg_29 : _T_2257; // @[Mux.scala 98:16]
  wire [1:0] _T_2259 = gw_config_reg_re_28 ? gw_config_reg_28 : _T_2258; // @[Mux.scala 98:16]
  wire [1:0] _T_2260 = gw_config_reg_re_27 ? gw_config_reg_27 : _T_2259; // @[Mux.scala 98:16]
  wire [1:0] _T_2261 = gw_config_reg_re_26 ? gw_config_reg_26 : _T_2260; // @[Mux.scala 98:16]
  wire [1:0] _T_2262 = gw_config_reg_re_25 ? gw_config_reg_25 : _T_2261; // @[Mux.scala 98:16]
  wire [1:0] _T_2263 = gw_config_reg_re_24 ? gw_config_reg_24 : _T_2262; // @[Mux.scala 98:16]
  wire [1:0] _T_2264 = gw_config_reg_re_23 ? gw_config_reg_23 : _T_2263; // @[Mux.scala 98:16]
  wire [1:0] _T_2265 = gw_config_reg_re_22 ? gw_config_reg_22 : _T_2264; // @[Mux.scala 98:16]
  wire [1:0] _T_2266 = gw_config_reg_re_21 ? gw_config_reg_21 : _T_2265; // @[Mux.scala 98:16]
  wire [1:0] _T_2267 = gw_config_reg_re_20 ? gw_config_reg_20 : _T_2266; // @[Mux.scala 98:16]
  wire [1:0] _T_2268 = gw_config_reg_re_19 ? gw_config_reg_19 : _T_2267; // @[Mux.scala 98:16]
  wire [1:0] _T_2269 = gw_config_reg_re_18 ? gw_config_reg_18 : _T_2268; // @[Mux.scala 98:16]
  wire [1:0] _T_2270 = gw_config_reg_re_17 ? gw_config_reg_17 : _T_2269; // @[Mux.scala 98:16]
  wire [1:0] _T_2271 = gw_config_reg_re_16 ? gw_config_reg_16 : _T_2270; // @[Mux.scala 98:16]
  wire [1:0] _T_2272 = gw_config_reg_re_15 ? gw_config_reg_15 : _T_2271; // @[Mux.scala 98:16]
  wire [1:0] _T_2273 = gw_config_reg_re_14 ? gw_config_reg_14 : _T_2272; // @[Mux.scala 98:16]
  wire [1:0] _T_2274 = gw_config_reg_re_13 ? gw_config_reg_13 : _T_2273; // @[Mux.scala 98:16]
  wire [1:0] _T_2275 = gw_config_reg_re_12 ? gw_config_reg_12 : _T_2274; // @[Mux.scala 98:16]
  wire [1:0] _T_2276 = gw_config_reg_re_11 ? gw_config_reg_11 : _T_2275; // @[Mux.scala 98:16]
  wire [1:0] _T_2277 = gw_config_reg_re_10 ? gw_config_reg_10 : _T_2276; // @[Mux.scala 98:16]
  wire [1:0] _T_2278 = gw_config_reg_re_9 ? gw_config_reg_9 : _T_2277; // @[Mux.scala 98:16]
  wire [1:0] _T_2279 = gw_config_reg_re_8 ? gw_config_reg_8 : _T_2278; // @[Mux.scala 98:16]
  wire [1:0] _T_2280 = gw_config_reg_re_7 ? gw_config_reg_7 : _T_2279; // @[Mux.scala 98:16]
  wire [1:0] _T_2281 = gw_config_reg_re_6 ? gw_config_reg_6 : _T_2280; // @[Mux.scala 98:16]
  wire [1:0] _T_2282 = gw_config_reg_re_5 ? gw_config_reg_5 : _T_2281; // @[Mux.scala 98:16]
  wire [1:0] _T_2283 = gw_config_reg_re_4 ? gw_config_reg_4 : _T_2282; // @[Mux.scala 98:16]
  wire [1:0] _T_2284 = gw_config_reg_re_3 ? gw_config_reg_3 : _T_2283; // @[Mux.scala 98:16]
  wire [1:0] _T_2285 = gw_config_reg_re_2 ? gw_config_reg_2 : _T_2284; // @[Mux.scala 98:16]
  wire [1:0] gw_config_rd_out = gw_config_reg_re_1 ? gw_config_reg_1 : _T_2285; // @[Mux.scala 98:16]
  wire [31:0] _T_2290 = {28'h0,intpriority_rd_out}; // @[Cat.scala 29:58]
  wire [31:0] _T_2293 = {31'h0,intenable_rd_out}; // @[Cat.scala 29:58]
  wire [31:0] _T_2296 = {30'h0,gw_config_rd_out}; // @[Cat.scala 29:58]
  wire [31:0] _T_2299 = {31'h0,config_reg}; // @[Cat.scala 29:58]
  wire [14:0] address = picm_raddr_ff[14:0]; // @[pic_ctrl.scala 322:30]
  wire  _T_2339 = 15'h3000 == address; // @[Conditional.scala 37:30]
  wire  _T_2340 = 15'h4004 == address; // @[Conditional.scala 37:30]
  wire  _T_2341 = 15'h4008 == address; // @[Conditional.scala 37:30]
  wire  _T_2342 = 15'h400c == address; // @[Conditional.scala 37:30]
  wire  _T_2343 = 15'h4010 == address; // @[Conditional.scala 37:30]
  wire  _T_2344 = 15'h4014 == address; // @[Conditional.scala 37:30]
  wire  _T_2345 = 15'h4018 == address; // @[Conditional.scala 37:30]
  wire  _T_2346 = 15'h401c == address; // @[Conditional.scala 37:30]
  wire  _T_2347 = 15'h4020 == address; // @[Conditional.scala 37:30]
  wire  _T_2348 = 15'h4024 == address; // @[Conditional.scala 37:30]
  wire  _T_2349 = 15'h4028 == address; // @[Conditional.scala 37:30]
  wire  _T_2350 = 15'h402c == address; // @[Conditional.scala 37:30]
  wire  _T_2351 = 15'h4030 == address; // @[Conditional.scala 37:30]
  wire  _T_2352 = 15'h4034 == address; // @[Conditional.scala 37:30]
  wire  _T_2353 = 15'h4038 == address; // @[Conditional.scala 37:30]
  wire  _T_2354 = 15'h403c == address; // @[Conditional.scala 37:30]
  wire  _T_2355 = 15'h4040 == address; // @[Conditional.scala 37:30]
  wire  _T_2356 = 15'h4044 == address; // @[Conditional.scala 37:30]
  wire  _T_2357 = 15'h4048 == address; // @[Conditional.scala 37:30]
  wire  _T_2358 = 15'h404c == address; // @[Conditional.scala 37:30]
  wire  _T_2359 = 15'h4050 == address; // @[Conditional.scala 37:30]
  wire  _T_2360 = 15'h4054 == address; // @[Conditional.scala 37:30]
  wire  _T_2361 = 15'h4058 == address; // @[Conditional.scala 37:30]
  wire  _T_2362 = 15'h405c == address; // @[Conditional.scala 37:30]
  wire  _T_2363 = 15'h4060 == address; // @[Conditional.scala 37:30]
  wire  _T_2364 = 15'h4064 == address; // @[Conditional.scala 37:30]
  wire  _T_2365 = 15'h4068 == address; // @[Conditional.scala 37:30]
  wire  _T_2366 = 15'h406c == address; // @[Conditional.scala 37:30]
  wire  _T_2367 = 15'h4070 == address; // @[Conditional.scala 37:30]
  wire  _T_2368 = 15'h4074 == address; // @[Conditional.scala 37:30]
  wire  _T_2369 = 15'h4078 == address; // @[Conditional.scala 37:30]
  wire  _T_2370 = 15'h407c == address; // @[Conditional.scala 37:30]
  wire  _T_2371 = 15'h2004 == address; // @[Conditional.scala 37:30]
  wire  _T_2372 = 15'h2008 == address; // @[Conditional.scala 37:30]
  wire  _T_2373 = 15'h200c == address; // @[Conditional.scala 37:30]
  wire  _T_2374 = 15'h2010 == address; // @[Conditional.scala 37:30]
  wire  _T_2375 = 15'h2014 == address; // @[Conditional.scala 37:30]
  wire  _T_2376 = 15'h2018 == address; // @[Conditional.scala 37:30]
  wire  _T_2377 = 15'h201c == address; // @[Conditional.scala 37:30]
  wire  _T_2378 = 15'h2020 == address; // @[Conditional.scala 37:30]
  wire  _T_2379 = 15'h2024 == address; // @[Conditional.scala 37:30]
  wire  _T_2380 = 15'h2028 == address; // @[Conditional.scala 37:30]
  wire  _T_2381 = 15'h202c == address; // @[Conditional.scala 37:30]
  wire  _T_2382 = 15'h2030 == address; // @[Conditional.scala 37:30]
  wire  _T_2383 = 15'h2034 == address; // @[Conditional.scala 37:30]
  wire  _T_2384 = 15'h2038 == address; // @[Conditional.scala 37:30]
  wire  _T_2385 = 15'h203c == address; // @[Conditional.scala 37:30]
  wire  _T_2386 = 15'h2040 == address; // @[Conditional.scala 37:30]
  wire  _T_2387 = 15'h2044 == address; // @[Conditional.scala 37:30]
  wire  _T_2388 = 15'h2048 == address; // @[Conditional.scala 37:30]
  wire  _T_2389 = 15'h204c == address; // @[Conditional.scala 37:30]
  wire  _T_2390 = 15'h2050 == address; // @[Conditional.scala 37:30]
  wire  _T_2391 = 15'h2054 == address; // @[Conditional.scala 37:30]
  wire  _T_2392 = 15'h2058 == address; // @[Conditional.scala 37:30]
  wire  _T_2393 = 15'h205c == address; // @[Conditional.scala 37:30]
  wire  _T_2394 = 15'h2060 == address; // @[Conditional.scala 37:30]
  wire  _T_2395 = 15'h2064 == address; // @[Conditional.scala 37:30]
  wire  _T_2396 = 15'h2068 == address; // @[Conditional.scala 37:30]
  wire  _T_2397 = 15'h206c == address; // @[Conditional.scala 37:30]
  wire  _T_2398 = 15'h2070 == address; // @[Conditional.scala 37:30]
  wire  _T_2399 = 15'h2074 == address; // @[Conditional.scala 37:30]
  wire  _T_2400 = 15'h2078 == address; // @[Conditional.scala 37:30]
  wire  _T_2401 = 15'h207c == address; // @[Conditional.scala 37:30]
  wire  _T_2402 = 15'h4 == address; // @[Conditional.scala 37:30]
  wire  _T_2403 = 15'h8 == address; // @[Conditional.scala 37:30]
  wire  _T_2404 = 15'hc == address; // @[Conditional.scala 37:30]
  wire  _T_2405 = 15'h10 == address; // @[Conditional.scala 37:30]
  wire  _T_2406 = 15'h14 == address; // @[Conditional.scala 37:30]
  wire  _T_2407 = 15'h18 == address; // @[Conditional.scala 37:30]
  wire  _T_2408 = 15'h1c == address; // @[Conditional.scala 37:30]
  wire  _T_2409 = 15'h20 == address; // @[Conditional.scala 37:30]
  wire  _T_2410 = 15'h24 == address; // @[Conditional.scala 37:30]
  wire  _T_2411 = 15'h28 == address; // @[Conditional.scala 37:30]
  wire  _T_2412 = 15'h2c == address; // @[Conditional.scala 37:30]
  wire  _T_2413 = 15'h30 == address; // @[Conditional.scala 37:30]
  wire  _T_2414 = 15'h34 == address; // @[Conditional.scala 37:30]
  wire  _T_2415 = 15'h38 == address; // @[Conditional.scala 37:30]
  wire  _T_2416 = 15'h3c == address; // @[Conditional.scala 37:30]
  wire  _T_2417 = 15'h40 == address; // @[Conditional.scala 37:30]
  wire  _T_2418 = 15'h44 == address; // @[Conditional.scala 37:30]
  wire  _T_2419 = 15'h48 == address; // @[Conditional.scala 37:30]
  wire  _T_2420 = 15'h4c == address; // @[Conditional.scala 37:30]
  wire  _T_2421 = 15'h50 == address; // @[Conditional.scala 37:30]
  wire  _T_2422 = 15'h54 == address; // @[Conditional.scala 37:30]
  wire  _T_2423 = 15'h58 == address; // @[Conditional.scala 37:30]
  wire  _T_2424 = 15'h5c == address; // @[Conditional.scala 37:30]
  wire  _T_2425 = 15'h60 == address; // @[Conditional.scala 37:30]
  wire  _T_2426 = 15'h64 == address; // @[Conditional.scala 37:30]
  wire  _T_2427 = 15'h68 == address; // @[Conditional.scala 37:30]
  wire  _T_2428 = 15'h6c == address; // @[Conditional.scala 37:30]
  wire  _T_2429 = 15'h70 == address; // @[Conditional.scala 37:30]
  wire  _T_2430 = 15'h74 == address; // @[Conditional.scala 37:30]
  wire  _T_2431 = 15'h78 == address; // @[Conditional.scala 37:30]
  wire  _T_2432 = 15'h7c == address; // @[Conditional.scala 37:30]
  wire [3:0] _GEN_187 = _T_2432 ? 4'h2 : 4'h1; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_188 = _T_2431 ? 4'h2 : _GEN_187; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_189 = _T_2430 ? 4'h2 : _GEN_188; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_190 = _T_2429 ? 4'h2 : _GEN_189; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_191 = _T_2428 ? 4'h2 : _GEN_190; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_192 = _T_2427 ? 4'h2 : _GEN_191; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_193 = _T_2426 ? 4'h2 : _GEN_192; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_194 = _T_2425 ? 4'h2 : _GEN_193; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_195 = _T_2424 ? 4'h2 : _GEN_194; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_196 = _T_2423 ? 4'h2 : _GEN_195; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_197 = _T_2422 ? 4'h2 : _GEN_196; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_198 = _T_2421 ? 4'h2 : _GEN_197; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_199 = _T_2420 ? 4'h2 : _GEN_198; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_200 = _T_2419 ? 4'h2 : _GEN_199; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_201 = _T_2418 ? 4'h2 : _GEN_200; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_202 = _T_2417 ? 4'h2 : _GEN_201; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_203 = _T_2416 ? 4'h2 : _GEN_202; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_204 = _T_2415 ? 4'h2 : _GEN_203; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_205 = _T_2414 ? 4'h2 : _GEN_204; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_206 = _T_2413 ? 4'h2 : _GEN_205; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_207 = _T_2412 ? 4'h2 : _GEN_206; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_208 = _T_2411 ? 4'h2 : _GEN_207; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_209 = _T_2410 ? 4'h2 : _GEN_208; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_210 = _T_2409 ? 4'h2 : _GEN_209; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_211 = _T_2408 ? 4'h2 : _GEN_210; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_212 = _T_2407 ? 4'h2 : _GEN_211; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_213 = _T_2406 ? 4'h2 : _GEN_212; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_214 = _T_2405 ? 4'h2 : _GEN_213; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_215 = _T_2404 ? 4'h2 : _GEN_214; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_216 = _T_2403 ? 4'h2 : _GEN_215; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_217 = _T_2402 ? 4'h2 : _GEN_216; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_218 = _T_2401 ? 4'h4 : _GEN_217; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_219 = _T_2400 ? 4'h4 : _GEN_218; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_220 = _T_2399 ? 4'h4 : _GEN_219; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_221 = _T_2398 ? 4'h4 : _GEN_220; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_222 = _T_2397 ? 4'h4 : _GEN_221; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_223 = _T_2396 ? 4'h4 : _GEN_222; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_224 = _T_2395 ? 4'h4 : _GEN_223; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_225 = _T_2394 ? 4'h4 : _GEN_224; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_226 = _T_2393 ? 4'h4 : _GEN_225; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_227 = _T_2392 ? 4'h4 : _GEN_226; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_228 = _T_2391 ? 4'h4 : _GEN_227; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_229 = _T_2390 ? 4'h4 : _GEN_228; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_230 = _T_2389 ? 4'h4 : _GEN_229; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_231 = _T_2388 ? 4'h4 : _GEN_230; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_232 = _T_2387 ? 4'h4 : _GEN_231; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_233 = _T_2386 ? 4'h4 : _GEN_232; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_234 = _T_2385 ? 4'h4 : _GEN_233; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_235 = _T_2384 ? 4'h4 : _GEN_234; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_236 = _T_2383 ? 4'h4 : _GEN_235; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_237 = _T_2382 ? 4'h4 : _GEN_236; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_238 = _T_2381 ? 4'h4 : _GEN_237; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_239 = _T_2380 ? 4'h4 : _GEN_238; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_240 = _T_2379 ? 4'h4 : _GEN_239; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_241 = _T_2378 ? 4'h4 : _GEN_240; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_242 = _T_2377 ? 4'h4 : _GEN_241; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_243 = _T_2376 ? 4'h4 : _GEN_242; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_244 = _T_2375 ? 4'h4 : _GEN_243; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_245 = _T_2374 ? 4'h4 : _GEN_244; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_246 = _T_2373 ? 4'h4 : _GEN_245; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_247 = _T_2372 ? 4'h4 : _GEN_246; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_248 = _T_2371 ? 4'h4 : _GEN_247; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_249 = _T_2370 ? 4'h8 : _GEN_248; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_250 = _T_2369 ? 4'h8 : _GEN_249; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_251 = _T_2368 ? 4'h8 : _GEN_250; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_252 = _T_2367 ? 4'h8 : _GEN_251; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_253 = _T_2366 ? 4'h8 : _GEN_252; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_254 = _T_2365 ? 4'h8 : _GEN_253; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_255 = _T_2364 ? 4'h8 : _GEN_254; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_256 = _T_2363 ? 4'h8 : _GEN_255; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_257 = _T_2362 ? 4'h8 : _GEN_256; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_258 = _T_2361 ? 4'h8 : _GEN_257; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_259 = _T_2360 ? 4'h8 : _GEN_258; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_260 = _T_2359 ? 4'h8 : _GEN_259; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_261 = _T_2358 ? 4'h8 : _GEN_260; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_262 = _T_2357 ? 4'h8 : _GEN_261; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_263 = _T_2356 ? 4'h8 : _GEN_262; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_264 = _T_2355 ? 4'h8 : _GEN_263; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_265 = _T_2354 ? 4'h8 : _GEN_264; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_266 = _T_2353 ? 4'h8 : _GEN_265; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_267 = _T_2352 ? 4'h8 : _GEN_266; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_268 = _T_2351 ? 4'h8 : _GEN_267; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_269 = _T_2350 ? 4'h8 : _GEN_268; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_270 = _T_2349 ? 4'h8 : _GEN_269; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_271 = _T_2348 ? 4'h8 : _GEN_270; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_272 = _T_2347 ? 4'h8 : _GEN_271; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_273 = _T_2346 ? 4'h8 : _GEN_272; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_274 = _T_2345 ? 4'h8 : _GEN_273; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_275 = _T_2344 ? 4'h8 : _GEN_274; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_276 = _T_2343 ? 4'h8 : _GEN_275; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_277 = _T_2342 ? 4'h8 : _GEN_276; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_278 = _T_2341 ? 4'h8 : _GEN_277; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_279 = _T_2340 ? 4'h8 : _GEN_278; // @[Conditional.scala 39:67]
  wire [3:0] mask = _T_2339 ? 4'h4 : _GEN_279; // @[Conditional.scala 40:58]
  wire  _T_2301 = picm_mken_ff & mask[3]; // @[pic_ctrl.scala 315:19]
  wire  _T_2306 = picm_mken_ff & mask[2]; // @[pic_ctrl.scala 316:19]
  wire  _T_2311 = picm_mken_ff & mask[1]; // @[pic_ctrl.scala 317:19]
  wire [31:0] _T_2319 = intpend_reg_read ? intpend_rd_out : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2320 = _T_53 ? _T_2290 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2321 = _T_56 ? _T_2293 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2322 = _T_59 ? _T_2296 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2323 = config_reg_re ? _T_2299 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2324 = _T_2301 ? 32'h3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2325 = _T_2306 ? 32'h1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2326 = _T_2311 ? 32'hf : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2328 = _T_2319 | _T_2320; // @[Mux.scala 27:72]
  wire [31:0] _T_2329 = _T_2328 | _T_2321; // @[Mux.scala 27:72]
  wire [31:0] _T_2330 = _T_2329 | _T_2322; // @[Mux.scala 27:72]
  wire [31:0] _T_2331 = _T_2330 | _T_2323; // @[Mux.scala 27:72]
  wire [31:0] _T_2332 = _T_2331 | _T_2324; // @[Mux.scala 27:72]
  wire [31:0] _T_2333 = _T_2332 | _T_2325; // @[Mux.scala 27:72]
  wire [31:0] picm_rd_data_in = _T_2333 | _T_2326; // @[Mux.scala 27:72]
  wire [7:0] level_intpend_id_5_0 = out_id_34; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30 pic_ctrl.scala 248:43]
  wire [7:0] level_intpend_id_1_18 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_1_19 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_1_20 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_1_21 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_1_22 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_1_23 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_1_24 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_1_25 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_1_26 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_1_27 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_1_28 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_1_29 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_1_30 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_1_31 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_1_32 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_1_33 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_2_10 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_2_11 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_2_12 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_2_13 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_2_14 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_2_15 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_2_16 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_2_17 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_2_18 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_2_19 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_2_20 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_2_21 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_2_22 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_2_23 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_2_24 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_2_25 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_2_26 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_2_27 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_2_28 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_2_29 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_2_30 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_2_31 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_2_32 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_2_33 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_3_6 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_3_7 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_3_8 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_3_9 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_3_10 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_3_11 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_3_12 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_3_13 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_3_14 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_3_15 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_3_16 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_3_17 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_3_18 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_3_19 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_3_20 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_3_21 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_3_22 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_3_23 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_3_24 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_3_25 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_3_26 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_3_27 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_3_28 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_3_29 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_3_30 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_3_31 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_3_32 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_3_33 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_4_4 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_4_5 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_4_6 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_4_7 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_4_8 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_4_9 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_4_10 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_4_11 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_4_12 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_4_13 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_4_14 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_4_15 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_4_16 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_4_17 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_4_18 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_4_19 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_4_20 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_4_21 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_4_22 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_4_23 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_4_24 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_4_25 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_4_26 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_4_27 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_4_28 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_4_29 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_4_30 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_4_31 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_4_32 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_4_33 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_5_1 = out_id_33; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30 pic_ctrl.scala 248:43]
  wire [7:0] level_intpend_id_5_2 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30 pic_ctrl.scala 245:46]
  wire [7:0] level_intpend_id_5_3 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_5_4 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_5_5 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_5_6 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_5_7 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_5_8 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_5_9 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_5_10 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_5_11 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_5_12 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_5_13 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_5_14 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_5_15 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_5_16 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_5_17 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_5_18 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_5_19 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_5_20 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_5_21 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_5_22 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_5_23 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_5_24 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_5_25 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_5_26 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_5_27 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_5_28 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_5_29 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_5_30 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_5_31 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_5_32 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  wire [7:0] level_intpend_id_5_33 = 8'h0; // @[pic_ctrl.scala 230:32 pic_ctrl.scala 234:30]
  assign io_lsu_pic_picm_rd_data = picm_bypass_ff ? picm_wr_data_ff : picm_rd_data_in; // @[pic_ctrl.scala 321:27]
  assign io_dec_pic_pic_claimid = _T_2042; // @[pic_ctrl.scala 278:49]
  assign io_dec_pic_pic_pl = _T_2043; // @[pic_ctrl.scala 279:44]
  assign io_dec_pic_mhwakeup = _T_2052; // @[pic_ctrl.scala 286:23]
  assign io_dec_pic_mexintpend = _T_2050; // @[pic_ctrl.scala 283:25]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  picm_raddr_ff = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  picm_waddr_ff = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  picm_wren_ff = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  picm_rden_ff = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  picm_mken_ff = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  picm_wr_data_ff = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  gw_config_reg_31 = _RAND_6[1:0];
  _RAND_7 = {1{`RANDOM}};
  intenable_reg_31 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  gw_config_reg_30 = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  intenable_reg_30 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  gw_config_reg_29 = _RAND_10[1:0];
  _RAND_11 = {1{`RANDOM}};
  intenable_reg_29 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  gw_config_reg_28 = _RAND_12[1:0];
  _RAND_13 = {1{`RANDOM}};
  intenable_reg_28 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  gw_config_reg_27 = _RAND_14[1:0];
  _RAND_15 = {1{`RANDOM}};
  intenable_reg_27 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  gw_config_reg_26 = _RAND_16[1:0];
  _RAND_17 = {1{`RANDOM}};
  intenable_reg_26 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  gw_config_reg_25 = _RAND_18[1:0];
  _RAND_19 = {1{`RANDOM}};
  intenable_reg_25 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  gw_config_reg_24 = _RAND_20[1:0];
  _RAND_21 = {1{`RANDOM}};
  intenable_reg_24 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  gw_config_reg_23 = _RAND_22[1:0];
  _RAND_23 = {1{`RANDOM}};
  intenable_reg_23 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  gw_config_reg_22 = _RAND_24[1:0];
  _RAND_25 = {1{`RANDOM}};
  intenable_reg_22 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  gw_config_reg_21 = _RAND_26[1:0];
  _RAND_27 = {1{`RANDOM}};
  intenable_reg_21 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  gw_config_reg_20 = _RAND_28[1:0];
  _RAND_29 = {1{`RANDOM}};
  intenable_reg_20 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  gw_config_reg_19 = _RAND_30[1:0];
  _RAND_31 = {1{`RANDOM}};
  intenable_reg_19 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  gw_config_reg_18 = _RAND_32[1:0];
  _RAND_33 = {1{`RANDOM}};
  intenable_reg_18 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  gw_config_reg_17 = _RAND_34[1:0];
  _RAND_35 = {1{`RANDOM}};
  intenable_reg_17 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  gw_config_reg_16 = _RAND_36[1:0];
  _RAND_37 = {1{`RANDOM}};
  intenable_reg_16 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  gw_config_reg_15 = _RAND_38[1:0];
  _RAND_39 = {1{`RANDOM}};
  intenable_reg_15 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  gw_config_reg_14 = _RAND_40[1:0];
  _RAND_41 = {1{`RANDOM}};
  intenable_reg_14 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  gw_config_reg_13 = _RAND_42[1:0];
  _RAND_43 = {1{`RANDOM}};
  intenable_reg_13 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  gw_config_reg_12 = _RAND_44[1:0];
  _RAND_45 = {1{`RANDOM}};
  intenable_reg_12 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  gw_config_reg_11 = _RAND_46[1:0];
  _RAND_47 = {1{`RANDOM}};
  intenable_reg_11 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  gw_config_reg_10 = _RAND_48[1:0];
  _RAND_49 = {1{`RANDOM}};
  intenable_reg_10 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  gw_config_reg_9 = _RAND_50[1:0];
  _RAND_51 = {1{`RANDOM}};
  intenable_reg_9 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  gw_config_reg_8 = _RAND_52[1:0];
  _RAND_53 = {1{`RANDOM}};
  intenable_reg_8 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  gw_config_reg_7 = _RAND_54[1:0];
  _RAND_55 = {1{`RANDOM}};
  intenable_reg_7 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  gw_config_reg_6 = _RAND_56[1:0];
  _RAND_57 = {1{`RANDOM}};
  intenable_reg_6 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  gw_config_reg_5 = _RAND_58[1:0];
  _RAND_59 = {1{`RANDOM}};
  intenable_reg_5 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  gw_config_reg_4 = _RAND_60[1:0];
  _RAND_61 = {1{`RANDOM}};
  intenable_reg_4 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  gw_config_reg_3 = _RAND_62[1:0];
  _RAND_63 = {1{`RANDOM}};
  intenable_reg_3 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  gw_config_reg_2 = _RAND_64[1:0];
  _RAND_65 = {1{`RANDOM}};
  intenable_reg_2 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  gw_config_reg_1 = _RAND_66[1:0];
  _RAND_67 = {1{`RANDOM}};
  intenable_reg_1 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  _T_66 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  extintsrc_req_sync_1 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  _T_70 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  extintsrc_req_sync_2 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  _T_74 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  extintsrc_req_sync_3 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  _T_78 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  extintsrc_req_sync_4 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  _T_82 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  extintsrc_req_sync_5 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  _T_86 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  extintsrc_req_sync_6 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  _T_90 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  extintsrc_req_sync_7 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  _T_94 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  extintsrc_req_sync_8 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  _T_98 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  extintsrc_req_sync_9 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  _T_102 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  extintsrc_req_sync_10 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  _T_106 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  extintsrc_req_sync_11 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  _T_110 = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  extintsrc_req_sync_12 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  _T_114 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  extintsrc_req_sync_13 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  _T_118 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  extintsrc_req_sync_14 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  _T_122 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  extintsrc_req_sync_15 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  _T_126 = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  extintsrc_req_sync_16 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  _T_130 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  extintsrc_req_sync_17 = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  _T_134 = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  extintsrc_req_sync_18 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  _T_138 = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  extintsrc_req_sync_19 = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  _T_142 = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  extintsrc_req_sync_20 = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  _T_146 = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  extintsrc_req_sync_21 = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  _T_150 = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  extintsrc_req_sync_22 = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  _T_154 = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  extintsrc_req_sync_23 = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  _T_158 = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  extintsrc_req_sync_24 = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  _T_162 = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  extintsrc_req_sync_25 = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  _T_166 = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  extintsrc_req_sync_26 = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  _T_170 = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  extintsrc_req_sync_27 = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  _T_174 = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  extintsrc_req_sync_28 = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  _T_178 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  extintsrc_req_sync_29 = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  _T_182 = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  extintsrc_req_sync_30 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  _T_186 = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  extintsrc_req_sync_31 = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  intpriority_reg_1 = _RAND_130[3:0];
  _RAND_131 = {1{`RANDOM}};
  intpriority_reg_2 = _RAND_131[3:0];
  _RAND_132 = {1{`RANDOM}};
  intpriority_reg_3 = _RAND_132[3:0];
  _RAND_133 = {1{`RANDOM}};
  intpriority_reg_4 = _RAND_133[3:0];
  _RAND_134 = {1{`RANDOM}};
  intpriority_reg_5 = _RAND_134[3:0];
  _RAND_135 = {1{`RANDOM}};
  intpriority_reg_6 = _RAND_135[3:0];
  _RAND_136 = {1{`RANDOM}};
  intpriority_reg_7 = _RAND_136[3:0];
  _RAND_137 = {1{`RANDOM}};
  intpriority_reg_8 = _RAND_137[3:0];
  _RAND_138 = {1{`RANDOM}};
  intpriority_reg_9 = _RAND_138[3:0];
  _RAND_139 = {1{`RANDOM}};
  intpriority_reg_10 = _RAND_139[3:0];
  _RAND_140 = {1{`RANDOM}};
  intpriority_reg_11 = _RAND_140[3:0];
  _RAND_141 = {1{`RANDOM}};
  intpriority_reg_12 = _RAND_141[3:0];
  _RAND_142 = {1{`RANDOM}};
  intpriority_reg_13 = _RAND_142[3:0];
  _RAND_143 = {1{`RANDOM}};
  intpriority_reg_14 = _RAND_143[3:0];
  _RAND_144 = {1{`RANDOM}};
  intpriority_reg_15 = _RAND_144[3:0];
  _RAND_145 = {1{`RANDOM}};
  intpriority_reg_16 = _RAND_145[3:0];
  _RAND_146 = {1{`RANDOM}};
  intpriority_reg_17 = _RAND_146[3:0];
  _RAND_147 = {1{`RANDOM}};
  intpriority_reg_18 = _RAND_147[3:0];
  _RAND_148 = {1{`RANDOM}};
  intpriority_reg_19 = _RAND_148[3:0];
  _RAND_149 = {1{`RANDOM}};
  intpriority_reg_20 = _RAND_149[3:0];
  _RAND_150 = {1{`RANDOM}};
  intpriority_reg_21 = _RAND_150[3:0];
  _RAND_151 = {1{`RANDOM}};
  intpriority_reg_22 = _RAND_151[3:0];
  _RAND_152 = {1{`RANDOM}};
  intpriority_reg_23 = _RAND_152[3:0];
  _RAND_153 = {1{`RANDOM}};
  intpriority_reg_24 = _RAND_153[3:0];
  _RAND_154 = {1{`RANDOM}};
  intpriority_reg_25 = _RAND_154[3:0];
  _RAND_155 = {1{`RANDOM}};
  intpriority_reg_26 = _RAND_155[3:0];
  _RAND_156 = {1{`RANDOM}};
  intpriority_reg_27 = _RAND_156[3:0];
  _RAND_157 = {1{`RANDOM}};
  intpriority_reg_28 = _RAND_157[3:0];
  _RAND_158 = {1{`RANDOM}};
  intpriority_reg_29 = _RAND_158[3:0];
  _RAND_159 = {1{`RANDOM}};
  intpriority_reg_30 = _RAND_159[3:0];
  _RAND_160 = {1{`RANDOM}};
  intpriority_reg_31 = _RAND_160[3:0];
  _RAND_161 = {1{`RANDOM}};
  _T_1283 = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  _T_1298 = _RAND_162[0:0];
  _RAND_163 = {1{`RANDOM}};
  _T_1313 = _RAND_163[0:0];
  _RAND_164 = {1{`RANDOM}};
  _T_1328 = _RAND_164[0:0];
  _RAND_165 = {1{`RANDOM}};
  _T_1343 = _RAND_165[0:0];
  _RAND_166 = {1{`RANDOM}};
  _T_1358 = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  _T_1373 = _RAND_167[0:0];
  _RAND_168 = {1{`RANDOM}};
  _T_1388 = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  _T_1403 = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  _T_1418 = _RAND_170[0:0];
  _RAND_171 = {1{`RANDOM}};
  _T_1433 = _RAND_171[0:0];
  _RAND_172 = {1{`RANDOM}};
  _T_1448 = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  _T_1463 = _RAND_173[0:0];
  _RAND_174 = {1{`RANDOM}};
  _T_1478 = _RAND_174[0:0];
  _RAND_175 = {1{`RANDOM}};
  _T_1493 = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  _T_1508 = _RAND_176[0:0];
  _RAND_177 = {1{`RANDOM}};
  _T_1523 = _RAND_177[0:0];
  _RAND_178 = {1{`RANDOM}};
  _T_1538 = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  _T_1553 = _RAND_179[0:0];
  _RAND_180 = {1{`RANDOM}};
  _T_1568 = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  _T_1583 = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  _T_1598 = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  _T_1613 = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  _T_1628 = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  _T_1643 = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  _T_1658 = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  _T_1673 = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  _T_1688 = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  _T_1703 = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  _T_1718 = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  _T_1733 = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  config_reg = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  _T_2042 = _RAND_193[7:0];
  _RAND_194 = {1{`RANDOM}};
  _T_2043 = _RAND_194[3:0];
  _RAND_195 = {1{`RANDOM}};
  _T_2050 = _RAND_195[0:0];
  _RAND_196 = {1{`RANDOM}};
  _T_2052 = _RAND_196[0:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    picm_raddr_ff = 32'h0;
  end
  if (reset) begin
    picm_waddr_ff = 32'h0;
  end
  if (reset) begin
    picm_wren_ff = 1'h0;
  end
  if (reset) begin
    picm_rden_ff = 1'h0;
  end
  if (reset) begin
    picm_mken_ff = 1'h0;
  end
  if (reset) begin
    picm_wr_data_ff = 32'h0;
  end
  if (reset) begin
    gw_config_reg_31 = 2'h0;
  end
  if (reset) begin
    intenable_reg_31 = 1'h0;
  end
  if (reset) begin
    gw_config_reg_30 = 2'h0;
  end
  if (reset) begin
    intenable_reg_30 = 1'h0;
  end
  if (reset) begin
    gw_config_reg_29 = 2'h0;
  end
  if (reset) begin
    intenable_reg_29 = 1'h0;
  end
  if (reset) begin
    gw_config_reg_28 = 2'h0;
  end
  if (reset) begin
    intenable_reg_28 = 1'h0;
  end
  if (reset) begin
    gw_config_reg_27 = 2'h0;
  end
  if (reset) begin
    intenable_reg_27 = 1'h0;
  end
  if (reset) begin
    gw_config_reg_26 = 2'h0;
  end
  if (reset) begin
    intenable_reg_26 = 1'h0;
  end
  if (reset) begin
    gw_config_reg_25 = 2'h0;
  end
  if (reset) begin
    intenable_reg_25 = 1'h0;
  end
  if (reset) begin
    gw_config_reg_24 = 2'h0;
  end
  if (reset) begin
    intenable_reg_24 = 1'h0;
  end
  if (reset) begin
    gw_config_reg_23 = 2'h0;
  end
  if (reset) begin
    intenable_reg_23 = 1'h0;
  end
  if (reset) begin
    gw_config_reg_22 = 2'h0;
  end
  if (reset) begin
    intenable_reg_22 = 1'h0;
  end
  if (reset) begin
    gw_config_reg_21 = 2'h0;
  end
  if (reset) begin
    intenable_reg_21 = 1'h0;
  end
  if (reset) begin
    gw_config_reg_20 = 2'h0;
  end
  if (reset) begin
    intenable_reg_20 = 1'h0;
  end
  if (reset) begin
    gw_config_reg_19 = 2'h0;
  end
  if (reset) begin
    intenable_reg_19 = 1'h0;
  end
  if (reset) begin
    gw_config_reg_18 = 2'h0;
  end
  if (reset) begin
    intenable_reg_18 = 1'h0;
  end
  if (reset) begin
    gw_config_reg_17 = 2'h0;
  end
  if (reset) begin
    intenable_reg_17 = 1'h0;
  end
  if (reset) begin
    gw_config_reg_16 = 2'h0;
  end
  if (reset) begin
    intenable_reg_16 = 1'h0;
  end
  if (reset) begin
    gw_config_reg_15 = 2'h0;
  end
  if (reset) begin
    intenable_reg_15 = 1'h0;
  end
  if (reset) begin
    gw_config_reg_14 = 2'h0;
  end
  if (reset) begin
    intenable_reg_14 = 1'h0;
  end
  if (reset) begin
    gw_config_reg_13 = 2'h0;
  end
  if (reset) begin
    intenable_reg_13 = 1'h0;
  end
  if (reset) begin
    gw_config_reg_12 = 2'h0;
  end
  if (reset) begin
    intenable_reg_12 = 1'h0;
  end
  if (reset) begin
    gw_config_reg_11 = 2'h0;
  end
  if (reset) begin
    intenable_reg_11 = 1'h0;
  end
  if (reset) begin
    gw_config_reg_10 = 2'h0;
  end
  if (reset) begin
    intenable_reg_10 = 1'h0;
  end
  if (reset) begin
    gw_config_reg_9 = 2'h0;
  end
  if (reset) begin
    intenable_reg_9 = 1'h0;
  end
  if (reset) begin
    gw_config_reg_8 = 2'h0;
  end
  if (reset) begin
    intenable_reg_8 = 1'h0;
  end
  if (reset) begin
    gw_config_reg_7 = 2'h0;
  end
  if (reset) begin
    intenable_reg_7 = 1'h0;
  end
  if (reset) begin
    gw_config_reg_6 = 2'h0;
  end
  if (reset) begin
    intenable_reg_6 = 1'h0;
  end
  if (reset) begin
    gw_config_reg_5 = 2'h0;
  end
  if (reset) begin
    intenable_reg_5 = 1'h0;
  end
  if (reset) begin
    gw_config_reg_4 = 2'h0;
  end
  if (reset) begin
    intenable_reg_4 = 1'h0;
  end
  if (reset) begin
    gw_config_reg_3 = 2'h0;
  end
  if (reset) begin
    intenable_reg_3 = 1'h0;
  end
  if (reset) begin
    gw_config_reg_2 = 2'h0;
  end
  if (reset) begin
    intenable_reg_2 = 1'h0;
  end
  if (reset) begin
    gw_config_reg_1 = 2'h0;
  end
  if (reset) begin
    intenable_reg_1 = 1'h0;
  end
  if (reset) begin
    _T_66 = 1'h0;
  end
  if (reset) begin
    extintsrc_req_sync_1 = 1'h0;
  end
  if (reset) begin
    _T_70 = 1'h0;
  end
  if (reset) begin
    extintsrc_req_sync_2 = 1'h0;
  end
  if (reset) begin
    _T_74 = 1'h0;
  end
  if (reset) begin
    extintsrc_req_sync_3 = 1'h0;
  end
  if (reset) begin
    _T_78 = 1'h0;
  end
  if (reset) begin
    extintsrc_req_sync_4 = 1'h0;
  end
  if (reset) begin
    _T_82 = 1'h0;
  end
  if (reset) begin
    extintsrc_req_sync_5 = 1'h0;
  end
  if (reset) begin
    _T_86 = 1'h0;
  end
  if (reset) begin
    extintsrc_req_sync_6 = 1'h0;
  end
  if (reset) begin
    _T_90 = 1'h0;
  end
  if (reset) begin
    extintsrc_req_sync_7 = 1'h0;
  end
  if (reset) begin
    _T_94 = 1'h0;
  end
  if (reset) begin
    extintsrc_req_sync_8 = 1'h0;
  end
  if (reset) begin
    _T_98 = 1'h0;
  end
  if (reset) begin
    extintsrc_req_sync_9 = 1'h0;
  end
  if (reset) begin
    _T_102 = 1'h0;
  end
  if (reset) begin
    extintsrc_req_sync_10 = 1'h0;
  end
  if (reset) begin
    _T_106 = 1'h0;
  end
  if (reset) begin
    extintsrc_req_sync_11 = 1'h0;
  end
  if (reset) begin
    _T_110 = 1'h0;
  end
  if (reset) begin
    extintsrc_req_sync_12 = 1'h0;
  end
  if (reset) begin
    _T_114 = 1'h0;
  end
  if (reset) begin
    extintsrc_req_sync_13 = 1'h0;
  end
  if (reset) begin
    _T_118 = 1'h0;
  end
  if (reset) begin
    extintsrc_req_sync_14 = 1'h0;
  end
  if (reset) begin
    _T_122 = 1'h0;
  end
  if (reset) begin
    extintsrc_req_sync_15 = 1'h0;
  end
  if (reset) begin
    _T_126 = 1'h0;
  end
  if (reset) begin
    extintsrc_req_sync_16 = 1'h0;
  end
  if (reset) begin
    _T_130 = 1'h0;
  end
  if (reset) begin
    extintsrc_req_sync_17 = 1'h0;
  end
  if (reset) begin
    _T_134 = 1'h0;
  end
  if (reset) begin
    extintsrc_req_sync_18 = 1'h0;
  end
  if (reset) begin
    _T_138 = 1'h0;
  end
  if (reset) begin
    extintsrc_req_sync_19 = 1'h0;
  end
  if (reset) begin
    _T_142 = 1'h0;
  end
  if (reset) begin
    extintsrc_req_sync_20 = 1'h0;
  end
  if (reset) begin
    _T_146 = 1'h0;
  end
  if (reset) begin
    extintsrc_req_sync_21 = 1'h0;
  end
  if (reset) begin
    _T_150 = 1'h0;
  end
  if (reset) begin
    extintsrc_req_sync_22 = 1'h0;
  end
  if (reset) begin
    _T_154 = 1'h0;
  end
  if (reset) begin
    extintsrc_req_sync_23 = 1'h0;
  end
  if (reset) begin
    _T_158 = 1'h0;
  end
  if (reset) begin
    extintsrc_req_sync_24 = 1'h0;
  end
  if (reset) begin
    _T_162 = 1'h0;
  end
  if (reset) begin
    extintsrc_req_sync_25 = 1'h0;
  end
  if (reset) begin
    _T_166 = 1'h0;
  end
  if (reset) begin
    extintsrc_req_sync_26 = 1'h0;
  end
  if (reset) begin
    _T_170 = 1'h0;
  end
  if (reset) begin
    extintsrc_req_sync_27 = 1'h0;
  end
  if (reset) begin
    _T_174 = 1'h0;
  end
  if (reset) begin
    extintsrc_req_sync_28 = 1'h0;
  end
  if (reset) begin
    _T_178 = 1'h0;
  end
  if (reset) begin
    extintsrc_req_sync_29 = 1'h0;
  end
  if (reset) begin
    _T_182 = 1'h0;
  end
  if (reset) begin
    extintsrc_req_sync_30 = 1'h0;
  end
  if (reset) begin
    _T_186 = 1'h0;
  end
  if (reset) begin
    extintsrc_req_sync_31 = 1'h0;
  end
  if (reset) begin
    intpriority_reg_1 = 4'h0;
  end
  if (reset) begin
    intpriority_reg_2 = 4'h0;
  end
  if (reset) begin
    intpriority_reg_3 = 4'h0;
  end
  if (reset) begin
    intpriority_reg_4 = 4'h0;
  end
  if (reset) begin
    intpriority_reg_5 = 4'h0;
  end
  if (reset) begin
    intpriority_reg_6 = 4'h0;
  end
  if (reset) begin
    intpriority_reg_7 = 4'h0;
  end
  if (reset) begin
    intpriority_reg_8 = 4'h0;
  end
  if (reset) begin
    intpriority_reg_9 = 4'h0;
  end
  if (reset) begin
    intpriority_reg_10 = 4'h0;
  end
  if (reset) begin
    intpriority_reg_11 = 4'h0;
  end
  if (reset) begin
    intpriority_reg_12 = 4'h0;
  end
  if (reset) begin
    intpriority_reg_13 = 4'h0;
  end
  if (reset) begin
    intpriority_reg_14 = 4'h0;
  end
  if (reset) begin
    intpriority_reg_15 = 4'h0;
  end
  if (reset) begin
    intpriority_reg_16 = 4'h0;
  end
  if (reset) begin
    intpriority_reg_17 = 4'h0;
  end
  if (reset) begin
    intpriority_reg_18 = 4'h0;
  end
  if (reset) begin
    intpriority_reg_19 = 4'h0;
  end
  if (reset) begin
    intpriority_reg_20 = 4'h0;
  end
  if (reset) begin
    intpriority_reg_21 = 4'h0;
  end
  if (reset) begin
    intpriority_reg_22 = 4'h0;
  end
  if (reset) begin
    intpriority_reg_23 = 4'h0;
  end
  if (reset) begin
    intpriority_reg_24 = 4'h0;
  end
  if (reset) begin
    intpriority_reg_25 = 4'h0;
  end
  if (reset) begin
    intpriority_reg_26 = 4'h0;
  end
  if (reset) begin
    intpriority_reg_27 = 4'h0;
  end
  if (reset) begin
    intpriority_reg_28 = 4'h0;
  end
  if (reset) begin
    intpriority_reg_29 = 4'h0;
  end
  if (reset) begin
    intpriority_reg_30 = 4'h0;
  end
  if (reset) begin
    intpriority_reg_31 = 4'h0;
  end
  if (reset) begin
    _T_1283 = 1'h0;
  end
  if (reset) begin
    _T_1298 = 1'h0;
  end
  if (reset) begin
    _T_1313 = 1'h0;
  end
  if (reset) begin
    _T_1328 = 1'h0;
  end
  if (reset) begin
    _T_1343 = 1'h0;
  end
  if (reset) begin
    _T_1358 = 1'h0;
  end
  if (reset) begin
    _T_1373 = 1'h0;
  end
  if (reset) begin
    _T_1388 = 1'h0;
  end
  if (reset) begin
    _T_1403 = 1'h0;
  end
  if (reset) begin
    _T_1418 = 1'h0;
  end
  if (reset) begin
    _T_1433 = 1'h0;
  end
  if (reset) begin
    _T_1448 = 1'h0;
  end
  if (reset) begin
    _T_1463 = 1'h0;
  end
  if (reset) begin
    _T_1478 = 1'h0;
  end
  if (reset) begin
    _T_1493 = 1'h0;
  end
  if (reset) begin
    _T_1508 = 1'h0;
  end
  if (reset) begin
    _T_1523 = 1'h0;
  end
  if (reset) begin
    _T_1538 = 1'h0;
  end
  if (reset) begin
    _T_1553 = 1'h0;
  end
  if (reset) begin
    _T_1568 = 1'h0;
  end
  if (reset) begin
    _T_1583 = 1'h0;
  end
  if (reset) begin
    _T_1598 = 1'h0;
  end
  if (reset) begin
    _T_1613 = 1'h0;
  end
  if (reset) begin
    _T_1628 = 1'h0;
  end
  if (reset) begin
    _T_1643 = 1'h0;
  end
  if (reset) begin
    _T_1658 = 1'h0;
  end
  if (reset) begin
    _T_1673 = 1'h0;
  end
  if (reset) begin
    _T_1688 = 1'h0;
  end
  if (reset) begin
    _T_1703 = 1'h0;
  end
  if (reset) begin
    _T_1718 = 1'h0;
  end
  if (reset) begin
    _T_1733 = 1'h0;
  end
  if (reset) begin
    config_reg = 1'h0;
  end
  if (reset) begin
    _T_2042 = 8'h0;
  end
  if (reset) begin
    _T_2043 = 4'h0;
  end
  if (reset) begin
    _T_2050 = 1'h0;
  end
  if (reset) begin
    _T_2052 = 1'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      picm_raddr_ff <= 32'h0;
    end else begin
      picm_raddr_ff <= io_lsu_pic_picm_rdaddr;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      picm_waddr_ff <= 32'h0;
    end else begin
      picm_waddr_ff <= io_lsu_pic_picm_wraddr;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      picm_wren_ff <= 1'h0;
    end else begin
      picm_wren_ff <= io_lsu_pic_picm_wren;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      picm_rden_ff <= 1'h0;
    end else begin
      picm_rden_ff <= io_lsu_pic_picm_rden;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      picm_mken_ff <= 1'h0;
    end else begin
      picm_mken_ff <= io_lsu_pic_picm_mken;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      picm_wr_data_ff <= 32'h0;
    end else begin
      picm_wr_data_ff <= io_lsu_pic_picm_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      gw_config_reg_31 <= 2'h0;
    end else if (gw_config_reg_we_31) begin
      gw_config_reg_31 <= picm_wr_data_ff[1:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      intenable_reg_31 <= 1'h0;
    end else if (intenable_reg_we_31) begin
      intenable_reg_31 <= picm_wr_data_ff[0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      gw_config_reg_30 <= 2'h0;
    end else if (gw_config_reg_we_30) begin
      gw_config_reg_30 <= picm_wr_data_ff[1:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      intenable_reg_30 <= 1'h0;
    end else if (intenable_reg_we_30) begin
      intenable_reg_30 <= picm_wr_data_ff[0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      gw_config_reg_29 <= 2'h0;
    end else if (gw_config_reg_we_29) begin
      gw_config_reg_29 <= picm_wr_data_ff[1:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      intenable_reg_29 <= 1'h0;
    end else if (intenable_reg_we_29) begin
      intenable_reg_29 <= picm_wr_data_ff[0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      gw_config_reg_28 <= 2'h0;
    end else if (gw_config_reg_we_28) begin
      gw_config_reg_28 <= picm_wr_data_ff[1:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      intenable_reg_28 <= 1'h0;
    end else if (intenable_reg_we_28) begin
      intenable_reg_28 <= picm_wr_data_ff[0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      gw_config_reg_27 <= 2'h0;
    end else if (gw_config_reg_we_27) begin
      gw_config_reg_27 <= picm_wr_data_ff[1:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      intenable_reg_27 <= 1'h0;
    end else if (intenable_reg_we_27) begin
      intenable_reg_27 <= picm_wr_data_ff[0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      gw_config_reg_26 <= 2'h0;
    end else if (gw_config_reg_we_26) begin
      gw_config_reg_26 <= picm_wr_data_ff[1:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      intenable_reg_26 <= 1'h0;
    end else if (intenable_reg_we_26) begin
      intenable_reg_26 <= picm_wr_data_ff[0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      gw_config_reg_25 <= 2'h0;
    end else if (gw_config_reg_we_25) begin
      gw_config_reg_25 <= picm_wr_data_ff[1:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      intenable_reg_25 <= 1'h0;
    end else if (intenable_reg_we_25) begin
      intenable_reg_25 <= picm_wr_data_ff[0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      gw_config_reg_24 <= 2'h0;
    end else if (gw_config_reg_we_24) begin
      gw_config_reg_24 <= picm_wr_data_ff[1:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      intenable_reg_24 <= 1'h0;
    end else if (intenable_reg_we_24) begin
      intenable_reg_24 <= picm_wr_data_ff[0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      gw_config_reg_23 <= 2'h0;
    end else if (gw_config_reg_we_23) begin
      gw_config_reg_23 <= picm_wr_data_ff[1:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      intenable_reg_23 <= 1'h0;
    end else if (intenable_reg_we_23) begin
      intenable_reg_23 <= picm_wr_data_ff[0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      gw_config_reg_22 <= 2'h0;
    end else if (gw_config_reg_we_22) begin
      gw_config_reg_22 <= picm_wr_data_ff[1:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      intenable_reg_22 <= 1'h0;
    end else if (intenable_reg_we_22) begin
      intenable_reg_22 <= picm_wr_data_ff[0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      gw_config_reg_21 <= 2'h0;
    end else if (gw_config_reg_we_21) begin
      gw_config_reg_21 <= picm_wr_data_ff[1:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      intenable_reg_21 <= 1'h0;
    end else if (intenable_reg_we_21) begin
      intenable_reg_21 <= picm_wr_data_ff[0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      gw_config_reg_20 <= 2'h0;
    end else if (gw_config_reg_we_20) begin
      gw_config_reg_20 <= picm_wr_data_ff[1:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      intenable_reg_20 <= 1'h0;
    end else if (intenable_reg_we_20) begin
      intenable_reg_20 <= picm_wr_data_ff[0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      gw_config_reg_19 <= 2'h0;
    end else if (gw_config_reg_we_19) begin
      gw_config_reg_19 <= picm_wr_data_ff[1:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      intenable_reg_19 <= 1'h0;
    end else if (intenable_reg_we_19) begin
      intenable_reg_19 <= picm_wr_data_ff[0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      gw_config_reg_18 <= 2'h0;
    end else if (gw_config_reg_we_18) begin
      gw_config_reg_18 <= picm_wr_data_ff[1:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      intenable_reg_18 <= 1'h0;
    end else if (intenable_reg_we_18) begin
      intenable_reg_18 <= picm_wr_data_ff[0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      gw_config_reg_17 <= 2'h0;
    end else if (gw_config_reg_we_17) begin
      gw_config_reg_17 <= picm_wr_data_ff[1:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      intenable_reg_17 <= 1'h0;
    end else if (intenable_reg_we_17) begin
      intenable_reg_17 <= picm_wr_data_ff[0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      gw_config_reg_16 <= 2'h0;
    end else if (gw_config_reg_we_16) begin
      gw_config_reg_16 <= picm_wr_data_ff[1:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      intenable_reg_16 <= 1'h0;
    end else if (intenable_reg_we_16) begin
      intenable_reg_16 <= picm_wr_data_ff[0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      gw_config_reg_15 <= 2'h0;
    end else if (gw_config_reg_we_15) begin
      gw_config_reg_15 <= picm_wr_data_ff[1:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      intenable_reg_15 <= 1'h0;
    end else if (intenable_reg_we_15) begin
      intenable_reg_15 <= picm_wr_data_ff[0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      gw_config_reg_14 <= 2'h0;
    end else if (gw_config_reg_we_14) begin
      gw_config_reg_14 <= picm_wr_data_ff[1:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      intenable_reg_14 <= 1'h0;
    end else if (intenable_reg_we_14) begin
      intenable_reg_14 <= picm_wr_data_ff[0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      gw_config_reg_13 <= 2'h0;
    end else if (gw_config_reg_we_13) begin
      gw_config_reg_13 <= picm_wr_data_ff[1:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      intenable_reg_13 <= 1'h0;
    end else if (intenable_reg_we_13) begin
      intenable_reg_13 <= picm_wr_data_ff[0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      gw_config_reg_12 <= 2'h0;
    end else if (gw_config_reg_we_12) begin
      gw_config_reg_12 <= picm_wr_data_ff[1:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      intenable_reg_12 <= 1'h0;
    end else if (intenable_reg_we_12) begin
      intenable_reg_12 <= picm_wr_data_ff[0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      gw_config_reg_11 <= 2'h0;
    end else if (gw_config_reg_we_11) begin
      gw_config_reg_11 <= picm_wr_data_ff[1:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      intenable_reg_11 <= 1'h0;
    end else if (intenable_reg_we_11) begin
      intenable_reg_11 <= picm_wr_data_ff[0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      gw_config_reg_10 <= 2'h0;
    end else if (gw_config_reg_we_10) begin
      gw_config_reg_10 <= picm_wr_data_ff[1:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      intenable_reg_10 <= 1'h0;
    end else if (intenable_reg_we_10) begin
      intenable_reg_10 <= picm_wr_data_ff[0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      gw_config_reg_9 <= 2'h0;
    end else if (gw_config_reg_we_9) begin
      gw_config_reg_9 <= picm_wr_data_ff[1:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      intenable_reg_9 <= 1'h0;
    end else if (intenable_reg_we_9) begin
      intenable_reg_9 <= picm_wr_data_ff[0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      gw_config_reg_8 <= 2'h0;
    end else if (gw_config_reg_we_8) begin
      gw_config_reg_8 <= picm_wr_data_ff[1:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      intenable_reg_8 <= 1'h0;
    end else if (intenable_reg_we_8) begin
      intenable_reg_8 <= picm_wr_data_ff[0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      gw_config_reg_7 <= 2'h0;
    end else if (gw_config_reg_we_7) begin
      gw_config_reg_7 <= picm_wr_data_ff[1:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      intenable_reg_7 <= 1'h0;
    end else if (intenable_reg_we_7) begin
      intenable_reg_7 <= picm_wr_data_ff[0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      gw_config_reg_6 <= 2'h0;
    end else if (gw_config_reg_we_6) begin
      gw_config_reg_6 <= picm_wr_data_ff[1:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      intenable_reg_6 <= 1'h0;
    end else if (intenable_reg_we_6) begin
      intenable_reg_6 <= picm_wr_data_ff[0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      gw_config_reg_5 <= 2'h0;
    end else if (gw_config_reg_we_5) begin
      gw_config_reg_5 <= picm_wr_data_ff[1:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      intenable_reg_5 <= 1'h0;
    end else if (intenable_reg_we_5) begin
      intenable_reg_5 <= picm_wr_data_ff[0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      gw_config_reg_4 <= 2'h0;
    end else if (gw_config_reg_we_4) begin
      gw_config_reg_4 <= picm_wr_data_ff[1:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      intenable_reg_4 <= 1'h0;
    end else if (intenable_reg_we_4) begin
      intenable_reg_4 <= picm_wr_data_ff[0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      gw_config_reg_3 <= 2'h0;
    end else if (gw_config_reg_we_3) begin
      gw_config_reg_3 <= picm_wr_data_ff[1:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      intenable_reg_3 <= 1'h0;
    end else if (intenable_reg_we_3) begin
      intenable_reg_3 <= picm_wr_data_ff[0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      gw_config_reg_2 <= 2'h0;
    end else if (gw_config_reg_we_2) begin
      gw_config_reg_2 <= picm_wr_data_ff[1:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      intenable_reg_2 <= 1'h0;
    end else if (intenable_reg_we_2) begin
      intenable_reg_2 <= picm_wr_data_ff[0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      gw_config_reg_1 <= 2'h0;
    end else if (gw_config_reg_we_1) begin
      gw_config_reg_1 <= picm_wr_data_ff[1:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      intenable_reg_1 <= 1'h0;
    end else if (intenable_reg_we_1) begin
      intenable_reg_1 <= picm_wr_data_ff[0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_66 <= 1'h0;
    end else if (intenable_clk_enable_grp_0) begin
      _T_66 <= io_extintsrc_req[1];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      extintsrc_req_sync_1 <= 1'h0;
    end else if (intenable_clk_enable_grp_0) begin
      extintsrc_req_sync_1 <= _T_66;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_70 <= 1'h0;
    end else if (intenable_clk_enable_grp_0) begin
      _T_70 <= io_extintsrc_req[2];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      extintsrc_req_sync_2 <= 1'h0;
    end else if (intenable_clk_enable_grp_0) begin
      extintsrc_req_sync_2 <= _T_70;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_74 <= 1'h0;
    end else if (intenable_clk_enable_grp_0) begin
      _T_74 <= io_extintsrc_req[3];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      extintsrc_req_sync_3 <= 1'h0;
    end else if (intenable_clk_enable_grp_0) begin
      extintsrc_req_sync_3 <= _T_74;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_78 <= 1'h0;
    end else if (intenable_clk_enable_grp_1) begin
      _T_78 <= io_extintsrc_req[4];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      extintsrc_req_sync_4 <= 1'h0;
    end else if (intenable_clk_enable_grp_1) begin
      extintsrc_req_sync_4 <= _T_78;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_82 <= 1'h0;
    end else if (intenable_clk_enable_grp_1) begin
      _T_82 <= io_extintsrc_req[5];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      extintsrc_req_sync_5 <= 1'h0;
    end else if (intenable_clk_enable_grp_1) begin
      extintsrc_req_sync_5 <= _T_82;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_86 <= 1'h0;
    end else if (intenable_clk_enable_grp_1) begin
      _T_86 <= io_extintsrc_req[6];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      extintsrc_req_sync_6 <= 1'h0;
    end else if (intenable_clk_enable_grp_1) begin
      extintsrc_req_sync_6 <= _T_86;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_90 <= 1'h0;
    end else if (intenable_clk_enable_grp_1) begin
      _T_90 <= io_extintsrc_req[7];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      extintsrc_req_sync_7 <= 1'h0;
    end else if (intenable_clk_enable_grp_1) begin
      extintsrc_req_sync_7 <= _T_90;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_94 <= 1'h0;
    end else if (intenable_clk_enable_grp_2) begin
      _T_94 <= io_extintsrc_req[8];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      extintsrc_req_sync_8 <= 1'h0;
    end else if (intenable_clk_enable_grp_2) begin
      extintsrc_req_sync_8 <= _T_94;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_98 <= 1'h0;
    end else if (intenable_clk_enable_grp_2) begin
      _T_98 <= io_extintsrc_req[9];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      extintsrc_req_sync_9 <= 1'h0;
    end else if (intenable_clk_enable_grp_2) begin
      extintsrc_req_sync_9 <= _T_98;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_102 <= 1'h0;
    end else if (intenable_clk_enable_grp_2) begin
      _T_102 <= io_extintsrc_req[10];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      extintsrc_req_sync_10 <= 1'h0;
    end else if (intenable_clk_enable_grp_2) begin
      extintsrc_req_sync_10 <= _T_102;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_106 <= 1'h0;
    end else if (intenable_clk_enable_grp_2) begin
      _T_106 <= io_extintsrc_req[11];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      extintsrc_req_sync_11 <= 1'h0;
    end else if (intenable_clk_enable_grp_2) begin
      extintsrc_req_sync_11 <= _T_106;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_110 <= 1'h0;
    end else if (intenable_clk_enable_grp_3) begin
      _T_110 <= io_extintsrc_req[12];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      extintsrc_req_sync_12 <= 1'h0;
    end else if (intenable_clk_enable_grp_3) begin
      extintsrc_req_sync_12 <= _T_110;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_114 <= 1'h0;
    end else if (intenable_clk_enable_grp_3) begin
      _T_114 <= io_extintsrc_req[13];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      extintsrc_req_sync_13 <= 1'h0;
    end else if (intenable_clk_enable_grp_3) begin
      extintsrc_req_sync_13 <= _T_114;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_118 <= 1'h0;
    end else if (intenable_clk_enable_grp_3) begin
      _T_118 <= io_extintsrc_req[14];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      extintsrc_req_sync_14 <= 1'h0;
    end else if (intenable_clk_enable_grp_3) begin
      extintsrc_req_sync_14 <= _T_118;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_122 <= 1'h0;
    end else if (intenable_clk_enable_grp_3) begin
      _T_122 <= io_extintsrc_req[15];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      extintsrc_req_sync_15 <= 1'h0;
    end else if (intenable_clk_enable_grp_3) begin
      extintsrc_req_sync_15 <= _T_122;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_126 <= 1'h0;
    end else if (intenable_clk_enable_grp_4) begin
      _T_126 <= io_extintsrc_req[16];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      extintsrc_req_sync_16 <= 1'h0;
    end else if (intenable_clk_enable_grp_4) begin
      extintsrc_req_sync_16 <= _T_126;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_130 <= 1'h0;
    end else if (intenable_clk_enable_grp_4) begin
      _T_130 <= io_extintsrc_req[17];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      extintsrc_req_sync_17 <= 1'h0;
    end else if (intenable_clk_enable_grp_4) begin
      extintsrc_req_sync_17 <= _T_130;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_134 <= 1'h0;
    end else if (intenable_clk_enable_grp_4) begin
      _T_134 <= io_extintsrc_req[18];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      extintsrc_req_sync_18 <= 1'h0;
    end else if (intenable_clk_enable_grp_4) begin
      extintsrc_req_sync_18 <= _T_134;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_138 <= 1'h0;
    end else if (intenable_clk_enable_grp_4) begin
      _T_138 <= io_extintsrc_req[19];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      extintsrc_req_sync_19 <= 1'h0;
    end else if (intenable_clk_enable_grp_4) begin
      extintsrc_req_sync_19 <= _T_138;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_142 <= 1'h0;
    end else if (intenable_clk_enable_grp_5) begin
      _T_142 <= io_extintsrc_req[20];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      extintsrc_req_sync_20 <= 1'h0;
    end else if (intenable_clk_enable_grp_5) begin
      extintsrc_req_sync_20 <= _T_142;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_146 <= 1'h0;
    end else if (intenable_clk_enable_grp_5) begin
      _T_146 <= io_extintsrc_req[21];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      extintsrc_req_sync_21 <= 1'h0;
    end else if (intenable_clk_enable_grp_5) begin
      extintsrc_req_sync_21 <= _T_146;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_150 <= 1'h0;
    end else if (intenable_clk_enable_grp_5) begin
      _T_150 <= io_extintsrc_req[22];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      extintsrc_req_sync_22 <= 1'h0;
    end else if (intenable_clk_enable_grp_5) begin
      extintsrc_req_sync_22 <= _T_150;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_154 <= 1'h0;
    end else if (intenable_clk_enable_grp_5) begin
      _T_154 <= io_extintsrc_req[23];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      extintsrc_req_sync_23 <= 1'h0;
    end else if (intenable_clk_enable_grp_5) begin
      extintsrc_req_sync_23 <= _T_154;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_158 <= 1'h0;
    end else if (intenable_clk_enable_grp_6) begin
      _T_158 <= io_extintsrc_req[24];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      extintsrc_req_sync_24 <= 1'h0;
    end else if (intenable_clk_enable_grp_6) begin
      extintsrc_req_sync_24 <= _T_158;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_162 <= 1'h0;
    end else if (intenable_clk_enable_grp_6) begin
      _T_162 <= io_extintsrc_req[25];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      extintsrc_req_sync_25 <= 1'h0;
    end else if (intenable_clk_enable_grp_6) begin
      extintsrc_req_sync_25 <= _T_162;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_166 <= 1'h0;
    end else if (intenable_clk_enable_grp_6) begin
      _T_166 <= io_extintsrc_req[26];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      extintsrc_req_sync_26 <= 1'h0;
    end else if (intenable_clk_enable_grp_6) begin
      extintsrc_req_sync_26 <= _T_166;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_170 <= 1'h0;
    end else if (intenable_clk_enable_grp_6) begin
      _T_170 <= io_extintsrc_req[27];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      extintsrc_req_sync_27 <= 1'h0;
    end else if (intenable_clk_enable_grp_6) begin
      extintsrc_req_sync_27 <= _T_170;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_174 <= 1'h0;
    end else if (intenable_clk_enable_grp_7) begin
      _T_174 <= io_extintsrc_req[28];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      extintsrc_req_sync_28 <= 1'h0;
    end else if (intenable_clk_enable_grp_7) begin
      extintsrc_req_sync_28 <= _T_174;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_178 <= 1'h0;
    end else if (intenable_clk_enable_grp_7) begin
      _T_178 <= io_extintsrc_req[29];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      extintsrc_req_sync_29 <= 1'h0;
    end else if (intenable_clk_enable_grp_7) begin
      extintsrc_req_sync_29 <= _T_178;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_182 <= 1'h0;
    end else if (intenable_clk_enable_grp_7) begin
      _T_182 <= io_extintsrc_req[30];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      extintsrc_req_sync_30 <= 1'h0;
    end else if (intenable_clk_enable_grp_7) begin
      extintsrc_req_sync_30 <= _T_182;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_186 <= 1'h0;
    end else if (intenable_clk_enable_grp_7) begin
      _T_186 <= io_extintsrc_req[31];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      extintsrc_req_sync_31 <= 1'h0;
    end else if (intenable_clk_enable_grp_7) begin
      extintsrc_req_sync_31 <= _T_186;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      intpriority_reg_1 <= 4'h0;
    end else if (intpriority_reg_we_1) begin
      intpriority_reg_1 <= picm_wr_data_ff[3:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      intpriority_reg_2 <= 4'h0;
    end else if (intpriority_reg_we_2) begin
      intpriority_reg_2 <= picm_wr_data_ff[3:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      intpriority_reg_3 <= 4'h0;
    end else if (intpriority_reg_we_3) begin
      intpriority_reg_3 <= picm_wr_data_ff[3:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      intpriority_reg_4 <= 4'h0;
    end else if (intpriority_reg_we_4) begin
      intpriority_reg_4 <= picm_wr_data_ff[3:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      intpriority_reg_5 <= 4'h0;
    end else if (intpriority_reg_we_5) begin
      intpriority_reg_5 <= picm_wr_data_ff[3:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      intpriority_reg_6 <= 4'h0;
    end else if (intpriority_reg_we_6) begin
      intpriority_reg_6 <= picm_wr_data_ff[3:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      intpriority_reg_7 <= 4'h0;
    end else if (intpriority_reg_we_7) begin
      intpriority_reg_7 <= picm_wr_data_ff[3:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      intpriority_reg_8 <= 4'h0;
    end else if (intpriority_reg_we_8) begin
      intpriority_reg_8 <= picm_wr_data_ff[3:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      intpriority_reg_9 <= 4'h0;
    end else if (intpriority_reg_we_9) begin
      intpriority_reg_9 <= picm_wr_data_ff[3:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      intpriority_reg_10 <= 4'h0;
    end else if (intpriority_reg_we_10) begin
      intpriority_reg_10 <= picm_wr_data_ff[3:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      intpriority_reg_11 <= 4'h0;
    end else if (intpriority_reg_we_11) begin
      intpriority_reg_11 <= picm_wr_data_ff[3:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      intpriority_reg_12 <= 4'h0;
    end else if (intpriority_reg_we_12) begin
      intpriority_reg_12 <= picm_wr_data_ff[3:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      intpriority_reg_13 <= 4'h0;
    end else if (intpriority_reg_we_13) begin
      intpriority_reg_13 <= picm_wr_data_ff[3:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      intpriority_reg_14 <= 4'h0;
    end else if (intpriority_reg_we_14) begin
      intpriority_reg_14 <= picm_wr_data_ff[3:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      intpriority_reg_15 <= 4'h0;
    end else if (intpriority_reg_we_15) begin
      intpriority_reg_15 <= picm_wr_data_ff[3:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      intpriority_reg_16 <= 4'h0;
    end else if (intpriority_reg_we_16) begin
      intpriority_reg_16 <= picm_wr_data_ff[3:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      intpriority_reg_17 <= 4'h0;
    end else if (intpriority_reg_we_17) begin
      intpriority_reg_17 <= picm_wr_data_ff[3:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      intpriority_reg_18 <= 4'h0;
    end else if (intpriority_reg_we_18) begin
      intpriority_reg_18 <= picm_wr_data_ff[3:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      intpriority_reg_19 <= 4'h0;
    end else if (intpriority_reg_we_19) begin
      intpriority_reg_19 <= picm_wr_data_ff[3:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      intpriority_reg_20 <= 4'h0;
    end else if (intpriority_reg_we_20) begin
      intpriority_reg_20 <= picm_wr_data_ff[3:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      intpriority_reg_21 <= 4'h0;
    end else if (intpriority_reg_we_21) begin
      intpriority_reg_21 <= picm_wr_data_ff[3:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      intpriority_reg_22 <= 4'h0;
    end else if (intpriority_reg_we_22) begin
      intpriority_reg_22 <= picm_wr_data_ff[3:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      intpriority_reg_23 <= 4'h0;
    end else if (intpriority_reg_we_23) begin
      intpriority_reg_23 <= picm_wr_data_ff[3:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      intpriority_reg_24 <= 4'h0;
    end else if (intpriority_reg_we_24) begin
      intpriority_reg_24 <= picm_wr_data_ff[3:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      intpriority_reg_25 <= 4'h0;
    end else if (intpriority_reg_we_25) begin
      intpriority_reg_25 <= picm_wr_data_ff[3:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      intpriority_reg_26 <= 4'h0;
    end else if (intpriority_reg_we_26) begin
      intpriority_reg_26 <= picm_wr_data_ff[3:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      intpriority_reg_27 <= 4'h0;
    end else if (intpriority_reg_we_27) begin
      intpriority_reg_27 <= picm_wr_data_ff[3:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      intpriority_reg_28 <= 4'h0;
    end else if (intpriority_reg_we_28) begin
      intpriority_reg_28 <= picm_wr_data_ff[3:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      intpriority_reg_29 <= 4'h0;
    end else if (intpriority_reg_we_29) begin
      intpriority_reg_29 <= picm_wr_data_ff[3:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      intpriority_reg_30 <= 4'h0;
    end else if (intpriority_reg_we_30) begin
      intpriority_reg_30 <= picm_wr_data_ff[3:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      intpriority_reg_31 <= 4'h0;
    end else if (intpriority_reg_we_31) begin
      intpriority_reg_31 <= picm_wr_data_ff[3:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1283 <= 1'h0;
    end else if (intenable_clk_enable_grp_0) begin
      _T_1283 <= _T_1282;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1298 <= 1'h0;
    end else if (intenable_clk_enable_grp_0) begin
      _T_1298 <= _T_1297;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1313 <= 1'h0;
    end else if (intenable_clk_enable_grp_0) begin
      _T_1313 <= _T_1312;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1328 <= 1'h0;
    end else if (intenable_clk_enable_grp_1) begin
      _T_1328 <= _T_1327;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1343 <= 1'h0;
    end else if (intenable_clk_enable_grp_1) begin
      _T_1343 <= _T_1342;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1358 <= 1'h0;
    end else if (intenable_clk_enable_grp_1) begin
      _T_1358 <= _T_1357;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1373 <= 1'h0;
    end else if (intenable_clk_enable_grp_1) begin
      _T_1373 <= _T_1372;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1388 <= 1'h0;
    end else if (intenable_clk_enable_grp_2) begin
      _T_1388 <= _T_1387;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1403 <= 1'h0;
    end else if (intenable_clk_enable_grp_2) begin
      _T_1403 <= _T_1402;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1418 <= 1'h0;
    end else if (intenable_clk_enable_grp_2) begin
      _T_1418 <= _T_1417;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1433 <= 1'h0;
    end else if (intenable_clk_enable_grp_2) begin
      _T_1433 <= _T_1432;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1448 <= 1'h0;
    end else if (intenable_clk_enable_grp_3) begin
      _T_1448 <= _T_1447;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1463 <= 1'h0;
    end else if (intenable_clk_enable_grp_3) begin
      _T_1463 <= _T_1462;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1478 <= 1'h0;
    end else if (intenable_clk_enable_grp_3) begin
      _T_1478 <= _T_1477;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1493 <= 1'h0;
    end else if (intenable_clk_enable_grp_3) begin
      _T_1493 <= _T_1492;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1508 <= 1'h0;
    end else if (intenable_clk_enable_grp_4) begin
      _T_1508 <= _T_1507;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1523 <= 1'h0;
    end else if (intenable_clk_enable_grp_4) begin
      _T_1523 <= _T_1522;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1538 <= 1'h0;
    end else if (intenable_clk_enable_grp_4) begin
      _T_1538 <= _T_1537;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1553 <= 1'h0;
    end else if (intenable_clk_enable_grp_4) begin
      _T_1553 <= _T_1552;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1568 <= 1'h0;
    end else if (intenable_clk_enable_grp_5) begin
      _T_1568 <= _T_1567;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1583 <= 1'h0;
    end else if (intenable_clk_enable_grp_5) begin
      _T_1583 <= _T_1582;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1598 <= 1'h0;
    end else if (intenable_clk_enable_grp_5) begin
      _T_1598 <= _T_1597;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1613 <= 1'h0;
    end else if (intenable_clk_enable_grp_5) begin
      _T_1613 <= _T_1612;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1628 <= 1'h0;
    end else if (intenable_clk_enable_grp_6) begin
      _T_1628 <= _T_1627;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1643 <= 1'h0;
    end else if (intenable_clk_enable_grp_6) begin
      _T_1643 <= _T_1642;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1658 <= 1'h0;
    end else if (intenable_clk_enable_grp_6) begin
      _T_1658 <= _T_1657;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1673 <= 1'h0;
    end else if (intenable_clk_enable_grp_6) begin
      _T_1673 <= _T_1672;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1688 <= 1'h0;
    end else if (intenable_clk_enable_grp_7) begin
      _T_1688 <= _T_1687;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1703 <= 1'h0;
    end else if (intenable_clk_enable_grp_7) begin
      _T_1703 <= _T_1702;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1718 <= 1'h0;
    end else if (intenable_clk_enable_grp_7) begin
      _T_1718 <= _T_1717;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      _T_1733 <= 1'h0;
    end else if (intenable_clk_enable_grp_7) begin
      _T_1733 <= _T_1732;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      config_reg <= 1'h0;
    end else if (config_reg_we) begin
      config_reg <= picm_wr_data_ff[0];
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      _T_2042 <= 8'h0;
    end else begin
      _T_2042 <= level_intpend_id_5_0;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      _T_2043 <= 4'h0;
    end else if (config_reg) begin
      _T_2043 <= _T_2041;
    end else begin
      _T_2043 <= level_intpend_w_prior_en_5_0;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      _T_2050 <= 1'h0;
    end else begin
      _T_2050 <= _T_2048 & _T_2049;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      _T_2052 <= 1'h0;
    end else begin
      _T_2052 <= pl_in_q == maxint;
    end
  end
endmodule
