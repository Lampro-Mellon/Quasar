module el2_ifu_mem_ctl(
  input         clock,
  input         reset,
  input         io_free_clk,
  input         io_active_clk,
  input         io_exu_flush_final,
  input         io_dec_tlu_flush_lower_wb,
  input         io_dec_tlu_flush_err_wb,
  input         io_dec_tlu_i0_commit_cmt,
  input         io_dec_tlu_force_halt,
  input  [30:0] io_ifc_fetch_addr_bf,
  input         io_ifc_fetch_uncacheable_bf,
  input         io_ifc_fetch_req_bf,
  input         io_ifc_fetch_req_bf_raw,
  input         io_ifc_iccm_access_bf,
  input         io_ifc_region_acc_fault_bf,
  input         io_ifc_dma_access_ok,
  input         io_dec_tlu_fence_i_wb,
  input         io_ifu_bp_hit_taken_f,
  input         io_ifu_bp_inst_mask_f,
  input         io_ifu_axi_arready,
  input         io_ifu_axi_rvalid,
  input  [2:0]  io_ifu_axi_rid,
  input  [63:0] io_ifu_axi_rdata,
  input  [1:0]  io_ifu_axi_rresp,
  input         io_ifu_bus_clk_en,
  input         io_dma_iccm_req,
  input  [31:0] io_dma_mem_addr,
  input  [2:0]  io_dma_mem_sz,
  input         io_dma_mem_write,
  input  [63:0] io_dma_mem_wdata,
  input  [2:0]  io_dma_mem_tag,
  input  [63:0] io_ic_rd_data,
  input  [70:0] io_ic_debug_rd_data,
  input  [25:0] io_ictag_debug_rd_data,
  input  [1:0]  io_ic_eccerr,
  input  [1:0]  io_ic_parerr,
  input  [1:0]  io_ic_rd_hit,
  input         io_ic_tag_perr,
  input  [63:0] io_iccm_rd_data,
  input  [77:0] io_iccm_rd_data_ecc,
  input  [1:0]  io_ifu_fetch_val,
  input  [70:0] io_dec_tlu_ic_diag_pkt_icache_wrdata,
  input  [16:0] io_dec_tlu_ic_diag_pkt_icache_dicawics,
  input         io_dec_tlu_ic_diag_pkt_icache_rd_valid,
  input         io_dec_tlu_ic_diag_pkt_icache_wr_valid,
  output        io_ifu_miss_state_idle,
  output        io_ifu_ic_mb_empty,
  output        io_ic_dma_active,
  output        io_ic_write_stall,
  output        io_ifu_pmu_ic_miss,
  output        io_ifu_pmu_ic_hit,
  output        io_ifu_pmu_bus_error,
  output        io_ifu_pmu_bus_busy,
  output        io_ifu_pmu_bus_trxn,
  output        io_ifu_axi_awvalid,
  output [2:0]  io_ifu_axi_awid,
  output [31:0] io_ifu_axi_awaddr,
  output [3:0]  io_ifu_axi_awregion,
  output [7:0]  io_ifu_axi_awlen,
  output [2:0]  io_ifu_axi_awsize,
  output [1:0]  io_ifu_axi_awburst,
  output        io_ifu_axi_awlock,
  output [3:0]  io_ifu_axi_awcache,
  output [2:0]  io_ifu_axi_awprot,
  output [3:0]  io_ifu_axi_awqos,
  output        io_ifu_axi_wvalid,
  output [63:0] io_ifu_axi_wdata,
  output [7:0]  io_ifu_axi_wstrb,
  output        io_ifu_axi_wlast,
  output        io_ifu_axi_bready,
  output        io_ifu_axi_arvalid,
  output [2:0]  io_ifu_axi_arid,
  output [31:0] io_ifu_axi_araddr,
  output [3:0]  io_ifu_axi_arregion,
  output [7:0]  io_ifu_axi_arlen,
  output [2:0]  io_ifu_axi_arsize,
  output [1:0]  io_ifu_axi_arburst,
  output        io_ifu_axi_arlock,
  output [3:0]  io_ifu_axi_arcache,
  output [2:0]  io_ifu_axi_arprot,
  output [3:0]  io_ifu_axi_arqos,
  output        io_ifu_axi_rready,
  output        io_iccm_dma_ecc_error,
  output        io_iccm_dma_rvalid,
  output [63:0] io_iccm_dma_rdata,
  output [2:0]  io_iccm_dma_rtag,
  output        io_iccm_ready,
  output [30:0] io_ic_rw_addr,
  output [1:0]  io_ic_wr_en,
  output        io_ic_rd_en,
  output [70:0] io_ic_wr_data_0,
  output [70:0] io_ic_wr_data_1,
  output [70:0] io_ic_debug_wr_data,
  output [70:0] io_ifu_ic_debug_rd_data,
  output [9:0]  io_ic_debug_addr,
  output        io_ic_debug_rd_en,
  output        io_ic_debug_wr_en,
  output        io_ic_debug_tag_array,
  output [1:0]  io_ic_debug_way,
  output [1:0]  io_ic_tag_valid,
  output [14:0] io_iccm_rw_addr,
  output        io_iccm_wren,
  output        io_iccm_rden,
  output [77:0] io_iccm_wr_data,
  output [2:0]  io_iccm_wr_size,
  output        io_ic_hit_f,
  output        io_ic_access_fault_f,
  output [1:0]  io_ic_access_fault_type_f,
  output        io_iccm_rd_ecc_single_err,
  output        io_iccm_rd_ecc_double_err,
  output        io_ic_error_start,
  output        io_ifu_async_error_start,
  output        io_iccm_dma_sb_error,
  output [1:0]  io_ic_fetch_val_f,
  output [31:0] io_ic_data_f,
  output [63:0] io_ic_premux_data,
  output        io_ic_sel_premux_data,
  input         io_dec_tlu_core_ecc_disable,
  output        io_ifu_ic_debug_rd_data_valid,
  output        io_iccm_buf_correct_ecc,
  output        io_iccm_correction_state,
  input         io_scan_mode
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [63:0] _RAND_163;
  reg [63:0] _RAND_164;
  reg [63:0] _RAND_165;
  reg [63:0] _RAND_166;
  reg [63:0] _RAND_167;
  reg [63:0] _RAND_168;
  reg [63:0] _RAND_169;
  reg [63:0] _RAND_170;
  reg [63:0] _RAND_171;
  reg [63:0] _RAND_172;
  reg [63:0] _RAND_173;
  reg [63:0] _RAND_174;
  reg [63:0] _RAND_175;
  reg [63:0] _RAND_176;
  reg [63:0] _RAND_177;
  reg [63:0] _RAND_178;
  reg [63:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [95:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [63:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [63:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
`endif // RANDOMIZE_REG_INIT
  reg  flush_final_f; // @[el2_ifu_mem_ctl.scala 180:30]
  reg  ifc_fetch_req_f_raw; // @[el2_ifu_mem_ctl.scala 315:36]
  wire  _T_318 = ~io_exu_flush_final; // @[el2_ifu_mem_ctl.scala 316:44]
  wire  ifc_fetch_req_f = ifc_fetch_req_f_raw & _T_318; // @[el2_ifu_mem_ctl.scala 316:42]
  reg [2:0] miss_state; // @[Reg.scala 27:20]
  wire  miss_pending = miss_state != 3'h0; // @[el2_ifu_mem_ctl.scala 248:30]
  reg  scnd_miss_req_q; // @[el2_ifu_mem_ctl.scala 540:52]
  wire  scnd_miss_req = scnd_miss_req_q & _T_318; // @[el2_ifu_mem_ctl.scala 542:36]
  wire  debug_c1_clken = io_ic_debug_rd_en | io_ic_debug_wr_en; // @[el2_ifu_mem_ctl.scala 182:42]
  wire [3:0] ic_fetch_val_int_f = {2'h0,io_ic_fetch_val_f}; // @[Cat.scala 29:58]
  reg [30:0] ifu_fetch_addr_int_f; // @[el2_ifu_mem_ctl.scala 303:34]
  wire [4:0] _GEN_463 = {{1'd0}, ic_fetch_val_int_f}; // @[el2_ifu_mem_ctl.scala 657:53]
  wire [4:0] ic_fetch_val_shift_right = _GEN_463 << ifu_fetch_addr_int_f[0]; // @[el2_ifu_mem_ctl.scala 657:53]
  wire [1:0] _GEN_464 = {{1'd0}, _T_318}; // @[el2_ifu_mem_ctl.scala 660:91]
  wire [1:0] _T_3070 = ic_fetch_val_shift_right[3:2] & _GEN_464; // @[el2_ifu_mem_ctl.scala 660:91]
  reg  ifc_iccm_access_f; // @[el2_ifu_mem_ctl.scala 317:31]
  wire  fetch_req_iccm_f = ifc_fetch_req_f & ifc_iccm_access_f; // @[el2_ifu_mem_ctl.scala 270:46]
  wire [1:0] _GEN_465 = {{1'd0}, fetch_req_iccm_f}; // @[el2_ifu_mem_ctl.scala 660:113]
  wire [1:0] _T_3071 = _T_3070 & _GEN_465; // @[el2_ifu_mem_ctl.scala 660:113]
  reg  iccm_dma_rvalid_in; // @[el2_ifu_mem_ctl.scala 646:59]
  wire [1:0] _GEN_466 = {{1'd0}, iccm_dma_rvalid_in}; // @[el2_ifu_mem_ctl.scala 660:130]
  wire [1:0] _T_3072 = _T_3071 | _GEN_466; // @[el2_ifu_mem_ctl.scala 660:130]
  wire  _T_3073 = ~io_dec_tlu_core_ecc_disable; // @[el2_ifu_mem_ctl.scala 660:154]
  wire [1:0] _GEN_467 = {{1'd0}, _T_3073}; // @[el2_ifu_mem_ctl.scala 660:152]
  wire [1:0] _T_3074 = _T_3072 & _GEN_467; // @[el2_ifu_mem_ctl.scala 660:152]
  wire [1:0] _T_3063 = ic_fetch_val_shift_right[1:0] & _GEN_464; // @[el2_ifu_mem_ctl.scala 660:91]
  wire [1:0] _T_3064 = _T_3063 & _GEN_465; // @[el2_ifu_mem_ctl.scala 660:113]
  wire [1:0] _T_3065 = _T_3064 | _GEN_466; // @[el2_ifu_mem_ctl.scala 660:130]
  wire [1:0] _T_3067 = _T_3065 & _GEN_467; // @[el2_ifu_mem_ctl.scala 660:152]
  wire [3:0] iccm_ecc_word_enable = {_T_3074,_T_3067}; // @[Cat.scala 29:58]
  wire  _T_3174 = ^io_iccm_rd_data_ecc[31:0]; // @[el2_lib.scala 301:30]
  wire  _T_3175 = ^io_iccm_rd_data_ecc[38:32]; // @[el2_lib.scala 301:44]
  wire  _T_3176 = _T_3174 ^ _T_3175; // @[el2_lib.scala 301:35]
  wire [5:0] _T_3184 = {io_iccm_rd_data_ecc[31],io_iccm_rd_data_ecc[30],io_iccm_rd_data_ecc[29],io_iccm_rd_data_ecc[28],io_iccm_rd_data_ecc[27],io_iccm_rd_data_ecc[26]}; // @[el2_lib.scala 301:76]
  wire  _T_3185 = ^_T_3184; // @[el2_lib.scala 301:83]
  wire  _T_3186 = io_iccm_rd_data_ecc[37] ^ _T_3185; // @[el2_lib.scala 301:71]
  wire [6:0] _T_3193 = {io_iccm_rd_data_ecc[17],io_iccm_rd_data_ecc[16],io_iccm_rd_data_ecc[15],io_iccm_rd_data_ecc[14],io_iccm_rd_data_ecc[13],io_iccm_rd_data_ecc[12],io_iccm_rd_data_ecc[11]}; // @[el2_lib.scala 301:103]
  wire [14:0] _T_3201 = {io_iccm_rd_data_ecc[25],io_iccm_rd_data_ecc[24],io_iccm_rd_data_ecc[23],io_iccm_rd_data_ecc[22],io_iccm_rd_data_ecc[21],io_iccm_rd_data_ecc[20],io_iccm_rd_data_ecc[19],io_iccm_rd_data_ecc[18],_T_3193}; // @[el2_lib.scala 301:103]
  wire  _T_3202 = ^_T_3201; // @[el2_lib.scala 301:110]
  wire  _T_3203 = io_iccm_rd_data_ecc[36] ^ _T_3202; // @[el2_lib.scala 301:98]
  wire [6:0] _T_3210 = {io_iccm_rd_data_ecc[10],io_iccm_rd_data_ecc[9],io_iccm_rd_data_ecc[8],io_iccm_rd_data_ecc[7],io_iccm_rd_data_ecc[6],io_iccm_rd_data_ecc[5],io_iccm_rd_data_ecc[4]}; // @[el2_lib.scala 301:130]
  wire [14:0] _T_3218 = {io_iccm_rd_data_ecc[25],io_iccm_rd_data_ecc[24],io_iccm_rd_data_ecc[23],io_iccm_rd_data_ecc[22],io_iccm_rd_data_ecc[21],io_iccm_rd_data_ecc[20],io_iccm_rd_data_ecc[19],io_iccm_rd_data_ecc[18],_T_3210}; // @[el2_lib.scala 301:130]
  wire  _T_3219 = ^_T_3218; // @[el2_lib.scala 301:137]
  wire  _T_3220 = io_iccm_rd_data_ecc[35] ^ _T_3219; // @[el2_lib.scala 301:125]
  wire [8:0] _T_3229 = {io_iccm_rd_data_ecc[15],io_iccm_rd_data_ecc[14],io_iccm_rd_data_ecc[10],io_iccm_rd_data_ecc[9],io_iccm_rd_data_ecc[8],io_iccm_rd_data_ecc[7],io_iccm_rd_data_ecc[3],io_iccm_rd_data_ecc[2],io_iccm_rd_data_ecc[1]}; // @[el2_lib.scala 301:157]
  wire [17:0] _T_3238 = {io_iccm_rd_data_ecc[31],io_iccm_rd_data_ecc[30],io_iccm_rd_data_ecc[29],io_iccm_rd_data_ecc[25],io_iccm_rd_data_ecc[24],io_iccm_rd_data_ecc[23],io_iccm_rd_data_ecc[22],io_iccm_rd_data_ecc[17],io_iccm_rd_data_ecc[16],_T_3229}; // @[el2_lib.scala 301:157]
  wire  _T_3239 = ^_T_3238; // @[el2_lib.scala 301:164]
  wire  _T_3240 = io_iccm_rd_data_ecc[34] ^ _T_3239; // @[el2_lib.scala 301:152]
  wire [8:0] _T_3249 = {io_iccm_rd_data_ecc[13],io_iccm_rd_data_ecc[12],io_iccm_rd_data_ecc[10],io_iccm_rd_data_ecc[9],io_iccm_rd_data_ecc[6],io_iccm_rd_data_ecc[5],io_iccm_rd_data_ecc[3],io_iccm_rd_data_ecc[2],io_iccm_rd_data_ecc[0]}; // @[el2_lib.scala 301:184]
  wire [17:0] _T_3258 = {io_iccm_rd_data_ecc[31],io_iccm_rd_data_ecc[28],io_iccm_rd_data_ecc[27],io_iccm_rd_data_ecc[25],io_iccm_rd_data_ecc[24],io_iccm_rd_data_ecc[21],io_iccm_rd_data_ecc[20],io_iccm_rd_data_ecc[17],io_iccm_rd_data_ecc[16],_T_3249}; // @[el2_lib.scala 301:184]
  wire  _T_3259 = ^_T_3258; // @[el2_lib.scala 301:191]
  wire  _T_3260 = io_iccm_rd_data_ecc[33] ^ _T_3259; // @[el2_lib.scala 301:179]
  wire [8:0] _T_3269 = {io_iccm_rd_data_ecc[13],io_iccm_rd_data_ecc[11],io_iccm_rd_data_ecc[10],io_iccm_rd_data_ecc[8],io_iccm_rd_data_ecc[6],io_iccm_rd_data_ecc[4],io_iccm_rd_data_ecc[3],io_iccm_rd_data_ecc[1],io_iccm_rd_data_ecc[0]}; // @[el2_lib.scala 301:211]
  wire [17:0] _T_3278 = {io_iccm_rd_data_ecc[30],io_iccm_rd_data_ecc[28],io_iccm_rd_data_ecc[26],io_iccm_rd_data_ecc[25],io_iccm_rd_data_ecc[23],io_iccm_rd_data_ecc[21],io_iccm_rd_data_ecc[19],io_iccm_rd_data_ecc[17],io_iccm_rd_data_ecc[15],_T_3269}; // @[el2_lib.scala 301:211]
  wire  _T_3279 = ^_T_3278; // @[el2_lib.scala 301:218]
  wire  _T_3280 = io_iccm_rd_data_ecc[32] ^ _T_3279; // @[el2_lib.scala 301:206]
  wire [6:0] _T_3286 = {_T_3176,_T_3186,_T_3203,_T_3220,_T_3240,_T_3260,_T_3280}; // @[Cat.scala 29:58]
  wire  _T_3287 = _T_3286 != 7'h0; // @[el2_lib.scala 302:44]
  wire  _T_3288 = iccm_ecc_word_enable[0] & _T_3287; // @[el2_lib.scala 302:32]
  wire  _T_3290 = _T_3288 & _T_3286[6]; // @[el2_lib.scala 302:53]
  wire  _T_3559 = ^io_iccm_rd_data_ecc[70:39]; // @[el2_lib.scala 301:30]
  wire  _T_3560 = ^io_iccm_rd_data_ecc[77:71]; // @[el2_lib.scala 301:44]
  wire  _T_3561 = _T_3559 ^ _T_3560; // @[el2_lib.scala 301:35]
  wire [5:0] _T_3569 = {io_iccm_rd_data_ecc[70],io_iccm_rd_data_ecc[69],io_iccm_rd_data_ecc[68],io_iccm_rd_data_ecc[67],io_iccm_rd_data_ecc[66],io_iccm_rd_data_ecc[65]}; // @[el2_lib.scala 301:76]
  wire  _T_3570 = ^_T_3569; // @[el2_lib.scala 301:83]
  wire  _T_3571 = io_iccm_rd_data_ecc[76] ^ _T_3570; // @[el2_lib.scala 301:71]
  wire [6:0] _T_3578 = {io_iccm_rd_data_ecc[56],io_iccm_rd_data_ecc[55],io_iccm_rd_data_ecc[54],io_iccm_rd_data_ecc[53],io_iccm_rd_data_ecc[52],io_iccm_rd_data_ecc[51],io_iccm_rd_data_ecc[50]}; // @[el2_lib.scala 301:103]
  wire [14:0] _T_3586 = {io_iccm_rd_data_ecc[64],io_iccm_rd_data_ecc[63],io_iccm_rd_data_ecc[62],io_iccm_rd_data_ecc[61],io_iccm_rd_data_ecc[60],io_iccm_rd_data_ecc[59],io_iccm_rd_data_ecc[58],io_iccm_rd_data_ecc[57],_T_3578}; // @[el2_lib.scala 301:103]
  wire  _T_3587 = ^_T_3586; // @[el2_lib.scala 301:110]
  wire  _T_3588 = io_iccm_rd_data_ecc[75] ^ _T_3587; // @[el2_lib.scala 301:98]
  wire [6:0] _T_3595 = {io_iccm_rd_data_ecc[49],io_iccm_rd_data_ecc[48],io_iccm_rd_data_ecc[47],io_iccm_rd_data_ecc[46],io_iccm_rd_data_ecc[45],io_iccm_rd_data_ecc[44],io_iccm_rd_data_ecc[43]}; // @[el2_lib.scala 301:130]
  wire [14:0] _T_3603 = {io_iccm_rd_data_ecc[64],io_iccm_rd_data_ecc[63],io_iccm_rd_data_ecc[62],io_iccm_rd_data_ecc[61],io_iccm_rd_data_ecc[60],io_iccm_rd_data_ecc[59],io_iccm_rd_data_ecc[58],io_iccm_rd_data_ecc[57],_T_3595}; // @[el2_lib.scala 301:130]
  wire  _T_3604 = ^_T_3603; // @[el2_lib.scala 301:137]
  wire  _T_3605 = io_iccm_rd_data_ecc[74] ^ _T_3604; // @[el2_lib.scala 301:125]
  wire [8:0] _T_3614 = {io_iccm_rd_data_ecc[54],io_iccm_rd_data_ecc[53],io_iccm_rd_data_ecc[49],io_iccm_rd_data_ecc[48],io_iccm_rd_data_ecc[47],io_iccm_rd_data_ecc[46],io_iccm_rd_data_ecc[42],io_iccm_rd_data_ecc[41],io_iccm_rd_data_ecc[40]}; // @[el2_lib.scala 301:157]
  wire [17:0] _T_3623 = {io_iccm_rd_data_ecc[70],io_iccm_rd_data_ecc[69],io_iccm_rd_data_ecc[68],io_iccm_rd_data_ecc[64],io_iccm_rd_data_ecc[63],io_iccm_rd_data_ecc[62],io_iccm_rd_data_ecc[61],io_iccm_rd_data_ecc[56],io_iccm_rd_data_ecc[55],_T_3614}; // @[el2_lib.scala 301:157]
  wire  _T_3624 = ^_T_3623; // @[el2_lib.scala 301:164]
  wire  _T_3625 = io_iccm_rd_data_ecc[73] ^ _T_3624; // @[el2_lib.scala 301:152]
  wire [8:0] _T_3634 = {io_iccm_rd_data_ecc[52],io_iccm_rd_data_ecc[51],io_iccm_rd_data_ecc[49],io_iccm_rd_data_ecc[48],io_iccm_rd_data_ecc[45],io_iccm_rd_data_ecc[44],io_iccm_rd_data_ecc[42],io_iccm_rd_data_ecc[41],io_iccm_rd_data_ecc[39]}; // @[el2_lib.scala 301:184]
  wire [17:0] _T_3643 = {io_iccm_rd_data_ecc[70],io_iccm_rd_data_ecc[67],io_iccm_rd_data_ecc[66],io_iccm_rd_data_ecc[64],io_iccm_rd_data_ecc[63],io_iccm_rd_data_ecc[60],io_iccm_rd_data_ecc[59],io_iccm_rd_data_ecc[56],io_iccm_rd_data_ecc[55],_T_3634}; // @[el2_lib.scala 301:184]
  wire  _T_3644 = ^_T_3643; // @[el2_lib.scala 301:191]
  wire  _T_3645 = io_iccm_rd_data_ecc[72] ^ _T_3644; // @[el2_lib.scala 301:179]
  wire [8:0] _T_3654 = {io_iccm_rd_data_ecc[52],io_iccm_rd_data_ecc[50],io_iccm_rd_data_ecc[49],io_iccm_rd_data_ecc[47],io_iccm_rd_data_ecc[45],io_iccm_rd_data_ecc[43],io_iccm_rd_data_ecc[42],io_iccm_rd_data_ecc[40],io_iccm_rd_data_ecc[39]}; // @[el2_lib.scala 301:211]
  wire [17:0] _T_3663 = {io_iccm_rd_data_ecc[69],io_iccm_rd_data_ecc[67],io_iccm_rd_data_ecc[65],io_iccm_rd_data_ecc[64],io_iccm_rd_data_ecc[62],io_iccm_rd_data_ecc[60],io_iccm_rd_data_ecc[58],io_iccm_rd_data_ecc[56],io_iccm_rd_data_ecc[54],_T_3654}; // @[el2_lib.scala 301:211]
  wire  _T_3664 = ^_T_3663; // @[el2_lib.scala 301:218]
  wire  _T_3665 = io_iccm_rd_data_ecc[71] ^ _T_3664; // @[el2_lib.scala 301:206]
  wire [6:0] _T_3671 = {_T_3561,_T_3571,_T_3588,_T_3605,_T_3625,_T_3645,_T_3665}; // @[Cat.scala 29:58]
  wire  _T_3672 = _T_3671 != 7'h0; // @[el2_lib.scala 302:44]
  wire  _T_3673 = iccm_ecc_word_enable[1] & _T_3672; // @[el2_lib.scala 302:32]
  wire  _T_3675 = _T_3673 & _T_3671[6]; // @[el2_lib.scala 302:53]
  wire [1:0] iccm_single_ecc_error = {_T_3290,_T_3675}; // @[Cat.scala 29:58]
  wire  _T_3 = |iccm_single_ecc_error; // @[el2_ifu_mem_ctl.scala 185:52]
  reg  dma_iccm_req_f; // @[el2_ifu_mem_ctl.scala 624:51]
  wire  _T_6 = io_iccm_rd_ecc_single_err | io_ic_error_start; // @[el2_ifu_mem_ctl.scala 186:57]
  reg [2:0] perr_state; // @[Reg.scala 27:20]
  wire  _T_7 = perr_state == 3'h4; // @[el2_ifu_mem_ctl.scala 187:54]
  wire  iccm_correct_ecc = perr_state == 3'h3; // @[el2_ifu_mem_ctl.scala 469:34]
  wire  _T_8 = iccm_correct_ecc | _T_7; // @[el2_ifu_mem_ctl.scala 187:40]
  reg [1:0] err_stop_state; // @[Reg.scala 27:20]
  wire  _T_9 = err_stop_state == 2'h3; // @[el2_ifu_mem_ctl.scala 187:90]
  wire  _T_10 = _T_8 | _T_9; // @[el2_ifu_mem_ctl.scala 187:72]
  wire  _T_2439 = 2'h0 == err_stop_state; // @[Conditional.scala 37:30]
  wire  _T_2444 = 2'h1 == err_stop_state; // @[Conditional.scala 37:30]
  wire  _T_2464 = io_ifu_fetch_val == 2'h3; // @[el2_ifu_mem_ctl.scala 519:48]
  wire  two_byte_instr = io_ic_data_f[1:0] != 2'h3; // @[el2_ifu_mem_ctl.scala 385:42]
  wire  _T_2466 = io_ifu_fetch_val[0] & two_byte_instr; // @[el2_ifu_mem_ctl.scala 519:79]
  wire  _T_2467 = _T_2464 | _T_2466; // @[el2_ifu_mem_ctl.scala 519:56]
  wire  _T_2468 = io_exu_flush_final | io_dec_tlu_i0_commit_cmt; // @[el2_ifu_mem_ctl.scala 519:122]
  wire  _T_2469 = ~_T_2468; // @[el2_ifu_mem_ctl.scala 519:101]
  wire  _T_2470 = _T_2467 & _T_2469; // @[el2_ifu_mem_ctl.scala 519:99]
  wire  _T_2471 = 2'h2 == err_stop_state; // @[Conditional.scala 37:30]
  wire  _T_2485 = io_ifu_fetch_val[0] & _T_318; // @[el2_ifu_mem_ctl.scala 526:45]
  wire  _T_2486 = ~io_dec_tlu_i0_commit_cmt; // @[el2_ifu_mem_ctl.scala 526:69]
  wire  _T_2487 = _T_2485 & _T_2486; // @[el2_ifu_mem_ctl.scala 526:67]
  wire  _T_2488 = 2'h3 == err_stop_state; // @[Conditional.scala 37:30]
  wire  _GEN_54 = _T_2471 ? _T_2487 : _T_2488; // @[Conditional.scala 39:67]
  wire  _GEN_58 = _T_2444 ? _T_2470 : _GEN_54; // @[Conditional.scala 39:67]
  wire  err_stop_fetch = _T_2439 ? 1'h0 : _GEN_58; // @[Conditional.scala 40:58]
  wire  _T_11 = _T_10 | err_stop_fetch; // @[el2_ifu_mem_ctl.scala 187:112]
  wire  _T_13 = io_ifu_axi_rvalid & io_ifu_bus_clk_en; // @[el2_ifu_mem_ctl.scala 188:44]
  wire  _T_14 = _T_13 & io_ifu_axi_rready; // @[el2_ifu_mem_ctl.scala 188:65]
  wire  _T_228 = |io_ic_rd_hit; // @[el2_ifu_mem_ctl.scala 278:37]
  wire  _T_229 = ~_T_228; // @[el2_ifu_mem_ctl.scala 278:23]
  reg  reset_all_tags; // @[el2_ifu_mem_ctl.scala 692:53]
  wire  _T_230 = _T_229 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 278:41]
  wire  _T_208 = ~ifc_iccm_access_f; // @[el2_ifu_mem_ctl.scala 269:48]
  wire  _T_209 = ifc_fetch_req_f & _T_208; // @[el2_ifu_mem_ctl.scala 269:46]
  reg  ifc_region_acc_fault_final_f; // @[el2_ifu_mem_ctl.scala 319:42]
  wire  _T_210 = ~ifc_region_acc_fault_final_f; // @[el2_ifu_mem_ctl.scala 269:69]
  wire  fetch_req_icache_f = _T_209 & _T_210; // @[el2_ifu_mem_ctl.scala 269:67]
  wire  _T_231 = _T_230 & fetch_req_icache_f; // @[el2_ifu_mem_ctl.scala 278:59]
  wire  _T_232 = ~miss_pending; // @[el2_ifu_mem_ctl.scala 278:82]
  wire  _T_233 = _T_231 & _T_232; // @[el2_ifu_mem_ctl.scala 278:80]
  wire  _T_234 = _T_233 | scnd_miss_req; // @[el2_ifu_mem_ctl.scala 278:97]
  wire  ic_act_miss_f = _T_234 & _T_210; // @[el2_ifu_mem_ctl.scala 278:114]
  reg  ifu_bus_rvalid_unq_ff; // @[Reg.scala 27:20]
  reg  bus_ifu_bus_clk_en_ff; // @[el2_ifu_mem_ctl.scala 539:61]
  wire  ifu_bus_rvalid_ff = ifu_bus_rvalid_unq_ff & bus_ifu_bus_clk_en_ff; // @[el2_ifu_mem_ctl.scala 581:49]
  wire  bus_ifu_wr_en_ff = ifu_bus_rvalid_ff & miss_pending; // @[el2_ifu_mem_ctl.scala 608:41]
  reg  uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 305:33]
  reg [2:0] bus_data_beat_count; // @[el2_ifu_mem_ctl.scala 589:56]
  wire  _T_2590 = bus_data_beat_count == 3'h1; // @[el2_ifu_mem_ctl.scala 606:69]
  wire  _T_2591 = &bus_data_beat_count; // @[el2_ifu_mem_ctl.scala 606:101]
  wire  bus_last_data_beat = uncacheable_miss_ff ? _T_2590 : _T_2591; // @[el2_ifu_mem_ctl.scala 606:28]
  wire  _T_2537 = bus_ifu_wr_en_ff & bus_last_data_beat; // @[el2_ifu_mem_ctl.scala 585:68]
  wire  _T_2538 = ic_act_miss_f | _T_2537; // @[el2_ifu_mem_ctl.scala 585:48]
  wire  bus_reset_data_beat_cnt = _T_2538 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 585:91]
  wire  _T_2534 = ~bus_last_data_beat; // @[el2_ifu_mem_ctl.scala 584:50]
  wire  _T_2535 = bus_ifu_wr_en_ff & _T_2534; // @[el2_ifu_mem_ctl.scala 584:48]
  wire  _T_2536 = ~io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 584:72]
  wire  bus_inc_data_beat_cnt = _T_2535 & _T_2536; // @[el2_ifu_mem_ctl.scala 584:70]
  wire [2:0] _T_2542 = bus_data_beat_count + 3'h1; // @[el2_ifu_mem_ctl.scala 588:115]
  wire [2:0] _T_2544 = bus_inc_data_beat_cnt ? _T_2542 : 3'h0; // @[Mux.scala 27:72]
  wire  _T_2539 = ~bus_inc_data_beat_cnt; // @[el2_ifu_mem_ctl.scala 586:32]
  wire  _T_2540 = ~bus_reset_data_beat_cnt; // @[el2_ifu_mem_ctl.scala 586:57]
  wire  bus_hold_data_beat_cnt = _T_2539 & _T_2540; // @[el2_ifu_mem_ctl.scala 586:55]
  wire [2:0] _T_2545 = bus_hold_data_beat_cnt ? bus_data_beat_count : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] bus_new_data_beat_count = _T_2544 | _T_2545; // @[Mux.scala 27:72]
  wire  _T_15 = &bus_new_data_beat_count; // @[el2_ifu_mem_ctl.scala 188:111]
  wire  _T_16 = _T_14 & _T_15; // @[el2_ifu_mem_ctl.scala 188:85]
  wire  _T_17 = miss_state == 3'h5; // @[el2_ifu_mem_ctl.scala 189:39]
  wire  _T_25 = 3'h0 == miss_state; // @[Conditional.scala 37:30]
  wire  _T_27 = ic_act_miss_f & _T_318; // @[el2_ifu_mem_ctl.scala 195:43]
  wire [2:0] _T_29 = _T_27 ? 3'h1 : 3'h2; // @[el2_ifu_mem_ctl.scala 195:27]
  wire  _T_32 = 3'h1 == miss_state; // @[Conditional.scala 37:30]
  wire [4:0] byp_fetch_index = ifu_fetch_addr_int_f[4:0]; // @[el2_ifu_mem_ctl.scala 421:45]
  wire  _T_2109 = byp_fetch_index[4:2] == 3'h0; // @[el2_ifu_mem_ctl.scala 442:127]
  reg [7:0] ic_miss_buff_data_valid; // @[el2_ifu_mem_ctl.scala 398:60]
  wire  _T_2140 = _T_2109 & ic_miss_buff_data_valid[0]; // @[Mux.scala 27:72]
  wire  _T_2113 = byp_fetch_index[4:2] == 3'h1; // @[el2_ifu_mem_ctl.scala 442:127]
  wire  _T_2141 = _T_2113 & ic_miss_buff_data_valid[1]; // @[Mux.scala 27:72]
  wire  _T_2148 = _T_2140 | _T_2141; // @[Mux.scala 27:72]
  wire  _T_2117 = byp_fetch_index[4:2] == 3'h2; // @[el2_ifu_mem_ctl.scala 442:127]
  wire  _T_2142 = _T_2117 & ic_miss_buff_data_valid[2]; // @[Mux.scala 27:72]
  wire  _T_2149 = _T_2148 | _T_2142; // @[Mux.scala 27:72]
  wire  _T_2121 = byp_fetch_index[4:2] == 3'h3; // @[el2_ifu_mem_ctl.scala 442:127]
  wire  _T_2143 = _T_2121 & ic_miss_buff_data_valid[3]; // @[Mux.scala 27:72]
  wire  _T_2150 = _T_2149 | _T_2143; // @[Mux.scala 27:72]
  wire  _T_2125 = byp_fetch_index[4:2] == 3'h4; // @[el2_ifu_mem_ctl.scala 442:127]
  wire  _T_2144 = _T_2125 & ic_miss_buff_data_valid[4]; // @[Mux.scala 27:72]
  wire  _T_2151 = _T_2150 | _T_2144; // @[Mux.scala 27:72]
  wire  _T_2129 = byp_fetch_index[4:2] == 3'h5; // @[el2_ifu_mem_ctl.scala 442:127]
  wire  _T_2145 = _T_2129 & ic_miss_buff_data_valid[5]; // @[Mux.scala 27:72]
  wire  _T_2152 = _T_2151 | _T_2145; // @[Mux.scala 27:72]
  wire  _T_2133 = byp_fetch_index[4:2] == 3'h6; // @[el2_ifu_mem_ctl.scala 442:127]
  wire  _T_2146 = _T_2133 & ic_miss_buff_data_valid[6]; // @[Mux.scala 27:72]
  wire  _T_2153 = _T_2152 | _T_2146; // @[Mux.scala 27:72]
  wire  _T_2137 = byp_fetch_index[4:2] == 3'h7; // @[el2_ifu_mem_ctl.scala 442:127]
  wire  _T_2147 = _T_2137 & ic_miss_buff_data_valid[7]; // @[Mux.scala 27:72]
  wire  ic_miss_buff_data_valid_bypass_index = _T_2153 | _T_2147; // @[Mux.scala 27:72]
  wire  _T_2195 = ~byp_fetch_index[1]; // @[el2_ifu_mem_ctl.scala 444:69]
  wire  _T_2196 = ic_miss_buff_data_valid_bypass_index & _T_2195; // @[el2_ifu_mem_ctl.scala 444:67]
  wire  _T_2198 = ~byp_fetch_index[0]; // @[el2_ifu_mem_ctl.scala 444:91]
  wire  _T_2199 = _T_2196 & _T_2198; // @[el2_ifu_mem_ctl.scala 444:89]
  wire  _T_2204 = _T_2196 & byp_fetch_index[0]; // @[el2_ifu_mem_ctl.scala 445:65]
  wire  _T_2205 = _T_2199 | _T_2204; // @[el2_ifu_mem_ctl.scala 444:112]
  wire  _T_2207 = ic_miss_buff_data_valid_bypass_index & byp_fetch_index[1]; // @[el2_ifu_mem_ctl.scala 446:43]
  wire  _T_2210 = _T_2207 & _T_2198; // @[el2_ifu_mem_ctl.scala 446:65]
  wire  _T_2211 = _T_2205 | _T_2210; // @[el2_ifu_mem_ctl.scala 445:88]
  wire  _T_2215 = _T_2207 & byp_fetch_index[0]; // @[el2_ifu_mem_ctl.scala 447:65]
  wire [2:0] byp_fetch_index_inc = ifu_fetch_addr_int_f[4:2] + 3'h1; // @[el2_ifu_mem_ctl.scala 424:75]
  wire  _T_2155 = byp_fetch_index_inc == 3'h0; // @[el2_ifu_mem_ctl.scala 443:110]
  wire  _T_2179 = _T_2155 & ic_miss_buff_data_valid[0]; // @[Mux.scala 27:72]
  wire  _T_2158 = byp_fetch_index_inc == 3'h1; // @[el2_ifu_mem_ctl.scala 443:110]
  wire  _T_2180 = _T_2158 & ic_miss_buff_data_valid[1]; // @[Mux.scala 27:72]
  wire  _T_2187 = _T_2179 | _T_2180; // @[Mux.scala 27:72]
  wire  _T_2161 = byp_fetch_index_inc == 3'h2; // @[el2_ifu_mem_ctl.scala 443:110]
  wire  _T_2181 = _T_2161 & ic_miss_buff_data_valid[2]; // @[Mux.scala 27:72]
  wire  _T_2188 = _T_2187 | _T_2181; // @[Mux.scala 27:72]
  wire  _T_2164 = byp_fetch_index_inc == 3'h3; // @[el2_ifu_mem_ctl.scala 443:110]
  wire  _T_2182 = _T_2164 & ic_miss_buff_data_valid[3]; // @[Mux.scala 27:72]
  wire  _T_2189 = _T_2188 | _T_2182; // @[Mux.scala 27:72]
  wire  _T_2167 = byp_fetch_index_inc == 3'h4; // @[el2_ifu_mem_ctl.scala 443:110]
  wire  _T_2183 = _T_2167 & ic_miss_buff_data_valid[4]; // @[Mux.scala 27:72]
  wire  _T_2190 = _T_2189 | _T_2183; // @[Mux.scala 27:72]
  wire  _T_2170 = byp_fetch_index_inc == 3'h5; // @[el2_ifu_mem_ctl.scala 443:110]
  wire  _T_2184 = _T_2170 & ic_miss_buff_data_valid[5]; // @[Mux.scala 27:72]
  wire  _T_2191 = _T_2190 | _T_2184; // @[Mux.scala 27:72]
  wire  _T_2173 = byp_fetch_index_inc == 3'h6; // @[el2_ifu_mem_ctl.scala 443:110]
  wire  _T_2185 = _T_2173 & ic_miss_buff_data_valid[6]; // @[Mux.scala 27:72]
  wire  _T_2192 = _T_2191 | _T_2185; // @[Mux.scala 27:72]
  wire  _T_2176 = byp_fetch_index_inc == 3'h7; // @[el2_ifu_mem_ctl.scala 443:110]
  wire  _T_2186 = _T_2176 & ic_miss_buff_data_valid[7]; // @[Mux.scala 27:72]
  wire  ic_miss_buff_data_valid_inc_bypass_index = _T_2192 | _T_2186; // @[Mux.scala 27:72]
  wire  _T_2216 = _T_2215 & ic_miss_buff_data_valid_inc_bypass_index; // @[el2_ifu_mem_ctl.scala 447:87]
  wire  _T_2217 = _T_2211 | _T_2216; // @[el2_ifu_mem_ctl.scala 446:88]
  wire  _T_2221 = ic_miss_buff_data_valid_bypass_index & _T_2137; // @[el2_ifu_mem_ctl.scala 448:43]
  wire  miss_buff_hit_unq_f = _T_2217 | _T_2221; // @[el2_ifu_mem_ctl.scala 447:131]
  wire  _T_2237 = miss_state == 3'h4; // @[el2_ifu_mem_ctl.scala 453:55]
  wire  _T_2238 = miss_state == 3'h1; // @[el2_ifu_mem_ctl.scala 453:87]
  wire  _T_2239 = _T_2237 | _T_2238; // @[el2_ifu_mem_ctl.scala 453:74]
  wire  crit_byp_hit_f = miss_buff_hit_unq_f & _T_2239; // @[el2_ifu_mem_ctl.scala 453:41]
  wire  _T_2222 = miss_state == 3'h6; // @[el2_ifu_mem_ctl.scala 450:30]
  reg [30:0] imb_ff; // @[el2_ifu_mem_ctl.scala 306:20]
  wire  miss_wrap_f = imb_ff[5] != ifu_fetch_addr_int_f[6]; // @[el2_ifu_mem_ctl.scala 441:51]
  wire  _T_2223 = ~miss_wrap_f; // @[el2_ifu_mem_ctl.scala 450:68]
  wire  _T_2224 = miss_buff_hit_unq_f & _T_2223; // @[el2_ifu_mem_ctl.scala 450:66]
  wire  stream_hit_f = _T_2222 & _T_2224; // @[el2_ifu_mem_ctl.scala 450:43]
  wire  _T_216 = crit_byp_hit_f | stream_hit_f; // @[el2_ifu_mem_ctl.scala 273:35]
  wire  _T_217 = _T_216 & fetch_req_icache_f; // @[el2_ifu_mem_ctl.scala 273:52]
  wire  ic_byp_hit_f = _T_217 & miss_pending; // @[el2_ifu_mem_ctl.scala 273:73]
  reg  last_data_recieved_ff; // @[el2_ifu_mem_ctl.scala 591:58]
  wire  last_beat = bus_last_data_beat & bus_ifu_wr_en_ff; // @[el2_ifu_mem_ctl.scala 618:35]
  wire  _T_33 = bus_ifu_wr_en_ff & last_beat; // @[el2_ifu_mem_ctl.scala 199:113]
  wire  _T_34 = last_data_recieved_ff | _T_33; // @[el2_ifu_mem_ctl.scala 199:93]
  wire  _T_35 = ic_byp_hit_f & _T_34; // @[el2_ifu_mem_ctl.scala 199:67]
  wire  _T_36 = _T_35 & uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 199:127]
  wire  _T_37 = io_dec_tlu_force_halt | _T_36; // @[el2_ifu_mem_ctl.scala 199:51]
  wire  _T_39 = ~last_data_recieved_ff; // @[el2_ifu_mem_ctl.scala 200:30]
  wire  _T_40 = ic_byp_hit_f & _T_39; // @[el2_ifu_mem_ctl.scala 200:27]
  wire  _T_41 = _T_40 & uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 200:53]
  wire  _T_43 = ~ic_byp_hit_f; // @[el2_ifu_mem_ctl.scala 201:16]
  wire  _T_45 = _T_43 & _T_318; // @[el2_ifu_mem_ctl.scala 201:30]
  wire  _T_47 = _T_45 & _T_33; // @[el2_ifu_mem_ctl.scala 201:52]
  wire  _T_48 = _T_47 & uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 201:85]
  wire  _T_51 = ~uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 202:51]
  wire  _T_52 = _T_33 & _T_51; // @[el2_ifu_mem_ctl.scala 202:49]
  wire  _T_55 = ic_byp_hit_f & _T_318; // @[el2_ifu_mem_ctl.scala 203:33]
  wire  _T_57 = ~_T_33; // @[el2_ifu_mem_ctl.scala 203:57]
  wire  _T_58 = _T_55 & _T_57; // @[el2_ifu_mem_ctl.scala 203:55]
  wire  ifu_bp_hit_taken_q_f = io_ifu_bp_hit_taken_f & io_ic_hit_f; // @[el2_ifu_mem_ctl.scala 191:52]
  wire  _T_59 = ~ifu_bp_hit_taken_q_f; // @[el2_ifu_mem_ctl.scala 203:91]
  wire  _T_60 = _T_58 & _T_59; // @[el2_ifu_mem_ctl.scala 203:89]
  wire  _T_62 = _T_60 & _T_51; // @[el2_ifu_mem_ctl.scala 203:113]
  wire  _T_65 = bus_ifu_wr_en_ff & _T_318; // @[el2_ifu_mem_ctl.scala 204:39]
  wire  _T_68 = _T_65 & _T_57; // @[el2_ifu_mem_ctl.scala 204:61]
  wire  _T_70 = _T_68 & _T_59; // @[el2_ifu_mem_ctl.scala 204:95]
  wire  _T_72 = _T_70 & _T_51; // @[el2_ifu_mem_ctl.scala 204:119]
  wire  _T_80 = _T_47 & _T_51; // @[el2_ifu_mem_ctl.scala 205:100]
  wire  _T_82 = io_exu_flush_final | ifu_bp_hit_taken_q_f; // @[el2_ifu_mem_ctl.scala 206:44]
  wire  _T_85 = _T_82 & _T_57; // @[el2_ifu_mem_ctl.scala 206:68]
  wire [2:0] _T_87 = _T_85 ? 3'h2 : 3'h0; // @[el2_ifu_mem_ctl.scala 206:22]
  wire [2:0] _T_88 = _T_80 ? 3'h0 : _T_87; // @[el2_ifu_mem_ctl.scala 205:20]
  wire [2:0] _T_89 = _T_72 ? 3'h6 : _T_88; // @[el2_ifu_mem_ctl.scala 204:20]
  wire [2:0] _T_90 = _T_62 ? 3'h6 : _T_89; // @[el2_ifu_mem_ctl.scala 203:18]
  wire [2:0] _T_91 = _T_52 ? 3'h0 : _T_90; // @[el2_ifu_mem_ctl.scala 202:16]
  wire [2:0] _T_92 = _T_48 ? 3'h4 : _T_91; // @[el2_ifu_mem_ctl.scala 201:14]
  wire [2:0] _T_93 = _T_41 ? 3'h3 : _T_92; // @[el2_ifu_mem_ctl.scala 200:12]
  wire [2:0] _T_94 = _T_37 ? 3'h0 : _T_93; // @[el2_ifu_mem_ctl.scala 199:27]
  wire  _T_103 = 3'h4 == miss_state; // @[Conditional.scala 37:30]
  wire  _T_107 = 3'h6 == miss_state; // @[Conditional.scala 37:30]
  wire  _T_2234 = byp_fetch_index[4:1] == 4'h7; // @[el2_ifu_mem_ctl.scala 452:60]
  wire  _T_2235 = _T_2234 & ifc_fetch_req_f; // @[el2_ifu_mem_ctl.scala 452:92]
  wire  stream_eol_f = _T_2235 & stream_hit_f; // @[el2_ifu_mem_ctl.scala 452:110]
  wire  _T_109 = _T_82 | stream_eol_f; // @[el2_ifu_mem_ctl.scala 214:72]
  wire  _T_112 = _T_109 & _T_57; // @[el2_ifu_mem_ctl.scala 214:87]
  wire  _T_114 = _T_112 & _T_2536; // @[el2_ifu_mem_ctl.scala 214:122]
  wire [2:0] _T_116 = _T_114 ? 3'h2 : 3'h0; // @[el2_ifu_mem_ctl.scala 214:27]
  wire  _T_122 = 3'h3 == miss_state; // @[Conditional.scala 37:30]
  wire  _T_125 = io_exu_flush_final & _T_57; // @[el2_ifu_mem_ctl.scala 218:48]
  wire  _T_127 = _T_125 & _T_2536; // @[el2_ifu_mem_ctl.scala 218:82]
  wire [2:0] _T_129 = _T_127 ? 3'h2 : 3'h0; // @[el2_ifu_mem_ctl.scala 218:27]
  wire  _T_133 = 3'h2 == miss_state; // @[Conditional.scala 37:30]
  wire  _T_237 = io_ic_rd_hit == 2'h0; // @[el2_ifu_mem_ctl.scala 279:28]
  wire  _T_238 = _T_237 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 279:42]
  wire  _T_239 = _T_238 & fetch_req_icache_f; // @[el2_ifu_mem_ctl.scala 279:60]
  wire  _T_240 = miss_state == 3'h2; // @[el2_ifu_mem_ctl.scala 279:94]
  wire  _T_241 = _T_239 & _T_240; // @[el2_ifu_mem_ctl.scala 279:81]
  wire  _T_244 = imb_ff[30:5] != ifu_fetch_addr_int_f[30:5]; // @[el2_ifu_mem_ctl.scala 280:39]
  wire  _T_245 = _T_241 & _T_244; // @[el2_ifu_mem_ctl.scala 279:111]
  wire  _T_247 = _T_245 & _T_51; // @[el2_ifu_mem_ctl.scala 280:91]
  reg  sel_mb_addr_ff; // @[el2_ifu_mem_ctl.scala 333:51]
  wire  _T_248 = ~sel_mb_addr_ff; // @[el2_ifu_mem_ctl.scala 280:116]
  wire  _T_249 = _T_247 & _T_248; // @[el2_ifu_mem_ctl.scala 280:114]
  wire  ic_miss_under_miss_f = _T_249 & _T_210; // @[el2_ifu_mem_ctl.scala 280:132]
  wire  _T_136 = ic_miss_under_miss_f & _T_57; // @[el2_ifu_mem_ctl.scala 222:50]
  wire  _T_138 = _T_136 & _T_2536; // @[el2_ifu_mem_ctl.scala 222:84]
  wire  _T_257 = _T_231 & _T_240; // @[el2_ifu_mem_ctl.scala 281:85]
  wire  _T_260 = imb_ff[30:5] == ifu_fetch_addr_int_f[30:5]; // @[el2_ifu_mem_ctl.scala 282:39]
  wire  _T_261 = _T_260 | uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 282:91]
  wire  ic_ignore_2nd_miss_f = _T_257 & _T_261; // @[el2_ifu_mem_ctl.scala 281:117]
  wire  _T_142 = ic_ignore_2nd_miss_f & _T_57; // @[el2_ifu_mem_ctl.scala 223:35]
  wire  _T_144 = _T_142 & _T_2536; // @[el2_ifu_mem_ctl.scala 223:69]
  wire [2:0] _T_146 = _T_144 ? 3'h7 : 3'h0; // @[el2_ifu_mem_ctl.scala 223:12]
  wire [2:0] _T_147 = _T_138 ? 3'h5 : _T_146; // @[el2_ifu_mem_ctl.scala 222:27]
  wire  _T_152 = 3'h5 == miss_state; // @[Conditional.scala 37:30]
  wire [2:0] _T_155 = _T_33 ? 3'h0 : 3'h2; // @[el2_ifu_mem_ctl.scala 228:12]
  wire [2:0] _T_156 = io_exu_flush_final ? _T_155 : 3'h1; // @[el2_ifu_mem_ctl.scala 227:62]
  wire [2:0] _T_157 = io_dec_tlu_force_halt ? 3'h0 : _T_156; // @[el2_ifu_mem_ctl.scala 227:27]
  wire  _T_161 = 3'h7 == miss_state; // @[Conditional.scala 37:30]
  wire [2:0] _T_165 = io_exu_flush_final ? _T_155 : 3'h0; // @[el2_ifu_mem_ctl.scala 232:62]
  wire [2:0] _T_166 = io_dec_tlu_force_halt ? 3'h0 : _T_165; // @[el2_ifu_mem_ctl.scala 232:27]
  wire [2:0] _GEN_0 = _T_161 ? _T_166 : 3'h0; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_2 = _T_152 ? _T_157 : _GEN_0; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_4 = _T_133 ? _T_147 : _GEN_2; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_6 = _T_122 ? _T_129 : _GEN_4; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_8 = _T_107 ? _T_116 : _GEN_6; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_10 = _T_103 ? 3'h0 : _GEN_8; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_12 = _T_32 ? _T_94 : _GEN_10; // @[Conditional.scala 39:67]
  wire [2:0] miss_nxtstate = _T_25 ? _T_29 : _GEN_12; // @[Conditional.scala 40:58]
  wire  _T_18 = miss_nxtstate == 3'h5; // @[el2_ifu_mem_ctl.scala 189:71]
  wire  _T_19 = _T_17 | _T_18; // @[el2_ifu_mem_ctl.scala 189:55]
  wire  _T_20 = uncacheable_miss_ff >> _T_19; // @[el2_ifu_mem_ctl.scala 189:26]
  wire  _T_22 = ~_T_20; // @[el2_ifu_mem_ctl.scala 189:5]
  wire  _T_23 = _T_16 & _T_22; // @[el2_ifu_mem_ctl.scala 188:116]
  wire  scnd_miss_req_in = _T_23 & _T_318; // @[el2_ifu_mem_ctl.scala 189:89]
  wire  _T_31 = ic_act_miss_f & _T_2536; // @[el2_ifu_mem_ctl.scala 196:38]
  wire  _T_95 = io_dec_tlu_force_halt | io_exu_flush_final; // @[el2_ifu_mem_ctl.scala 207:46]
  wire  _T_96 = _T_95 | ic_byp_hit_f; // @[el2_ifu_mem_ctl.scala 207:67]
  wire  _T_97 = _T_96 | ifu_bp_hit_taken_q_f; // @[el2_ifu_mem_ctl.scala 207:82]
  wire  _T_99 = _T_97 | _T_33; // @[el2_ifu_mem_ctl.scala 207:105]
  wire  _T_101 = bus_ifu_wr_en_ff & _T_51; // @[el2_ifu_mem_ctl.scala 207:158]
  wire  _T_102 = _T_99 | _T_101; // @[el2_ifu_mem_ctl.scala 207:138]
  wire  _T_104 = io_exu_flush_final | flush_final_f; // @[el2_ifu_mem_ctl.scala 211:43]
  wire  _T_105 = _T_104 | ic_byp_hit_f; // @[el2_ifu_mem_ctl.scala 211:59]
  wire  _T_106 = _T_105 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 211:74]
  wire  _T_120 = _T_109 | _T_33; // @[el2_ifu_mem_ctl.scala 215:84]
  wire  _T_121 = _T_120 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 215:118]
  wire  _T_131 = io_exu_flush_final | _T_33; // @[el2_ifu_mem_ctl.scala 219:43]
  wire  _T_132 = _T_131 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 219:76]
  wire  _T_149 = _T_33 | ic_miss_under_miss_f; // @[el2_ifu_mem_ctl.scala 224:55]
  wire  _T_150 = _T_149 | ic_ignore_2nd_miss_f; // @[el2_ifu_mem_ctl.scala 224:78]
  wire  _T_151 = _T_150 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 224:101]
  wire  _T_159 = _T_33 | io_exu_flush_final; // @[el2_ifu_mem_ctl.scala 229:55]
  wire  _T_160 = _T_159 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 229:76]
  wire  _GEN_1 = _T_161 & _T_160; // @[Conditional.scala 39:67]
  wire  _GEN_3 = _T_152 ? _T_160 : _GEN_1; // @[Conditional.scala 39:67]
  wire  _GEN_5 = _T_133 ? _T_151 : _GEN_3; // @[Conditional.scala 39:67]
  wire  _GEN_7 = _T_122 ? _T_132 : _GEN_5; // @[Conditional.scala 39:67]
  wire  _GEN_9 = _T_107 ? _T_121 : _GEN_7; // @[Conditional.scala 39:67]
  wire  _GEN_11 = _T_103 ? _T_106 : _GEN_9; // @[Conditional.scala 39:67]
  wire  _GEN_13 = _T_32 ? _T_102 : _GEN_11; // @[Conditional.scala 39:67]
  wire  miss_state_en = _T_25 ? _T_31 : _GEN_13; // @[Conditional.scala 40:58]
  wire  _T_175 = ~flush_final_f; // @[el2_ifu_mem_ctl.scala 249:95]
  wire  _T_176 = _T_2237 & _T_175; // @[el2_ifu_mem_ctl.scala 249:93]
  wire  crit_wd_byp_ok_ff = _T_2238 | _T_176; // @[el2_ifu_mem_ctl.scala 249:58]
  wire  _T_179 = miss_pending & _T_57; // @[el2_ifu_mem_ctl.scala 250:36]
  wire  _T_181 = _T_2237 & io_exu_flush_final; // @[el2_ifu_mem_ctl.scala 250:106]
  wire  _T_182 = ~_T_181; // @[el2_ifu_mem_ctl.scala 250:72]
  wire  _T_183 = _T_179 & _T_182; // @[el2_ifu_mem_ctl.scala 250:70]
  wire  _T_185 = _T_2237 & crit_byp_hit_f; // @[el2_ifu_mem_ctl.scala 251:57]
  wire  _T_186 = ~_T_185; // @[el2_ifu_mem_ctl.scala 251:23]
  wire  _T_187 = _T_183 & _T_186; // @[el2_ifu_mem_ctl.scala 250:128]
  wire  _T_188 = _T_187 | ic_act_miss_f; // @[el2_ifu_mem_ctl.scala 251:77]
  wire  _T_189 = miss_nxtstate == 3'h4; // @[el2_ifu_mem_ctl.scala 252:36]
  wire  _T_190 = miss_pending & _T_189; // @[el2_ifu_mem_ctl.scala 252:19]
  wire  sel_hold_imb = _T_188 | _T_190; // @[el2_ifu_mem_ctl.scala 251:93]
  wire  _T_192 = _T_17 | ic_miss_under_miss_f; // @[el2_ifu_mem_ctl.scala 254:57]
  wire  sel_hold_imb_scnd = _T_192 & _T_175; // @[el2_ifu_mem_ctl.scala 254:81]
  reg  way_status_mb_scnd_ff; // @[el2_ifu_mem_ctl.scala 262:35]
  reg [6:0] _T_5115; // @[el2_ifu_mem_ctl.scala 720:14]
  wire [5:0] ifu_ic_rw_int_addr_ff = _T_5115[5:0]; // @[el2_ifu_mem_ctl.scala 719:27]
  wire [6:0] _GEN_472 = {{1'd0}, ifu_ic_rw_int_addr_ff}; // @[el2_ifu_mem_ctl.scala 716:121]
  wire  _T_4980 = _GEN_472 == 7'h7f; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4982 = _T_4980 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4471; // @[Reg.scala 27:20]
  wire  way_status_out_127 = _T_4471[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_473 = {{5'd0}, way_status_out_127}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4983 = _T_4982 & _GEN_473; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4976 = _GEN_472 == 7'h7e; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4978 = _T_4976 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4467; // @[Reg.scala 27:20]
  wire  way_status_out_126 = _T_4467[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_475 = {{5'd0}, way_status_out_126}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4979 = _T_4978 & _GEN_475; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4972 = _GEN_472 == 7'h7d; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4974 = _T_4972 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4463; // @[Reg.scala 27:20]
  wire  way_status_out_125 = _T_4463[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_477 = {{5'd0}, way_status_out_125}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4975 = _T_4974 & _GEN_477; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4968 = _GEN_472 == 7'h7c; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4970 = _T_4968 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4459; // @[Reg.scala 27:20]
  wire  way_status_out_124 = _T_4459[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_479 = {{5'd0}, way_status_out_124}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4971 = _T_4970 & _GEN_479; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4964 = _GEN_472 == 7'h7b; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4966 = _T_4964 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4455; // @[Reg.scala 27:20]
  wire  way_status_out_123 = _T_4455[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_481 = {{5'd0}, way_status_out_123}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4967 = _T_4966 & _GEN_481; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4960 = _GEN_472 == 7'h7a; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4962 = _T_4960 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4451; // @[Reg.scala 27:20]
  wire  way_status_out_122 = _T_4451[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_483 = {{5'd0}, way_status_out_122}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4963 = _T_4962 & _GEN_483; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4956 = _GEN_472 == 7'h79; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4958 = _T_4956 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4447; // @[Reg.scala 27:20]
  wire  way_status_out_121 = _T_4447[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_485 = {{5'd0}, way_status_out_121}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4959 = _T_4958 & _GEN_485; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4952 = _GEN_472 == 7'h78; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4954 = _T_4952 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4443; // @[Reg.scala 27:20]
  wire  way_status_out_120 = _T_4443[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_487 = {{5'd0}, way_status_out_120}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4955 = _T_4954 & _GEN_487; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4948 = _GEN_472 == 7'h77; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4950 = _T_4948 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4439; // @[Reg.scala 27:20]
  wire  way_status_out_119 = _T_4439[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_489 = {{5'd0}, way_status_out_119}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4951 = _T_4950 & _GEN_489; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4944 = _GEN_472 == 7'h76; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4946 = _T_4944 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4435; // @[Reg.scala 27:20]
  wire  way_status_out_118 = _T_4435[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_491 = {{5'd0}, way_status_out_118}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4947 = _T_4946 & _GEN_491; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [59:0] _T_4992 = {_T_4983,_T_4979,_T_4975,_T_4971,_T_4967,_T_4963,_T_4959,_T_4955,_T_4951,_T_4947}; // @[Cat.scala 29:58]
  wire  _T_4940 = _GEN_472 == 7'h75; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4942 = _T_4940 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4431; // @[Reg.scala 27:20]
  wire  way_status_out_117 = _T_4431[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_493 = {{5'd0}, way_status_out_117}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4943 = _T_4942 & _GEN_493; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4936 = _GEN_472 == 7'h74; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4938 = _T_4936 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4427; // @[Reg.scala 27:20]
  wire  way_status_out_116 = _T_4427[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_495 = {{5'd0}, way_status_out_116}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4939 = _T_4938 & _GEN_495; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4932 = _GEN_472 == 7'h73; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4934 = _T_4932 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4423; // @[Reg.scala 27:20]
  wire  way_status_out_115 = _T_4423[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_497 = {{5'd0}, way_status_out_115}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4935 = _T_4934 & _GEN_497; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4928 = _GEN_472 == 7'h72; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4930 = _T_4928 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4419; // @[Reg.scala 27:20]
  wire  way_status_out_114 = _T_4419[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_499 = {{5'd0}, way_status_out_114}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4931 = _T_4930 & _GEN_499; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4924 = _GEN_472 == 7'h71; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4926 = _T_4924 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4415; // @[Reg.scala 27:20]
  wire  way_status_out_113 = _T_4415[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_501 = {{5'd0}, way_status_out_113}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4927 = _T_4926 & _GEN_501; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4920 = _GEN_472 == 7'h70; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4922 = _T_4920 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4411; // @[Reg.scala 27:20]
  wire  way_status_out_112 = _T_4411[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_503 = {{5'd0}, way_status_out_112}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4923 = _T_4922 & _GEN_503; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4916 = _GEN_472 == 7'h6f; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4918 = _T_4916 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4407; // @[Reg.scala 27:20]
  wire  way_status_out_111 = _T_4407[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_505 = {{5'd0}, way_status_out_111}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4919 = _T_4918 & _GEN_505; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4912 = _GEN_472 == 7'h6e; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4914 = _T_4912 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4403; // @[Reg.scala 27:20]
  wire  way_status_out_110 = _T_4403[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_507 = {{5'd0}, way_status_out_110}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4915 = _T_4914 & _GEN_507; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4908 = _GEN_472 == 7'h6d; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4910 = _T_4908 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4399; // @[Reg.scala 27:20]
  wire  way_status_out_109 = _T_4399[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_509 = {{5'd0}, way_status_out_109}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4911 = _T_4910 & _GEN_509; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [113:0] _T_5001 = {_T_4992,_T_4943,_T_4939,_T_4935,_T_4931,_T_4927,_T_4923,_T_4919,_T_4915,_T_4911}; // @[Cat.scala 29:58]
  wire  _T_4904 = _GEN_472 == 7'h6c; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4906 = _T_4904 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4395; // @[Reg.scala 27:20]
  wire  way_status_out_108 = _T_4395[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_511 = {{5'd0}, way_status_out_108}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4907 = _T_4906 & _GEN_511; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4900 = _GEN_472 == 7'h6b; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4902 = _T_4900 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4391; // @[Reg.scala 27:20]
  wire  way_status_out_107 = _T_4391[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_513 = {{5'd0}, way_status_out_107}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4903 = _T_4902 & _GEN_513; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4896 = _GEN_472 == 7'h6a; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4898 = _T_4896 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4387; // @[Reg.scala 27:20]
  wire  way_status_out_106 = _T_4387[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_515 = {{5'd0}, way_status_out_106}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4899 = _T_4898 & _GEN_515; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4892 = _GEN_472 == 7'h69; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4894 = _T_4892 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4383; // @[Reg.scala 27:20]
  wire  way_status_out_105 = _T_4383[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_517 = {{5'd0}, way_status_out_105}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4895 = _T_4894 & _GEN_517; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4888 = _GEN_472 == 7'h68; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4890 = _T_4888 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4379; // @[Reg.scala 27:20]
  wire  way_status_out_104 = _T_4379[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_519 = {{5'd0}, way_status_out_104}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4891 = _T_4890 & _GEN_519; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4884 = _GEN_472 == 7'h67; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4886 = _T_4884 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4375; // @[Reg.scala 27:20]
  wire  way_status_out_103 = _T_4375[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_521 = {{5'd0}, way_status_out_103}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4887 = _T_4886 & _GEN_521; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4880 = _GEN_472 == 7'h66; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4882 = _T_4880 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4371; // @[Reg.scala 27:20]
  wire  way_status_out_102 = _T_4371[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_523 = {{5'd0}, way_status_out_102}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4883 = _T_4882 & _GEN_523; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4876 = _GEN_472 == 7'h65; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4878 = _T_4876 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4367; // @[Reg.scala 27:20]
  wire  way_status_out_101 = _T_4367[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_525 = {{5'd0}, way_status_out_101}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4879 = _T_4878 & _GEN_525; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4872 = _GEN_472 == 7'h64; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4874 = _T_4872 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4363; // @[Reg.scala 27:20]
  wire  way_status_out_100 = _T_4363[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_527 = {{5'd0}, way_status_out_100}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4875 = _T_4874 & _GEN_527; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [167:0] _T_5010 = {_T_5001,_T_4907,_T_4903,_T_4899,_T_4895,_T_4891,_T_4887,_T_4883,_T_4879,_T_4875}; // @[Cat.scala 29:58]
  wire  _T_4868 = _GEN_472 == 7'h63; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4870 = _T_4868 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4359; // @[Reg.scala 27:20]
  wire  way_status_out_99 = _T_4359[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_529 = {{5'd0}, way_status_out_99}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4871 = _T_4870 & _GEN_529; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4864 = _GEN_472 == 7'h62; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4866 = _T_4864 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4355; // @[Reg.scala 27:20]
  wire  way_status_out_98 = _T_4355[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_531 = {{5'd0}, way_status_out_98}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4867 = _T_4866 & _GEN_531; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4860 = _GEN_472 == 7'h61; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4862 = _T_4860 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4351; // @[Reg.scala 27:20]
  wire  way_status_out_97 = _T_4351[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_533 = {{5'd0}, way_status_out_97}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4863 = _T_4862 & _GEN_533; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4856 = _GEN_472 == 7'h60; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4858 = _T_4856 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4347; // @[Reg.scala 27:20]
  wire  way_status_out_96 = _T_4347[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_535 = {{5'd0}, way_status_out_96}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4859 = _T_4858 & _GEN_535; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4852 = _GEN_472 == 7'h5f; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4854 = _T_4852 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4343; // @[Reg.scala 27:20]
  wire  way_status_out_95 = _T_4343[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_537 = {{5'd0}, way_status_out_95}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4855 = _T_4854 & _GEN_537; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4848 = _GEN_472 == 7'h5e; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4850 = _T_4848 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4339; // @[Reg.scala 27:20]
  wire  way_status_out_94 = _T_4339[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_539 = {{5'd0}, way_status_out_94}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4851 = _T_4850 & _GEN_539; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4844 = _GEN_472 == 7'h5d; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4846 = _T_4844 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4335; // @[Reg.scala 27:20]
  wire  way_status_out_93 = _T_4335[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_541 = {{5'd0}, way_status_out_93}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4847 = _T_4846 & _GEN_541; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4840 = _GEN_472 == 7'h5c; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4842 = _T_4840 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4331; // @[Reg.scala 27:20]
  wire  way_status_out_92 = _T_4331[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_543 = {{5'd0}, way_status_out_92}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4843 = _T_4842 & _GEN_543; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4836 = _GEN_472 == 7'h5b; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4838 = _T_4836 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4327; // @[Reg.scala 27:20]
  wire  way_status_out_91 = _T_4327[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_545 = {{5'd0}, way_status_out_91}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4839 = _T_4838 & _GEN_545; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [221:0] _T_5019 = {_T_5010,_T_4871,_T_4867,_T_4863,_T_4859,_T_4855,_T_4851,_T_4847,_T_4843,_T_4839}; // @[Cat.scala 29:58]
  wire  _T_4832 = _GEN_472 == 7'h5a; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4834 = _T_4832 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4323; // @[Reg.scala 27:20]
  wire  way_status_out_90 = _T_4323[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_547 = {{5'd0}, way_status_out_90}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4835 = _T_4834 & _GEN_547; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4828 = _GEN_472 == 7'h59; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4830 = _T_4828 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4319; // @[Reg.scala 27:20]
  wire  way_status_out_89 = _T_4319[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_549 = {{5'd0}, way_status_out_89}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4831 = _T_4830 & _GEN_549; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4824 = _GEN_472 == 7'h58; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4826 = _T_4824 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4315; // @[Reg.scala 27:20]
  wire  way_status_out_88 = _T_4315[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_551 = {{5'd0}, way_status_out_88}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4827 = _T_4826 & _GEN_551; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4820 = _GEN_472 == 7'h57; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4822 = _T_4820 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4311; // @[Reg.scala 27:20]
  wire  way_status_out_87 = _T_4311[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_553 = {{5'd0}, way_status_out_87}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4823 = _T_4822 & _GEN_553; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4816 = _GEN_472 == 7'h56; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4818 = _T_4816 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4307; // @[Reg.scala 27:20]
  wire  way_status_out_86 = _T_4307[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_555 = {{5'd0}, way_status_out_86}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4819 = _T_4818 & _GEN_555; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4812 = _GEN_472 == 7'h55; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4814 = _T_4812 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4303; // @[Reg.scala 27:20]
  wire  way_status_out_85 = _T_4303[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_557 = {{5'd0}, way_status_out_85}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4815 = _T_4814 & _GEN_557; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4808 = _GEN_472 == 7'h54; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4810 = _T_4808 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4299; // @[Reg.scala 27:20]
  wire  way_status_out_84 = _T_4299[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_559 = {{5'd0}, way_status_out_84}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4811 = _T_4810 & _GEN_559; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4804 = _GEN_472 == 7'h53; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4806 = _T_4804 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4295; // @[Reg.scala 27:20]
  wire  way_status_out_83 = _T_4295[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_561 = {{5'd0}, way_status_out_83}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4807 = _T_4806 & _GEN_561; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4800 = _GEN_472 == 7'h52; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4802 = _T_4800 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4291; // @[Reg.scala 27:20]
  wire  way_status_out_82 = _T_4291[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_563 = {{5'd0}, way_status_out_82}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4803 = _T_4802 & _GEN_563; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [275:0] _T_5028 = {_T_5019,_T_4835,_T_4831,_T_4827,_T_4823,_T_4819,_T_4815,_T_4811,_T_4807,_T_4803}; // @[Cat.scala 29:58]
  wire  _T_4796 = _GEN_472 == 7'h51; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4798 = _T_4796 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4287; // @[Reg.scala 27:20]
  wire  way_status_out_81 = _T_4287[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_565 = {{5'd0}, way_status_out_81}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4799 = _T_4798 & _GEN_565; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4792 = _GEN_472 == 7'h50; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4794 = _T_4792 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4283; // @[Reg.scala 27:20]
  wire  way_status_out_80 = _T_4283[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_567 = {{5'd0}, way_status_out_80}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4795 = _T_4794 & _GEN_567; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4788 = _GEN_472 == 7'h4f; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4790 = _T_4788 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4279; // @[Reg.scala 27:20]
  wire  way_status_out_79 = _T_4279[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_569 = {{5'd0}, way_status_out_79}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4791 = _T_4790 & _GEN_569; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4784 = _GEN_472 == 7'h4e; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4786 = _T_4784 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4275; // @[Reg.scala 27:20]
  wire  way_status_out_78 = _T_4275[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_571 = {{5'd0}, way_status_out_78}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4787 = _T_4786 & _GEN_571; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4780 = _GEN_472 == 7'h4d; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4782 = _T_4780 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4271; // @[Reg.scala 27:20]
  wire  way_status_out_77 = _T_4271[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_573 = {{5'd0}, way_status_out_77}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4783 = _T_4782 & _GEN_573; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4776 = _GEN_472 == 7'h4c; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4778 = _T_4776 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4267; // @[Reg.scala 27:20]
  wire  way_status_out_76 = _T_4267[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_575 = {{5'd0}, way_status_out_76}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4779 = _T_4778 & _GEN_575; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4772 = _GEN_472 == 7'h4b; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4774 = _T_4772 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4263; // @[Reg.scala 27:20]
  wire  way_status_out_75 = _T_4263[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_577 = {{5'd0}, way_status_out_75}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4775 = _T_4774 & _GEN_577; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4768 = _GEN_472 == 7'h4a; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4770 = _T_4768 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4259; // @[Reg.scala 27:20]
  wire  way_status_out_74 = _T_4259[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_579 = {{5'd0}, way_status_out_74}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4771 = _T_4770 & _GEN_579; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4764 = _GEN_472 == 7'h49; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4766 = _T_4764 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4255; // @[Reg.scala 27:20]
  wire  way_status_out_73 = _T_4255[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_581 = {{5'd0}, way_status_out_73}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4767 = _T_4766 & _GEN_581; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [329:0] _T_5037 = {_T_5028,_T_4799,_T_4795,_T_4791,_T_4787,_T_4783,_T_4779,_T_4775,_T_4771,_T_4767}; // @[Cat.scala 29:58]
  wire  _T_4760 = _GEN_472 == 7'h48; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4762 = _T_4760 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4251; // @[Reg.scala 27:20]
  wire  way_status_out_72 = _T_4251[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_583 = {{5'd0}, way_status_out_72}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4763 = _T_4762 & _GEN_583; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4756 = _GEN_472 == 7'h47; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4758 = _T_4756 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4247; // @[Reg.scala 27:20]
  wire  way_status_out_71 = _T_4247[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_585 = {{5'd0}, way_status_out_71}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4759 = _T_4758 & _GEN_585; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4752 = _GEN_472 == 7'h46; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4754 = _T_4752 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4243; // @[Reg.scala 27:20]
  wire  way_status_out_70 = _T_4243[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_587 = {{5'd0}, way_status_out_70}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4755 = _T_4754 & _GEN_587; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4748 = _GEN_472 == 7'h45; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4750 = _T_4748 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4239; // @[Reg.scala 27:20]
  wire  way_status_out_69 = _T_4239[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_589 = {{5'd0}, way_status_out_69}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4751 = _T_4750 & _GEN_589; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4744 = _GEN_472 == 7'h44; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4746 = _T_4744 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4235; // @[Reg.scala 27:20]
  wire  way_status_out_68 = _T_4235[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_591 = {{5'd0}, way_status_out_68}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4747 = _T_4746 & _GEN_591; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4740 = _GEN_472 == 7'h43; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4742 = _T_4740 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4231; // @[Reg.scala 27:20]
  wire  way_status_out_67 = _T_4231[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_593 = {{5'd0}, way_status_out_67}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4743 = _T_4742 & _GEN_593; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4736 = _GEN_472 == 7'h42; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4738 = _T_4736 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4227; // @[Reg.scala 27:20]
  wire  way_status_out_66 = _T_4227[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_595 = {{5'd0}, way_status_out_66}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4739 = _T_4738 & _GEN_595; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4732 = _GEN_472 == 7'h41; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4734 = _T_4732 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4223; // @[Reg.scala 27:20]
  wire  way_status_out_65 = _T_4223[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_597 = {{5'd0}, way_status_out_65}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4735 = _T_4734 & _GEN_597; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4728 = _GEN_472 == 7'h40; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4730 = _T_4728 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4219; // @[Reg.scala 27:20]
  wire  way_status_out_64 = _T_4219[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_599 = {{5'd0}, way_status_out_64}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4731 = _T_4730 & _GEN_599; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [383:0] _T_5046 = {_T_5037,_T_4763,_T_4759,_T_4755,_T_4751,_T_4747,_T_4743,_T_4739,_T_4735,_T_4731}; // @[Cat.scala 29:58]
  wire  _T_4724 = ifu_ic_rw_int_addr_ff == 6'h3f; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4726 = _T_4724 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4215; // @[Reg.scala 27:20]
  wire  way_status_out_63 = _T_4215[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_600 = {{5'd0}, way_status_out_63}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4727 = _T_4726 & _GEN_600; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4720 = ifu_ic_rw_int_addr_ff == 6'h3e; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4722 = _T_4720 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4211; // @[Reg.scala 27:20]
  wire  way_status_out_62 = _T_4211[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_601 = {{5'd0}, way_status_out_62}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4723 = _T_4722 & _GEN_601; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4716 = ifu_ic_rw_int_addr_ff == 6'h3d; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4718 = _T_4716 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4207; // @[Reg.scala 27:20]
  wire  way_status_out_61 = _T_4207[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_602 = {{5'd0}, way_status_out_61}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4719 = _T_4718 & _GEN_602; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4712 = ifu_ic_rw_int_addr_ff == 6'h3c; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4714 = _T_4712 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4203; // @[Reg.scala 27:20]
  wire  way_status_out_60 = _T_4203[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_603 = {{5'd0}, way_status_out_60}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4715 = _T_4714 & _GEN_603; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4708 = ifu_ic_rw_int_addr_ff == 6'h3b; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4710 = _T_4708 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4199; // @[Reg.scala 27:20]
  wire  way_status_out_59 = _T_4199[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_604 = {{5'd0}, way_status_out_59}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4711 = _T_4710 & _GEN_604; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4704 = ifu_ic_rw_int_addr_ff == 6'h3a; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4706 = _T_4704 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4195; // @[Reg.scala 27:20]
  wire  way_status_out_58 = _T_4195[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_605 = {{5'd0}, way_status_out_58}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4707 = _T_4706 & _GEN_605; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4700 = ifu_ic_rw_int_addr_ff == 6'h39; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4702 = _T_4700 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4191; // @[Reg.scala 27:20]
  wire  way_status_out_57 = _T_4191[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_606 = {{5'd0}, way_status_out_57}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4703 = _T_4702 & _GEN_606; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4696 = ifu_ic_rw_int_addr_ff == 6'h38; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4698 = _T_4696 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4187; // @[Reg.scala 27:20]
  wire  way_status_out_56 = _T_4187[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_607 = {{5'd0}, way_status_out_56}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4699 = _T_4698 & _GEN_607; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4692 = ifu_ic_rw_int_addr_ff == 6'h37; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4694 = _T_4692 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4183; // @[Reg.scala 27:20]
  wire  way_status_out_55 = _T_4183[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_608 = {{5'd0}, way_status_out_55}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4695 = _T_4694 & _GEN_608; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [437:0] _T_5055 = {_T_5046,_T_4727,_T_4723,_T_4719,_T_4715,_T_4711,_T_4707,_T_4703,_T_4699,_T_4695}; // @[Cat.scala 29:58]
  wire  _T_4688 = ifu_ic_rw_int_addr_ff == 6'h36; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4690 = _T_4688 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4179; // @[Reg.scala 27:20]
  wire  way_status_out_54 = _T_4179[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_609 = {{5'd0}, way_status_out_54}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4691 = _T_4690 & _GEN_609; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4684 = ifu_ic_rw_int_addr_ff == 6'h35; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4686 = _T_4684 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4175; // @[Reg.scala 27:20]
  wire  way_status_out_53 = _T_4175[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_610 = {{5'd0}, way_status_out_53}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4687 = _T_4686 & _GEN_610; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4680 = ifu_ic_rw_int_addr_ff == 6'h34; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4682 = _T_4680 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4171; // @[Reg.scala 27:20]
  wire  way_status_out_52 = _T_4171[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_611 = {{5'd0}, way_status_out_52}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4683 = _T_4682 & _GEN_611; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4676 = ifu_ic_rw_int_addr_ff == 6'h33; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4678 = _T_4676 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4167; // @[Reg.scala 27:20]
  wire  way_status_out_51 = _T_4167[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_612 = {{5'd0}, way_status_out_51}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4679 = _T_4678 & _GEN_612; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4672 = ifu_ic_rw_int_addr_ff == 6'h32; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4674 = _T_4672 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4163; // @[Reg.scala 27:20]
  wire  way_status_out_50 = _T_4163[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_613 = {{5'd0}, way_status_out_50}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4675 = _T_4674 & _GEN_613; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4668 = ifu_ic_rw_int_addr_ff == 6'h31; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4670 = _T_4668 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4159; // @[Reg.scala 27:20]
  wire  way_status_out_49 = _T_4159[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_614 = {{5'd0}, way_status_out_49}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4671 = _T_4670 & _GEN_614; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4664 = ifu_ic_rw_int_addr_ff == 6'h30; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4666 = _T_4664 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4155; // @[Reg.scala 27:20]
  wire  way_status_out_48 = _T_4155[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_615 = {{5'd0}, way_status_out_48}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4667 = _T_4666 & _GEN_615; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4660 = ifu_ic_rw_int_addr_ff == 6'h2f; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4662 = _T_4660 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4151; // @[Reg.scala 27:20]
  wire  way_status_out_47 = _T_4151[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_616 = {{5'd0}, way_status_out_47}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4663 = _T_4662 & _GEN_616; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4656 = ifu_ic_rw_int_addr_ff == 6'h2e; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4658 = _T_4656 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4147; // @[Reg.scala 27:20]
  wire  way_status_out_46 = _T_4147[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_617 = {{5'd0}, way_status_out_46}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4659 = _T_4658 & _GEN_617; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [491:0] _T_5064 = {_T_5055,_T_4691,_T_4687,_T_4683,_T_4679,_T_4675,_T_4671,_T_4667,_T_4663,_T_4659}; // @[Cat.scala 29:58]
  wire  _T_4652 = ifu_ic_rw_int_addr_ff == 6'h2d; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4654 = _T_4652 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4143; // @[Reg.scala 27:20]
  wire  way_status_out_45 = _T_4143[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_618 = {{5'd0}, way_status_out_45}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4655 = _T_4654 & _GEN_618; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4648 = ifu_ic_rw_int_addr_ff == 6'h2c; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4650 = _T_4648 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4139; // @[Reg.scala 27:20]
  wire  way_status_out_44 = _T_4139[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_619 = {{5'd0}, way_status_out_44}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4651 = _T_4650 & _GEN_619; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4644 = ifu_ic_rw_int_addr_ff == 6'h2b; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4646 = _T_4644 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4135; // @[Reg.scala 27:20]
  wire  way_status_out_43 = _T_4135[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_620 = {{5'd0}, way_status_out_43}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4647 = _T_4646 & _GEN_620; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4640 = ifu_ic_rw_int_addr_ff == 6'h2a; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4642 = _T_4640 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4131; // @[Reg.scala 27:20]
  wire  way_status_out_42 = _T_4131[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_621 = {{5'd0}, way_status_out_42}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4643 = _T_4642 & _GEN_621; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4636 = ifu_ic_rw_int_addr_ff == 6'h29; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4638 = _T_4636 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4127; // @[Reg.scala 27:20]
  wire  way_status_out_41 = _T_4127[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_622 = {{5'd0}, way_status_out_41}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4639 = _T_4638 & _GEN_622; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4632 = ifu_ic_rw_int_addr_ff == 6'h28; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4634 = _T_4632 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4123; // @[Reg.scala 27:20]
  wire  way_status_out_40 = _T_4123[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_623 = {{5'd0}, way_status_out_40}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4635 = _T_4634 & _GEN_623; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4628 = ifu_ic_rw_int_addr_ff == 6'h27; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4630 = _T_4628 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4119; // @[Reg.scala 27:20]
  wire  way_status_out_39 = _T_4119[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_624 = {{5'd0}, way_status_out_39}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4631 = _T_4630 & _GEN_624; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4624 = ifu_ic_rw_int_addr_ff == 6'h26; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4626 = _T_4624 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4115; // @[Reg.scala 27:20]
  wire  way_status_out_38 = _T_4115[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_625 = {{5'd0}, way_status_out_38}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4627 = _T_4626 & _GEN_625; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4620 = ifu_ic_rw_int_addr_ff == 6'h25; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4622 = _T_4620 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4111; // @[Reg.scala 27:20]
  wire  way_status_out_37 = _T_4111[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_626 = {{5'd0}, way_status_out_37}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4623 = _T_4622 & _GEN_626; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [545:0] _T_5073 = {_T_5064,_T_4655,_T_4651,_T_4647,_T_4643,_T_4639,_T_4635,_T_4631,_T_4627,_T_4623}; // @[Cat.scala 29:58]
  wire  _T_4616 = ifu_ic_rw_int_addr_ff == 6'h24; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4618 = _T_4616 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4107; // @[Reg.scala 27:20]
  wire  way_status_out_36 = _T_4107[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_627 = {{5'd0}, way_status_out_36}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4619 = _T_4618 & _GEN_627; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4612 = ifu_ic_rw_int_addr_ff == 6'h23; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4614 = _T_4612 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4103; // @[Reg.scala 27:20]
  wire  way_status_out_35 = _T_4103[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_628 = {{5'd0}, way_status_out_35}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4615 = _T_4614 & _GEN_628; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4608 = ifu_ic_rw_int_addr_ff == 6'h22; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4610 = _T_4608 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4099; // @[Reg.scala 27:20]
  wire  way_status_out_34 = _T_4099[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_629 = {{5'd0}, way_status_out_34}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4611 = _T_4610 & _GEN_629; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4604 = ifu_ic_rw_int_addr_ff == 6'h21; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4606 = _T_4604 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4095; // @[Reg.scala 27:20]
  wire  way_status_out_33 = _T_4095[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_630 = {{5'd0}, way_status_out_33}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4607 = _T_4606 & _GEN_630; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4600 = ifu_ic_rw_int_addr_ff == 6'h20; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4602 = _T_4600 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4091; // @[Reg.scala 27:20]
  wire  way_status_out_32 = _T_4091[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_631 = {{5'd0}, way_status_out_32}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4603 = _T_4602 & _GEN_631; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4596 = ifu_ic_rw_int_addr_ff == 6'h1f; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4598 = _T_4596 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4087; // @[Reg.scala 27:20]
  wire  way_status_out_31 = _T_4087[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_632 = {{5'd0}, way_status_out_31}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4599 = _T_4598 & _GEN_632; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4592 = ifu_ic_rw_int_addr_ff == 6'h1e; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4594 = _T_4592 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4083; // @[Reg.scala 27:20]
  wire  way_status_out_30 = _T_4083[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_633 = {{5'd0}, way_status_out_30}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4595 = _T_4594 & _GEN_633; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4588 = ifu_ic_rw_int_addr_ff == 6'h1d; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4590 = _T_4588 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4079; // @[Reg.scala 27:20]
  wire  way_status_out_29 = _T_4079[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_634 = {{5'd0}, way_status_out_29}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4591 = _T_4590 & _GEN_634; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4584 = ifu_ic_rw_int_addr_ff == 6'h1c; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4586 = _T_4584 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4075; // @[Reg.scala 27:20]
  wire  way_status_out_28 = _T_4075[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_635 = {{5'd0}, way_status_out_28}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4587 = _T_4586 & _GEN_635; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [599:0] _T_5082 = {_T_5073,_T_4619,_T_4615,_T_4611,_T_4607,_T_4603,_T_4599,_T_4595,_T_4591,_T_4587}; // @[Cat.scala 29:58]
  wire  _T_4580 = ifu_ic_rw_int_addr_ff == 6'h1b; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4582 = _T_4580 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4071; // @[Reg.scala 27:20]
  wire  way_status_out_27 = _T_4071[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_636 = {{5'd0}, way_status_out_27}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4583 = _T_4582 & _GEN_636; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4576 = ifu_ic_rw_int_addr_ff == 6'h1a; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4578 = _T_4576 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4067; // @[Reg.scala 27:20]
  wire  way_status_out_26 = _T_4067[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_637 = {{5'd0}, way_status_out_26}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4579 = _T_4578 & _GEN_637; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4572 = ifu_ic_rw_int_addr_ff == 6'h19; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4574 = _T_4572 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4063; // @[Reg.scala 27:20]
  wire  way_status_out_25 = _T_4063[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_638 = {{5'd0}, way_status_out_25}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4575 = _T_4574 & _GEN_638; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4568 = ifu_ic_rw_int_addr_ff == 6'h18; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4570 = _T_4568 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4059; // @[Reg.scala 27:20]
  wire  way_status_out_24 = _T_4059[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_639 = {{5'd0}, way_status_out_24}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4571 = _T_4570 & _GEN_639; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4564 = ifu_ic_rw_int_addr_ff == 6'h17; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4566 = _T_4564 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4055; // @[Reg.scala 27:20]
  wire  way_status_out_23 = _T_4055[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_640 = {{5'd0}, way_status_out_23}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4567 = _T_4566 & _GEN_640; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4560 = ifu_ic_rw_int_addr_ff == 6'h16; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4562 = _T_4560 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4051; // @[Reg.scala 27:20]
  wire  way_status_out_22 = _T_4051[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_641 = {{5'd0}, way_status_out_22}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4563 = _T_4562 & _GEN_641; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4556 = ifu_ic_rw_int_addr_ff == 6'h15; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4558 = _T_4556 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4047; // @[Reg.scala 27:20]
  wire  way_status_out_21 = _T_4047[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_642 = {{5'd0}, way_status_out_21}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4559 = _T_4558 & _GEN_642; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4552 = ifu_ic_rw_int_addr_ff == 6'h14; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4554 = _T_4552 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4043; // @[Reg.scala 27:20]
  wire  way_status_out_20 = _T_4043[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_643 = {{5'd0}, way_status_out_20}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4555 = _T_4554 & _GEN_643; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4548 = ifu_ic_rw_int_addr_ff == 6'h13; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4550 = _T_4548 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4039; // @[Reg.scala 27:20]
  wire  way_status_out_19 = _T_4039[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_644 = {{5'd0}, way_status_out_19}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4551 = _T_4550 & _GEN_644; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [653:0] _T_5091 = {_T_5082,_T_4583,_T_4579,_T_4575,_T_4571,_T_4567,_T_4563,_T_4559,_T_4555,_T_4551}; // @[Cat.scala 29:58]
  wire  _T_4544 = ifu_ic_rw_int_addr_ff == 6'h12; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4546 = _T_4544 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4035; // @[Reg.scala 27:20]
  wire  way_status_out_18 = _T_4035[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_645 = {{5'd0}, way_status_out_18}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4547 = _T_4546 & _GEN_645; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4540 = ifu_ic_rw_int_addr_ff == 6'h11; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4542 = _T_4540 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4031; // @[Reg.scala 27:20]
  wire  way_status_out_17 = _T_4031[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_646 = {{5'd0}, way_status_out_17}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4543 = _T_4542 & _GEN_646; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4536 = ifu_ic_rw_int_addr_ff == 6'h10; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4538 = _T_4536 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4027; // @[Reg.scala 27:20]
  wire  way_status_out_16 = _T_4027[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_647 = {{5'd0}, way_status_out_16}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4539 = _T_4538 & _GEN_647; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4532 = ifu_ic_rw_int_addr_ff == 6'hf; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4534 = _T_4532 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4023; // @[Reg.scala 27:20]
  wire  way_status_out_15 = _T_4023[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_648 = {{5'd0}, way_status_out_15}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4535 = _T_4534 & _GEN_648; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4528 = ifu_ic_rw_int_addr_ff == 6'he; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4530 = _T_4528 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4019; // @[Reg.scala 27:20]
  wire  way_status_out_14 = _T_4019[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_649 = {{5'd0}, way_status_out_14}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4531 = _T_4530 & _GEN_649; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4524 = ifu_ic_rw_int_addr_ff == 6'hd; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4526 = _T_4524 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4015; // @[Reg.scala 27:20]
  wire  way_status_out_13 = _T_4015[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_650 = {{5'd0}, way_status_out_13}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4527 = _T_4526 & _GEN_650; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4520 = ifu_ic_rw_int_addr_ff == 6'hc; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4522 = _T_4520 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4011; // @[Reg.scala 27:20]
  wire  way_status_out_12 = _T_4011[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_651 = {{5'd0}, way_status_out_12}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4523 = _T_4522 & _GEN_651; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4516 = ifu_ic_rw_int_addr_ff == 6'hb; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4518 = _T_4516 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4007; // @[Reg.scala 27:20]
  wire  way_status_out_11 = _T_4007[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_652 = {{5'd0}, way_status_out_11}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4519 = _T_4518 & _GEN_652; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4512 = ifu_ic_rw_int_addr_ff == 6'ha; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4514 = _T_4512 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4003; // @[Reg.scala 27:20]
  wire  way_status_out_10 = _T_4003[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_653 = {{5'd0}, way_status_out_10}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4515 = _T_4514 & _GEN_653; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [707:0] _T_5100 = {_T_5091,_T_4547,_T_4543,_T_4539,_T_4535,_T_4531,_T_4527,_T_4523,_T_4519,_T_4515}; // @[Cat.scala 29:58]
  wire  _T_4508 = ifu_ic_rw_int_addr_ff == 6'h9; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4510 = _T_4508 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3999; // @[Reg.scala 27:20]
  wire  way_status_out_9 = _T_3999[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_654 = {{5'd0}, way_status_out_9}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4511 = _T_4510 & _GEN_654; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4504 = ifu_ic_rw_int_addr_ff == 6'h8; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4506 = _T_4504 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3995; // @[Reg.scala 27:20]
  wire  way_status_out_8 = _T_3995[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_655 = {{5'd0}, way_status_out_8}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4507 = _T_4506 & _GEN_655; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4500 = ifu_ic_rw_int_addr_ff == 6'h7; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4502 = _T_4500 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3991; // @[Reg.scala 27:20]
  wire  way_status_out_7 = _T_3991[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_656 = {{5'd0}, way_status_out_7}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4503 = _T_4502 & _GEN_656; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4496 = ifu_ic_rw_int_addr_ff == 6'h6; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4498 = _T_4496 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3987; // @[Reg.scala 27:20]
  wire  way_status_out_6 = _T_3987[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_657 = {{5'd0}, way_status_out_6}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4499 = _T_4498 & _GEN_657; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4492 = ifu_ic_rw_int_addr_ff == 6'h5; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4494 = _T_4492 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3983; // @[Reg.scala 27:20]
  wire  way_status_out_5 = _T_3983[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_658 = {{5'd0}, way_status_out_5}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4495 = _T_4494 & _GEN_658; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4488 = ifu_ic_rw_int_addr_ff == 6'h4; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4490 = _T_4488 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3979; // @[Reg.scala 27:20]
  wire  way_status_out_4 = _T_3979[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_659 = {{5'd0}, way_status_out_4}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4491 = _T_4490 & _GEN_659; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4484 = ifu_ic_rw_int_addr_ff == 6'h3; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4486 = _T_4484 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3975; // @[Reg.scala 27:20]
  wire  way_status_out_3 = _T_3975[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_660 = {{5'd0}, way_status_out_3}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4487 = _T_4486 & _GEN_660; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4480 = ifu_ic_rw_int_addr_ff == 6'h2; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4482 = _T_4480 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3971; // @[Reg.scala 27:20]
  wire  way_status_out_2 = _T_3971[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_661 = {{5'd0}, way_status_out_2}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4483 = _T_4482 & _GEN_661; // @[el2_ifu_mem_ctl.scala 716:130]
  wire  _T_4476 = ifu_ic_rw_int_addr_ff == 6'h1; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4478 = _T_4476 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3967; // @[Reg.scala 27:20]
  wire  way_status_out_1 = _T_3967[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_662 = {{5'd0}, way_status_out_1}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4479 = _T_4478 & _GEN_662; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [761:0] _T_5109 = {_T_5100,_T_4511,_T_4507,_T_4503,_T_4499,_T_4495,_T_4491,_T_4487,_T_4483,_T_4479}; // @[Cat.scala 29:58]
  wire  _T_4472 = ifu_ic_rw_int_addr_ff == 6'h0; // @[el2_ifu_mem_ctl.scala 716:121]
  wire [5:0] _T_4474 = _T_4472 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3963; // @[Reg.scala 27:20]
  wire  way_status_out_0 = _T_3963[0]; // @[el2_ifu_mem_ctl.scala 713:30 el2_ifu_mem_ctl.scala 715:33]
  wire [5:0] _GEN_663 = {{5'd0}, way_status_out_0}; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [5:0] _T_4475 = _T_4474 & _GEN_663; // @[el2_ifu_mem_ctl.scala 716:130]
  wire [767:0] _T_5110 = {_T_5109,_T_4475}; // @[Cat.scala 29:58]
  wire  way_status = _T_5110[0]; // @[el2_ifu_mem_ctl.scala 716:16]
  wire  _T_196 = ~reset_all_tags; // @[el2_ifu_mem_ctl.scala 257:96]
  reg  uncacheable_miss_scnd_ff; // @[el2_ifu_mem_ctl.scala 259:38]
  reg [30:0] imb_scnd_ff; // @[el2_ifu_mem_ctl.scala 261:25]
  wire [2:0] _T_207 = bus_ifu_wr_en_ff ? 3'h7 : 3'h0; // @[Bitwise.scala 72:12]
  reg [2:0] ifu_bus_rid_ff; // @[Reg.scala 27:20]
  wire [2:0] ic_wr_addr_bits_hi_3 = ifu_bus_rid_ff & _T_207; // @[el2_ifu_mem_ctl.scala 266:45]
  wire  _T_213 = _T_232 | _T_240; // @[el2_ifu_mem_ctl.scala 271:59]
  wire  _T_215 = _T_213 | _T_2222; // @[el2_ifu_mem_ctl.scala 271:91]
  wire  ic_iccm_hit_f = fetch_req_iccm_f & _T_215; // @[el2_ifu_mem_ctl.scala 271:41]
  wire  _T_220 = _T_228 & fetch_req_icache_f; // @[el2_ifu_mem_ctl.scala 277:39]
  wire  _T_222 = _T_220 & _T_196; // @[el2_ifu_mem_ctl.scala 277:60]
  wire  _T_226 = _T_222 & _T_213; // @[el2_ifu_mem_ctl.scala 277:78]
  wire  ic_act_hit_f = _T_226 & _T_248; // @[el2_ifu_mem_ctl.scala 277:126]
  wire  _T_263 = ic_act_hit_f | ic_byp_hit_f; // @[el2_ifu_mem_ctl.scala 284:31]
  wire  _T_264 = _T_263 | ic_iccm_hit_f; // @[el2_ifu_mem_ctl.scala 284:46]
  wire  _T_265 = ifc_region_acc_fault_final_f & ifc_fetch_req_f; // @[el2_ifu_mem_ctl.scala 284:94]
  wire  _T_269 = sel_hold_imb ? uncacheable_miss_ff : io_ifc_fetch_uncacheable_bf; // @[el2_ifu_mem_ctl.scala 285:84]
  wire  uncacheable_miss_in = scnd_miss_req ? uncacheable_miss_scnd_ff : _T_269; // @[el2_ifu_mem_ctl.scala 285:32]
  wire  _T_275 = imb_ff[12:6] == imb_scnd_ff[12:6]; // @[el2_ifu_mem_ctl.scala 288:75]
  wire  _T_276 = _T_275 & scnd_miss_req; // @[el2_ifu_mem_ctl.scala 288:127]
  reg [1:0] ifu_bus_rresp_ff; // @[Reg.scala 27:20]
  wire  _T_2611 = |ifu_bus_rresp_ff; // @[el2_ifu_mem_ctl.scala 614:48]
  wire  _T_2612 = _T_2611 & ifu_bus_rvalid_ff; // @[el2_ifu_mem_ctl.scala 614:52]
  wire  bus_ifu_wr_data_error_ff = _T_2612 & miss_pending; // @[el2_ifu_mem_ctl.scala 614:73]
  reg  ifu_wr_data_comb_err_ff; // @[el2_ifu_mem_ctl.scala 360:61]
  wire  ifu_wr_cumulative_err_data = bus_ifu_wr_data_error_ff | ifu_wr_data_comb_err_ff; // @[el2_ifu_mem_ctl.scala 359:55]
  wire  _T_277 = ~ifu_wr_cumulative_err_data; // @[el2_ifu_mem_ctl.scala 288:145]
  wire  scnd_miss_index_match = _T_276 & _T_277; // @[el2_ifu_mem_ctl.scala 288:143]
  wire  _T_278 = ~scnd_miss_index_match; // @[el2_ifu_mem_ctl.scala 291:47]
  wire  _T_279 = scnd_miss_req & _T_278; // @[el2_ifu_mem_ctl.scala 291:45]
  wire  _T_281 = scnd_miss_req & scnd_miss_index_match; // @[el2_ifu_mem_ctl.scala 292:26]
  reg  way_status_mb_ff; // @[el2_ifu_mem_ctl.scala 311:30]
  wire  _T_10060 = ~way_status_mb_ff; // @[el2_ifu_mem_ctl.scala 769:33]
  reg [1:0] tagv_mb_ff; // @[el2_ifu_mem_ctl.scala 312:24]
  wire  _T_10062 = _T_10060 & tagv_mb_ff[0]; // @[el2_ifu_mem_ctl.scala 769:51]
  wire  _T_10064 = _T_10062 & tagv_mb_ff[1]; // @[el2_ifu_mem_ctl.scala 769:67]
  wire  _T_10066 = ~tagv_mb_ff[0]; // @[el2_ifu_mem_ctl.scala 769:86]
  wire  replace_way_mb_any_0 = _T_10064 | _T_10066; // @[el2_ifu_mem_ctl.scala 769:84]
  wire [1:0] _T_288 = scnd_miss_index_match ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire  _T_10069 = way_status_mb_ff & tagv_mb_ff[0]; // @[el2_ifu_mem_ctl.scala 770:50]
  wire  _T_10071 = _T_10069 & tagv_mb_ff[1]; // @[el2_ifu_mem_ctl.scala 770:66]
  wire  _T_10073 = ~tagv_mb_ff[1]; // @[el2_ifu_mem_ctl.scala 770:85]
  wire  _T_10075 = _T_10073 & tagv_mb_ff[0]; // @[el2_ifu_mem_ctl.scala 770:100]
  wire  replace_way_mb_any_1 = _T_10071 | _T_10075; // @[el2_ifu_mem_ctl.scala 770:83]
  wire [1:0] _T_289 = {replace_way_mb_any_1,replace_way_mb_any_0}; // @[Cat.scala 29:58]
  wire [1:0] _T_290 = _T_288 & _T_289; // @[el2_ifu_mem_ctl.scala 296:110]
  wire  _T_298 = ~scnd_miss_req_q; // @[el2_ifu_mem_ctl.scala 300:36]
  wire  _T_299 = miss_pending & _T_298; // @[el2_ifu_mem_ctl.scala 300:34]
  reg  reset_ic_ff; // @[el2_ifu_mem_ctl.scala 301:25]
  wire  _T_300 = reset_all_tags | reset_ic_ff; // @[el2_ifu_mem_ctl.scala 300:72]
  wire  reset_ic_in = _T_299 & _T_300; // @[el2_ifu_mem_ctl.scala 300:53]
  reg  fetch_uncacheable_ff; // @[el2_ifu_mem_ctl.scala 302:37]
  reg [25:0] miss_addr; // @[el2_ifu_mem_ctl.scala 310:23]
  wire  _T_314 = _T_2237 & flush_final_f; // @[el2_ifu_mem_ctl.scala 314:87]
  wire  _T_315 = ~_T_314; // @[el2_ifu_mem_ctl.scala 314:55]
  wire  _T_316 = io_ifc_fetch_req_bf & _T_315; // @[el2_ifu_mem_ctl.scala 314:53]
  wire  _T_2229 = ~_T_2224; // @[el2_ifu_mem_ctl.scala 451:46]
  wire  _T_2230 = _T_2222 & _T_2229; // @[el2_ifu_mem_ctl.scala 451:44]
  wire  stream_miss_f = _T_2230 & ifc_fetch_req_f; // @[el2_ifu_mem_ctl.scala 451:84]
  wire  _T_317 = ~stream_miss_f; // @[el2_ifu_mem_ctl.scala 314:106]
  wire  ifc_fetch_req_qual_bf = _T_316 & _T_317; // @[el2_ifu_mem_ctl.scala 314:104]
  reg  ifc_region_acc_fault_f; // @[el2_ifu_mem_ctl.scala 320:39]
  reg [2:0] bus_rd_addr_count; // @[Reg.scala 27:20]
  wire [28:0] ifu_ic_req_addr_f = {miss_addr,bus_rd_addr_count}; // @[Cat.scala 29:58]
  wire  _T_324 = _T_240 | _T_2222; // @[el2_ifu_mem_ctl.scala 322:55]
  wire  _T_327 = _T_324 & _T_57; // @[el2_ifu_mem_ctl.scala 322:82]
  wire  _T_2243 = ~ifu_bus_rid_ff[0]; // @[el2_ifu_mem_ctl.scala 456:55]
  wire [2:0] other_tag = {ifu_bus_rid_ff[2:1],_T_2243}; // @[Cat.scala 29:58]
  wire  _T_2244 = other_tag == 3'h0; // @[el2_ifu_mem_ctl.scala 457:81]
  wire  _T_2268 = _T_2244 & ic_miss_buff_data_valid[0]; // @[Mux.scala 27:72]
  wire  _T_2247 = other_tag == 3'h1; // @[el2_ifu_mem_ctl.scala 457:81]
  wire  _T_2269 = _T_2247 & ic_miss_buff_data_valid[1]; // @[Mux.scala 27:72]
  wire  _T_2276 = _T_2268 | _T_2269; // @[Mux.scala 27:72]
  wire  _T_2250 = other_tag == 3'h2; // @[el2_ifu_mem_ctl.scala 457:81]
  wire  _T_2270 = _T_2250 & ic_miss_buff_data_valid[2]; // @[Mux.scala 27:72]
  wire  _T_2277 = _T_2276 | _T_2270; // @[Mux.scala 27:72]
  wire  _T_2253 = other_tag == 3'h3; // @[el2_ifu_mem_ctl.scala 457:81]
  wire  _T_2271 = _T_2253 & ic_miss_buff_data_valid[3]; // @[Mux.scala 27:72]
  wire  _T_2278 = _T_2277 | _T_2271; // @[Mux.scala 27:72]
  wire  _T_2256 = other_tag == 3'h4; // @[el2_ifu_mem_ctl.scala 457:81]
  wire  _T_2272 = _T_2256 & ic_miss_buff_data_valid[4]; // @[Mux.scala 27:72]
  wire  _T_2279 = _T_2278 | _T_2272; // @[Mux.scala 27:72]
  wire  _T_2259 = other_tag == 3'h5; // @[el2_ifu_mem_ctl.scala 457:81]
  wire  _T_2273 = _T_2259 & ic_miss_buff_data_valid[5]; // @[Mux.scala 27:72]
  wire  _T_2280 = _T_2279 | _T_2273; // @[Mux.scala 27:72]
  wire  _T_2262 = other_tag == 3'h6; // @[el2_ifu_mem_ctl.scala 457:81]
  wire  _T_2274 = _T_2262 & ic_miss_buff_data_valid[6]; // @[Mux.scala 27:72]
  wire  _T_2281 = _T_2280 | _T_2274; // @[Mux.scala 27:72]
  wire  _T_2265 = other_tag == 3'h7; // @[el2_ifu_mem_ctl.scala 457:81]
  wire  _T_2275 = _T_2265 & ic_miss_buff_data_valid[7]; // @[Mux.scala 27:72]
  wire  second_half_available = _T_2281 | _T_2275; // @[Mux.scala 27:72]
  wire  write_ic_16_bytes = second_half_available & bus_ifu_wr_en_ff; // @[el2_ifu_mem_ctl.scala 458:46]
  wire  _T_331 = miss_pending & write_ic_16_bytes; // @[el2_ifu_mem_ctl.scala 326:35]
  wire  _T_333 = _T_331 & _T_51; // @[el2_ifu_mem_ctl.scala 326:55]
  reg  ic_act_miss_f_delayed; // @[el2_ifu_mem_ctl.scala 611:61]
  wire  _T_2605 = ic_act_miss_f_delayed & _T_2238; // @[el2_ifu_mem_ctl.scala 612:53]
  wire  reset_tag_valid_for_miss = _T_2605 & _T_51; // @[el2_ifu_mem_ctl.scala 612:84]
  wire  sel_mb_addr = _T_333 | reset_tag_valid_for_miss; // @[el2_ifu_mem_ctl.scala 326:79]
  wire [30:0] _T_338 = {imb_ff[30:5],ic_wr_addr_bits_hi_3,imb_ff[1:0]}; // @[Cat.scala 29:58]
  wire  _T_340 = ~sel_mb_addr; // @[el2_ifu_mem_ctl.scala 328:37]
  wire [30:0] _T_341 = sel_mb_addr ? _T_338 : 31'h0; // @[Mux.scala 27:72]
  wire [30:0] _T_342 = _T_340 ? ifu_fetch_addr_int_f : 31'h0; // @[Mux.scala 27:72]
  wire [30:0] ifu_ic_rw_int_addr = _T_341 | _T_342; // @[Mux.scala 27:72]
  wire  _T_347 = _T_333 & last_beat; // @[el2_ifu_mem_ctl.scala 330:84]
  wire  _T_2599 = ~_T_2611; // @[el2_ifu_mem_ctl.scala 609:84]
  wire  _T_2600 = _T_101 & _T_2599; // @[el2_ifu_mem_ctl.scala 609:82]
  wire  bus_ifu_wr_en_ff_q = _T_2600 & write_ic_16_bytes; // @[el2_ifu_mem_ctl.scala 609:108]
  wire  sel_mb_status_addr = _T_347 & bus_ifu_wr_en_ff_q; // @[el2_ifu_mem_ctl.scala 330:96]
  wire [30:0] ifu_status_wr_addr = sel_mb_status_addr ? _T_338 : ifu_fetch_addr_int_f; // @[el2_ifu_mem_ctl.scala 331:31]
  reg [63:0] ifu_bus_rdata_ff; // @[Reg.scala 27:20]
  wire [7:0] _T_571 = {ifu_bus_rdata_ff[11],ifu_bus_rdata_ff[10],ifu_bus_rdata_ff[8],ifu_bus_rdata_ff[6],ifu_bus_rdata_ff[4],ifu_bus_rdata_ff[3],ifu_bus_rdata_ff[1],ifu_bus_rdata_ff[0]}; // @[el2_lib.scala 348:27]
  wire [16:0] _T_580 = {ifu_bus_rdata_ff[28],ifu_bus_rdata_ff[26],ifu_bus_rdata_ff[25],ifu_bus_rdata_ff[23],ifu_bus_rdata_ff[21],ifu_bus_rdata_ff[19],ifu_bus_rdata_ff[17],ifu_bus_rdata_ff[15],ifu_bus_rdata_ff[13],_T_571}; // @[el2_lib.scala 348:27]
  wire [8:0] _T_588 = {ifu_bus_rdata_ff[46],ifu_bus_rdata_ff[44],ifu_bus_rdata_ff[42],ifu_bus_rdata_ff[40],ifu_bus_rdata_ff[38],ifu_bus_rdata_ff[36],ifu_bus_rdata_ff[34],ifu_bus_rdata_ff[32],ifu_bus_rdata_ff[30]}; // @[el2_lib.scala 348:27]
  wire [17:0] _T_597 = {ifu_bus_rdata_ff[63],ifu_bus_rdata_ff[61],ifu_bus_rdata_ff[59],ifu_bus_rdata_ff[57],ifu_bus_rdata_ff[56],ifu_bus_rdata_ff[54],ifu_bus_rdata_ff[52],ifu_bus_rdata_ff[50],ifu_bus_rdata_ff[48],_T_588}; // @[el2_lib.scala 348:27]
  wire [34:0] _T_598 = {_T_597,_T_580}; // @[el2_lib.scala 348:27]
  wire  _T_599 = ^_T_598; // @[el2_lib.scala 348:34]
  wire [7:0] _T_606 = {ifu_bus_rdata_ff[12],ifu_bus_rdata_ff[10],ifu_bus_rdata_ff[9],ifu_bus_rdata_ff[6],ifu_bus_rdata_ff[5],ifu_bus_rdata_ff[3],ifu_bus_rdata_ff[2],ifu_bus_rdata_ff[0]}; // @[el2_lib.scala 348:44]
  wire [16:0] _T_615 = {ifu_bus_rdata_ff[28],ifu_bus_rdata_ff[27],ifu_bus_rdata_ff[25],ifu_bus_rdata_ff[24],ifu_bus_rdata_ff[21],ifu_bus_rdata_ff[20],ifu_bus_rdata_ff[17],ifu_bus_rdata_ff[16],ifu_bus_rdata_ff[13],_T_606}; // @[el2_lib.scala 348:44]
  wire [8:0] _T_623 = {ifu_bus_rdata_ff[47],ifu_bus_rdata_ff[44],ifu_bus_rdata_ff[43],ifu_bus_rdata_ff[40],ifu_bus_rdata_ff[39],ifu_bus_rdata_ff[36],ifu_bus_rdata_ff[35],ifu_bus_rdata_ff[32],ifu_bus_rdata_ff[31]}; // @[el2_lib.scala 348:44]
  wire [17:0] _T_632 = {ifu_bus_rdata_ff[63],ifu_bus_rdata_ff[62],ifu_bus_rdata_ff[59],ifu_bus_rdata_ff[58],ifu_bus_rdata_ff[56],ifu_bus_rdata_ff[55],ifu_bus_rdata_ff[52],ifu_bus_rdata_ff[51],ifu_bus_rdata_ff[48],_T_623}; // @[el2_lib.scala 348:44]
  wire [34:0] _T_633 = {_T_632,_T_615}; // @[el2_lib.scala 348:44]
  wire  _T_634 = ^_T_633; // @[el2_lib.scala 348:51]
  wire [7:0] _T_641 = {ifu_bus_rdata_ff[14],ifu_bus_rdata_ff[10],ifu_bus_rdata_ff[9],ifu_bus_rdata_ff[8],ifu_bus_rdata_ff[7],ifu_bus_rdata_ff[3],ifu_bus_rdata_ff[2],ifu_bus_rdata_ff[1]}; // @[el2_lib.scala 348:61]
  wire [16:0] _T_650 = {ifu_bus_rdata_ff[30],ifu_bus_rdata_ff[29],ifu_bus_rdata_ff[25],ifu_bus_rdata_ff[24],ifu_bus_rdata_ff[23],ifu_bus_rdata_ff[22],ifu_bus_rdata_ff[17],ifu_bus_rdata_ff[16],ifu_bus_rdata_ff[15],_T_641}; // @[el2_lib.scala 348:61]
  wire [8:0] _T_658 = {ifu_bus_rdata_ff[47],ifu_bus_rdata_ff[46],ifu_bus_rdata_ff[45],ifu_bus_rdata_ff[40],ifu_bus_rdata_ff[39],ifu_bus_rdata_ff[38],ifu_bus_rdata_ff[37],ifu_bus_rdata_ff[32],ifu_bus_rdata_ff[31]}; // @[el2_lib.scala 348:61]
  wire [17:0] _T_667 = {ifu_bus_rdata_ff[63],ifu_bus_rdata_ff[62],ifu_bus_rdata_ff[61],ifu_bus_rdata_ff[60],ifu_bus_rdata_ff[56],ifu_bus_rdata_ff[55],ifu_bus_rdata_ff[54],ifu_bus_rdata_ff[53],ifu_bus_rdata_ff[48],_T_658}; // @[el2_lib.scala 348:61]
  wire [34:0] _T_668 = {_T_667,_T_650}; // @[el2_lib.scala 348:61]
  wire  _T_669 = ^_T_668; // @[el2_lib.scala 348:68]
  wire [6:0] _T_675 = {ifu_bus_rdata_ff[10],ifu_bus_rdata_ff[9],ifu_bus_rdata_ff[8],ifu_bus_rdata_ff[7],ifu_bus_rdata_ff[6],ifu_bus_rdata_ff[5],ifu_bus_rdata_ff[4]}; // @[el2_lib.scala 348:78]
  wire [14:0] _T_683 = {ifu_bus_rdata_ff[25],ifu_bus_rdata_ff[24],ifu_bus_rdata_ff[23],ifu_bus_rdata_ff[22],ifu_bus_rdata_ff[21],ifu_bus_rdata_ff[20],ifu_bus_rdata_ff[19],ifu_bus_rdata_ff[18],_T_675}; // @[el2_lib.scala 348:78]
  wire [7:0] _T_690 = {ifu_bus_rdata_ff[40],ifu_bus_rdata_ff[39],ifu_bus_rdata_ff[38],ifu_bus_rdata_ff[37],ifu_bus_rdata_ff[36],ifu_bus_rdata_ff[35],ifu_bus_rdata_ff[34],ifu_bus_rdata_ff[33]}; // @[el2_lib.scala 348:78]
  wire [30:0] _T_699 = {ifu_bus_rdata_ff[56],ifu_bus_rdata_ff[55],ifu_bus_rdata_ff[54],ifu_bus_rdata_ff[53],ifu_bus_rdata_ff[52],ifu_bus_rdata_ff[51],ifu_bus_rdata_ff[50],ifu_bus_rdata_ff[49],_T_690,_T_683}; // @[el2_lib.scala 348:78]
  wire  _T_700 = ^_T_699; // @[el2_lib.scala 348:85]
  wire [6:0] _T_706 = {ifu_bus_rdata_ff[17],ifu_bus_rdata_ff[16],ifu_bus_rdata_ff[15],ifu_bus_rdata_ff[14],ifu_bus_rdata_ff[13],ifu_bus_rdata_ff[12],ifu_bus_rdata_ff[11]}; // @[el2_lib.scala 348:95]
  wire [14:0] _T_714 = {ifu_bus_rdata_ff[25],ifu_bus_rdata_ff[24],ifu_bus_rdata_ff[23],ifu_bus_rdata_ff[22],ifu_bus_rdata_ff[21],ifu_bus_rdata_ff[20],ifu_bus_rdata_ff[19],ifu_bus_rdata_ff[18],_T_706}; // @[el2_lib.scala 348:95]
  wire [7:0] _T_721 = {ifu_bus_rdata_ff[48],ifu_bus_rdata_ff[47],ifu_bus_rdata_ff[46],ifu_bus_rdata_ff[45],ifu_bus_rdata_ff[44],ifu_bus_rdata_ff[43],ifu_bus_rdata_ff[42],ifu_bus_rdata_ff[41]}; // @[el2_lib.scala 348:95]
  wire [30:0] _T_730 = {ifu_bus_rdata_ff[56],ifu_bus_rdata_ff[55],ifu_bus_rdata_ff[54],ifu_bus_rdata_ff[53],ifu_bus_rdata_ff[52],ifu_bus_rdata_ff[51],ifu_bus_rdata_ff[50],ifu_bus_rdata_ff[49],_T_721,_T_714}; // @[el2_lib.scala 348:95]
  wire  _T_731 = ^_T_730; // @[el2_lib.scala 348:102]
  wire [6:0] _T_737 = {ifu_bus_rdata_ff[32],ifu_bus_rdata_ff[31],ifu_bus_rdata_ff[30],ifu_bus_rdata_ff[29],ifu_bus_rdata_ff[28],ifu_bus_rdata_ff[27],ifu_bus_rdata_ff[26]}; // @[el2_lib.scala 348:112]
  wire [14:0] _T_745 = {ifu_bus_rdata_ff[40],ifu_bus_rdata_ff[39],ifu_bus_rdata_ff[38],ifu_bus_rdata_ff[37],ifu_bus_rdata_ff[36],ifu_bus_rdata_ff[35],ifu_bus_rdata_ff[34],ifu_bus_rdata_ff[33],_T_737}; // @[el2_lib.scala 348:112]
  wire [30:0] _T_761 = {ifu_bus_rdata_ff[56],ifu_bus_rdata_ff[55],ifu_bus_rdata_ff[54],ifu_bus_rdata_ff[53],ifu_bus_rdata_ff[52],ifu_bus_rdata_ff[51],ifu_bus_rdata_ff[50],ifu_bus_rdata_ff[49],_T_721,_T_745}; // @[el2_lib.scala 348:112]
  wire  _T_762 = ^_T_761; // @[el2_lib.scala 348:119]
  wire [6:0] _T_768 = {ifu_bus_rdata_ff[63],ifu_bus_rdata_ff[62],ifu_bus_rdata_ff[61],ifu_bus_rdata_ff[60],ifu_bus_rdata_ff[59],ifu_bus_rdata_ff[58],ifu_bus_rdata_ff[57]}; // @[el2_lib.scala 348:129]
  wire  _T_769 = ^_T_768; // @[el2_lib.scala 348:136]
  wire [3:0] _T_2284 = {ifu_bus_rid_ff[2:1],_T_2243,1'h1}; // @[Cat.scala 29:58]
  wire  _T_2285 = _T_2284 == 4'h0; // @[el2_ifu_mem_ctl.scala 459:89]
  reg [63:0] _T_1296; // @[Reg.scala 27:20]
  wire [31:0] ic_miss_buff_data_0 = _T_1296[31:0]; // @[el2_ifu_mem_ctl.scala 392:31 el2_ifu_mem_ctl.scala 394:26]
  wire [31:0] _T_2332 = _T_2285 ? ic_miss_buff_data_0 : 32'h0; // @[Mux.scala 27:72]
  wire  _T_2288 = _T_2284 == 4'h1; // @[el2_ifu_mem_ctl.scala 459:89]
  reg [63:0] _T_1298; // @[Reg.scala 27:20]
  wire [31:0] ic_miss_buff_data_1 = _T_1298[31:0]; // @[el2_ifu_mem_ctl.scala 392:31 el2_ifu_mem_ctl.scala 395:28]
  wire [31:0] _T_2333 = _T_2288 ? ic_miss_buff_data_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2348 = _T_2332 | _T_2333; // @[Mux.scala 27:72]
  wire  _T_2291 = _T_2284 == 4'h2; // @[el2_ifu_mem_ctl.scala 459:89]
  reg [63:0] _T_1300; // @[Reg.scala 27:20]
  wire [31:0] ic_miss_buff_data_2 = _T_1300[31:0]; // @[el2_ifu_mem_ctl.scala 392:31 el2_ifu_mem_ctl.scala 394:26]
  wire [31:0] _T_2334 = _T_2291 ? ic_miss_buff_data_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2349 = _T_2348 | _T_2334; // @[Mux.scala 27:72]
  wire  _T_2294 = _T_2284 == 4'h3; // @[el2_ifu_mem_ctl.scala 459:89]
  reg [63:0] _T_1302; // @[Reg.scala 27:20]
  wire [31:0] ic_miss_buff_data_3 = _T_1302[31:0]; // @[el2_ifu_mem_ctl.scala 392:31 el2_ifu_mem_ctl.scala 395:28]
  wire [31:0] _T_2335 = _T_2294 ? ic_miss_buff_data_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2350 = _T_2349 | _T_2335; // @[Mux.scala 27:72]
  wire  _T_2297 = _T_2284 == 4'h4; // @[el2_ifu_mem_ctl.scala 459:89]
  reg [63:0] _T_1304; // @[Reg.scala 27:20]
  wire [31:0] ic_miss_buff_data_4 = _T_1304[31:0]; // @[el2_ifu_mem_ctl.scala 392:31 el2_ifu_mem_ctl.scala 394:26]
  wire [31:0] _T_2336 = _T_2297 ? ic_miss_buff_data_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2351 = _T_2350 | _T_2336; // @[Mux.scala 27:72]
  wire  _T_2300 = _T_2284 == 4'h5; // @[el2_ifu_mem_ctl.scala 459:89]
  reg [63:0] _T_1306; // @[Reg.scala 27:20]
  wire [31:0] ic_miss_buff_data_5 = _T_1306[31:0]; // @[el2_ifu_mem_ctl.scala 392:31 el2_ifu_mem_ctl.scala 395:28]
  wire [31:0] _T_2337 = _T_2300 ? ic_miss_buff_data_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2352 = _T_2351 | _T_2337; // @[Mux.scala 27:72]
  wire  _T_2303 = _T_2284 == 4'h6; // @[el2_ifu_mem_ctl.scala 459:89]
  reg [63:0] _T_1308; // @[Reg.scala 27:20]
  wire [31:0] ic_miss_buff_data_6 = _T_1308[31:0]; // @[el2_ifu_mem_ctl.scala 392:31 el2_ifu_mem_ctl.scala 394:26]
  wire [31:0] _T_2338 = _T_2303 ? ic_miss_buff_data_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2353 = _T_2352 | _T_2338; // @[Mux.scala 27:72]
  wire  _T_2306 = _T_2284 == 4'h7; // @[el2_ifu_mem_ctl.scala 459:89]
  reg [63:0] _T_1310; // @[Reg.scala 27:20]
  wire [31:0] ic_miss_buff_data_7 = _T_1310[31:0]; // @[el2_ifu_mem_ctl.scala 392:31 el2_ifu_mem_ctl.scala 395:28]
  wire [31:0] _T_2339 = _T_2306 ? ic_miss_buff_data_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2354 = _T_2353 | _T_2339; // @[Mux.scala 27:72]
  wire  _T_2309 = _T_2284 == 4'h8; // @[el2_ifu_mem_ctl.scala 459:89]
  reg [63:0] _T_1312; // @[Reg.scala 27:20]
  wire [31:0] ic_miss_buff_data_8 = _T_1312[31:0]; // @[el2_ifu_mem_ctl.scala 392:31 el2_ifu_mem_ctl.scala 394:26]
  wire [31:0] _T_2340 = _T_2309 ? ic_miss_buff_data_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2355 = _T_2354 | _T_2340; // @[Mux.scala 27:72]
  wire  _T_2312 = _T_2284 == 4'h9; // @[el2_ifu_mem_ctl.scala 459:89]
  reg [63:0] _T_1314; // @[Reg.scala 27:20]
  wire [31:0] ic_miss_buff_data_9 = _T_1314[31:0]; // @[el2_ifu_mem_ctl.scala 392:31 el2_ifu_mem_ctl.scala 395:28]
  wire [31:0] _T_2341 = _T_2312 ? ic_miss_buff_data_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2356 = _T_2355 | _T_2341; // @[Mux.scala 27:72]
  wire  _T_2315 = _T_2284 == 4'ha; // @[el2_ifu_mem_ctl.scala 459:89]
  reg [63:0] _T_1316; // @[Reg.scala 27:20]
  wire [31:0] ic_miss_buff_data_10 = _T_1316[31:0]; // @[el2_ifu_mem_ctl.scala 392:31 el2_ifu_mem_ctl.scala 394:26]
  wire [31:0] _T_2342 = _T_2315 ? ic_miss_buff_data_10 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2357 = _T_2356 | _T_2342; // @[Mux.scala 27:72]
  wire  _T_2318 = _T_2284 == 4'hb; // @[el2_ifu_mem_ctl.scala 459:89]
  reg [63:0] _T_1318; // @[Reg.scala 27:20]
  wire [31:0] ic_miss_buff_data_11 = _T_1318[31:0]; // @[el2_ifu_mem_ctl.scala 392:31 el2_ifu_mem_ctl.scala 395:28]
  wire [31:0] _T_2343 = _T_2318 ? ic_miss_buff_data_11 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2358 = _T_2357 | _T_2343; // @[Mux.scala 27:72]
  wire  _T_2321 = _T_2284 == 4'hc; // @[el2_ifu_mem_ctl.scala 459:89]
  reg [63:0] _T_1320; // @[Reg.scala 27:20]
  wire [31:0] ic_miss_buff_data_12 = _T_1320[31:0]; // @[el2_ifu_mem_ctl.scala 392:31 el2_ifu_mem_ctl.scala 394:26]
  wire [31:0] _T_2344 = _T_2321 ? ic_miss_buff_data_12 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2359 = _T_2358 | _T_2344; // @[Mux.scala 27:72]
  wire  _T_2324 = _T_2284 == 4'hd; // @[el2_ifu_mem_ctl.scala 459:89]
  reg [63:0] _T_1322; // @[Reg.scala 27:20]
  wire [31:0] ic_miss_buff_data_13 = _T_1322[31:0]; // @[el2_ifu_mem_ctl.scala 392:31 el2_ifu_mem_ctl.scala 395:28]
  wire [31:0] _T_2345 = _T_2324 ? ic_miss_buff_data_13 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2360 = _T_2359 | _T_2345; // @[Mux.scala 27:72]
  wire  _T_2327 = _T_2284 == 4'he; // @[el2_ifu_mem_ctl.scala 459:89]
  reg [63:0] _T_1324; // @[Reg.scala 27:20]
  wire [31:0] ic_miss_buff_data_14 = _T_1324[31:0]; // @[el2_ifu_mem_ctl.scala 392:31 el2_ifu_mem_ctl.scala 394:26]
  wire [31:0] _T_2346 = _T_2327 ? ic_miss_buff_data_14 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2361 = _T_2360 | _T_2346; // @[Mux.scala 27:72]
  wire  _T_2330 = _T_2284 == 4'hf; // @[el2_ifu_mem_ctl.scala 459:89]
  reg [63:0] _T_1326; // @[Reg.scala 27:20]
  wire [31:0] ic_miss_buff_data_15 = _T_1326[31:0]; // @[el2_ifu_mem_ctl.scala 392:31 el2_ifu_mem_ctl.scala 395:28]
  wire [31:0] _T_2347 = _T_2330 ? ic_miss_buff_data_15 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2362 = _T_2361 | _T_2347; // @[Mux.scala 27:72]
  wire [3:0] _T_2364 = {ifu_bus_rid_ff[2:1],_T_2243,1'h0}; // @[Cat.scala 29:58]
  wire  _T_2365 = _T_2364 == 4'h0; // @[el2_ifu_mem_ctl.scala 460:64]
  wire [31:0] _T_2388 = _T_2365 ? ic_miss_buff_data_0 : 32'h0; // @[Mux.scala 27:72]
  wire  _T_2368 = _T_2364 == 4'h1; // @[el2_ifu_mem_ctl.scala 460:64]
  wire [31:0] _T_2389 = _T_2368 ? ic_miss_buff_data_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2396 = _T_2388 | _T_2389; // @[Mux.scala 27:72]
  wire  _T_2371 = _T_2364 == 4'h2; // @[el2_ifu_mem_ctl.scala 460:64]
  wire [31:0] _T_2390 = _T_2371 ? ic_miss_buff_data_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2397 = _T_2396 | _T_2390; // @[Mux.scala 27:72]
  wire  _T_2374 = _T_2364 == 4'h3; // @[el2_ifu_mem_ctl.scala 460:64]
  wire [31:0] _T_2391 = _T_2374 ? ic_miss_buff_data_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2398 = _T_2397 | _T_2391; // @[Mux.scala 27:72]
  wire  _T_2377 = _T_2364 == 4'h4; // @[el2_ifu_mem_ctl.scala 460:64]
  wire [31:0] _T_2392 = _T_2377 ? ic_miss_buff_data_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2399 = _T_2398 | _T_2392; // @[Mux.scala 27:72]
  wire  _T_2380 = _T_2364 == 4'h5; // @[el2_ifu_mem_ctl.scala 460:64]
  wire [31:0] _T_2393 = _T_2380 ? ic_miss_buff_data_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2400 = _T_2399 | _T_2393; // @[Mux.scala 27:72]
  wire  _T_2383 = _T_2364 == 4'h6; // @[el2_ifu_mem_ctl.scala 460:64]
  wire [31:0] _T_2394 = _T_2383 ? ic_miss_buff_data_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2401 = _T_2400 | _T_2394; // @[Mux.scala 27:72]
  wire  _T_2386 = _T_2364 == 4'h7; // @[el2_ifu_mem_ctl.scala 460:64]
  wire [31:0] _T_2395 = _T_2386 ? ic_miss_buff_data_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2402 = _T_2401 | _T_2395; // @[Mux.scala 27:72]
  wire [63:0] ic_miss_buff_half = {_T_2362,_T_2402}; // @[Cat.scala 29:58]
  wire [7:0] _T_993 = {ic_miss_buff_half[11],ic_miss_buff_half[10],ic_miss_buff_half[8],ic_miss_buff_half[6],ic_miss_buff_half[4],ic_miss_buff_half[3],ic_miss_buff_half[1],ic_miss_buff_half[0]}; // @[el2_lib.scala 348:27]
  wire [16:0] _T_1002 = {ic_miss_buff_half[28],ic_miss_buff_half[26],ic_miss_buff_half[25],ic_miss_buff_half[23],ic_miss_buff_half[21],ic_miss_buff_half[19],ic_miss_buff_half[17],ic_miss_buff_half[15],ic_miss_buff_half[13],_T_993}; // @[el2_lib.scala 348:27]
  wire [8:0] _T_1010 = {ic_miss_buff_half[46],ic_miss_buff_half[44],ic_miss_buff_half[42],ic_miss_buff_half[40],ic_miss_buff_half[38],ic_miss_buff_half[36],ic_miss_buff_half[34],ic_miss_buff_half[32],ic_miss_buff_half[30]}; // @[el2_lib.scala 348:27]
  wire [17:0] _T_1019 = {ic_miss_buff_half[63],ic_miss_buff_half[61],ic_miss_buff_half[59],ic_miss_buff_half[57],ic_miss_buff_half[56],ic_miss_buff_half[54],ic_miss_buff_half[52],ic_miss_buff_half[50],ic_miss_buff_half[48],_T_1010}; // @[el2_lib.scala 348:27]
  wire [34:0] _T_1020 = {_T_1019,_T_1002}; // @[el2_lib.scala 348:27]
  wire  _T_1021 = ^_T_1020; // @[el2_lib.scala 348:34]
  wire [7:0] _T_1028 = {ic_miss_buff_half[12],ic_miss_buff_half[10],ic_miss_buff_half[9],ic_miss_buff_half[6],ic_miss_buff_half[5],ic_miss_buff_half[3],ic_miss_buff_half[2],ic_miss_buff_half[0]}; // @[el2_lib.scala 348:44]
  wire [16:0] _T_1037 = {ic_miss_buff_half[28],ic_miss_buff_half[27],ic_miss_buff_half[25],ic_miss_buff_half[24],ic_miss_buff_half[21],ic_miss_buff_half[20],ic_miss_buff_half[17],ic_miss_buff_half[16],ic_miss_buff_half[13],_T_1028}; // @[el2_lib.scala 348:44]
  wire [8:0] _T_1045 = {ic_miss_buff_half[47],ic_miss_buff_half[44],ic_miss_buff_half[43],ic_miss_buff_half[40],ic_miss_buff_half[39],ic_miss_buff_half[36],ic_miss_buff_half[35],ic_miss_buff_half[32],ic_miss_buff_half[31]}; // @[el2_lib.scala 348:44]
  wire [17:0] _T_1054 = {ic_miss_buff_half[63],ic_miss_buff_half[62],ic_miss_buff_half[59],ic_miss_buff_half[58],ic_miss_buff_half[56],ic_miss_buff_half[55],ic_miss_buff_half[52],ic_miss_buff_half[51],ic_miss_buff_half[48],_T_1045}; // @[el2_lib.scala 348:44]
  wire [34:0] _T_1055 = {_T_1054,_T_1037}; // @[el2_lib.scala 348:44]
  wire  _T_1056 = ^_T_1055; // @[el2_lib.scala 348:51]
  wire [7:0] _T_1063 = {ic_miss_buff_half[14],ic_miss_buff_half[10],ic_miss_buff_half[9],ic_miss_buff_half[8],ic_miss_buff_half[7],ic_miss_buff_half[3],ic_miss_buff_half[2],ic_miss_buff_half[1]}; // @[el2_lib.scala 348:61]
  wire [16:0] _T_1072 = {ic_miss_buff_half[30],ic_miss_buff_half[29],ic_miss_buff_half[25],ic_miss_buff_half[24],ic_miss_buff_half[23],ic_miss_buff_half[22],ic_miss_buff_half[17],ic_miss_buff_half[16],ic_miss_buff_half[15],_T_1063}; // @[el2_lib.scala 348:61]
  wire [8:0] _T_1080 = {ic_miss_buff_half[47],ic_miss_buff_half[46],ic_miss_buff_half[45],ic_miss_buff_half[40],ic_miss_buff_half[39],ic_miss_buff_half[38],ic_miss_buff_half[37],ic_miss_buff_half[32],ic_miss_buff_half[31]}; // @[el2_lib.scala 348:61]
  wire [17:0] _T_1089 = {ic_miss_buff_half[63],ic_miss_buff_half[62],ic_miss_buff_half[61],ic_miss_buff_half[60],ic_miss_buff_half[56],ic_miss_buff_half[55],ic_miss_buff_half[54],ic_miss_buff_half[53],ic_miss_buff_half[48],_T_1080}; // @[el2_lib.scala 348:61]
  wire [34:0] _T_1090 = {_T_1089,_T_1072}; // @[el2_lib.scala 348:61]
  wire  _T_1091 = ^_T_1090; // @[el2_lib.scala 348:68]
  wire [6:0] _T_1097 = {ic_miss_buff_half[10],ic_miss_buff_half[9],ic_miss_buff_half[8],ic_miss_buff_half[7],ic_miss_buff_half[6],ic_miss_buff_half[5],ic_miss_buff_half[4]}; // @[el2_lib.scala 348:78]
  wire [14:0] _T_1105 = {ic_miss_buff_half[25],ic_miss_buff_half[24],ic_miss_buff_half[23],ic_miss_buff_half[22],ic_miss_buff_half[21],ic_miss_buff_half[20],ic_miss_buff_half[19],ic_miss_buff_half[18],_T_1097}; // @[el2_lib.scala 348:78]
  wire [7:0] _T_1112 = {ic_miss_buff_half[40],ic_miss_buff_half[39],ic_miss_buff_half[38],ic_miss_buff_half[37],ic_miss_buff_half[36],ic_miss_buff_half[35],ic_miss_buff_half[34],ic_miss_buff_half[33]}; // @[el2_lib.scala 348:78]
  wire [30:0] _T_1121 = {ic_miss_buff_half[56],ic_miss_buff_half[55],ic_miss_buff_half[54],ic_miss_buff_half[53],ic_miss_buff_half[52],ic_miss_buff_half[51],ic_miss_buff_half[50],ic_miss_buff_half[49],_T_1112,_T_1105}; // @[el2_lib.scala 348:78]
  wire  _T_1122 = ^_T_1121; // @[el2_lib.scala 348:85]
  wire [6:0] _T_1128 = {ic_miss_buff_half[17],ic_miss_buff_half[16],ic_miss_buff_half[15],ic_miss_buff_half[14],ic_miss_buff_half[13],ic_miss_buff_half[12],ic_miss_buff_half[11]}; // @[el2_lib.scala 348:95]
  wire [14:0] _T_1136 = {ic_miss_buff_half[25],ic_miss_buff_half[24],ic_miss_buff_half[23],ic_miss_buff_half[22],ic_miss_buff_half[21],ic_miss_buff_half[20],ic_miss_buff_half[19],ic_miss_buff_half[18],_T_1128}; // @[el2_lib.scala 348:95]
  wire [7:0] _T_1143 = {ic_miss_buff_half[48],ic_miss_buff_half[47],ic_miss_buff_half[46],ic_miss_buff_half[45],ic_miss_buff_half[44],ic_miss_buff_half[43],ic_miss_buff_half[42],ic_miss_buff_half[41]}; // @[el2_lib.scala 348:95]
  wire [30:0] _T_1152 = {ic_miss_buff_half[56],ic_miss_buff_half[55],ic_miss_buff_half[54],ic_miss_buff_half[53],ic_miss_buff_half[52],ic_miss_buff_half[51],ic_miss_buff_half[50],ic_miss_buff_half[49],_T_1143,_T_1136}; // @[el2_lib.scala 348:95]
  wire  _T_1153 = ^_T_1152; // @[el2_lib.scala 348:102]
  wire [6:0] _T_1159 = {ic_miss_buff_half[32],ic_miss_buff_half[31],ic_miss_buff_half[30],ic_miss_buff_half[29],ic_miss_buff_half[28],ic_miss_buff_half[27],ic_miss_buff_half[26]}; // @[el2_lib.scala 348:112]
  wire [14:0] _T_1167 = {ic_miss_buff_half[40],ic_miss_buff_half[39],ic_miss_buff_half[38],ic_miss_buff_half[37],ic_miss_buff_half[36],ic_miss_buff_half[35],ic_miss_buff_half[34],ic_miss_buff_half[33],_T_1159}; // @[el2_lib.scala 348:112]
  wire [30:0] _T_1183 = {ic_miss_buff_half[56],ic_miss_buff_half[55],ic_miss_buff_half[54],ic_miss_buff_half[53],ic_miss_buff_half[52],ic_miss_buff_half[51],ic_miss_buff_half[50],ic_miss_buff_half[49],_T_1143,_T_1167}; // @[el2_lib.scala 348:112]
  wire  _T_1184 = ^_T_1183; // @[el2_lib.scala 348:119]
  wire [6:0] _T_1190 = {ic_miss_buff_half[63],ic_miss_buff_half[62],ic_miss_buff_half[61],ic_miss_buff_half[60],ic_miss_buff_half[59],ic_miss_buff_half[58],ic_miss_buff_half[57]}; // @[el2_lib.scala 348:129]
  wire  _T_1191 = ^_T_1190; // @[el2_lib.scala 348:136]
  wire [70:0] _T_1238 = {_T_599,_T_634,_T_669,_T_700,_T_731,_T_762,_T_769,ifu_bus_rdata_ff}; // @[Cat.scala 29:58]
  wire [70:0] _T_1237 = {_T_1021,_T_1056,_T_1091,_T_1122,_T_1153,_T_1184,_T_1191,_T_2362,_T_2402}; // @[Cat.scala 29:58]
  wire [141:0] _T_1239 = {_T_599,_T_634,_T_669,_T_700,_T_731,_T_762,_T_769,ifu_bus_rdata_ff,_T_1237}; // @[Cat.scala 29:58]
  wire [141:0] _T_1242 = {_T_1021,_T_1056,_T_1091,_T_1122,_T_1153,_T_1184,_T_1191,_T_2362,_T_2402,_T_1238}; // @[Cat.scala 29:58]
  wire [141:0] ic_wr_16bytes_data = ifu_bus_rid_ff[0] ? _T_1239 : _T_1242; // @[el2_ifu_mem_ctl.scala 352:28]
  wire  _T_1199 = |io_ic_eccerr; // @[el2_ifu_mem_ctl.scala 342:56]
  wire  _T_1200 = _T_1199 & ic_act_hit_f; // @[el2_ifu_mem_ctl.scala 342:83]
  wire [4:0] bypass_index = imb_ff[4:0]; // @[el2_ifu_mem_ctl.scala 406:28]
  wire  _T_1402 = bypass_index[4:2] == 3'h0; // @[el2_ifu_mem_ctl.scala 408:114]
  wire  bus_ifu_wr_en = _T_13 & miss_pending; // @[el2_ifu_mem_ctl.scala 607:35]
  wire  _T_1287 = io_ifu_axi_rid == 3'h0; // @[el2_ifu_mem_ctl.scala 391:91]
  wire  write_fill_data_0 = bus_ifu_wr_en & _T_1287; // @[el2_ifu_mem_ctl.scala 391:73]
  wire  _T_1328 = ~ic_act_miss_f; // @[el2_ifu_mem_ctl.scala 397:118]
  wire  _T_1329 = ic_miss_buff_data_valid[0] & _T_1328; // @[el2_ifu_mem_ctl.scala 397:116]
  wire  ic_miss_buff_data_valid_in_0 = write_fill_data_0 | _T_1329; // @[el2_ifu_mem_ctl.scala 397:88]
  wire  _T_1425 = _T_1402 & ic_miss_buff_data_valid_in_0; // @[Mux.scala 27:72]
  wire  _T_1405 = bypass_index[4:2] == 3'h1; // @[el2_ifu_mem_ctl.scala 408:114]
  wire  _T_1288 = io_ifu_axi_rid == 3'h1; // @[el2_ifu_mem_ctl.scala 391:91]
  wire  write_fill_data_1 = bus_ifu_wr_en & _T_1288; // @[el2_ifu_mem_ctl.scala 391:73]
  wire  _T_1332 = ic_miss_buff_data_valid[1] & _T_1328; // @[el2_ifu_mem_ctl.scala 397:116]
  wire  ic_miss_buff_data_valid_in_1 = write_fill_data_1 | _T_1332; // @[el2_ifu_mem_ctl.scala 397:88]
  wire  _T_1426 = _T_1405 & ic_miss_buff_data_valid_in_1; // @[Mux.scala 27:72]
  wire  _T_1433 = _T_1425 | _T_1426; // @[Mux.scala 27:72]
  wire  _T_1408 = bypass_index[4:2] == 3'h2; // @[el2_ifu_mem_ctl.scala 408:114]
  wire  _T_1289 = io_ifu_axi_rid == 3'h2; // @[el2_ifu_mem_ctl.scala 391:91]
  wire  write_fill_data_2 = bus_ifu_wr_en & _T_1289; // @[el2_ifu_mem_ctl.scala 391:73]
  wire  _T_1335 = ic_miss_buff_data_valid[2] & _T_1328; // @[el2_ifu_mem_ctl.scala 397:116]
  wire  ic_miss_buff_data_valid_in_2 = write_fill_data_2 | _T_1335; // @[el2_ifu_mem_ctl.scala 397:88]
  wire  _T_1427 = _T_1408 & ic_miss_buff_data_valid_in_2; // @[Mux.scala 27:72]
  wire  _T_1434 = _T_1433 | _T_1427; // @[Mux.scala 27:72]
  wire  _T_1411 = bypass_index[4:2] == 3'h3; // @[el2_ifu_mem_ctl.scala 408:114]
  wire  _T_1290 = io_ifu_axi_rid == 3'h3; // @[el2_ifu_mem_ctl.scala 391:91]
  wire  write_fill_data_3 = bus_ifu_wr_en & _T_1290; // @[el2_ifu_mem_ctl.scala 391:73]
  wire  _T_1338 = ic_miss_buff_data_valid[3] & _T_1328; // @[el2_ifu_mem_ctl.scala 397:116]
  wire  ic_miss_buff_data_valid_in_3 = write_fill_data_3 | _T_1338; // @[el2_ifu_mem_ctl.scala 397:88]
  wire  _T_1428 = _T_1411 & ic_miss_buff_data_valid_in_3; // @[Mux.scala 27:72]
  wire  _T_1435 = _T_1434 | _T_1428; // @[Mux.scala 27:72]
  wire  _T_1414 = bypass_index[4:2] == 3'h4; // @[el2_ifu_mem_ctl.scala 408:114]
  wire  _T_1291 = io_ifu_axi_rid == 3'h4; // @[el2_ifu_mem_ctl.scala 391:91]
  wire  write_fill_data_4 = bus_ifu_wr_en & _T_1291; // @[el2_ifu_mem_ctl.scala 391:73]
  wire  _T_1341 = ic_miss_buff_data_valid[4] & _T_1328; // @[el2_ifu_mem_ctl.scala 397:116]
  wire  ic_miss_buff_data_valid_in_4 = write_fill_data_4 | _T_1341; // @[el2_ifu_mem_ctl.scala 397:88]
  wire  _T_1429 = _T_1414 & ic_miss_buff_data_valid_in_4; // @[Mux.scala 27:72]
  wire  _T_1436 = _T_1435 | _T_1429; // @[Mux.scala 27:72]
  wire  _T_1417 = bypass_index[4:2] == 3'h5; // @[el2_ifu_mem_ctl.scala 408:114]
  wire  _T_1292 = io_ifu_axi_rid == 3'h5; // @[el2_ifu_mem_ctl.scala 391:91]
  wire  write_fill_data_5 = bus_ifu_wr_en & _T_1292; // @[el2_ifu_mem_ctl.scala 391:73]
  wire  _T_1344 = ic_miss_buff_data_valid[5] & _T_1328; // @[el2_ifu_mem_ctl.scala 397:116]
  wire  ic_miss_buff_data_valid_in_5 = write_fill_data_5 | _T_1344; // @[el2_ifu_mem_ctl.scala 397:88]
  wire  _T_1430 = _T_1417 & ic_miss_buff_data_valid_in_5; // @[Mux.scala 27:72]
  wire  _T_1437 = _T_1436 | _T_1430; // @[Mux.scala 27:72]
  wire  _T_1420 = bypass_index[4:2] == 3'h6; // @[el2_ifu_mem_ctl.scala 408:114]
  wire  _T_1293 = io_ifu_axi_rid == 3'h6; // @[el2_ifu_mem_ctl.scala 391:91]
  wire  write_fill_data_6 = bus_ifu_wr_en & _T_1293; // @[el2_ifu_mem_ctl.scala 391:73]
  wire  _T_1347 = ic_miss_buff_data_valid[6] & _T_1328; // @[el2_ifu_mem_ctl.scala 397:116]
  wire  ic_miss_buff_data_valid_in_6 = write_fill_data_6 | _T_1347; // @[el2_ifu_mem_ctl.scala 397:88]
  wire  _T_1431 = _T_1420 & ic_miss_buff_data_valid_in_6; // @[Mux.scala 27:72]
  wire  _T_1438 = _T_1437 | _T_1431; // @[Mux.scala 27:72]
  wire  _T_1423 = bypass_index[4:2] == 3'h7; // @[el2_ifu_mem_ctl.scala 408:114]
  wire  _T_1294 = io_ifu_axi_rid == 3'h7; // @[el2_ifu_mem_ctl.scala 391:91]
  wire  write_fill_data_7 = bus_ifu_wr_en & _T_1294; // @[el2_ifu_mem_ctl.scala 391:73]
  wire  _T_1350 = ic_miss_buff_data_valid[7] & _T_1328; // @[el2_ifu_mem_ctl.scala 397:116]
  wire  ic_miss_buff_data_valid_in_7 = write_fill_data_7 | _T_1350; // @[el2_ifu_mem_ctl.scala 397:88]
  wire  _T_1432 = _T_1423 & ic_miss_buff_data_valid_in_7; // @[Mux.scala 27:72]
  wire  bypass_valid_value_check = _T_1438 | _T_1432; // @[Mux.scala 27:72]
  wire  _T_1441 = ~bypass_index[1]; // @[el2_ifu_mem_ctl.scala 409:58]
  wire  _T_1442 = bypass_valid_value_check & _T_1441; // @[el2_ifu_mem_ctl.scala 409:56]
  wire  _T_1444 = ~bypass_index[0]; // @[el2_ifu_mem_ctl.scala 409:77]
  wire  _T_1445 = _T_1442 & _T_1444; // @[el2_ifu_mem_ctl.scala 409:75]
  wire  _T_1450 = _T_1442 & bypass_index[0]; // @[el2_ifu_mem_ctl.scala 410:75]
  wire  _T_1451 = _T_1445 | _T_1450; // @[el2_ifu_mem_ctl.scala 409:95]
  wire  _T_1453 = bypass_valid_value_check & bypass_index[1]; // @[el2_ifu_mem_ctl.scala 411:56]
  wire  _T_1456 = _T_1453 & _T_1444; // @[el2_ifu_mem_ctl.scala 411:74]
  wire  _T_1457 = _T_1451 | _T_1456; // @[el2_ifu_mem_ctl.scala 410:94]
  wire  _T_1461 = _T_1453 & bypass_index[0]; // @[el2_ifu_mem_ctl.scala 412:51]
  wire [2:0] bypass_index_5_3_inc = bypass_index[4:2] + 3'h1; // @[el2_ifu_mem_ctl.scala 407:70]
  wire  _T_1462 = bypass_index_5_3_inc == 3'h0; // @[el2_ifu_mem_ctl.scala 412:132]
  wire  _T_1478 = _T_1462 & ic_miss_buff_data_valid_in_0; // @[Mux.scala 27:72]
  wire  _T_1464 = bypass_index_5_3_inc == 3'h1; // @[el2_ifu_mem_ctl.scala 412:132]
  wire  _T_1479 = _T_1464 & ic_miss_buff_data_valid_in_1; // @[Mux.scala 27:72]
  wire  _T_1486 = _T_1478 | _T_1479; // @[Mux.scala 27:72]
  wire  _T_1466 = bypass_index_5_3_inc == 3'h2; // @[el2_ifu_mem_ctl.scala 412:132]
  wire  _T_1480 = _T_1466 & ic_miss_buff_data_valid_in_2; // @[Mux.scala 27:72]
  wire  _T_1487 = _T_1486 | _T_1480; // @[Mux.scala 27:72]
  wire  _T_1468 = bypass_index_5_3_inc == 3'h3; // @[el2_ifu_mem_ctl.scala 412:132]
  wire  _T_1481 = _T_1468 & ic_miss_buff_data_valid_in_3; // @[Mux.scala 27:72]
  wire  _T_1488 = _T_1487 | _T_1481; // @[Mux.scala 27:72]
  wire  _T_1470 = bypass_index_5_3_inc == 3'h4; // @[el2_ifu_mem_ctl.scala 412:132]
  wire  _T_1482 = _T_1470 & ic_miss_buff_data_valid_in_4; // @[Mux.scala 27:72]
  wire  _T_1489 = _T_1488 | _T_1482; // @[Mux.scala 27:72]
  wire  _T_1472 = bypass_index_5_3_inc == 3'h5; // @[el2_ifu_mem_ctl.scala 412:132]
  wire  _T_1483 = _T_1472 & ic_miss_buff_data_valid_in_5; // @[Mux.scala 27:72]
  wire  _T_1490 = _T_1489 | _T_1483; // @[Mux.scala 27:72]
  wire  _T_1474 = bypass_index_5_3_inc == 3'h6; // @[el2_ifu_mem_ctl.scala 412:132]
  wire  _T_1484 = _T_1474 & ic_miss_buff_data_valid_in_6; // @[Mux.scala 27:72]
  wire  _T_1491 = _T_1490 | _T_1484; // @[Mux.scala 27:72]
  wire  _T_1476 = bypass_index_5_3_inc == 3'h7; // @[el2_ifu_mem_ctl.scala 412:132]
  wire  _T_1485 = _T_1476 & ic_miss_buff_data_valid_in_7; // @[Mux.scala 27:72]
  wire  _T_1492 = _T_1491 | _T_1485; // @[Mux.scala 27:72]
  wire  _T_1494 = _T_1461 & _T_1492; // @[el2_ifu_mem_ctl.scala 412:69]
  wire  _T_1495 = _T_1457 | _T_1494; // @[el2_ifu_mem_ctl.scala 411:94]
  wire [4:0] _GEN_664 = {{2'd0}, bypass_index[4:2]}; // @[el2_ifu_mem_ctl.scala 413:95]
  wire  _T_1498 = _GEN_664 == 5'h1f; // @[el2_ifu_mem_ctl.scala 413:95]
  wire  _T_1499 = bypass_valid_value_check & _T_1498; // @[el2_ifu_mem_ctl.scala 413:56]
  wire  bypass_data_ready_in = _T_1495 | _T_1499; // @[el2_ifu_mem_ctl.scala 412:181]
  wire  _T_1500 = bypass_data_ready_in & crit_wd_byp_ok_ff; // @[el2_ifu_mem_ctl.scala 417:53]
  wire  _T_1501 = _T_1500 & uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 417:73]
  wire  _T_1503 = _T_1501 & _T_318; // @[el2_ifu_mem_ctl.scala 417:96]
  wire  _T_1505 = _T_1503 & _T_59; // @[el2_ifu_mem_ctl.scala 417:118]
  wire  _T_1507 = crit_wd_byp_ok_ff & _T_51; // @[el2_ifu_mem_ctl.scala 418:73]
  wire  _T_1509 = _T_1507 & _T_318; // @[el2_ifu_mem_ctl.scala 418:96]
  wire  _T_1511 = _T_1509 & _T_59; // @[el2_ifu_mem_ctl.scala 418:118]
  wire  _T_1512 = _T_1505 | _T_1511; // @[el2_ifu_mem_ctl.scala 417:143]
  reg  ic_crit_wd_rdy_new_ff; // @[el2_ifu_mem_ctl.scala 420:58]
  wire  _T_1513 = ic_crit_wd_rdy_new_ff & crit_wd_byp_ok_ff; // @[el2_ifu_mem_ctl.scala 419:54]
  wire  _T_1514 = ~fetch_req_icache_f; // @[el2_ifu_mem_ctl.scala 419:76]
  wire  _T_1515 = _T_1513 & _T_1514; // @[el2_ifu_mem_ctl.scala 419:74]
  wire  _T_1517 = _T_1515 & _T_318; // @[el2_ifu_mem_ctl.scala 419:96]
  wire  ic_crit_wd_rdy_new_in = _T_1512 | _T_1517; // @[el2_ifu_mem_ctl.scala 418:143]
  wire  ic_crit_wd_rdy = ic_crit_wd_rdy_new_in | ic_crit_wd_rdy_new_ff; // @[el2_ifu_mem_ctl.scala 617:43]
  wire  _T_1254 = ic_crit_wd_rdy | _T_2222; // @[el2_ifu_mem_ctl.scala 364:38]
  wire  _T_1256 = _T_1254 | _T_2238; // @[el2_ifu_mem_ctl.scala 364:64]
  wire  _T_1257 = ~_T_1256; // @[el2_ifu_mem_ctl.scala 364:21]
  wire  _T_1258 = ~fetch_req_iccm_f; // @[el2_ifu_mem_ctl.scala 364:98]
  wire  sel_ic_data = _T_1257 & _T_1258; // @[el2_ifu_mem_ctl.scala 364:96]
  wire  _T_2405 = io_ic_tag_perr & sel_ic_data; // @[el2_ifu_mem_ctl.scala 462:44]
  wire  _T_1611 = ifu_fetch_addr_int_f[1] & ifu_fetch_addr_int_f[0]; // @[el2_ifu_mem_ctl.scala 431:31]
  reg [7:0] ic_miss_buff_data_error; // @[el2_ifu_mem_ctl.scala 403:60]
  wire  _T_1555 = _T_1402 & ic_miss_buff_data_error[0]; // @[Mux.scala 27:72]
  wire  _T_1556 = _T_1405 & ic_miss_buff_data_error[1]; // @[Mux.scala 27:72]
  wire  _T_1563 = _T_1555 | _T_1556; // @[Mux.scala 27:72]
  wire  _T_1557 = _T_1408 & ic_miss_buff_data_error[2]; // @[Mux.scala 27:72]
  wire  _T_1564 = _T_1563 | _T_1557; // @[Mux.scala 27:72]
  wire  _T_1558 = _T_1411 & ic_miss_buff_data_error[3]; // @[Mux.scala 27:72]
  wire  _T_1565 = _T_1564 | _T_1558; // @[Mux.scala 27:72]
  wire  _T_1559 = _T_1414 & ic_miss_buff_data_error[4]; // @[Mux.scala 27:72]
  wire  _T_1566 = _T_1565 | _T_1559; // @[Mux.scala 27:72]
  wire  _T_1560 = _T_1417 & ic_miss_buff_data_error[5]; // @[Mux.scala 27:72]
  wire  _T_1567 = _T_1566 | _T_1560; // @[Mux.scala 27:72]
  wire  _T_1561 = _T_1420 & ic_miss_buff_data_error[6]; // @[Mux.scala 27:72]
  wire  _T_1568 = _T_1567 | _T_1561; // @[Mux.scala 27:72]
  wire  _T_1562 = _T_1423 & ic_miss_buff_data_error[7]; // @[Mux.scala 27:72]
  wire  ic_miss_buff_data_error_bypass = _T_1568 | _T_1562; // @[Mux.scala 27:72]
  wire  _T_1594 = _T_2155 & ic_miss_buff_data_error[0]; // @[Mux.scala 27:72]
  wire  _T_1595 = _T_2158 & ic_miss_buff_data_error[1]; // @[Mux.scala 27:72]
  wire  _T_1602 = _T_1594 | _T_1595; // @[Mux.scala 27:72]
  wire  _T_1596 = _T_2161 & ic_miss_buff_data_error[2]; // @[Mux.scala 27:72]
  wire  _T_1603 = _T_1602 | _T_1596; // @[Mux.scala 27:72]
  wire  _T_1597 = _T_2164 & ic_miss_buff_data_error[3]; // @[Mux.scala 27:72]
  wire  _T_1604 = _T_1603 | _T_1597; // @[Mux.scala 27:72]
  wire  _T_1598 = _T_2167 & ic_miss_buff_data_error[4]; // @[Mux.scala 27:72]
  wire  _T_1605 = _T_1604 | _T_1598; // @[Mux.scala 27:72]
  wire  _T_1599 = _T_2170 & ic_miss_buff_data_error[5]; // @[Mux.scala 27:72]
  wire  _T_1606 = _T_1605 | _T_1599; // @[Mux.scala 27:72]
  wire  _T_1600 = _T_2173 & ic_miss_buff_data_error[6]; // @[Mux.scala 27:72]
  wire  _T_1607 = _T_1606 | _T_1600; // @[Mux.scala 27:72]
  wire  _T_1601 = _T_2176 & ic_miss_buff_data_error[7]; // @[Mux.scala 27:72]
  wire  ic_miss_buff_data_error_bypass_inc = _T_1607 | _T_1601; // @[Mux.scala 27:72]
  wire  _T_1612 = ic_miss_buff_data_error_bypass | ic_miss_buff_data_error_bypass_inc; // @[el2_ifu_mem_ctl.scala 433:70]
  wire  ifu_byp_data_err_new = _T_1611 ? ic_miss_buff_data_error_bypass : _T_1612; // @[el2_ifu_mem_ctl.scala 431:56]
  wire  ifc_bus_acc_fault_f = ic_byp_hit_f & ifu_byp_data_err_new; // @[el2_ifu_mem_ctl.scala 375:42]
  wire  _T_2406 = ifc_region_acc_fault_final_f | ifc_bus_acc_fault_f; // @[el2_ifu_mem_ctl.scala 462:91]
  wire  _T_2407 = ~_T_2406; // @[el2_ifu_mem_ctl.scala 462:60]
  wire  ic_rd_parity_final_err = _T_2405 & _T_2407; // @[el2_ifu_mem_ctl.scala 462:58]
  reg  ic_debug_ict_array_sel_ff; // @[Reg.scala 27:20]
  reg  ic_tag_valid_out_1_0; // @[Reg.scala 27:20]
  wire  _T_9678 = _T_4472 ? 1'h0 : ic_tag_valid_out_1_0; // @[el2_ifu_mem_ctl.scala 744:10]
  reg  ic_tag_valid_out_1_1; // @[Reg.scala 27:20]
  wire  _T_9680 = _T_4476 ? 1'h0 : ic_tag_valid_out_1_1; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9933 = _T_9678 | _T_9680; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_2; // @[Reg.scala 27:20]
  wire  _T_9682 = _T_4480 ? 1'h0 : ic_tag_valid_out_1_2; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9934 = _T_9933 | _T_9682; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_3; // @[Reg.scala 27:20]
  wire  _T_9684 = _T_4484 ? 1'h0 : ic_tag_valid_out_1_3; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9935 = _T_9934 | _T_9684; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_4; // @[Reg.scala 27:20]
  wire  _T_9686 = _T_4488 ? 1'h0 : ic_tag_valid_out_1_4; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9936 = _T_9935 | _T_9686; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_5; // @[Reg.scala 27:20]
  wire  _T_9688 = _T_4492 ? 1'h0 : ic_tag_valid_out_1_5; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9937 = _T_9936 | _T_9688; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_6; // @[Reg.scala 27:20]
  wire  _T_9690 = _T_4496 ? 1'h0 : ic_tag_valid_out_1_6; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9938 = _T_9937 | _T_9690; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_7; // @[Reg.scala 27:20]
  wire  _T_9692 = _T_4500 ? 1'h0 : ic_tag_valid_out_1_7; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9939 = _T_9938 | _T_9692; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_8; // @[Reg.scala 27:20]
  wire  _T_9694 = _T_4504 ? 1'h0 : ic_tag_valid_out_1_8; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9940 = _T_9939 | _T_9694; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_9; // @[Reg.scala 27:20]
  wire  _T_9696 = _T_4508 ? 1'h0 : ic_tag_valid_out_1_9; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9941 = _T_9940 | _T_9696; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_10; // @[Reg.scala 27:20]
  wire  _T_9698 = _T_4512 ? 1'h0 : ic_tag_valid_out_1_10; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9942 = _T_9941 | _T_9698; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_11; // @[Reg.scala 27:20]
  wire  _T_9700 = _T_4516 ? 1'h0 : ic_tag_valid_out_1_11; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9943 = _T_9942 | _T_9700; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_12; // @[Reg.scala 27:20]
  wire  _T_9702 = _T_4520 ? 1'h0 : ic_tag_valid_out_1_12; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9944 = _T_9943 | _T_9702; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_13; // @[Reg.scala 27:20]
  wire  _T_9704 = _T_4524 ? 1'h0 : ic_tag_valid_out_1_13; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9945 = _T_9944 | _T_9704; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_14; // @[Reg.scala 27:20]
  wire  _T_9706 = _T_4528 ? 1'h0 : ic_tag_valid_out_1_14; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9946 = _T_9945 | _T_9706; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_15; // @[Reg.scala 27:20]
  wire  _T_9708 = _T_4532 ? 1'h0 : ic_tag_valid_out_1_15; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9947 = _T_9946 | _T_9708; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_16; // @[Reg.scala 27:20]
  wire  _T_9710 = _T_4536 ? 1'h0 : ic_tag_valid_out_1_16; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9948 = _T_9947 | _T_9710; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_17; // @[Reg.scala 27:20]
  wire  _T_9712 = _T_4540 ? 1'h0 : ic_tag_valid_out_1_17; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9949 = _T_9948 | _T_9712; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_18; // @[Reg.scala 27:20]
  wire  _T_9714 = _T_4544 ? 1'h0 : ic_tag_valid_out_1_18; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9950 = _T_9949 | _T_9714; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_19; // @[Reg.scala 27:20]
  wire  _T_9716 = _T_4548 ? 1'h0 : ic_tag_valid_out_1_19; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9951 = _T_9950 | _T_9716; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_20; // @[Reg.scala 27:20]
  wire  _T_9718 = _T_4552 ? 1'h0 : ic_tag_valid_out_1_20; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9952 = _T_9951 | _T_9718; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_21; // @[Reg.scala 27:20]
  wire  _T_9720 = _T_4556 ? 1'h0 : ic_tag_valid_out_1_21; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9953 = _T_9952 | _T_9720; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_22; // @[Reg.scala 27:20]
  wire  _T_9722 = _T_4560 ? 1'h0 : ic_tag_valid_out_1_22; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9954 = _T_9953 | _T_9722; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_23; // @[Reg.scala 27:20]
  wire  _T_9724 = _T_4564 ? 1'h0 : ic_tag_valid_out_1_23; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9955 = _T_9954 | _T_9724; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_24; // @[Reg.scala 27:20]
  wire  _T_9726 = _T_4568 ? 1'h0 : ic_tag_valid_out_1_24; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9956 = _T_9955 | _T_9726; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_25; // @[Reg.scala 27:20]
  wire  _T_9728 = _T_4572 ? 1'h0 : ic_tag_valid_out_1_25; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9957 = _T_9956 | _T_9728; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_26; // @[Reg.scala 27:20]
  wire  _T_9730 = _T_4576 ? 1'h0 : ic_tag_valid_out_1_26; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9958 = _T_9957 | _T_9730; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_27; // @[Reg.scala 27:20]
  wire  _T_9732 = _T_4580 ? 1'h0 : ic_tag_valid_out_1_27; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9959 = _T_9958 | _T_9732; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_28; // @[Reg.scala 27:20]
  wire  _T_9734 = _T_4584 ? 1'h0 : ic_tag_valid_out_1_28; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9960 = _T_9959 | _T_9734; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_29; // @[Reg.scala 27:20]
  wire  _T_9736 = _T_4588 ? 1'h0 : ic_tag_valid_out_1_29; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9961 = _T_9960 | _T_9736; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_30; // @[Reg.scala 27:20]
  wire  _T_9738 = _T_4592 ? 1'h0 : ic_tag_valid_out_1_30; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9962 = _T_9961 | _T_9738; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_31; // @[Reg.scala 27:20]
  wire  _T_9740 = _T_4596 ? 1'h0 : ic_tag_valid_out_1_31; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9963 = _T_9962 | _T_9740; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_32; // @[Reg.scala 27:20]
  wire  _T_9742 = _T_4600 ? 1'h0 : ic_tag_valid_out_1_32; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9964 = _T_9963 | _T_9742; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_33; // @[Reg.scala 27:20]
  wire  _T_9744 = _T_4604 ? 1'h0 : ic_tag_valid_out_1_33; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9965 = _T_9964 | _T_9744; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_34; // @[Reg.scala 27:20]
  wire  _T_9746 = _T_4608 ? 1'h0 : ic_tag_valid_out_1_34; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9966 = _T_9965 | _T_9746; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_35; // @[Reg.scala 27:20]
  wire  _T_9748 = _T_4612 ? 1'h0 : ic_tag_valid_out_1_35; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9967 = _T_9966 | _T_9748; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_36; // @[Reg.scala 27:20]
  wire  _T_9750 = _T_4616 ? 1'h0 : ic_tag_valid_out_1_36; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9968 = _T_9967 | _T_9750; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_37; // @[Reg.scala 27:20]
  wire  _T_9752 = _T_4620 ? 1'h0 : ic_tag_valid_out_1_37; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9969 = _T_9968 | _T_9752; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_38; // @[Reg.scala 27:20]
  wire  _T_9754 = _T_4624 ? 1'h0 : ic_tag_valid_out_1_38; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9970 = _T_9969 | _T_9754; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_39; // @[Reg.scala 27:20]
  wire  _T_9756 = _T_4628 ? 1'h0 : ic_tag_valid_out_1_39; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9971 = _T_9970 | _T_9756; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_40; // @[Reg.scala 27:20]
  wire  _T_9758 = _T_4632 ? 1'h0 : ic_tag_valid_out_1_40; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9972 = _T_9971 | _T_9758; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_41; // @[Reg.scala 27:20]
  wire  _T_9760 = _T_4636 ? 1'h0 : ic_tag_valid_out_1_41; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9973 = _T_9972 | _T_9760; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_42; // @[Reg.scala 27:20]
  wire  _T_9762 = _T_4640 ? 1'h0 : ic_tag_valid_out_1_42; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9974 = _T_9973 | _T_9762; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_43; // @[Reg.scala 27:20]
  wire  _T_9764 = _T_4644 ? 1'h0 : ic_tag_valid_out_1_43; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9975 = _T_9974 | _T_9764; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_44; // @[Reg.scala 27:20]
  wire  _T_9766 = _T_4648 ? 1'h0 : ic_tag_valid_out_1_44; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9976 = _T_9975 | _T_9766; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_45; // @[Reg.scala 27:20]
  wire  _T_9768 = _T_4652 ? 1'h0 : ic_tag_valid_out_1_45; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9977 = _T_9976 | _T_9768; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_46; // @[Reg.scala 27:20]
  wire  _T_9770 = _T_4656 ? 1'h0 : ic_tag_valid_out_1_46; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9978 = _T_9977 | _T_9770; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_47; // @[Reg.scala 27:20]
  wire  _T_9772 = _T_4660 ? 1'h0 : ic_tag_valid_out_1_47; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9979 = _T_9978 | _T_9772; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_48; // @[Reg.scala 27:20]
  wire  _T_9774 = _T_4664 ? 1'h0 : ic_tag_valid_out_1_48; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9980 = _T_9979 | _T_9774; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_49; // @[Reg.scala 27:20]
  wire  _T_9776 = _T_4668 ? 1'h0 : ic_tag_valid_out_1_49; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9981 = _T_9980 | _T_9776; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_50; // @[Reg.scala 27:20]
  wire  _T_9778 = _T_4672 ? 1'h0 : ic_tag_valid_out_1_50; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9982 = _T_9981 | _T_9778; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_51; // @[Reg.scala 27:20]
  wire  _T_9780 = _T_4676 ? 1'h0 : ic_tag_valid_out_1_51; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9983 = _T_9982 | _T_9780; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_52; // @[Reg.scala 27:20]
  wire  _T_9782 = _T_4680 ? 1'h0 : ic_tag_valid_out_1_52; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9984 = _T_9983 | _T_9782; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_53; // @[Reg.scala 27:20]
  wire  _T_9784 = _T_4684 ? 1'h0 : ic_tag_valid_out_1_53; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9985 = _T_9984 | _T_9784; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_54; // @[Reg.scala 27:20]
  wire  _T_9786 = _T_4688 ? 1'h0 : ic_tag_valid_out_1_54; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9986 = _T_9985 | _T_9786; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_55; // @[Reg.scala 27:20]
  wire  _T_9788 = _T_4692 ? 1'h0 : ic_tag_valid_out_1_55; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9987 = _T_9986 | _T_9788; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_56; // @[Reg.scala 27:20]
  wire  _T_9790 = _T_4696 ? 1'h0 : ic_tag_valid_out_1_56; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9988 = _T_9987 | _T_9790; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_57; // @[Reg.scala 27:20]
  wire  _T_9792 = _T_4700 ? 1'h0 : ic_tag_valid_out_1_57; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9989 = _T_9988 | _T_9792; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_58; // @[Reg.scala 27:20]
  wire  _T_9794 = _T_4704 ? 1'h0 : ic_tag_valid_out_1_58; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9990 = _T_9989 | _T_9794; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_59; // @[Reg.scala 27:20]
  wire  _T_9796 = _T_4708 ? 1'h0 : ic_tag_valid_out_1_59; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9991 = _T_9990 | _T_9796; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_60; // @[Reg.scala 27:20]
  wire  _T_9798 = _T_4712 ? 1'h0 : ic_tag_valid_out_1_60; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9992 = _T_9991 | _T_9798; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_61; // @[Reg.scala 27:20]
  wire  _T_9800 = _T_4716 ? 1'h0 : ic_tag_valid_out_1_61; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9993 = _T_9992 | _T_9800; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_62; // @[Reg.scala 27:20]
  wire  _T_9802 = _T_4720 ? 1'h0 : ic_tag_valid_out_1_62; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9994 = _T_9993 | _T_9802; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_63; // @[Reg.scala 27:20]
  wire  _T_9804 = _T_4724 ? 1'h0 : ic_tag_valid_out_1_63; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9995 = _T_9994 | _T_9804; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_64; // @[Reg.scala 27:20]
  wire  _T_9806 = _T_4728 ? 1'h0 : ic_tag_valid_out_1_64; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9996 = _T_9995 | _T_9806; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_65; // @[Reg.scala 27:20]
  wire  _T_9808 = _T_4732 ? 1'h0 : ic_tag_valid_out_1_65; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9997 = _T_9996 | _T_9808; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_66; // @[Reg.scala 27:20]
  wire  _T_9810 = _T_4736 ? 1'h0 : ic_tag_valid_out_1_66; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9998 = _T_9997 | _T_9810; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_67; // @[Reg.scala 27:20]
  wire  _T_9812 = _T_4740 ? 1'h0 : ic_tag_valid_out_1_67; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9999 = _T_9998 | _T_9812; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_68; // @[Reg.scala 27:20]
  wire  _T_9814 = _T_4744 ? 1'h0 : ic_tag_valid_out_1_68; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_10000 = _T_9999 | _T_9814; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_69; // @[Reg.scala 27:20]
  wire  _T_9816 = _T_4748 ? 1'h0 : ic_tag_valid_out_1_69; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_10001 = _T_10000 | _T_9816; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_70; // @[Reg.scala 27:20]
  wire  _T_9818 = _T_4752 ? 1'h0 : ic_tag_valid_out_1_70; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_10002 = _T_10001 | _T_9818; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_71; // @[Reg.scala 27:20]
  wire  _T_9820 = _T_4756 ? 1'h0 : ic_tag_valid_out_1_71; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_10003 = _T_10002 | _T_9820; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_72; // @[Reg.scala 27:20]
  wire  _T_9822 = _T_4760 ? 1'h0 : ic_tag_valid_out_1_72; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_10004 = _T_10003 | _T_9822; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_73; // @[Reg.scala 27:20]
  wire  _T_9824 = _T_4764 ? 1'h0 : ic_tag_valid_out_1_73; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_10005 = _T_10004 | _T_9824; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_74; // @[Reg.scala 27:20]
  wire  _T_9826 = _T_4768 ? 1'h0 : ic_tag_valid_out_1_74; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_10006 = _T_10005 | _T_9826; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_75; // @[Reg.scala 27:20]
  wire  _T_9828 = _T_4772 ? 1'h0 : ic_tag_valid_out_1_75; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_10007 = _T_10006 | _T_9828; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_76; // @[Reg.scala 27:20]
  wire  _T_9830 = _T_4776 ? 1'h0 : ic_tag_valid_out_1_76; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_10008 = _T_10007 | _T_9830; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_77; // @[Reg.scala 27:20]
  wire  _T_9832 = _T_4780 ? 1'h0 : ic_tag_valid_out_1_77; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_10009 = _T_10008 | _T_9832; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_78; // @[Reg.scala 27:20]
  wire  _T_9834 = _T_4784 ? 1'h0 : ic_tag_valid_out_1_78; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_10010 = _T_10009 | _T_9834; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_79; // @[Reg.scala 27:20]
  wire  _T_9836 = _T_4788 ? 1'h0 : ic_tag_valid_out_1_79; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_10011 = _T_10010 | _T_9836; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_80; // @[Reg.scala 27:20]
  wire  _T_9838 = _T_4792 ? 1'h0 : ic_tag_valid_out_1_80; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_10012 = _T_10011 | _T_9838; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_81; // @[Reg.scala 27:20]
  wire  _T_9840 = _T_4796 ? 1'h0 : ic_tag_valid_out_1_81; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_10013 = _T_10012 | _T_9840; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_82; // @[Reg.scala 27:20]
  wire  _T_9842 = _T_4800 ? 1'h0 : ic_tag_valid_out_1_82; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_10014 = _T_10013 | _T_9842; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_83; // @[Reg.scala 27:20]
  wire  _T_9844 = _T_4804 ? 1'h0 : ic_tag_valid_out_1_83; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_10015 = _T_10014 | _T_9844; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_84; // @[Reg.scala 27:20]
  wire  _T_9846 = _T_4808 ? 1'h0 : ic_tag_valid_out_1_84; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_10016 = _T_10015 | _T_9846; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_85; // @[Reg.scala 27:20]
  wire  _T_9848 = _T_4812 ? 1'h0 : ic_tag_valid_out_1_85; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_10017 = _T_10016 | _T_9848; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_86; // @[Reg.scala 27:20]
  wire  _T_9850 = _T_4816 ? 1'h0 : ic_tag_valid_out_1_86; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_10018 = _T_10017 | _T_9850; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_87; // @[Reg.scala 27:20]
  wire  _T_9852 = _T_4820 ? 1'h0 : ic_tag_valid_out_1_87; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_10019 = _T_10018 | _T_9852; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_88; // @[Reg.scala 27:20]
  wire  _T_9854 = _T_4824 ? 1'h0 : ic_tag_valid_out_1_88; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_10020 = _T_10019 | _T_9854; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_89; // @[Reg.scala 27:20]
  wire  _T_9856 = _T_4828 ? 1'h0 : ic_tag_valid_out_1_89; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_10021 = _T_10020 | _T_9856; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_90; // @[Reg.scala 27:20]
  wire  _T_9858 = _T_4832 ? 1'h0 : ic_tag_valid_out_1_90; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_10022 = _T_10021 | _T_9858; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_91; // @[Reg.scala 27:20]
  wire  _T_9860 = _T_4836 ? 1'h0 : ic_tag_valid_out_1_91; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_10023 = _T_10022 | _T_9860; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_92; // @[Reg.scala 27:20]
  wire  _T_9862 = _T_4840 ? 1'h0 : ic_tag_valid_out_1_92; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_10024 = _T_10023 | _T_9862; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_93; // @[Reg.scala 27:20]
  wire  _T_9864 = _T_4844 ? 1'h0 : ic_tag_valid_out_1_93; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_10025 = _T_10024 | _T_9864; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_94; // @[Reg.scala 27:20]
  wire  _T_9866 = _T_4848 ? 1'h0 : ic_tag_valid_out_1_94; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_10026 = _T_10025 | _T_9866; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_95; // @[Reg.scala 27:20]
  wire  _T_9868 = _T_4852 ? 1'h0 : ic_tag_valid_out_1_95; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_10027 = _T_10026 | _T_9868; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_96; // @[Reg.scala 27:20]
  wire  _T_9870 = _T_4856 ? 1'h0 : ic_tag_valid_out_1_96; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_10028 = _T_10027 | _T_9870; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_97; // @[Reg.scala 27:20]
  wire  _T_9872 = _T_4860 ? 1'h0 : ic_tag_valid_out_1_97; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_10029 = _T_10028 | _T_9872; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_98; // @[Reg.scala 27:20]
  wire  _T_9874 = _T_4864 ? 1'h0 : ic_tag_valid_out_1_98; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_10030 = _T_10029 | _T_9874; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_99; // @[Reg.scala 27:20]
  wire  _T_9876 = _T_4868 ? 1'h0 : ic_tag_valid_out_1_99; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_10031 = _T_10030 | _T_9876; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_100; // @[Reg.scala 27:20]
  wire  _T_9878 = _T_4872 ? 1'h0 : ic_tag_valid_out_1_100; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_10032 = _T_10031 | _T_9878; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_101; // @[Reg.scala 27:20]
  wire  _T_9880 = _T_4876 ? 1'h0 : ic_tag_valid_out_1_101; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_10033 = _T_10032 | _T_9880; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_102; // @[Reg.scala 27:20]
  wire  _T_9882 = _T_4880 ? 1'h0 : ic_tag_valid_out_1_102; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_10034 = _T_10033 | _T_9882; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_103; // @[Reg.scala 27:20]
  wire  _T_9884 = _T_4884 ? 1'h0 : ic_tag_valid_out_1_103; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_10035 = _T_10034 | _T_9884; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_104; // @[Reg.scala 27:20]
  wire  _T_9886 = _T_4888 ? 1'h0 : ic_tag_valid_out_1_104; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_10036 = _T_10035 | _T_9886; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_105; // @[Reg.scala 27:20]
  wire  _T_9888 = _T_4892 ? 1'h0 : ic_tag_valid_out_1_105; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_10037 = _T_10036 | _T_9888; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_106; // @[Reg.scala 27:20]
  wire  _T_9890 = _T_4896 ? 1'h0 : ic_tag_valid_out_1_106; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_10038 = _T_10037 | _T_9890; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_107; // @[Reg.scala 27:20]
  wire  _T_9892 = _T_4900 ? 1'h0 : ic_tag_valid_out_1_107; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_10039 = _T_10038 | _T_9892; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_108; // @[Reg.scala 27:20]
  wire  _T_9894 = _T_4904 ? 1'h0 : ic_tag_valid_out_1_108; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_10040 = _T_10039 | _T_9894; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_109; // @[Reg.scala 27:20]
  wire  _T_9896 = _T_4908 ? 1'h0 : ic_tag_valid_out_1_109; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_10041 = _T_10040 | _T_9896; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_110; // @[Reg.scala 27:20]
  wire  _T_9898 = _T_4912 ? 1'h0 : ic_tag_valid_out_1_110; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_10042 = _T_10041 | _T_9898; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_111; // @[Reg.scala 27:20]
  wire  _T_9900 = _T_4916 ? 1'h0 : ic_tag_valid_out_1_111; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_10043 = _T_10042 | _T_9900; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_112; // @[Reg.scala 27:20]
  wire  _T_9902 = _T_4920 ? 1'h0 : ic_tag_valid_out_1_112; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_10044 = _T_10043 | _T_9902; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_113; // @[Reg.scala 27:20]
  wire  _T_9904 = _T_4924 ? 1'h0 : ic_tag_valid_out_1_113; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_10045 = _T_10044 | _T_9904; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_114; // @[Reg.scala 27:20]
  wire  _T_9906 = _T_4928 ? 1'h0 : ic_tag_valid_out_1_114; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_10046 = _T_10045 | _T_9906; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_115; // @[Reg.scala 27:20]
  wire  _T_9908 = _T_4932 ? 1'h0 : ic_tag_valid_out_1_115; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_10047 = _T_10046 | _T_9908; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_116; // @[Reg.scala 27:20]
  wire  _T_9910 = _T_4936 ? 1'h0 : ic_tag_valid_out_1_116; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_10048 = _T_10047 | _T_9910; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_117; // @[Reg.scala 27:20]
  wire  _T_9912 = _T_4940 ? 1'h0 : ic_tag_valid_out_1_117; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_10049 = _T_10048 | _T_9912; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_118; // @[Reg.scala 27:20]
  wire  _T_9914 = _T_4944 ? 1'h0 : ic_tag_valid_out_1_118; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_10050 = _T_10049 | _T_9914; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_119; // @[Reg.scala 27:20]
  wire  _T_9916 = _T_4948 ? 1'h0 : ic_tag_valid_out_1_119; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_10051 = _T_10050 | _T_9916; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_120; // @[Reg.scala 27:20]
  wire  _T_9918 = _T_4952 ? 1'h0 : ic_tag_valid_out_1_120; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_10052 = _T_10051 | _T_9918; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_121; // @[Reg.scala 27:20]
  wire  _T_9920 = _T_4956 ? 1'h0 : ic_tag_valid_out_1_121; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_10053 = _T_10052 | _T_9920; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_122; // @[Reg.scala 27:20]
  wire  _T_9922 = _T_4960 ? 1'h0 : ic_tag_valid_out_1_122; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_10054 = _T_10053 | _T_9922; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_123; // @[Reg.scala 27:20]
  wire  _T_9924 = _T_4964 ? 1'h0 : ic_tag_valid_out_1_123; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_10055 = _T_10054 | _T_9924; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_124; // @[Reg.scala 27:20]
  wire  _T_9926 = _T_4968 ? 1'h0 : ic_tag_valid_out_1_124; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_10056 = _T_10055 | _T_9926; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_125; // @[Reg.scala 27:20]
  wire  _T_9928 = _T_4972 ? 1'h0 : ic_tag_valid_out_1_125; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_10057 = _T_10056 | _T_9928; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_126; // @[Reg.scala 27:20]
  wire  _T_9930 = _T_4976 ? 1'h0 : ic_tag_valid_out_1_126; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_10058 = _T_10057 | _T_9930; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_1_127; // @[Reg.scala 27:20]
  wire  _T_9932 = _T_4980 ? 1'h0 : ic_tag_valid_out_1_127; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_10059 = _T_10058 | _T_9932; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_0; // @[Reg.scala 27:20]
  wire  _T_9295 = _T_4472 ? 1'h0 : ic_tag_valid_out_0_0; // @[el2_ifu_mem_ctl.scala 744:10]
  reg  ic_tag_valid_out_0_1; // @[Reg.scala 27:20]
  wire  _T_9297 = _T_4476 ? 1'h0 : ic_tag_valid_out_0_1; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9550 = _T_9295 | _T_9297; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_2; // @[Reg.scala 27:20]
  wire  _T_9299 = _T_4480 ? 1'h0 : ic_tag_valid_out_0_2; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9551 = _T_9550 | _T_9299; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_3; // @[Reg.scala 27:20]
  wire  _T_9301 = _T_4484 ? 1'h0 : ic_tag_valid_out_0_3; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9552 = _T_9551 | _T_9301; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_4; // @[Reg.scala 27:20]
  wire  _T_9303 = _T_4488 ? 1'h0 : ic_tag_valid_out_0_4; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9553 = _T_9552 | _T_9303; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_5; // @[Reg.scala 27:20]
  wire  _T_9305 = _T_4492 ? 1'h0 : ic_tag_valid_out_0_5; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9554 = _T_9553 | _T_9305; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_6; // @[Reg.scala 27:20]
  wire  _T_9307 = _T_4496 ? 1'h0 : ic_tag_valid_out_0_6; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9555 = _T_9554 | _T_9307; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_7; // @[Reg.scala 27:20]
  wire  _T_9309 = _T_4500 ? 1'h0 : ic_tag_valid_out_0_7; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9556 = _T_9555 | _T_9309; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_8; // @[Reg.scala 27:20]
  wire  _T_9311 = _T_4504 ? 1'h0 : ic_tag_valid_out_0_8; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9557 = _T_9556 | _T_9311; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_9; // @[Reg.scala 27:20]
  wire  _T_9313 = _T_4508 ? 1'h0 : ic_tag_valid_out_0_9; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9558 = _T_9557 | _T_9313; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_10; // @[Reg.scala 27:20]
  wire  _T_9315 = _T_4512 ? 1'h0 : ic_tag_valid_out_0_10; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9559 = _T_9558 | _T_9315; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_11; // @[Reg.scala 27:20]
  wire  _T_9317 = _T_4516 ? 1'h0 : ic_tag_valid_out_0_11; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9560 = _T_9559 | _T_9317; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_12; // @[Reg.scala 27:20]
  wire  _T_9319 = _T_4520 ? 1'h0 : ic_tag_valid_out_0_12; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9561 = _T_9560 | _T_9319; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_13; // @[Reg.scala 27:20]
  wire  _T_9321 = _T_4524 ? 1'h0 : ic_tag_valid_out_0_13; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9562 = _T_9561 | _T_9321; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_14; // @[Reg.scala 27:20]
  wire  _T_9323 = _T_4528 ? 1'h0 : ic_tag_valid_out_0_14; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9563 = _T_9562 | _T_9323; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_15; // @[Reg.scala 27:20]
  wire  _T_9325 = _T_4532 ? 1'h0 : ic_tag_valid_out_0_15; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9564 = _T_9563 | _T_9325; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_16; // @[Reg.scala 27:20]
  wire  _T_9327 = _T_4536 ? 1'h0 : ic_tag_valid_out_0_16; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9565 = _T_9564 | _T_9327; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_17; // @[Reg.scala 27:20]
  wire  _T_9329 = _T_4540 ? 1'h0 : ic_tag_valid_out_0_17; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9566 = _T_9565 | _T_9329; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_18; // @[Reg.scala 27:20]
  wire  _T_9331 = _T_4544 ? 1'h0 : ic_tag_valid_out_0_18; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9567 = _T_9566 | _T_9331; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_19; // @[Reg.scala 27:20]
  wire  _T_9333 = _T_4548 ? 1'h0 : ic_tag_valid_out_0_19; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9568 = _T_9567 | _T_9333; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_20; // @[Reg.scala 27:20]
  wire  _T_9335 = _T_4552 ? 1'h0 : ic_tag_valid_out_0_20; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9569 = _T_9568 | _T_9335; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_21; // @[Reg.scala 27:20]
  wire  _T_9337 = _T_4556 ? 1'h0 : ic_tag_valid_out_0_21; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9570 = _T_9569 | _T_9337; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_22; // @[Reg.scala 27:20]
  wire  _T_9339 = _T_4560 ? 1'h0 : ic_tag_valid_out_0_22; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9571 = _T_9570 | _T_9339; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_23; // @[Reg.scala 27:20]
  wire  _T_9341 = _T_4564 ? 1'h0 : ic_tag_valid_out_0_23; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9572 = _T_9571 | _T_9341; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_24; // @[Reg.scala 27:20]
  wire  _T_9343 = _T_4568 ? 1'h0 : ic_tag_valid_out_0_24; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9573 = _T_9572 | _T_9343; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_25; // @[Reg.scala 27:20]
  wire  _T_9345 = _T_4572 ? 1'h0 : ic_tag_valid_out_0_25; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9574 = _T_9573 | _T_9345; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_26; // @[Reg.scala 27:20]
  wire  _T_9347 = _T_4576 ? 1'h0 : ic_tag_valid_out_0_26; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9575 = _T_9574 | _T_9347; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_27; // @[Reg.scala 27:20]
  wire  _T_9349 = _T_4580 ? 1'h0 : ic_tag_valid_out_0_27; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9576 = _T_9575 | _T_9349; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_28; // @[Reg.scala 27:20]
  wire  _T_9351 = _T_4584 ? 1'h0 : ic_tag_valid_out_0_28; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9577 = _T_9576 | _T_9351; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_29; // @[Reg.scala 27:20]
  wire  _T_9353 = _T_4588 ? 1'h0 : ic_tag_valid_out_0_29; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9578 = _T_9577 | _T_9353; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_30; // @[Reg.scala 27:20]
  wire  _T_9355 = _T_4592 ? 1'h0 : ic_tag_valid_out_0_30; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9579 = _T_9578 | _T_9355; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_31; // @[Reg.scala 27:20]
  wire  _T_9357 = _T_4596 ? 1'h0 : ic_tag_valid_out_0_31; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9580 = _T_9579 | _T_9357; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_32; // @[Reg.scala 27:20]
  wire  _T_9359 = _T_4600 ? 1'h0 : ic_tag_valid_out_0_32; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9581 = _T_9580 | _T_9359; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_33; // @[Reg.scala 27:20]
  wire  _T_9361 = _T_4604 ? 1'h0 : ic_tag_valid_out_0_33; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9582 = _T_9581 | _T_9361; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_34; // @[Reg.scala 27:20]
  wire  _T_9363 = _T_4608 ? 1'h0 : ic_tag_valid_out_0_34; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9583 = _T_9582 | _T_9363; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_35; // @[Reg.scala 27:20]
  wire  _T_9365 = _T_4612 ? 1'h0 : ic_tag_valid_out_0_35; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9584 = _T_9583 | _T_9365; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_36; // @[Reg.scala 27:20]
  wire  _T_9367 = _T_4616 ? 1'h0 : ic_tag_valid_out_0_36; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9585 = _T_9584 | _T_9367; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_37; // @[Reg.scala 27:20]
  wire  _T_9369 = _T_4620 ? 1'h0 : ic_tag_valid_out_0_37; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9586 = _T_9585 | _T_9369; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_38; // @[Reg.scala 27:20]
  wire  _T_9371 = _T_4624 ? 1'h0 : ic_tag_valid_out_0_38; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9587 = _T_9586 | _T_9371; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_39; // @[Reg.scala 27:20]
  wire  _T_9373 = _T_4628 ? 1'h0 : ic_tag_valid_out_0_39; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9588 = _T_9587 | _T_9373; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_40; // @[Reg.scala 27:20]
  wire  _T_9375 = _T_4632 ? 1'h0 : ic_tag_valid_out_0_40; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9589 = _T_9588 | _T_9375; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_41; // @[Reg.scala 27:20]
  wire  _T_9377 = _T_4636 ? 1'h0 : ic_tag_valid_out_0_41; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9590 = _T_9589 | _T_9377; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_42; // @[Reg.scala 27:20]
  wire  _T_9379 = _T_4640 ? 1'h0 : ic_tag_valid_out_0_42; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9591 = _T_9590 | _T_9379; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_43; // @[Reg.scala 27:20]
  wire  _T_9381 = _T_4644 ? 1'h0 : ic_tag_valid_out_0_43; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9592 = _T_9591 | _T_9381; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_44; // @[Reg.scala 27:20]
  wire  _T_9383 = _T_4648 ? 1'h0 : ic_tag_valid_out_0_44; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9593 = _T_9592 | _T_9383; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_45; // @[Reg.scala 27:20]
  wire  _T_9385 = _T_4652 ? 1'h0 : ic_tag_valid_out_0_45; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9594 = _T_9593 | _T_9385; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_46; // @[Reg.scala 27:20]
  wire  _T_9387 = _T_4656 ? 1'h0 : ic_tag_valid_out_0_46; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9595 = _T_9594 | _T_9387; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_47; // @[Reg.scala 27:20]
  wire  _T_9389 = _T_4660 ? 1'h0 : ic_tag_valid_out_0_47; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9596 = _T_9595 | _T_9389; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_48; // @[Reg.scala 27:20]
  wire  _T_9391 = _T_4664 ? 1'h0 : ic_tag_valid_out_0_48; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9597 = _T_9596 | _T_9391; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_49; // @[Reg.scala 27:20]
  wire  _T_9393 = _T_4668 ? 1'h0 : ic_tag_valid_out_0_49; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9598 = _T_9597 | _T_9393; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_50; // @[Reg.scala 27:20]
  wire  _T_9395 = _T_4672 ? 1'h0 : ic_tag_valid_out_0_50; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9599 = _T_9598 | _T_9395; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_51; // @[Reg.scala 27:20]
  wire  _T_9397 = _T_4676 ? 1'h0 : ic_tag_valid_out_0_51; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9600 = _T_9599 | _T_9397; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_52; // @[Reg.scala 27:20]
  wire  _T_9399 = _T_4680 ? 1'h0 : ic_tag_valid_out_0_52; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9601 = _T_9600 | _T_9399; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_53; // @[Reg.scala 27:20]
  wire  _T_9401 = _T_4684 ? 1'h0 : ic_tag_valid_out_0_53; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9602 = _T_9601 | _T_9401; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_54; // @[Reg.scala 27:20]
  wire  _T_9403 = _T_4688 ? 1'h0 : ic_tag_valid_out_0_54; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9603 = _T_9602 | _T_9403; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_55; // @[Reg.scala 27:20]
  wire  _T_9405 = _T_4692 ? 1'h0 : ic_tag_valid_out_0_55; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9604 = _T_9603 | _T_9405; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_56; // @[Reg.scala 27:20]
  wire  _T_9407 = _T_4696 ? 1'h0 : ic_tag_valid_out_0_56; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9605 = _T_9604 | _T_9407; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_57; // @[Reg.scala 27:20]
  wire  _T_9409 = _T_4700 ? 1'h0 : ic_tag_valid_out_0_57; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9606 = _T_9605 | _T_9409; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_58; // @[Reg.scala 27:20]
  wire  _T_9411 = _T_4704 ? 1'h0 : ic_tag_valid_out_0_58; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9607 = _T_9606 | _T_9411; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_59; // @[Reg.scala 27:20]
  wire  _T_9413 = _T_4708 ? 1'h0 : ic_tag_valid_out_0_59; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9608 = _T_9607 | _T_9413; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_60; // @[Reg.scala 27:20]
  wire  _T_9415 = _T_4712 ? 1'h0 : ic_tag_valid_out_0_60; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9609 = _T_9608 | _T_9415; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_61; // @[Reg.scala 27:20]
  wire  _T_9417 = _T_4716 ? 1'h0 : ic_tag_valid_out_0_61; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9610 = _T_9609 | _T_9417; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_62; // @[Reg.scala 27:20]
  wire  _T_9419 = _T_4720 ? 1'h0 : ic_tag_valid_out_0_62; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9611 = _T_9610 | _T_9419; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_63; // @[Reg.scala 27:20]
  wire  _T_9421 = _T_4724 ? 1'h0 : ic_tag_valid_out_0_63; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9612 = _T_9611 | _T_9421; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_64; // @[Reg.scala 27:20]
  wire  _T_9423 = _T_4728 ? 1'h0 : ic_tag_valid_out_0_64; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9613 = _T_9612 | _T_9423; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_65; // @[Reg.scala 27:20]
  wire  _T_9425 = _T_4732 ? 1'h0 : ic_tag_valid_out_0_65; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9614 = _T_9613 | _T_9425; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_66; // @[Reg.scala 27:20]
  wire  _T_9427 = _T_4736 ? 1'h0 : ic_tag_valid_out_0_66; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9615 = _T_9614 | _T_9427; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_67; // @[Reg.scala 27:20]
  wire  _T_9429 = _T_4740 ? 1'h0 : ic_tag_valid_out_0_67; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9616 = _T_9615 | _T_9429; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_68; // @[Reg.scala 27:20]
  wire  _T_9431 = _T_4744 ? 1'h0 : ic_tag_valid_out_0_68; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9617 = _T_9616 | _T_9431; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_69; // @[Reg.scala 27:20]
  wire  _T_9433 = _T_4748 ? 1'h0 : ic_tag_valid_out_0_69; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9618 = _T_9617 | _T_9433; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_70; // @[Reg.scala 27:20]
  wire  _T_9435 = _T_4752 ? 1'h0 : ic_tag_valid_out_0_70; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9619 = _T_9618 | _T_9435; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_71; // @[Reg.scala 27:20]
  wire  _T_9437 = _T_4756 ? 1'h0 : ic_tag_valid_out_0_71; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9620 = _T_9619 | _T_9437; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_72; // @[Reg.scala 27:20]
  wire  _T_9439 = _T_4760 ? 1'h0 : ic_tag_valid_out_0_72; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9621 = _T_9620 | _T_9439; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_73; // @[Reg.scala 27:20]
  wire  _T_9441 = _T_4764 ? 1'h0 : ic_tag_valid_out_0_73; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9622 = _T_9621 | _T_9441; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_74; // @[Reg.scala 27:20]
  wire  _T_9443 = _T_4768 ? 1'h0 : ic_tag_valid_out_0_74; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9623 = _T_9622 | _T_9443; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_75; // @[Reg.scala 27:20]
  wire  _T_9445 = _T_4772 ? 1'h0 : ic_tag_valid_out_0_75; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9624 = _T_9623 | _T_9445; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_76; // @[Reg.scala 27:20]
  wire  _T_9447 = _T_4776 ? 1'h0 : ic_tag_valid_out_0_76; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9625 = _T_9624 | _T_9447; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_77; // @[Reg.scala 27:20]
  wire  _T_9449 = _T_4780 ? 1'h0 : ic_tag_valid_out_0_77; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9626 = _T_9625 | _T_9449; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_78; // @[Reg.scala 27:20]
  wire  _T_9451 = _T_4784 ? 1'h0 : ic_tag_valid_out_0_78; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9627 = _T_9626 | _T_9451; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_79; // @[Reg.scala 27:20]
  wire  _T_9453 = _T_4788 ? 1'h0 : ic_tag_valid_out_0_79; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9628 = _T_9627 | _T_9453; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_80; // @[Reg.scala 27:20]
  wire  _T_9455 = _T_4792 ? 1'h0 : ic_tag_valid_out_0_80; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9629 = _T_9628 | _T_9455; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_81; // @[Reg.scala 27:20]
  wire  _T_9457 = _T_4796 ? 1'h0 : ic_tag_valid_out_0_81; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9630 = _T_9629 | _T_9457; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_82; // @[Reg.scala 27:20]
  wire  _T_9459 = _T_4800 ? 1'h0 : ic_tag_valid_out_0_82; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9631 = _T_9630 | _T_9459; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_83; // @[Reg.scala 27:20]
  wire  _T_9461 = _T_4804 ? 1'h0 : ic_tag_valid_out_0_83; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9632 = _T_9631 | _T_9461; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_84; // @[Reg.scala 27:20]
  wire  _T_9463 = _T_4808 ? 1'h0 : ic_tag_valid_out_0_84; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9633 = _T_9632 | _T_9463; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_85; // @[Reg.scala 27:20]
  wire  _T_9465 = _T_4812 ? 1'h0 : ic_tag_valid_out_0_85; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9634 = _T_9633 | _T_9465; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_86; // @[Reg.scala 27:20]
  wire  _T_9467 = _T_4816 ? 1'h0 : ic_tag_valid_out_0_86; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9635 = _T_9634 | _T_9467; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_87; // @[Reg.scala 27:20]
  wire  _T_9469 = _T_4820 ? 1'h0 : ic_tag_valid_out_0_87; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9636 = _T_9635 | _T_9469; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_88; // @[Reg.scala 27:20]
  wire  _T_9471 = _T_4824 ? 1'h0 : ic_tag_valid_out_0_88; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9637 = _T_9636 | _T_9471; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_89; // @[Reg.scala 27:20]
  wire  _T_9473 = _T_4828 ? 1'h0 : ic_tag_valid_out_0_89; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9638 = _T_9637 | _T_9473; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_90; // @[Reg.scala 27:20]
  wire  _T_9475 = _T_4832 ? 1'h0 : ic_tag_valid_out_0_90; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9639 = _T_9638 | _T_9475; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_91; // @[Reg.scala 27:20]
  wire  _T_9477 = _T_4836 ? 1'h0 : ic_tag_valid_out_0_91; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9640 = _T_9639 | _T_9477; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_92; // @[Reg.scala 27:20]
  wire  _T_9479 = _T_4840 ? 1'h0 : ic_tag_valid_out_0_92; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9641 = _T_9640 | _T_9479; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_93; // @[Reg.scala 27:20]
  wire  _T_9481 = _T_4844 ? 1'h0 : ic_tag_valid_out_0_93; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9642 = _T_9641 | _T_9481; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_94; // @[Reg.scala 27:20]
  wire  _T_9483 = _T_4848 ? 1'h0 : ic_tag_valid_out_0_94; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9643 = _T_9642 | _T_9483; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_95; // @[Reg.scala 27:20]
  wire  _T_9485 = _T_4852 ? 1'h0 : ic_tag_valid_out_0_95; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9644 = _T_9643 | _T_9485; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_96; // @[Reg.scala 27:20]
  wire  _T_9487 = _T_4856 ? 1'h0 : ic_tag_valid_out_0_96; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9645 = _T_9644 | _T_9487; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_97; // @[Reg.scala 27:20]
  wire  _T_9489 = _T_4860 ? 1'h0 : ic_tag_valid_out_0_97; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9646 = _T_9645 | _T_9489; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_98; // @[Reg.scala 27:20]
  wire  _T_9491 = _T_4864 ? 1'h0 : ic_tag_valid_out_0_98; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9647 = _T_9646 | _T_9491; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_99; // @[Reg.scala 27:20]
  wire  _T_9493 = _T_4868 ? 1'h0 : ic_tag_valid_out_0_99; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9648 = _T_9647 | _T_9493; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_100; // @[Reg.scala 27:20]
  wire  _T_9495 = _T_4872 ? 1'h0 : ic_tag_valid_out_0_100; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9649 = _T_9648 | _T_9495; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_101; // @[Reg.scala 27:20]
  wire  _T_9497 = _T_4876 ? 1'h0 : ic_tag_valid_out_0_101; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9650 = _T_9649 | _T_9497; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_102; // @[Reg.scala 27:20]
  wire  _T_9499 = _T_4880 ? 1'h0 : ic_tag_valid_out_0_102; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9651 = _T_9650 | _T_9499; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_103; // @[Reg.scala 27:20]
  wire  _T_9501 = _T_4884 ? 1'h0 : ic_tag_valid_out_0_103; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9652 = _T_9651 | _T_9501; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_104; // @[Reg.scala 27:20]
  wire  _T_9503 = _T_4888 ? 1'h0 : ic_tag_valid_out_0_104; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9653 = _T_9652 | _T_9503; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_105; // @[Reg.scala 27:20]
  wire  _T_9505 = _T_4892 ? 1'h0 : ic_tag_valid_out_0_105; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9654 = _T_9653 | _T_9505; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_106; // @[Reg.scala 27:20]
  wire  _T_9507 = _T_4896 ? 1'h0 : ic_tag_valid_out_0_106; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9655 = _T_9654 | _T_9507; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_107; // @[Reg.scala 27:20]
  wire  _T_9509 = _T_4900 ? 1'h0 : ic_tag_valid_out_0_107; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9656 = _T_9655 | _T_9509; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_108; // @[Reg.scala 27:20]
  wire  _T_9511 = _T_4904 ? 1'h0 : ic_tag_valid_out_0_108; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9657 = _T_9656 | _T_9511; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_109; // @[Reg.scala 27:20]
  wire  _T_9513 = _T_4908 ? 1'h0 : ic_tag_valid_out_0_109; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9658 = _T_9657 | _T_9513; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_110; // @[Reg.scala 27:20]
  wire  _T_9515 = _T_4912 ? 1'h0 : ic_tag_valid_out_0_110; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9659 = _T_9658 | _T_9515; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_111; // @[Reg.scala 27:20]
  wire  _T_9517 = _T_4916 ? 1'h0 : ic_tag_valid_out_0_111; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9660 = _T_9659 | _T_9517; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_112; // @[Reg.scala 27:20]
  wire  _T_9519 = _T_4920 ? 1'h0 : ic_tag_valid_out_0_112; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9661 = _T_9660 | _T_9519; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_113; // @[Reg.scala 27:20]
  wire  _T_9521 = _T_4924 ? 1'h0 : ic_tag_valid_out_0_113; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9662 = _T_9661 | _T_9521; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_114; // @[Reg.scala 27:20]
  wire  _T_9523 = _T_4928 ? 1'h0 : ic_tag_valid_out_0_114; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9663 = _T_9662 | _T_9523; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_115; // @[Reg.scala 27:20]
  wire  _T_9525 = _T_4932 ? 1'h0 : ic_tag_valid_out_0_115; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9664 = _T_9663 | _T_9525; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_116; // @[Reg.scala 27:20]
  wire  _T_9527 = _T_4936 ? 1'h0 : ic_tag_valid_out_0_116; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9665 = _T_9664 | _T_9527; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_117; // @[Reg.scala 27:20]
  wire  _T_9529 = _T_4940 ? 1'h0 : ic_tag_valid_out_0_117; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9666 = _T_9665 | _T_9529; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_118; // @[Reg.scala 27:20]
  wire  _T_9531 = _T_4944 ? 1'h0 : ic_tag_valid_out_0_118; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9667 = _T_9666 | _T_9531; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_119; // @[Reg.scala 27:20]
  wire  _T_9533 = _T_4948 ? 1'h0 : ic_tag_valid_out_0_119; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9668 = _T_9667 | _T_9533; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_120; // @[Reg.scala 27:20]
  wire  _T_9535 = _T_4952 ? 1'h0 : ic_tag_valid_out_0_120; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9669 = _T_9668 | _T_9535; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_121; // @[Reg.scala 27:20]
  wire  _T_9537 = _T_4956 ? 1'h0 : ic_tag_valid_out_0_121; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9670 = _T_9669 | _T_9537; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_122; // @[Reg.scala 27:20]
  wire  _T_9539 = _T_4960 ? 1'h0 : ic_tag_valid_out_0_122; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9671 = _T_9670 | _T_9539; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_123; // @[Reg.scala 27:20]
  wire  _T_9541 = _T_4964 ? 1'h0 : ic_tag_valid_out_0_123; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9672 = _T_9671 | _T_9541; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_124; // @[Reg.scala 27:20]
  wire  _T_9543 = _T_4968 ? 1'h0 : ic_tag_valid_out_0_124; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9673 = _T_9672 | _T_9543; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_125; // @[Reg.scala 27:20]
  wire  _T_9545 = _T_4972 ? 1'h0 : ic_tag_valid_out_0_125; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9674 = _T_9673 | _T_9545; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_126; // @[Reg.scala 27:20]
  wire  _T_9547 = _T_4976 ? 1'h0 : ic_tag_valid_out_0_126; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9675 = _T_9674 | _T_9547; // @[el2_ifu_mem_ctl.scala 744:91]
  reg  ic_tag_valid_out_0_127; // @[Reg.scala 27:20]
  wire  _T_9549 = _T_4980 ? 1'h0 : ic_tag_valid_out_0_127; // @[el2_ifu_mem_ctl.scala 744:10]
  wire  _T_9676 = _T_9675 | _T_9549; // @[el2_ifu_mem_ctl.scala 744:91]
  wire [1:0] ic_tag_valid_unq = {_T_10059,_T_9676}; // @[Cat.scala 29:58]
  reg [1:0] ic_debug_way_ff; // @[Reg.scala 27:20]
  reg  ic_debug_rd_en_ff; // @[el2_ifu_mem_ctl.scala 817:54]
  wire [1:0] _T_10098 = ic_debug_rd_en_ff ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [1:0] _T_10099 = ic_debug_way_ff & _T_10098; // @[el2_ifu_mem_ctl.scala 798:67]
  wire [1:0] _T_10100 = ic_tag_valid_unq & _T_10099; // @[el2_ifu_mem_ctl.scala 798:48]
  wire  ic_debug_tag_val_rd_out = |_T_10100; // @[el2_ifu_mem_ctl.scala 798:115]
  wire [65:0] _T_1211 = {2'h0,io_ictag_debug_rd_data[25:21],32'h0,io_ictag_debug_rd_data[20:0],1'h0,way_status,3'h0,ic_debug_tag_val_rd_out}; // @[Cat.scala 29:58]
  reg [70:0] _T_1212; // @[el2_ifu_mem_ctl.scala 348:37]
  wire  ifu_wr_cumulative_err = ifu_wr_cumulative_err_data & _T_2540; // @[el2_ifu_mem_ctl.scala 358:80]
  wire  _T_1252 = ~ifu_byp_data_err_new; // @[el2_ifu_mem_ctl.scala 363:98]
  wire  sel_byp_data = _T_1256 & _T_1252; // @[el2_ifu_mem_ctl.scala 363:96]
  wire [63:0] _T_1263 = fetch_req_iccm_f ? 64'hffffffffffffffff : 64'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_1264 = _T_1263 & io_iccm_rd_data; // @[el2_ifu_mem_ctl.scala 370:64]
  wire [63:0] _T_1266 = sel_byp_data ? 64'hffffffffffffffff : 64'h0; // @[Bitwise.scala 72:12]
  wire  _T_2102 = ~ifu_fetch_addr_int_f[0]; // @[el2_ifu_mem_ctl.scala 439:31]
  wire [3:0] byp_fetch_index_inc_0 = {byp_fetch_index_inc,1'h0}; // @[Cat.scala 29:58]
  wire  _T_1616 = byp_fetch_index_inc_0 == 4'h0; // @[el2_ifu_mem_ctl.scala 436:73]
  wire [15:0] _T_1664 = _T_1616 ? ic_miss_buff_data_0[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire  _T_1619 = byp_fetch_index_inc_0 == 4'h1; // @[el2_ifu_mem_ctl.scala 436:73]
  wire [15:0] _T_1665 = _T_1619 ? ic_miss_buff_data_1[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1680 = _T_1664 | _T_1665; // @[Mux.scala 27:72]
  wire  _T_1622 = byp_fetch_index_inc_0 == 4'h2; // @[el2_ifu_mem_ctl.scala 436:73]
  wire [15:0] _T_1666 = _T_1622 ? ic_miss_buff_data_2[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1681 = _T_1680 | _T_1666; // @[Mux.scala 27:72]
  wire  _T_1625 = byp_fetch_index_inc_0 == 4'h3; // @[el2_ifu_mem_ctl.scala 436:73]
  wire [15:0] _T_1667 = _T_1625 ? ic_miss_buff_data_3[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1682 = _T_1681 | _T_1667; // @[Mux.scala 27:72]
  wire  _T_1628 = byp_fetch_index_inc_0 == 4'h4; // @[el2_ifu_mem_ctl.scala 436:73]
  wire [15:0] _T_1668 = _T_1628 ? ic_miss_buff_data_4[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1683 = _T_1682 | _T_1668; // @[Mux.scala 27:72]
  wire  _T_1631 = byp_fetch_index_inc_0 == 4'h5; // @[el2_ifu_mem_ctl.scala 436:73]
  wire [15:0] _T_1669 = _T_1631 ? ic_miss_buff_data_5[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1684 = _T_1683 | _T_1669; // @[Mux.scala 27:72]
  wire  _T_1634 = byp_fetch_index_inc_0 == 4'h6; // @[el2_ifu_mem_ctl.scala 436:73]
  wire [15:0] _T_1670 = _T_1634 ? ic_miss_buff_data_6[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1685 = _T_1684 | _T_1670; // @[Mux.scala 27:72]
  wire  _T_1637 = byp_fetch_index_inc_0 == 4'h7; // @[el2_ifu_mem_ctl.scala 436:73]
  wire [15:0] _T_1671 = _T_1637 ? ic_miss_buff_data_7[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1686 = _T_1685 | _T_1671; // @[Mux.scala 27:72]
  wire  _T_1640 = byp_fetch_index_inc_0 == 4'h8; // @[el2_ifu_mem_ctl.scala 436:73]
  wire [15:0] _T_1672 = _T_1640 ? ic_miss_buff_data_8[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1687 = _T_1686 | _T_1672; // @[Mux.scala 27:72]
  wire  _T_1643 = byp_fetch_index_inc_0 == 4'h9; // @[el2_ifu_mem_ctl.scala 436:73]
  wire [15:0] _T_1673 = _T_1643 ? ic_miss_buff_data_9[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1688 = _T_1687 | _T_1673; // @[Mux.scala 27:72]
  wire  _T_1646 = byp_fetch_index_inc_0 == 4'ha; // @[el2_ifu_mem_ctl.scala 436:73]
  wire [15:0] _T_1674 = _T_1646 ? ic_miss_buff_data_10[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1689 = _T_1688 | _T_1674; // @[Mux.scala 27:72]
  wire  _T_1649 = byp_fetch_index_inc_0 == 4'hb; // @[el2_ifu_mem_ctl.scala 436:73]
  wire [15:0] _T_1675 = _T_1649 ? ic_miss_buff_data_11[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1690 = _T_1689 | _T_1675; // @[Mux.scala 27:72]
  wire  _T_1652 = byp_fetch_index_inc_0 == 4'hc; // @[el2_ifu_mem_ctl.scala 436:73]
  wire [15:0] _T_1676 = _T_1652 ? ic_miss_buff_data_12[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1691 = _T_1690 | _T_1676; // @[Mux.scala 27:72]
  wire  _T_1655 = byp_fetch_index_inc_0 == 4'hd; // @[el2_ifu_mem_ctl.scala 436:73]
  wire [15:0] _T_1677 = _T_1655 ? ic_miss_buff_data_13[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1692 = _T_1691 | _T_1677; // @[Mux.scala 27:72]
  wire  _T_1658 = byp_fetch_index_inc_0 == 4'he; // @[el2_ifu_mem_ctl.scala 436:73]
  wire [15:0] _T_1678 = _T_1658 ? ic_miss_buff_data_14[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1693 = _T_1692 | _T_1678; // @[Mux.scala 27:72]
  wire  _T_1661 = byp_fetch_index_inc_0 == 4'hf; // @[el2_ifu_mem_ctl.scala 436:73]
  wire [15:0] _T_1679 = _T_1661 ? ic_miss_buff_data_15[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1694 = _T_1693 | _T_1679; // @[Mux.scala 27:72]
  wire [3:0] byp_fetch_index_1 = {ifu_fetch_addr_int_f[4:2],1'h1}; // @[Cat.scala 29:58]
  wire  _T_1696 = byp_fetch_index_1 == 4'h0; // @[el2_ifu_mem_ctl.scala 436:179]
  wire [31:0] _T_1744 = _T_1696 ? ic_miss_buff_data_0 : 32'h0; // @[Mux.scala 27:72]
  wire  _T_1699 = byp_fetch_index_1 == 4'h1; // @[el2_ifu_mem_ctl.scala 436:179]
  wire [31:0] _T_1745 = _T_1699 ? ic_miss_buff_data_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1760 = _T_1744 | _T_1745; // @[Mux.scala 27:72]
  wire  _T_1702 = byp_fetch_index_1 == 4'h2; // @[el2_ifu_mem_ctl.scala 436:179]
  wire [31:0] _T_1746 = _T_1702 ? ic_miss_buff_data_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1761 = _T_1760 | _T_1746; // @[Mux.scala 27:72]
  wire  _T_1705 = byp_fetch_index_1 == 4'h3; // @[el2_ifu_mem_ctl.scala 436:179]
  wire [31:0] _T_1747 = _T_1705 ? ic_miss_buff_data_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1762 = _T_1761 | _T_1747; // @[Mux.scala 27:72]
  wire  _T_1708 = byp_fetch_index_1 == 4'h4; // @[el2_ifu_mem_ctl.scala 436:179]
  wire [31:0] _T_1748 = _T_1708 ? ic_miss_buff_data_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1763 = _T_1762 | _T_1748; // @[Mux.scala 27:72]
  wire  _T_1711 = byp_fetch_index_1 == 4'h5; // @[el2_ifu_mem_ctl.scala 436:179]
  wire [31:0] _T_1749 = _T_1711 ? ic_miss_buff_data_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1764 = _T_1763 | _T_1749; // @[Mux.scala 27:72]
  wire  _T_1714 = byp_fetch_index_1 == 4'h6; // @[el2_ifu_mem_ctl.scala 436:179]
  wire [31:0] _T_1750 = _T_1714 ? ic_miss_buff_data_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1765 = _T_1764 | _T_1750; // @[Mux.scala 27:72]
  wire  _T_1717 = byp_fetch_index_1 == 4'h7; // @[el2_ifu_mem_ctl.scala 436:179]
  wire [31:0] _T_1751 = _T_1717 ? ic_miss_buff_data_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1766 = _T_1765 | _T_1751; // @[Mux.scala 27:72]
  wire  _T_1720 = byp_fetch_index_1 == 4'h8; // @[el2_ifu_mem_ctl.scala 436:179]
  wire [31:0] _T_1752 = _T_1720 ? ic_miss_buff_data_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1767 = _T_1766 | _T_1752; // @[Mux.scala 27:72]
  wire  _T_1723 = byp_fetch_index_1 == 4'h9; // @[el2_ifu_mem_ctl.scala 436:179]
  wire [31:0] _T_1753 = _T_1723 ? ic_miss_buff_data_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1768 = _T_1767 | _T_1753; // @[Mux.scala 27:72]
  wire  _T_1726 = byp_fetch_index_1 == 4'ha; // @[el2_ifu_mem_ctl.scala 436:179]
  wire [31:0] _T_1754 = _T_1726 ? ic_miss_buff_data_10 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1769 = _T_1768 | _T_1754; // @[Mux.scala 27:72]
  wire  _T_1729 = byp_fetch_index_1 == 4'hb; // @[el2_ifu_mem_ctl.scala 436:179]
  wire [31:0] _T_1755 = _T_1729 ? ic_miss_buff_data_11 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1770 = _T_1769 | _T_1755; // @[Mux.scala 27:72]
  wire  _T_1732 = byp_fetch_index_1 == 4'hc; // @[el2_ifu_mem_ctl.scala 436:179]
  wire [31:0] _T_1756 = _T_1732 ? ic_miss_buff_data_12 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1771 = _T_1770 | _T_1756; // @[Mux.scala 27:72]
  wire  _T_1735 = byp_fetch_index_1 == 4'hd; // @[el2_ifu_mem_ctl.scala 436:179]
  wire [31:0] _T_1757 = _T_1735 ? ic_miss_buff_data_13 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1772 = _T_1771 | _T_1757; // @[Mux.scala 27:72]
  wire  _T_1738 = byp_fetch_index_1 == 4'he; // @[el2_ifu_mem_ctl.scala 436:179]
  wire [31:0] _T_1758 = _T_1738 ? ic_miss_buff_data_14 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1773 = _T_1772 | _T_1758; // @[Mux.scala 27:72]
  wire  _T_1741 = byp_fetch_index_1 == 4'hf; // @[el2_ifu_mem_ctl.scala 436:179]
  wire [31:0] _T_1759 = _T_1741 ? ic_miss_buff_data_15 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1774 = _T_1773 | _T_1759; // @[Mux.scala 27:72]
  wire [3:0] byp_fetch_index_0 = {ifu_fetch_addr_int_f[4:2],1'h0}; // @[Cat.scala 29:58]
  wire  _T_1776 = byp_fetch_index_0 == 4'h0; // @[el2_ifu_mem_ctl.scala 436:285]
  wire [31:0] _T_1824 = _T_1776 ? ic_miss_buff_data_0 : 32'h0; // @[Mux.scala 27:72]
  wire  _T_1779 = byp_fetch_index_0 == 4'h1; // @[el2_ifu_mem_ctl.scala 436:285]
  wire [31:0] _T_1825 = _T_1779 ? ic_miss_buff_data_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1840 = _T_1824 | _T_1825; // @[Mux.scala 27:72]
  wire  _T_1782 = byp_fetch_index_0 == 4'h2; // @[el2_ifu_mem_ctl.scala 436:285]
  wire [31:0] _T_1826 = _T_1782 ? ic_miss_buff_data_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1841 = _T_1840 | _T_1826; // @[Mux.scala 27:72]
  wire  _T_1785 = byp_fetch_index_0 == 4'h3; // @[el2_ifu_mem_ctl.scala 436:285]
  wire [31:0] _T_1827 = _T_1785 ? ic_miss_buff_data_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1842 = _T_1841 | _T_1827; // @[Mux.scala 27:72]
  wire  _T_1788 = byp_fetch_index_0 == 4'h4; // @[el2_ifu_mem_ctl.scala 436:285]
  wire [31:0] _T_1828 = _T_1788 ? ic_miss_buff_data_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1843 = _T_1842 | _T_1828; // @[Mux.scala 27:72]
  wire  _T_1791 = byp_fetch_index_0 == 4'h5; // @[el2_ifu_mem_ctl.scala 436:285]
  wire [31:0] _T_1829 = _T_1791 ? ic_miss_buff_data_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1844 = _T_1843 | _T_1829; // @[Mux.scala 27:72]
  wire  _T_1794 = byp_fetch_index_0 == 4'h6; // @[el2_ifu_mem_ctl.scala 436:285]
  wire [31:0] _T_1830 = _T_1794 ? ic_miss_buff_data_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1845 = _T_1844 | _T_1830; // @[Mux.scala 27:72]
  wire  _T_1797 = byp_fetch_index_0 == 4'h7; // @[el2_ifu_mem_ctl.scala 436:285]
  wire [31:0] _T_1831 = _T_1797 ? ic_miss_buff_data_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1846 = _T_1845 | _T_1831; // @[Mux.scala 27:72]
  wire  _T_1800 = byp_fetch_index_0 == 4'h8; // @[el2_ifu_mem_ctl.scala 436:285]
  wire [31:0] _T_1832 = _T_1800 ? ic_miss_buff_data_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1847 = _T_1846 | _T_1832; // @[Mux.scala 27:72]
  wire  _T_1803 = byp_fetch_index_0 == 4'h9; // @[el2_ifu_mem_ctl.scala 436:285]
  wire [31:0] _T_1833 = _T_1803 ? ic_miss_buff_data_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1848 = _T_1847 | _T_1833; // @[Mux.scala 27:72]
  wire  _T_1806 = byp_fetch_index_0 == 4'ha; // @[el2_ifu_mem_ctl.scala 436:285]
  wire [31:0] _T_1834 = _T_1806 ? ic_miss_buff_data_10 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1849 = _T_1848 | _T_1834; // @[Mux.scala 27:72]
  wire  _T_1809 = byp_fetch_index_0 == 4'hb; // @[el2_ifu_mem_ctl.scala 436:285]
  wire [31:0] _T_1835 = _T_1809 ? ic_miss_buff_data_11 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1850 = _T_1849 | _T_1835; // @[Mux.scala 27:72]
  wire  _T_1812 = byp_fetch_index_0 == 4'hc; // @[el2_ifu_mem_ctl.scala 436:285]
  wire [31:0] _T_1836 = _T_1812 ? ic_miss_buff_data_12 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1851 = _T_1850 | _T_1836; // @[Mux.scala 27:72]
  wire  _T_1815 = byp_fetch_index_0 == 4'hd; // @[el2_ifu_mem_ctl.scala 436:285]
  wire [31:0] _T_1837 = _T_1815 ? ic_miss_buff_data_13 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1852 = _T_1851 | _T_1837; // @[Mux.scala 27:72]
  wire  _T_1818 = byp_fetch_index_0 == 4'he; // @[el2_ifu_mem_ctl.scala 436:285]
  wire [31:0] _T_1838 = _T_1818 ? ic_miss_buff_data_14 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1853 = _T_1852 | _T_1838; // @[Mux.scala 27:72]
  wire  _T_1821 = byp_fetch_index_0 == 4'hf; // @[el2_ifu_mem_ctl.scala 436:285]
  wire [31:0] _T_1839 = _T_1821 ? ic_miss_buff_data_15 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1854 = _T_1853 | _T_1839; // @[Mux.scala 27:72]
  wire [79:0] _T_1857 = {_T_1694,_T_1774,_T_1854}; // @[Cat.scala 29:58]
  wire [3:0] byp_fetch_index_inc_1 = {byp_fetch_index_inc,1'h1}; // @[Cat.scala 29:58]
  wire  _T_1858 = byp_fetch_index_inc_1 == 4'h0; // @[el2_ifu_mem_ctl.scala 437:73]
  wire [15:0] _T_1906 = _T_1858 ? ic_miss_buff_data_0[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire  _T_1861 = byp_fetch_index_inc_1 == 4'h1; // @[el2_ifu_mem_ctl.scala 437:73]
  wire [15:0] _T_1907 = _T_1861 ? ic_miss_buff_data_1[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1922 = _T_1906 | _T_1907; // @[Mux.scala 27:72]
  wire  _T_1864 = byp_fetch_index_inc_1 == 4'h2; // @[el2_ifu_mem_ctl.scala 437:73]
  wire [15:0] _T_1908 = _T_1864 ? ic_miss_buff_data_2[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1923 = _T_1922 | _T_1908; // @[Mux.scala 27:72]
  wire  _T_1867 = byp_fetch_index_inc_1 == 4'h3; // @[el2_ifu_mem_ctl.scala 437:73]
  wire [15:0] _T_1909 = _T_1867 ? ic_miss_buff_data_3[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1924 = _T_1923 | _T_1909; // @[Mux.scala 27:72]
  wire  _T_1870 = byp_fetch_index_inc_1 == 4'h4; // @[el2_ifu_mem_ctl.scala 437:73]
  wire [15:0] _T_1910 = _T_1870 ? ic_miss_buff_data_4[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1925 = _T_1924 | _T_1910; // @[Mux.scala 27:72]
  wire  _T_1873 = byp_fetch_index_inc_1 == 4'h5; // @[el2_ifu_mem_ctl.scala 437:73]
  wire [15:0] _T_1911 = _T_1873 ? ic_miss_buff_data_5[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1926 = _T_1925 | _T_1911; // @[Mux.scala 27:72]
  wire  _T_1876 = byp_fetch_index_inc_1 == 4'h6; // @[el2_ifu_mem_ctl.scala 437:73]
  wire [15:0] _T_1912 = _T_1876 ? ic_miss_buff_data_6[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1927 = _T_1926 | _T_1912; // @[Mux.scala 27:72]
  wire  _T_1879 = byp_fetch_index_inc_1 == 4'h7; // @[el2_ifu_mem_ctl.scala 437:73]
  wire [15:0] _T_1913 = _T_1879 ? ic_miss_buff_data_7[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1928 = _T_1927 | _T_1913; // @[Mux.scala 27:72]
  wire  _T_1882 = byp_fetch_index_inc_1 == 4'h8; // @[el2_ifu_mem_ctl.scala 437:73]
  wire [15:0] _T_1914 = _T_1882 ? ic_miss_buff_data_8[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1929 = _T_1928 | _T_1914; // @[Mux.scala 27:72]
  wire  _T_1885 = byp_fetch_index_inc_1 == 4'h9; // @[el2_ifu_mem_ctl.scala 437:73]
  wire [15:0] _T_1915 = _T_1885 ? ic_miss_buff_data_9[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1930 = _T_1929 | _T_1915; // @[Mux.scala 27:72]
  wire  _T_1888 = byp_fetch_index_inc_1 == 4'ha; // @[el2_ifu_mem_ctl.scala 437:73]
  wire [15:0] _T_1916 = _T_1888 ? ic_miss_buff_data_10[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1931 = _T_1930 | _T_1916; // @[Mux.scala 27:72]
  wire  _T_1891 = byp_fetch_index_inc_1 == 4'hb; // @[el2_ifu_mem_ctl.scala 437:73]
  wire [15:0] _T_1917 = _T_1891 ? ic_miss_buff_data_11[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1932 = _T_1931 | _T_1917; // @[Mux.scala 27:72]
  wire  _T_1894 = byp_fetch_index_inc_1 == 4'hc; // @[el2_ifu_mem_ctl.scala 437:73]
  wire [15:0] _T_1918 = _T_1894 ? ic_miss_buff_data_12[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1933 = _T_1932 | _T_1918; // @[Mux.scala 27:72]
  wire  _T_1897 = byp_fetch_index_inc_1 == 4'hd; // @[el2_ifu_mem_ctl.scala 437:73]
  wire [15:0] _T_1919 = _T_1897 ? ic_miss_buff_data_13[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1934 = _T_1933 | _T_1919; // @[Mux.scala 27:72]
  wire  _T_1900 = byp_fetch_index_inc_1 == 4'he; // @[el2_ifu_mem_ctl.scala 437:73]
  wire [15:0] _T_1920 = _T_1900 ? ic_miss_buff_data_14[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1935 = _T_1934 | _T_1920; // @[Mux.scala 27:72]
  wire  _T_1903 = byp_fetch_index_inc_1 == 4'hf; // @[el2_ifu_mem_ctl.scala 437:73]
  wire [15:0] _T_1921 = _T_1903 ? ic_miss_buff_data_15[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1936 = _T_1935 | _T_1921; // @[Mux.scala 27:72]
  wire [31:0] _T_1986 = _T_1616 ? ic_miss_buff_data_0 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1987 = _T_1619 ? ic_miss_buff_data_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2002 = _T_1986 | _T_1987; // @[Mux.scala 27:72]
  wire [31:0] _T_1988 = _T_1622 ? ic_miss_buff_data_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2003 = _T_2002 | _T_1988; // @[Mux.scala 27:72]
  wire [31:0] _T_1989 = _T_1625 ? ic_miss_buff_data_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2004 = _T_2003 | _T_1989; // @[Mux.scala 27:72]
  wire [31:0] _T_1990 = _T_1628 ? ic_miss_buff_data_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2005 = _T_2004 | _T_1990; // @[Mux.scala 27:72]
  wire [31:0] _T_1991 = _T_1631 ? ic_miss_buff_data_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2006 = _T_2005 | _T_1991; // @[Mux.scala 27:72]
  wire [31:0] _T_1992 = _T_1634 ? ic_miss_buff_data_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2007 = _T_2006 | _T_1992; // @[Mux.scala 27:72]
  wire [31:0] _T_1993 = _T_1637 ? ic_miss_buff_data_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2008 = _T_2007 | _T_1993; // @[Mux.scala 27:72]
  wire [31:0] _T_1994 = _T_1640 ? ic_miss_buff_data_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2009 = _T_2008 | _T_1994; // @[Mux.scala 27:72]
  wire [31:0] _T_1995 = _T_1643 ? ic_miss_buff_data_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2010 = _T_2009 | _T_1995; // @[Mux.scala 27:72]
  wire [31:0] _T_1996 = _T_1646 ? ic_miss_buff_data_10 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2011 = _T_2010 | _T_1996; // @[Mux.scala 27:72]
  wire [31:0] _T_1997 = _T_1649 ? ic_miss_buff_data_11 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2012 = _T_2011 | _T_1997; // @[Mux.scala 27:72]
  wire [31:0] _T_1998 = _T_1652 ? ic_miss_buff_data_12 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2013 = _T_2012 | _T_1998; // @[Mux.scala 27:72]
  wire [31:0] _T_1999 = _T_1655 ? ic_miss_buff_data_13 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2014 = _T_2013 | _T_1999; // @[Mux.scala 27:72]
  wire [31:0] _T_2000 = _T_1658 ? ic_miss_buff_data_14 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2015 = _T_2014 | _T_2000; // @[Mux.scala 27:72]
  wire [31:0] _T_2001 = _T_1661 ? ic_miss_buff_data_15 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2016 = _T_2015 | _T_2001; // @[Mux.scala 27:72]
  wire [79:0] _T_2099 = {_T_1936,_T_2016,_T_1774}; // @[Cat.scala 29:58]
  wire [79:0] ic_byp_data_only_pre_new = _T_2102 ? _T_1857 : _T_2099; // @[el2_ifu_mem_ctl.scala 435:37]
  wire [79:0] _T_2104 = {16'h0,ic_byp_data_only_pre_new[79:16]}; // @[Cat.scala 29:58]
  wire [79:0] ic_byp_data_only_new = _T_2102 ? ic_byp_data_only_pre_new : _T_2104; // @[el2_ifu_mem_ctl.scala 439:30]
  wire [79:0] _GEN_793 = {{16'd0}, _T_1266}; // @[el2_ifu_mem_ctl.scala 370:109]
  wire [79:0] _T_1267 = _GEN_793 & ic_byp_data_only_new; // @[el2_ifu_mem_ctl.scala 370:109]
  wire [79:0] _GEN_794 = {{16'd0}, _T_1264}; // @[el2_ifu_mem_ctl.scala 370:83]
  wire [79:0] ic_premux_data = _GEN_794 | _T_1267; // @[el2_ifu_mem_ctl.scala 370:83]
  wire  fetch_req_f_qual = io_ic_hit_f & _T_318; // @[el2_ifu_mem_ctl.scala 377:38]
  wire [1:0] _T_1276 = ifc_region_acc_fault_f ? 2'h2 : 2'h0; // @[el2_ifu_mem_ctl.scala 381:8]
  wire [7:0] _T_1357 = {ic_miss_buff_data_valid_in_7,ic_miss_buff_data_valid_in_6,ic_miss_buff_data_valid_in_5,ic_miss_buff_data_valid_in_4,ic_miss_buff_data_valid_in_3,ic_miss_buff_data_valid_in_2,ic_miss_buff_data_valid_in_1,ic_miss_buff_data_valid_in_0}; // @[Cat.scala 29:58]
  wire  _T_1362 = ic_miss_buff_data_error[0] & _T_1328; // @[el2_ifu_mem_ctl.scala 402:32]
  wire  _T_2608 = |io_ifu_axi_rresp; // @[el2_ifu_mem_ctl.scala 613:47]
  wire  _T_2609 = _T_2608 & _T_13; // @[el2_ifu_mem_ctl.scala 613:50]
  wire  bus_ifu_wr_data_error = _T_2609 & miss_pending; // @[el2_ifu_mem_ctl.scala 613:68]
  wire  ic_miss_buff_data_error_in_0 = write_fill_data_0 ? bus_ifu_wr_data_error : _T_1362; // @[el2_ifu_mem_ctl.scala 401:72]
  wire  _T_1366 = ic_miss_buff_data_error[1] & _T_1328; // @[el2_ifu_mem_ctl.scala 402:32]
  wire  ic_miss_buff_data_error_in_1 = write_fill_data_1 ? bus_ifu_wr_data_error : _T_1366; // @[el2_ifu_mem_ctl.scala 401:72]
  wire  _T_1370 = ic_miss_buff_data_error[2] & _T_1328; // @[el2_ifu_mem_ctl.scala 402:32]
  wire  ic_miss_buff_data_error_in_2 = write_fill_data_2 ? bus_ifu_wr_data_error : _T_1370; // @[el2_ifu_mem_ctl.scala 401:72]
  wire  _T_1374 = ic_miss_buff_data_error[3] & _T_1328; // @[el2_ifu_mem_ctl.scala 402:32]
  wire  ic_miss_buff_data_error_in_3 = write_fill_data_3 ? bus_ifu_wr_data_error : _T_1374; // @[el2_ifu_mem_ctl.scala 401:72]
  wire  _T_1378 = ic_miss_buff_data_error[4] & _T_1328; // @[el2_ifu_mem_ctl.scala 402:32]
  wire  ic_miss_buff_data_error_in_4 = write_fill_data_4 ? bus_ifu_wr_data_error : _T_1378; // @[el2_ifu_mem_ctl.scala 401:72]
  wire  _T_1382 = ic_miss_buff_data_error[5] & _T_1328; // @[el2_ifu_mem_ctl.scala 402:32]
  wire  ic_miss_buff_data_error_in_5 = write_fill_data_5 ? bus_ifu_wr_data_error : _T_1382; // @[el2_ifu_mem_ctl.scala 401:72]
  wire  _T_1386 = ic_miss_buff_data_error[6] & _T_1328; // @[el2_ifu_mem_ctl.scala 402:32]
  wire  ic_miss_buff_data_error_in_6 = write_fill_data_6 ? bus_ifu_wr_data_error : _T_1386; // @[el2_ifu_mem_ctl.scala 401:72]
  wire  _T_1390 = ic_miss_buff_data_error[7] & _T_1328; // @[el2_ifu_mem_ctl.scala 402:32]
  wire  ic_miss_buff_data_error_in_7 = write_fill_data_7 ? bus_ifu_wr_data_error : _T_1390; // @[el2_ifu_mem_ctl.scala 401:72]
  wire [7:0] _T_1397 = {ic_miss_buff_data_error_in_7,ic_miss_buff_data_error_in_6,ic_miss_buff_data_error_in_5,ic_miss_buff_data_error_in_4,ic_miss_buff_data_error_in_3,ic_miss_buff_data_error_in_2,ic_miss_buff_data_error_in_1,ic_miss_buff_data_error_in_0}; // @[Cat.scala 29:58]
  reg [5:0] perr_ic_index_ff; // @[Reg.scala 27:20]
  wire  _T_2414 = 3'h0 == perr_state; // @[Conditional.scala 37:30]
  wire  _T_2422 = _T_6 & _T_318; // @[el2_ifu_mem_ctl.scala 482:65]
  wire  _T_2423 = _T_2422 | io_iccm_dma_sb_error; // @[el2_ifu_mem_ctl.scala 482:88]
  wire  _T_2425 = _T_2423 & _T_2536; // @[el2_ifu_mem_ctl.scala 482:112]
  wire  _T_2426 = 3'h1 == perr_state; // @[Conditional.scala 37:30]
  wire  _T_2427 = io_dec_tlu_flush_lower_wb | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 487:50]
  wire  _T_2429 = 3'h2 == perr_state; // @[Conditional.scala 37:30]
  wire  _T_2435 = 3'h4 == perr_state; // @[Conditional.scala 37:30]
  wire  _T_2437 = 3'h3 == perr_state; // @[Conditional.scala 37:30]
  wire  _GEN_38 = _T_2435 | _T_2437; // @[Conditional.scala 39:67]
  wire  _GEN_40 = _T_2429 ? _T_2427 : _GEN_38; // @[Conditional.scala 39:67]
  wire  _GEN_42 = _T_2426 ? _T_2427 : _GEN_40; // @[Conditional.scala 39:67]
  wire  perr_state_en = _T_2414 ? _T_2425 : _GEN_42; // @[Conditional.scala 40:58]
  wire  perr_sb_write_status = _T_2414 & perr_state_en; // @[Conditional.scala 40:58]
  wire  _T_2428 = io_dec_tlu_flush_lower_wb & io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 488:56]
  wire  _GEN_43 = _T_2426 & _T_2428; // @[Conditional.scala 39:67]
  wire  perr_sel_invalidate = _T_2414 ? 1'h0 : _GEN_43; // @[Conditional.scala 40:58]
  wire [1:0] perr_err_inv_way = perr_sel_invalidate ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  reg  dma_sb_err_state_ff; // @[el2_ifu_mem_ctl.scala 473:58]
  wire  _T_2411 = ~dma_sb_err_state_ff; // @[el2_ifu_mem_ctl.scala 472:49]
  wire  _T_2416 = io_ic_error_start & _T_318; // @[el2_ifu_mem_ctl.scala 481:87]
  wire  _T_2430 = io_dec_tlu_flush_err_wb & io_dec_tlu_flush_lower_wb; // @[el2_ifu_mem_ctl.scala 491:54]
  wire  _T_2431 = _T_2430 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 491:84]
  wire  _T_2440 = perr_state == 3'h2; // @[el2_ifu_mem_ctl.scala 512:66]
  wire  _T_2441 = io_dec_tlu_flush_err_wb & _T_2440; // @[el2_ifu_mem_ctl.scala 512:52]
  wire  _T_2443 = _T_2441 & _T_2536; // @[el2_ifu_mem_ctl.scala 512:81]
  wire  _T_2445 = io_dec_tlu_flush_lower_wb | io_dec_tlu_i0_commit_cmt; // @[el2_ifu_mem_ctl.scala 515:59]
  wire  _T_2446 = _T_2445 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 515:86]
  wire  _T_2460 = _T_2445 | io_ifu_fetch_val[0]; // @[el2_ifu_mem_ctl.scala 518:81]
  wire  _T_2461 = _T_2460 | ifu_bp_hit_taken_q_f; // @[el2_ifu_mem_ctl.scala 518:103]
  wire  _T_2462 = _T_2461 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 518:126]
  wire  _T_2482 = _T_2460 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 525:103]
  wire  _T_2489 = ~io_dec_tlu_flush_err_wb; // @[el2_ifu_mem_ctl.scala 530:62]
  wire  _T_2490 = io_dec_tlu_flush_lower_wb & _T_2489; // @[el2_ifu_mem_ctl.scala 530:60]
  wire  _T_2491 = _T_2490 | io_dec_tlu_i0_commit_cmt; // @[el2_ifu_mem_ctl.scala 530:88]
  wire  _T_2492 = _T_2491 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 530:115]
  wire  _GEN_50 = _T_2488 & _T_2446; // @[Conditional.scala 39:67]
  wire  _GEN_53 = _T_2471 ? _T_2482 : _GEN_50; // @[Conditional.scala 39:67]
  wire  _GEN_55 = _T_2471 | _T_2488; // @[Conditional.scala 39:67]
  wire  _GEN_57 = _T_2444 ? _T_2462 : _GEN_53; // @[Conditional.scala 39:67]
  wire  _GEN_59 = _T_2444 | _GEN_55; // @[Conditional.scala 39:67]
  wire  err_stop_state_en = _T_2439 ? _T_2443 : _GEN_57; // @[Conditional.scala 40:58]
  reg  ifu_bus_cmd_valid; // @[Reg.scala 27:20]
  wire  _T_2504 = ic_act_miss_f | ifu_bus_cmd_valid; // @[el2_ifu_mem_ctl.scala 547:64]
  wire  _T_2506 = _T_2504 & _T_2536; // @[el2_ifu_mem_ctl.scala 547:85]
  reg [2:0] bus_cmd_beat_count; // @[Reg.scala 27:20]
  wire  _T_2508 = bus_cmd_beat_count == 3'h7; // @[el2_ifu_mem_ctl.scala 547:133]
  wire  _T_2509 = _T_2508 & ifu_bus_cmd_valid; // @[el2_ifu_mem_ctl.scala 547:164]
  wire  _T_2510 = _T_2509 & io_ifu_axi_arready; // @[el2_ifu_mem_ctl.scala 547:184]
  wire  _T_2511 = _T_2510 & miss_pending; // @[el2_ifu_mem_ctl.scala 547:204]
  wire  _T_2512 = ~_T_2511; // @[el2_ifu_mem_ctl.scala 547:112]
  wire  ifc_bus_ic_req_ff_in = _T_2506 & _T_2512; // @[el2_ifu_mem_ctl.scala 547:110]
  wire  _T_2513 = io_ifu_bus_clk_en | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 548:80]
  wire  ifu_bus_arready = io_ifu_axi_arready & io_ifu_bus_clk_en; // @[el2_ifu_mem_ctl.scala 579:45]
  wire  _T_2530 = io_ifu_axi_arvalid & ifu_bus_arready; // @[el2_ifu_mem_ctl.scala 582:35]
  wire  _T_2531 = _T_2530 & miss_pending; // @[el2_ifu_mem_ctl.scala 582:53]
  wire  bus_cmd_sent = _T_2531 & _T_2536; // @[el2_ifu_mem_ctl.scala 582:68]
  wire [2:0] _T_2521 = ifu_bus_cmd_valid ? 3'h7 : 3'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_2523 = {miss_addr,bus_rd_addr_count,3'h0}; // @[Cat.scala 29:58]
  wire [31:0] _T_2525 = ifu_bus_cmd_valid ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  reg  ifu_bus_arready_unq_ff; // @[Reg.scala 27:20]
  reg  ifu_bus_arvalid_ff; // @[Reg.scala 27:20]
  wire  ifu_bus_arready_ff = ifu_bus_arready_unq_ff & bus_ifu_bus_clk_en_ff; // @[el2_ifu_mem_ctl.scala 580:51]
  wire  _T_2551 = ~scnd_miss_req; // @[el2_ifu_mem_ctl.scala 590:73]
  wire  _T_2552 = _T_2537 & _T_2551; // @[el2_ifu_mem_ctl.scala 590:71]
  wire  _T_2554 = last_data_recieved_ff & _T_1328; // @[el2_ifu_mem_ctl.scala 590:114]
  wire  last_data_recieved_in = _T_2552 | _T_2554; // @[el2_ifu_mem_ctl.scala 590:89]
  wire [2:0] _T_2560 = bus_rd_addr_count + 3'h1; // @[el2_ifu_mem_ctl.scala 595:45]
  wire  _T_2563 = io_ifu_bus_clk_en | ic_act_miss_f; // @[el2_ifu_mem_ctl.scala 596:81]
  wire  _T_2564 = _T_2563 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 596:97]
  wire  _T_2566 = ifu_bus_cmd_valid & io_ifu_axi_arready; // @[el2_ifu_mem_ctl.scala 598:48]
  wire  _T_2567 = _T_2566 & miss_pending; // @[el2_ifu_mem_ctl.scala 598:68]
  wire  bus_inc_cmd_beat_cnt = _T_2567 & _T_2536; // @[el2_ifu_mem_ctl.scala 598:83]
  wire  bus_reset_cmd_beat_cnt_secondlast = ic_act_miss_f & uncacheable_miss_in; // @[el2_ifu_mem_ctl.scala 600:57]
  wire  _T_2571 = ~bus_inc_cmd_beat_cnt; // @[el2_ifu_mem_ctl.scala 601:31]
  wire  _T_2572 = ic_act_miss_f | scnd_miss_req; // @[el2_ifu_mem_ctl.scala 601:71]
  wire  _T_2573 = _T_2572 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 601:87]
  wire  _T_2574 = ~_T_2573; // @[el2_ifu_mem_ctl.scala 601:55]
  wire  bus_hold_cmd_beat_cnt = _T_2571 & _T_2574; // @[el2_ifu_mem_ctl.scala 601:53]
  wire  _T_2575 = bus_inc_cmd_beat_cnt | ic_act_miss_f; // @[el2_ifu_mem_ctl.scala 602:46]
  wire  bus_cmd_beat_en = _T_2575 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 602:62]
  wire [2:0] _T_2578 = bus_cmd_beat_count + 3'h1; // @[el2_ifu_mem_ctl.scala 604:46]
  wire [2:0] _T_2580 = bus_reset_cmd_beat_cnt_secondlast ? 3'h6 : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_2581 = bus_inc_cmd_beat_cnt ? _T_2578 : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_2582 = bus_hold_cmd_beat_cnt ? bus_cmd_beat_count : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_2584 = _T_2580 | _T_2581; // @[Mux.scala 27:72]
  wire [2:0] bus_new_cmd_beat_count = _T_2584 | _T_2582; // @[Mux.scala 27:72]
  wire  _T_2588 = _T_2564 & bus_cmd_beat_en; // @[el2_ifu_mem_ctl.scala 605:125]
  reg  ifc_dma_access_ok_prev; // @[el2_ifu_mem_ctl.scala 616:62]
  wire  _T_2616 = ~iccm_correct_ecc; // @[el2_ifu_mem_ctl.scala 621:50]
  wire  _T_2617 = io_ifc_dma_access_ok & _T_2616; // @[el2_ifu_mem_ctl.scala 621:47]
  wire  _T_2618 = ~io_iccm_dma_sb_error; // @[el2_ifu_mem_ctl.scala 621:70]
  wire  ifc_dma_access_ok_d = _T_2617 & _T_2618; // @[el2_ifu_mem_ctl.scala 621:68]
  wire  _T_2622 = _T_2617 & ifc_dma_access_ok_prev; // @[el2_ifu_mem_ctl.scala 622:72]
  wire  _T_2623 = perr_state == 3'h0; // @[el2_ifu_mem_ctl.scala 622:111]
  wire  _T_2624 = _T_2622 & _T_2623; // @[el2_ifu_mem_ctl.scala 622:97]
  wire  ifc_dma_access_q_ok = _T_2624 & _T_2618; // @[el2_ifu_mem_ctl.scala 622:127]
  wire  _T_2627 = ifc_dma_access_q_ok & io_dma_iccm_req; // @[el2_ifu_mem_ctl.scala 625:40]
  wire  _T_2628 = _T_2627 & io_dma_mem_write; // @[el2_ifu_mem_ctl.scala 625:58]
  wire  _T_2631 = ~io_dma_mem_write; // @[el2_ifu_mem_ctl.scala 626:60]
  wire  _T_2632 = _T_2627 & _T_2631; // @[el2_ifu_mem_ctl.scala 626:58]
  wire  _T_2633 = io_ifc_iccm_access_bf & io_ifc_fetch_req_bf; // @[el2_ifu_mem_ctl.scala 626:104]
  wire [2:0] _T_2638 = io_dma_iccm_req ? 3'h7 : 3'h0; // @[Bitwise.scala 72:12]
  wire [8:0] _T_2744 = {io_dma_mem_wdata[48],io_dma_mem_wdata[46],io_dma_mem_wdata[44],io_dma_mem_wdata[42],io_dma_mem_wdata[40],io_dma_mem_wdata[38],io_dma_mem_wdata[37],io_dma_mem_wdata[35],io_dma_mem_wdata[33]}; // @[el2_lib.scala 268:22]
  wire [17:0] _T_2753 = {io_dma_mem_wdata[63],io_dma_mem_wdata[62],io_dma_mem_wdata[60],io_dma_mem_wdata[59],io_dma_mem_wdata[57],io_dma_mem_wdata[55],io_dma_mem_wdata[53],io_dma_mem_wdata[52],io_dma_mem_wdata[50],_T_2744}; // @[el2_lib.scala 268:22]
  wire  _T_2754 = ^_T_2753; // @[el2_lib.scala 268:29]
  wire [8:0] _T_2762 = {io_dma_mem_wdata[47],io_dma_mem_wdata[46],io_dma_mem_wdata[43],io_dma_mem_wdata[42],io_dma_mem_wdata[39],io_dma_mem_wdata[38],io_dma_mem_wdata[36],io_dma_mem_wdata[35],io_dma_mem_wdata[32]}; // @[el2_lib.scala 268:39]
  wire [17:0] _T_2771 = {io_dma_mem_wdata[63],io_dma_mem_wdata[61],io_dma_mem_wdata[60],io_dma_mem_wdata[58],io_dma_mem_wdata[57],io_dma_mem_wdata[54],io_dma_mem_wdata[53],io_dma_mem_wdata[51],io_dma_mem_wdata[50],_T_2762}; // @[el2_lib.scala 268:39]
  wire  _T_2772 = ^_T_2771; // @[el2_lib.scala 268:46]
  wire [8:0] _T_2780 = {io_dma_mem_wdata[47],io_dma_mem_wdata[46],io_dma_mem_wdata[41],io_dma_mem_wdata[40],io_dma_mem_wdata[39],io_dma_mem_wdata[38],io_dma_mem_wdata[34],io_dma_mem_wdata[33],io_dma_mem_wdata[32]}; // @[el2_lib.scala 268:56]
  wire [17:0] _T_2789 = {io_dma_mem_wdata[62],io_dma_mem_wdata[61],io_dma_mem_wdata[60],io_dma_mem_wdata[56],io_dma_mem_wdata[55],io_dma_mem_wdata[54],io_dma_mem_wdata[53],io_dma_mem_wdata[49],io_dma_mem_wdata[48],_T_2780}; // @[el2_lib.scala 268:56]
  wire  _T_2790 = ^_T_2789; // @[el2_lib.scala 268:63]
  wire [6:0] _T_2796 = {io_dma_mem_wdata[44],io_dma_mem_wdata[43],io_dma_mem_wdata[42],io_dma_mem_wdata[41],io_dma_mem_wdata[40],io_dma_mem_wdata[39],io_dma_mem_wdata[38]}; // @[el2_lib.scala 268:73]
  wire [14:0] _T_2804 = {io_dma_mem_wdata[59],io_dma_mem_wdata[58],io_dma_mem_wdata[57],io_dma_mem_wdata[56],io_dma_mem_wdata[55],io_dma_mem_wdata[54],io_dma_mem_wdata[53],io_dma_mem_wdata[45],_T_2796}; // @[el2_lib.scala 268:73]
  wire  _T_2805 = ^_T_2804; // @[el2_lib.scala 268:80]
  wire [14:0] _T_2819 = {io_dma_mem_wdata[52],io_dma_mem_wdata[51],io_dma_mem_wdata[50],io_dma_mem_wdata[49],io_dma_mem_wdata[48],io_dma_mem_wdata[47],io_dma_mem_wdata[46],io_dma_mem_wdata[45],_T_2796}; // @[el2_lib.scala 268:90]
  wire  _T_2820 = ^_T_2819; // @[el2_lib.scala 268:97]
  wire [5:0] _T_2825 = {io_dma_mem_wdata[37],io_dma_mem_wdata[36],io_dma_mem_wdata[35],io_dma_mem_wdata[34],io_dma_mem_wdata[33],io_dma_mem_wdata[32]}; // @[el2_lib.scala 268:107]
  wire  _T_2826 = ^_T_2825; // @[el2_lib.scala 268:114]
  wire [5:0] _T_2831 = {_T_2754,_T_2772,_T_2790,_T_2805,_T_2820,_T_2826}; // @[Cat.scala 29:58]
  wire  _T_2832 = ^io_dma_mem_wdata[63:32]; // @[el2_lib.scala 269:13]
  wire  _T_2833 = ^_T_2831; // @[el2_lib.scala 269:23]
  wire  _T_2834 = _T_2832 ^ _T_2833; // @[el2_lib.scala 269:18]
  wire [8:0] _T_2940 = {io_dma_mem_wdata[16],io_dma_mem_wdata[14],io_dma_mem_wdata[12],io_dma_mem_wdata[10],io_dma_mem_wdata[8],io_dma_mem_wdata[6],io_dma_mem_wdata[5],io_dma_mem_wdata[3],io_dma_mem_wdata[1]}; // @[el2_lib.scala 268:22]
  wire [17:0] _T_2949 = {io_dma_mem_wdata[31],io_dma_mem_wdata[30],io_dma_mem_wdata[28],io_dma_mem_wdata[27],io_dma_mem_wdata[25],io_dma_mem_wdata[23],io_dma_mem_wdata[21],io_dma_mem_wdata[20],io_dma_mem_wdata[18],_T_2940}; // @[el2_lib.scala 268:22]
  wire  _T_2950 = ^_T_2949; // @[el2_lib.scala 268:29]
  wire [8:0] _T_2958 = {io_dma_mem_wdata[15],io_dma_mem_wdata[14],io_dma_mem_wdata[11],io_dma_mem_wdata[10],io_dma_mem_wdata[7],io_dma_mem_wdata[6],io_dma_mem_wdata[4],io_dma_mem_wdata[3],io_dma_mem_wdata[0]}; // @[el2_lib.scala 268:39]
  wire [17:0] _T_2967 = {io_dma_mem_wdata[31],io_dma_mem_wdata[29],io_dma_mem_wdata[28],io_dma_mem_wdata[26],io_dma_mem_wdata[25],io_dma_mem_wdata[22],io_dma_mem_wdata[21],io_dma_mem_wdata[19],io_dma_mem_wdata[18],_T_2958}; // @[el2_lib.scala 268:39]
  wire  _T_2968 = ^_T_2967; // @[el2_lib.scala 268:46]
  wire [8:0] _T_2976 = {io_dma_mem_wdata[15],io_dma_mem_wdata[14],io_dma_mem_wdata[9],io_dma_mem_wdata[8],io_dma_mem_wdata[7],io_dma_mem_wdata[6],io_dma_mem_wdata[2],io_dma_mem_wdata[1],io_dma_mem_wdata[0]}; // @[el2_lib.scala 268:56]
  wire [17:0] _T_2985 = {io_dma_mem_wdata[30],io_dma_mem_wdata[29],io_dma_mem_wdata[28],io_dma_mem_wdata[24],io_dma_mem_wdata[23],io_dma_mem_wdata[22],io_dma_mem_wdata[21],io_dma_mem_wdata[17],io_dma_mem_wdata[16],_T_2976}; // @[el2_lib.scala 268:56]
  wire  _T_2986 = ^_T_2985; // @[el2_lib.scala 268:63]
  wire [6:0] _T_2992 = {io_dma_mem_wdata[12],io_dma_mem_wdata[11],io_dma_mem_wdata[10],io_dma_mem_wdata[9],io_dma_mem_wdata[8],io_dma_mem_wdata[7],io_dma_mem_wdata[6]}; // @[el2_lib.scala 268:73]
  wire [14:0] _T_3000 = {io_dma_mem_wdata[27],io_dma_mem_wdata[26],io_dma_mem_wdata[25],io_dma_mem_wdata[24],io_dma_mem_wdata[23],io_dma_mem_wdata[22],io_dma_mem_wdata[21],io_dma_mem_wdata[13],_T_2992}; // @[el2_lib.scala 268:73]
  wire  _T_3001 = ^_T_3000; // @[el2_lib.scala 268:80]
  wire [14:0] _T_3015 = {io_dma_mem_wdata[20],io_dma_mem_wdata[19],io_dma_mem_wdata[18],io_dma_mem_wdata[17],io_dma_mem_wdata[16],io_dma_mem_wdata[15],io_dma_mem_wdata[14],io_dma_mem_wdata[13],_T_2992}; // @[el2_lib.scala 268:90]
  wire  _T_3016 = ^_T_3015; // @[el2_lib.scala 268:97]
  wire [5:0] _T_3021 = {io_dma_mem_wdata[5],io_dma_mem_wdata[4],io_dma_mem_wdata[3],io_dma_mem_wdata[2],io_dma_mem_wdata[1],io_dma_mem_wdata[0]}; // @[el2_lib.scala 268:107]
  wire  _T_3022 = ^_T_3021; // @[el2_lib.scala 268:114]
  wire [5:0] _T_3027 = {_T_2950,_T_2968,_T_2986,_T_3001,_T_3016,_T_3022}; // @[Cat.scala 29:58]
  wire  _T_3028 = ^io_dma_mem_wdata[31:0]; // @[el2_lib.scala 269:13]
  wire  _T_3029 = ^_T_3027; // @[el2_lib.scala 269:23]
  wire  _T_3030 = _T_3028 ^ _T_3029; // @[el2_lib.scala 269:18]
  wire [6:0] _T_3031 = {_T_3030,_T_2950,_T_2968,_T_2986,_T_3001,_T_3016,_T_3022}; // @[Cat.scala 29:58]
  wire [13:0] dma_mem_ecc = {_T_2834,_T_2754,_T_2772,_T_2790,_T_2805,_T_2820,_T_2826,_T_3031}; // @[Cat.scala 29:58]
  wire  _T_3033 = ~_T_2627; // @[el2_ifu_mem_ctl.scala 631:45]
  wire  _T_3034 = iccm_correct_ecc & _T_3033; // @[el2_ifu_mem_ctl.scala 631:43]
  reg [38:0] iccm_ecc_corr_data_ff; // @[Reg.scala 27:20]
  wire [77:0] _T_3035 = {iccm_ecc_corr_data_ff,iccm_ecc_corr_data_ff}; // @[Cat.scala 29:58]
  wire [77:0] _T_3042 = {dma_mem_ecc[13:7],io_dma_mem_wdata[63:32],dma_mem_ecc[6:0],io_dma_mem_wdata[31:0]}; // @[Cat.scala 29:58]
  reg [1:0] dma_mem_addr_ff; // @[el2_ifu_mem_ctl.scala 645:53]
  wire  _T_3374 = _T_3286[5:0] == 6'h27; // @[el2_lib.scala 307:41]
  wire  _T_3372 = _T_3286[5:0] == 6'h26; // @[el2_lib.scala 307:41]
  wire  _T_3370 = _T_3286[5:0] == 6'h25; // @[el2_lib.scala 307:41]
  wire  _T_3368 = _T_3286[5:0] == 6'h24; // @[el2_lib.scala 307:41]
  wire  _T_3366 = _T_3286[5:0] == 6'h23; // @[el2_lib.scala 307:41]
  wire  _T_3364 = _T_3286[5:0] == 6'h22; // @[el2_lib.scala 307:41]
  wire  _T_3362 = _T_3286[5:0] == 6'h21; // @[el2_lib.scala 307:41]
  wire  _T_3360 = _T_3286[5:0] == 6'h20; // @[el2_lib.scala 307:41]
  wire  _T_3358 = _T_3286[5:0] == 6'h1f; // @[el2_lib.scala 307:41]
  wire  _T_3356 = _T_3286[5:0] == 6'h1e; // @[el2_lib.scala 307:41]
  wire [9:0] _T_3432 = {_T_3374,_T_3372,_T_3370,_T_3368,_T_3366,_T_3364,_T_3362,_T_3360,_T_3358,_T_3356}; // @[el2_lib.scala 310:69]
  wire  _T_3354 = _T_3286[5:0] == 6'h1d; // @[el2_lib.scala 307:41]
  wire  _T_3352 = _T_3286[5:0] == 6'h1c; // @[el2_lib.scala 307:41]
  wire  _T_3350 = _T_3286[5:0] == 6'h1b; // @[el2_lib.scala 307:41]
  wire  _T_3348 = _T_3286[5:0] == 6'h1a; // @[el2_lib.scala 307:41]
  wire  _T_3346 = _T_3286[5:0] == 6'h19; // @[el2_lib.scala 307:41]
  wire  _T_3344 = _T_3286[5:0] == 6'h18; // @[el2_lib.scala 307:41]
  wire  _T_3342 = _T_3286[5:0] == 6'h17; // @[el2_lib.scala 307:41]
  wire  _T_3340 = _T_3286[5:0] == 6'h16; // @[el2_lib.scala 307:41]
  wire  _T_3338 = _T_3286[5:0] == 6'h15; // @[el2_lib.scala 307:41]
  wire  _T_3336 = _T_3286[5:0] == 6'h14; // @[el2_lib.scala 307:41]
  wire [9:0] _T_3423 = {_T_3354,_T_3352,_T_3350,_T_3348,_T_3346,_T_3344,_T_3342,_T_3340,_T_3338,_T_3336}; // @[el2_lib.scala 310:69]
  wire  _T_3334 = _T_3286[5:0] == 6'h13; // @[el2_lib.scala 307:41]
  wire  _T_3332 = _T_3286[5:0] == 6'h12; // @[el2_lib.scala 307:41]
  wire  _T_3330 = _T_3286[5:0] == 6'h11; // @[el2_lib.scala 307:41]
  wire  _T_3328 = _T_3286[5:0] == 6'h10; // @[el2_lib.scala 307:41]
  wire  _T_3326 = _T_3286[5:0] == 6'hf; // @[el2_lib.scala 307:41]
  wire  _T_3324 = _T_3286[5:0] == 6'he; // @[el2_lib.scala 307:41]
  wire  _T_3322 = _T_3286[5:0] == 6'hd; // @[el2_lib.scala 307:41]
  wire  _T_3320 = _T_3286[5:0] == 6'hc; // @[el2_lib.scala 307:41]
  wire  _T_3318 = _T_3286[5:0] == 6'hb; // @[el2_lib.scala 307:41]
  wire  _T_3316 = _T_3286[5:0] == 6'ha; // @[el2_lib.scala 307:41]
  wire [9:0] _T_3413 = {_T_3334,_T_3332,_T_3330,_T_3328,_T_3326,_T_3324,_T_3322,_T_3320,_T_3318,_T_3316}; // @[el2_lib.scala 310:69]
  wire  _T_3314 = _T_3286[5:0] == 6'h9; // @[el2_lib.scala 307:41]
  wire  _T_3312 = _T_3286[5:0] == 6'h8; // @[el2_lib.scala 307:41]
  wire  _T_3310 = _T_3286[5:0] == 6'h7; // @[el2_lib.scala 307:41]
  wire  _T_3308 = _T_3286[5:0] == 6'h6; // @[el2_lib.scala 307:41]
  wire  _T_3306 = _T_3286[5:0] == 6'h5; // @[el2_lib.scala 307:41]
  wire  _T_3304 = _T_3286[5:0] == 6'h4; // @[el2_lib.scala 307:41]
  wire  _T_3302 = _T_3286[5:0] == 6'h3; // @[el2_lib.scala 307:41]
  wire  _T_3300 = _T_3286[5:0] == 6'h2; // @[el2_lib.scala 307:41]
  wire  _T_3298 = _T_3286[5:0] == 6'h1; // @[el2_lib.scala 307:41]
  wire [18:0] _T_3414 = {_T_3413,_T_3314,_T_3312,_T_3310,_T_3308,_T_3306,_T_3304,_T_3302,_T_3300,_T_3298}; // @[el2_lib.scala 310:69]
  wire [38:0] _T_3434 = {_T_3432,_T_3423,_T_3414}; // @[el2_lib.scala 310:69]
  wire [7:0] _T_3389 = {io_iccm_rd_data_ecc[35],io_iccm_rd_data_ecc[3:1],io_iccm_rd_data_ecc[34],io_iccm_rd_data_ecc[0],io_iccm_rd_data_ecc[33:32]}; // @[Cat.scala 29:58]
  wire [38:0] _T_3395 = {io_iccm_rd_data_ecc[38],io_iccm_rd_data_ecc[31:26],io_iccm_rd_data_ecc[37],io_iccm_rd_data_ecc[25:11],io_iccm_rd_data_ecc[36],io_iccm_rd_data_ecc[10:4],_T_3389}; // @[Cat.scala 29:58]
  wire [38:0] _T_3435 = _T_3434 ^ _T_3395; // @[el2_lib.scala 310:76]
  wire [38:0] _T_3436 = _T_3290 ? _T_3435 : _T_3395; // @[el2_lib.scala 310:31]
  wire [31:0] iccm_corrected_data_0 = {_T_3436[37:32],_T_3436[30:16],_T_3436[14:8],_T_3436[6:4],_T_3436[2]}; // @[Cat.scala 29:58]
  wire  _T_3759 = _T_3671[5:0] == 6'h27; // @[el2_lib.scala 307:41]
  wire  _T_3757 = _T_3671[5:0] == 6'h26; // @[el2_lib.scala 307:41]
  wire  _T_3755 = _T_3671[5:0] == 6'h25; // @[el2_lib.scala 307:41]
  wire  _T_3753 = _T_3671[5:0] == 6'h24; // @[el2_lib.scala 307:41]
  wire  _T_3751 = _T_3671[5:0] == 6'h23; // @[el2_lib.scala 307:41]
  wire  _T_3749 = _T_3671[5:0] == 6'h22; // @[el2_lib.scala 307:41]
  wire  _T_3747 = _T_3671[5:0] == 6'h21; // @[el2_lib.scala 307:41]
  wire  _T_3745 = _T_3671[5:0] == 6'h20; // @[el2_lib.scala 307:41]
  wire  _T_3743 = _T_3671[5:0] == 6'h1f; // @[el2_lib.scala 307:41]
  wire  _T_3741 = _T_3671[5:0] == 6'h1e; // @[el2_lib.scala 307:41]
  wire [9:0] _T_3817 = {_T_3759,_T_3757,_T_3755,_T_3753,_T_3751,_T_3749,_T_3747,_T_3745,_T_3743,_T_3741}; // @[el2_lib.scala 310:69]
  wire  _T_3739 = _T_3671[5:0] == 6'h1d; // @[el2_lib.scala 307:41]
  wire  _T_3737 = _T_3671[5:0] == 6'h1c; // @[el2_lib.scala 307:41]
  wire  _T_3735 = _T_3671[5:0] == 6'h1b; // @[el2_lib.scala 307:41]
  wire  _T_3733 = _T_3671[5:0] == 6'h1a; // @[el2_lib.scala 307:41]
  wire  _T_3731 = _T_3671[5:0] == 6'h19; // @[el2_lib.scala 307:41]
  wire  _T_3729 = _T_3671[5:0] == 6'h18; // @[el2_lib.scala 307:41]
  wire  _T_3727 = _T_3671[5:0] == 6'h17; // @[el2_lib.scala 307:41]
  wire  _T_3725 = _T_3671[5:0] == 6'h16; // @[el2_lib.scala 307:41]
  wire  _T_3723 = _T_3671[5:0] == 6'h15; // @[el2_lib.scala 307:41]
  wire  _T_3721 = _T_3671[5:0] == 6'h14; // @[el2_lib.scala 307:41]
  wire [9:0] _T_3808 = {_T_3739,_T_3737,_T_3735,_T_3733,_T_3731,_T_3729,_T_3727,_T_3725,_T_3723,_T_3721}; // @[el2_lib.scala 310:69]
  wire  _T_3719 = _T_3671[5:0] == 6'h13; // @[el2_lib.scala 307:41]
  wire  _T_3717 = _T_3671[5:0] == 6'h12; // @[el2_lib.scala 307:41]
  wire  _T_3715 = _T_3671[5:0] == 6'h11; // @[el2_lib.scala 307:41]
  wire  _T_3713 = _T_3671[5:0] == 6'h10; // @[el2_lib.scala 307:41]
  wire  _T_3711 = _T_3671[5:0] == 6'hf; // @[el2_lib.scala 307:41]
  wire  _T_3709 = _T_3671[5:0] == 6'he; // @[el2_lib.scala 307:41]
  wire  _T_3707 = _T_3671[5:0] == 6'hd; // @[el2_lib.scala 307:41]
  wire  _T_3705 = _T_3671[5:0] == 6'hc; // @[el2_lib.scala 307:41]
  wire  _T_3703 = _T_3671[5:0] == 6'hb; // @[el2_lib.scala 307:41]
  wire  _T_3701 = _T_3671[5:0] == 6'ha; // @[el2_lib.scala 307:41]
  wire [9:0] _T_3798 = {_T_3719,_T_3717,_T_3715,_T_3713,_T_3711,_T_3709,_T_3707,_T_3705,_T_3703,_T_3701}; // @[el2_lib.scala 310:69]
  wire  _T_3699 = _T_3671[5:0] == 6'h9; // @[el2_lib.scala 307:41]
  wire  _T_3697 = _T_3671[5:0] == 6'h8; // @[el2_lib.scala 307:41]
  wire  _T_3695 = _T_3671[5:0] == 6'h7; // @[el2_lib.scala 307:41]
  wire  _T_3693 = _T_3671[5:0] == 6'h6; // @[el2_lib.scala 307:41]
  wire  _T_3691 = _T_3671[5:0] == 6'h5; // @[el2_lib.scala 307:41]
  wire  _T_3689 = _T_3671[5:0] == 6'h4; // @[el2_lib.scala 307:41]
  wire  _T_3687 = _T_3671[5:0] == 6'h3; // @[el2_lib.scala 307:41]
  wire  _T_3685 = _T_3671[5:0] == 6'h2; // @[el2_lib.scala 307:41]
  wire  _T_3683 = _T_3671[5:0] == 6'h1; // @[el2_lib.scala 307:41]
  wire [18:0] _T_3799 = {_T_3798,_T_3699,_T_3697,_T_3695,_T_3693,_T_3691,_T_3689,_T_3687,_T_3685,_T_3683}; // @[el2_lib.scala 310:69]
  wire [38:0] _T_3819 = {_T_3817,_T_3808,_T_3799}; // @[el2_lib.scala 310:69]
  wire [7:0] _T_3774 = {io_iccm_rd_data_ecc[74],io_iccm_rd_data_ecc[42:40],io_iccm_rd_data_ecc[73],io_iccm_rd_data_ecc[39],io_iccm_rd_data_ecc[72:71]}; // @[Cat.scala 29:58]
  wire [38:0] _T_3780 = {io_iccm_rd_data_ecc[77],io_iccm_rd_data_ecc[70:65],io_iccm_rd_data_ecc[76],io_iccm_rd_data_ecc[64:50],io_iccm_rd_data_ecc[75],io_iccm_rd_data_ecc[49:43],_T_3774}; // @[Cat.scala 29:58]
  wire [38:0] _T_3820 = _T_3819 ^ _T_3780; // @[el2_lib.scala 310:76]
  wire [38:0] _T_3821 = _T_3675 ? _T_3820 : _T_3780; // @[el2_lib.scala 310:31]
  wire [31:0] iccm_corrected_data_1 = {_T_3821[37:32],_T_3821[30:16],_T_3821[14:8],_T_3821[6:4],_T_3821[2]}; // @[Cat.scala 29:58]
  wire [31:0] iccm_dma_rdata_1_muxed = dma_mem_addr_ff[0] ? iccm_corrected_data_0 : iccm_corrected_data_1; // @[el2_ifu_mem_ctl.scala 637:35]
  wire  _T_3294 = ~_T_3286[6]; // @[el2_lib.scala 303:55]
  wire  _T_3295 = _T_3288 & _T_3294; // @[el2_lib.scala 303:53]
  wire  _T_3679 = ~_T_3671[6]; // @[el2_lib.scala 303:55]
  wire  _T_3680 = _T_3673 & _T_3679; // @[el2_lib.scala 303:53]
  wire [1:0] iccm_double_ecc_error = {_T_3295,_T_3680}; // @[Cat.scala 29:58]
  wire  iccm_dma_ecc_error_in = |iccm_double_ecc_error; // @[el2_ifu_mem_ctl.scala 639:53]
  wire [63:0] _T_3046 = {io_dma_mem_addr,io_dma_mem_addr}; // @[Cat.scala 29:58]
  wire [63:0] _T_3047 = {iccm_dma_rdata_1_muxed,_T_3436[37:32],_T_3436[30:16],_T_3436[14:8],_T_3436[6:4],_T_3436[2]}; // @[Cat.scala 29:58]
  reg [2:0] dma_mem_tag_ff; // @[el2_ifu_mem_ctl.scala 641:54]
  reg [2:0] iccm_dma_rtag; // @[el2_ifu_mem_ctl.scala 642:69]
  reg  iccm_dma_rvalid; // @[el2_ifu_mem_ctl.scala 647:71]
  reg [63:0] iccm_dma_rdata; // @[el2_ifu_mem_ctl.scala 651:70]
  wire  _T_3052 = _T_2627 & _T_2616; // @[el2_ifu_mem_ctl.scala 654:65]
  wire  _T_3055 = _T_3033 & iccm_correct_ecc; // @[el2_ifu_mem_ctl.scala 655:50]
  reg [13:0] iccm_ecc_corr_index_ff; // @[Reg.scala 27:20]
  wire [14:0] _T_3056 = {iccm_ecc_corr_index_ff,1'h0}; // @[Cat.scala 29:58]
  wire [15:0] _T_3058 = _T_3055 ? {{1'd0}, _T_3056} : io_ifc_fetch_addr_bf[15:0]; // @[el2_ifu_mem_ctl.scala 655:8]
  wire [31:0] _T_3059 = _T_3052 ? io_dma_mem_addr : {{16'd0}, _T_3058}; // @[el2_ifu_mem_ctl.scala 654:25]
  wire  _T_3448 = _T_3286 == 7'h40; // @[el2_lib.scala 313:62]
  wire  _T_3449 = _T_3436[38] ^ _T_3448; // @[el2_lib.scala 313:44]
  wire [6:0] iccm_corrected_ecc_0 = {_T_3449,_T_3436[31],_T_3436[15],_T_3436[7],_T_3436[3],_T_3436[1:0]}; // @[Cat.scala 29:58]
  wire  _T_3833 = _T_3671 == 7'h40; // @[el2_lib.scala 313:62]
  wire  _T_3834 = _T_3821[38] ^ _T_3833; // @[el2_lib.scala 313:44]
  wire [6:0] iccm_corrected_ecc_1 = {_T_3834,_T_3821[31],_T_3821[15],_T_3821[7],_T_3821[3],_T_3821[1:0]}; // @[Cat.scala 29:58]
  wire  _T_3850 = _T_3 & ifc_iccm_access_f; // @[el2_ifu_mem_ctl.scala 667:58]
  wire [31:0] iccm_corrected_data_f_mux = iccm_single_ecc_error[0] ? iccm_corrected_data_0 : iccm_corrected_data_1; // @[el2_ifu_mem_ctl.scala 669:38]
  wire [6:0] iccm_corrected_ecc_f_mux = iccm_single_ecc_error[0] ? iccm_corrected_ecc_0 : iccm_corrected_ecc_1; // @[el2_ifu_mem_ctl.scala 670:37]
  reg  iccm_rd_ecc_single_err_ff; // @[el2_ifu_mem_ctl.scala 678:62]
  wire  _T_3858 = ~iccm_rd_ecc_single_err_ff; // @[el2_ifu_mem_ctl.scala 672:76]
  wire  _T_3859 = io_iccm_rd_ecc_single_err & _T_3858; // @[el2_ifu_mem_ctl.scala 672:74]
  wire  _T_3861 = _T_3859 & _T_318; // @[el2_ifu_mem_ctl.scala 672:104]
  wire  iccm_ecc_write_status = _T_3861 | io_iccm_dma_sb_error; // @[el2_ifu_mem_ctl.scala 672:127]
  wire  _T_3862 = io_iccm_rd_ecc_single_err | iccm_rd_ecc_single_err_ff; // @[el2_ifu_mem_ctl.scala 673:67]
  wire  iccm_rd_ecc_single_err_hold_in = _T_3862 & _T_318; // @[el2_ifu_mem_ctl.scala 673:96]
  reg [13:0] iccm_rw_addr_f; // @[el2_ifu_mem_ctl.scala 677:51]
  wire [13:0] _T_3867 = iccm_rw_addr_f + 14'h1; // @[el2_ifu_mem_ctl.scala 676:102]
  wire [38:0] _T_3871 = {iccm_corrected_ecc_f_mux,iccm_corrected_data_f_mux}; // @[Cat.scala 29:58]
  wire  _T_3876 = ~io_ifc_fetch_uncacheable_bf; // @[el2_ifu_mem_ctl.scala 681:41]
  wire  _T_3877 = io_ifc_fetch_req_bf & _T_3876; // @[el2_ifu_mem_ctl.scala 681:39]
  wire  _T_3878 = ~io_ifc_iccm_access_bf; // @[el2_ifu_mem_ctl.scala 681:72]
  wire  _T_3879 = _T_3877 & _T_3878; // @[el2_ifu_mem_ctl.scala 681:70]
  wire  _T_3881 = ~miss_state_en; // @[el2_ifu_mem_ctl.scala 682:34]
  wire  _T_3882 = _T_2222 & _T_3881; // @[el2_ifu_mem_ctl.scala 682:32]
  wire  _T_3885 = _T_2238 & _T_3881; // @[el2_ifu_mem_ctl.scala 683:37]
  wire  _T_3886 = _T_3882 | _T_3885; // @[el2_ifu_mem_ctl.scala 682:88]
  wire  _T_3887 = miss_state == 3'h7; // @[el2_ifu_mem_ctl.scala 684:19]
  wire  _T_3889 = _T_3887 & _T_3881; // @[el2_ifu_mem_ctl.scala 684:41]
  wire  _T_3890 = _T_3886 | _T_3889; // @[el2_ifu_mem_ctl.scala 683:88]
  wire  _T_3891 = miss_state == 3'h3; // @[el2_ifu_mem_ctl.scala 685:19]
  wire  _T_3893 = _T_3891 & _T_3881; // @[el2_ifu_mem_ctl.scala 685:35]
  wire  _T_3894 = _T_3890 | _T_3893; // @[el2_ifu_mem_ctl.scala 684:88]
  wire  _T_3897 = _T_2237 & _T_3881; // @[el2_ifu_mem_ctl.scala 686:38]
  wire  _T_3898 = _T_3894 | _T_3897; // @[el2_ifu_mem_ctl.scala 685:88]
  wire  _T_3900 = _T_2238 & miss_state_en; // @[el2_ifu_mem_ctl.scala 687:37]
  wire  _T_3901 = miss_nxtstate == 3'h3; // @[el2_ifu_mem_ctl.scala 687:71]
  wire  _T_3902 = _T_3900 & _T_3901; // @[el2_ifu_mem_ctl.scala 687:54]
  wire  _T_3903 = _T_3898 | _T_3902; // @[el2_ifu_mem_ctl.scala 686:57]
  wire  _T_3904 = ~_T_3903; // @[el2_ifu_mem_ctl.scala 682:5]
  wire  _T_3905 = _T_3879 & _T_3904; // @[el2_ifu_mem_ctl.scala 681:96]
  wire  _T_3906 = io_ifc_fetch_req_bf & io_exu_flush_final; // @[el2_ifu_mem_ctl.scala 688:28]
  wire  _T_3908 = _T_3906 & _T_3876; // @[el2_ifu_mem_ctl.scala 688:50]
  wire  _T_3910 = _T_3908 & _T_3878; // @[el2_ifu_mem_ctl.scala 688:81]
  wire  _T_3919 = ~_T_109; // @[el2_ifu_mem_ctl.scala 691:106]
  wire  _T_3920 = _T_2222 & _T_3919; // @[el2_ifu_mem_ctl.scala 691:104]
  wire  _T_3921 = _T_2238 | _T_3920; // @[el2_ifu_mem_ctl.scala 691:77]
  wire  _T_3925 = ~_T_52; // @[el2_ifu_mem_ctl.scala 691:172]
  wire  _T_3926 = _T_3921 & _T_3925; // @[el2_ifu_mem_ctl.scala 691:170]
  wire  _T_3927 = ~_T_3926; // @[el2_ifu_mem_ctl.scala 691:44]
  wire  _T_3931 = reset_ic_in | reset_ic_ff; // @[el2_ifu_mem_ctl.scala 694:64]
  wire  _T_3932 = ~_T_3931; // @[el2_ifu_mem_ctl.scala 694:50]
  wire  _T_3933 = _T_277 & _T_3932; // @[el2_ifu_mem_ctl.scala 694:48]
  wire  _T_3934 = ~reset_tag_valid_for_miss; // @[el2_ifu_mem_ctl.scala 694:81]
  wire  ic_valid = _T_3933 & _T_3934; // @[el2_ifu_mem_ctl.scala 694:79]
  wire  _T_3936 = debug_c1_clken & io_ic_debug_tag_array; // @[el2_ifu_mem_ctl.scala 695:82]
  reg [6:0] ifu_status_wr_addr_ff; // @[el2_ifu_mem_ctl.scala 698:14]
  wire  _T_3939 = io_ic_debug_wr_en & io_ic_debug_tag_array; // @[el2_ifu_mem_ctl.scala 701:74]
  wire  _T_10081 = bus_ifu_wr_en_ff_q & last_beat; // @[el2_ifu_mem_ctl.scala 775:45]
  wire  way_status_wr_en = _T_10081 | ic_act_hit_f; // @[el2_ifu_mem_ctl.scala 775:58]
  wire  way_status_wr_en_w_debug = way_status_wr_en | _T_3939; // @[el2_ifu_mem_ctl.scala 701:53]
  reg  way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 703:14]
  wire [2:0] _T_3943 = {{2'd0}, io_ic_debug_wr_data[4]}; // @[el2_ifu_mem_ctl.scala 707:10]
  wire  way_status_hit_new = io_ic_rd_hit[0]; // @[el2_ifu_mem_ctl.scala 771:41]
  wire  way_status_new = _T_10081 ? replace_way_mb_any_0 : way_status_hit_new; // @[el2_ifu_mem_ctl.scala 774:26]
  reg [2:0] way_status_new_ff; // @[el2_ifu_mem_ctl.scala 709:14]
  wire  way_status_clken_0 = ifu_status_wr_addr_ff[6:3] == 4'h0; // @[el2_ifu_mem_ctl.scala 711:132]
  wire  way_status_clken_1 = ifu_status_wr_addr_ff[6:3] == 4'h1; // @[el2_ifu_mem_ctl.scala 711:132]
  wire  way_status_clken_2 = ifu_status_wr_addr_ff[6:3] == 4'h2; // @[el2_ifu_mem_ctl.scala 711:132]
  wire  way_status_clken_3 = ifu_status_wr_addr_ff[6:3] == 4'h3; // @[el2_ifu_mem_ctl.scala 711:132]
  wire  way_status_clken_4 = ifu_status_wr_addr_ff[6:3] == 4'h4; // @[el2_ifu_mem_ctl.scala 711:132]
  wire  way_status_clken_5 = ifu_status_wr_addr_ff[6:3] == 4'h5; // @[el2_ifu_mem_ctl.scala 711:132]
  wire  way_status_clken_6 = ifu_status_wr_addr_ff[6:3] == 4'h6; // @[el2_ifu_mem_ctl.scala 711:132]
  wire  way_status_clken_7 = ifu_status_wr_addr_ff[6:3] == 4'h7; // @[el2_ifu_mem_ctl.scala 711:132]
  wire  way_status_clken_8 = ifu_status_wr_addr_ff[6:3] == 4'h8; // @[el2_ifu_mem_ctl.scala 711:132]
  wire  way_status_clken_9 = ifu_status_wr_addr_ff[6:3] == 4'h9; // @[el2_ifu_mem_ctl.scala 711:132]
  wire  way_status_clken_10 = ifu_status_wr_addr_ff[6:3] == 4'ha; // @[el2_ifu_mem_ctl.scala 711:132]
  wire  way_status_clken_11 = ifu_status_wr_addr_ff[6:3] == 4'hb; // @[el2_ifu_mem_ctl.scala 711:132]
  wire  way_status_clken_12 = ifu_status_wr_addr_ff[6:3] == 4'hc; // @[el2_ifu_mem_ctl.scala 711:132]
  wire  way_status_clken_13 = ifu_status_wr_addr_ff[6:3] == 4'hd; // @[el2_ifu_mem_ctl.scala 711:132]
  wire  way_status_clken_14 = ifu_status_wr_addr_ff[6:3] == 4'he; // @[el2_ifu_mem_ctl.scala 711:132]
  wire  way_status_clken_15 = ifu_status_wr_addr_ff[6:3] == 4'hf; // @[el2_ifu_mem_ctl.scala 711:132]
  wire  _T_3960 = ifu_status_wr_addr_ff == 7'h0; // @[el2_ifu_mem_ctl.scala 715:93]
  wire  _T_3961 = _T_3960 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 715:102]
  wire  _T_3962 = _T_3961 & way_status_clken_0; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_3964 = ifu_status_wr_addr_ff == 7'h1; // @[el2_ifu_mem_ctl.scala 715:93]
  wire  _T_3965 = _T_3964 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 715:102]
  wire  _T_3966 = _T_3965 & way_status_clken_0; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_3968 = ifu_status_wr_addr_ff == 7'h2; // @[el2_ifu_mem_ctl.scala 715:93]
  wire  _T_3969 = _T_3968 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 715:102]
  wire  _T_3970 = _T_3969 & way_status_clken_0; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_3972 = ifu_status_wr_addr_ff == 7'h3; // @[el2_ifu_mem_ctl.scala 715:93]
  wire  _T_3973 = _T_3972 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 715:102]
  wire  _T_3974 = _T_3973 & way_status_clken_0; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_3976 = ifu_status_wr_addr_ff == 7'h4; // @[el2_ifu_mem_ctl.scala 715:93]
  wire  _T_3977 = _T_3976 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 715:102]
  wire  _T_3978 = _T_3977 & way_status_clken_0; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_3980 = ifu_status_wr_addr_ff == 7'h5; // @[el2_ifu_mem_ctl.scala 715:93]
  wire  _T_3981 = _T_3980 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 715:102]
  wire  _T_3982 = _T_3981 & way_status_clken_0; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_3984 = ifu_status_wr_addr_ff == 7'h6; // @[el2_ifu_mem_ctl.scala 715:93]
  wire  _T_3985 = _T_3984 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 715:102]
  wire  _T_3986 = _T_3985 & way_status_clken_0; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_3988 = ifu_status_wr_addr_ff == 7'h7; // @[el2_ifu_mem_ctl.scala 715:93]
  wire  _T_3989 = _T_3988 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 715:102]
  wire  _T_3990 = _T_3989 & way_status_clken_0; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_3994 = _T_3961 & way_status_clken_1; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_3998 = _T_3965 & way_status_clken_1; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4002 = _T_3969 & way_status_clken_1; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4006 = _T_3973 & way_status_clken_1; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4010 = _T_3977 & way_status_clken_1; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4014 = _T_3981 & way_status_clken_1; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4018 = _T_3985 & way_status_clken_1; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4022 = _T_3989 & way_status_clken_1; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4026 = _T_3961 & way_status_clken_2; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4030 = _T_3965 & way_status_clken_2; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4034 = _T_3969 & way_status_clken_2; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4038 = _T_3973 & way_status_clken_2; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4042 = _T_3977 & way_status_clken_2; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4046 = _T_3981 & way_status_clken_2; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4050 = _T_3985 & way_status_clken_2; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4054 = _T_3989 & way_status_clken_2; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4058 = _T_3961 & way_status_clken_3; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4062 = _T_3965 & way_status_clken_3; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4066 = _T_3969 & way_status_clken_3; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4070 = _T_3973 & way_status_clken_3; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4074 = _T_3977 & way_status_clken_3; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4078 = _T_3981 & way_status_clken_3; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4082 = _T_3985 & way_status_clken_3; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4086 = _T_3989 & way_status_clken_3; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4090 = _T_3961 & way_status_clken_4; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4094 = _T_3965 & way_status_clken_4; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4098 = _T_3969 & way_status_clken_4; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4102 = _T_3973 & way_status_clken_4; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4106 = _T_3977 & way_status_clken_4; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4110 = _T_3981 & way_status_clken_4; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4114 = _T_3985 & way_status_clken_4; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4118 = _T_3989 & way_status_clken_4; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4122 = _T_3961 & way_status_clken_5; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4126 = _T_3965 & way_status_clken_5; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4130 = _T_3969 & way_status_clken_5; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4134 = _T_3973 & way_status_clken_5; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4138 = _T_3977 & way_status_clken_5; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4142 = _T_3981 & way_status_clken_5; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4146 = _T_3985 & way_status_clken_5; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4150 = _T_3989 & way_status_clken_5; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4154 = _T_3961 & way_status_clken_6; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4158 = _T_3965 & way_status_clken_6; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4162 = _T_3969 & way_status_clken_6; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4166 = _T_3973 & way_status_clken_6; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4170 = _T_3977 & way_status_clken_6; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4174 = _T_3981 & way_status_clken_6; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4178 = _T_3985 & way_status_clken_6; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4182 = _T_3989 & way_status_clken_6; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4186 = _T_3961 & way_status_clken_7; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4190 = _T_3965 & way_status_clken_7; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4194 = _T_3969 & way_status_clken_7; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4198 = _T_3973 & way_status_clken_7; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4202 = _T_3977 & way_status_clken_7; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4206 = _T_3981 & way_status_clken_7; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4210 = _T_3985 & way_status_clken_7; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4214 = _T_3989 & way_status_clken_7; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4218 = _T_3961 & way_status_clken_8; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4222 = _T_3965 & way_status_clken_8; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4226 = _T_3969 & way_status_clken_8; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4230 = _T_3973 & way_status_clken_8; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4234 = _T_3977 & way_status_clken_8; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4238 = _T_3981 & way_status_clken_8; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4242 = _T_3985 & way_status_clken_8; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4246 = _T_3989 & way_status_clken_8; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4250 = _T_3961 & way_status_clken_9; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4254 = _T_3965 & way_status_clken_9; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4258 = _T_3969 & way_status_clken_9; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4262 = _T_3973 & way_status_clken_9; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4266 = _T_3977 & way_status_clken_9; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4270 = _T_3981 & way_status_clken_9; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4274 = _T_3985 & way_status_clken_9; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4278 = _T_3989 & way_status_clken_9; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4282 = _T_3961 & way_status_clken_10; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4286 = _T_3965 & way_status_clken_10; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4290 = _T_3969 & way_status_clken_10; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4294 = _T_3973 & way_status_clken_10; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4298 = _T_3977 & way_status_clken_10; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4302 = _T_3981 & way_status_clken_10; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4306 = _T_3985 & way_status_clken_10; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4310 = _T_3989 & way_status_clken_10; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4314 = _T_3961 & way_status_clken_11; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4318 = _T_3965 & way_status_clken_11; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4322 = _T_3969 & way_status_clken_11; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4326 = _T_3973 & way_status_clken_11; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4330 = _T_3977 & way_status_clken_11; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4334 = _T_3981 & way_status_clken_11; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4338 = _T_3985 & way_status_clken_11; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4342 = _T_3989 & way_status_clken_11; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4346 = _T_3961 & way_status_clken_12; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4350 = _T_3965 & way_status_clken_12; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4354 = _T_3969 & way_status_clken_12; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4358 = _T_3973 & way_status_clken_12; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4362 = _T_3977 & way_status_clken_12; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4366 = _T_3981 & way_status_clken_12; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4370 = _T_3985 & way_status_clken_12; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4374 = _T_3989 & way_status_clken_12; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4378 = _T_3961 & way_status_clken_13; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4382 = _T_3965 & way_status_clken_13; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4386 = _T_3969 & way_status_clken_13; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4390 = _T_3973 & way_status_clken_13; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4394 = _T_3977 & way_status_clken_13; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4398 = _T_3981 & way_status_clken_13; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4402 = _T_3985 & way_status_clken_13; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4406 = _T_3989 & way_status_clken_13; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4410 = _T_3961 & way_status_clken_14; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4414 = _T_3965 & way_status_clken_14; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4418 = _T_3969 & way_status_clken_14; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4422 = _T_3973 & way_status_clken_14; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4426 = _T_3977 & way_status_clken_14; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4430 = _T_3981 & way_status_clken_14; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4434 = _T_3985 & way_status_clken_14; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4438 = _T_3989 & way_status_clken_14; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4442 = _T_3961 & way_status_clken_15; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4446 = _T_3965 & way_status_clken_15; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4450 = _T_3969 & way_status_clken_15; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4454 = _T_3973 & way_status_clken_15; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4458 = _T_3977 & way_status_clken_15; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4462 = _T_3981 & way_status_clken_15; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4466 = _T_3985 & way_status_clken_15; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_4470 = _T_3989 & way_status_clken_15; // @[el2_ifu_mem_ctl.scala 715:124]
  wire  _T_10087 = _T_101 & replace_way_mb_any_1; // @[el2_ifu_mem_ctl.scala 778:84]
  wire  _T_10088 = _T_10087 & miss_pending; // @[el2_ifu_mem_ctl.scala 778:108]
  wire  bus_wren_last_1 = _T_10088 & bus_last_data_beat; // @[el2_ifu_mem_ctl.scala 778:123]
  wire  wren_reset_miss_1 = replace_way_mb_any_1 & reset_tag_valid_for_miss; // @[el2_ifu_mem_ctl.scala 779:84]
  wire  _T_10090 = bus_wren_last_1 | wren_reset_miss_1; // @[el2_ifu_mem_ctl.scala 780:73]
  wire  _T_10085 = _T_101 & replace_way_mb_any_0; // @[el2_ifu_mem_ctl.scala 778:84]
  wire  _T_10086 = _T_10085 & miss_pending; // @[el2_ifu_mem_ctl.scala 778:108]
  wire  bus_wren_last_0 = _T_10086 & bus_last_data_beat; // @[el2_ifu_mem_ctl.scala 778:123]
  wire  wren_reset_miss_0 = replace_way_mb_any_0 & reset_tag_valid_for_miss; // @[el2_ifu_mem_ctl.scala 779:84]
  wire  _T_10089 = bus_wren_last_0 | wren_reset_miss_0; // @[el2_ifu_mem_ctl.scala 780:73]
  wire [1:0] ifu_tag_wren = {_T_10090,_T_10089}; // @[Cat.scala 29:58]
  wire [1:0] _T_10124 = _T_3939 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [1:0] ic_debug_tag_wr_en = _T_10124 & io_ic_debug_way; // @[el2_ifu_mem_ctl.scala 813:90]
  wire [1:0] ifu_tag_wren_w_debug = ifu_tag_wren | ic_debug_tag_wr_en; // @[el2_ifu_mem_ctl.scala 724:45]
  reg [1:0] ifu_tag_wren_ff; // @[el2_ifu_mem_ctl.scala 726:14]
  reg  ic_valid_ff; // @[el2_ifu_mem_ctl.scala 730:14]
  wire  _T_5119 = ifu_ic_rw_int_addr_ff[5:4] == 2'h0; // @[el2_ifu_mem_ctl.scala 734:82]
  wire  _T_5121 = _T_5119 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 734:91]
  wire  _T_5123 = perr_ic_index_ff[5:4] == 2'h0; // @[el2_ifu_mem_ctl.scala 735:74]
  wire  _T_5125 = _T_5123 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 735:83]
  wire  _T_5126 = _T_5121 | _T_5125; // @[el2_ifu_mem_ctl.scala 734:113]
  wire  _T_5127 = _T_5126 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 735:106]
  wire  _T_5131 = _T_5119 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 734:91]
  wire  _T_5135 = _T_5123 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 735:83]
  wire  _T_5136 = _T_5131 | _T_5135; // @[el2_ifu_mem_ctl.scala 734:113]
  wire  _T_5137 = _T_5136 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 735:106]
  wire [1:0] tag_valid_clken_0 = {_T_5127,_T_5137}; // @[Cat.scala 29:58]
  wire  _T_5139 = ifu_ic_rw_int_addr_ff[5:4] == 2'h1; // @[el2_ifu_mem_ctl.scala 734:82]
  wire  _T_5141 = _T_5139 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 734:91]
  wire  _T_5143 = perr_ic_index_ff[5:4] == 2'h1; // @[el2_ifu_mem_ctl.scala 735:74]
  wire  _T_5145 = _T_5143 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 735:83]
  wire  _T_5146 = _T_5141 | _T_5145; // @[el2_ifu_mem_ctl.scala 734:113]
  wire  _T_5147 = _T_5146 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 735:106]
  wire  _T_5151 = _T_5139 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 734:91]
  wire  _T_5155 = _T_5143 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 735:83]
  wire  _T_5156 = _T_5151 | _T_5155; // @[el2_ifu_mem_ctl.scala 734:113]
  wire  _T_5157 = _T_5156 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 735:106]
  wire [1:0] tag_valid_clken_1 = {_T_5147,_T_5157}; // @[Cat.scala 29:58]
  wire  _T_5159 = ifu_ic_rw_int_addr_ff[5:4] == 2'h2; // @[el2_ifu_mem_ctl.scala 734:82]
  wire  _T_5161 = _T_5159 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 734:91]
  wire  _T_5163 = perr_ic_index_ff[5:4] == 2'h2; // @[el2_ifu_mem_ctl.scala 735:74]
  wire  _T_5165 = _T_5163 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 735:83]
  wire  _T_5166 = _T_5161 | _T_5165; // @[el2_ifu_mem_ctl.scala 734:113]
  wire  _T_5167 = _T_5166 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 735:106]
  wire  _T_5171 = _T_5159 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 734:91]
  wire  _T_5175 = _T_5163 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 735:83]
  wire  _T_5176 = _T_5171 | _T_5175; // @[el2_ifu_mem_ctl.scala 734:113]
  wire  _T_5177 = _T_5176 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 735:106]
  wire [1:0] tag_valid_clken_2 = {_T_5167,_T_5177}; // @[Cat.scala 29:58]
  wire  _T_5179 = ifu_ic_rw_int_addr_ff[5:4] == 2'h3; // @[el2_ifu_mem_ctl.scala 734:82]
  wire  _T_5181 = _T_5179 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 734:91]
  wire  _T_5183 = perr_ic_index_ff[5:4] == 2'h3; // @[el2_ifu_mem_ctl.scala 735:74]
  wire  _T_5185 = _T_5183 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 735:83]
  wire  _T_5186 = _T_5181 | _T_5185; // @[el2_ifu_mem_ctl.scala 734:113]
  wire  _T_5187 = _T_5186 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 735:106]
  wire  _T_5191 = _T_5179 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 734:91]
  wire  _T_5195 = _T_5183 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 735:83]
  wire  _T_5196 = _T_5191 | _T_5195; // @[el2_ifu_mem_ctl.scala 734:113]
  wire  _T_5197 = _T_5196 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 735:106]
  wire [1:0] tag_valid_clken_3 = {_T_5187,_T_5197}; // @[Cat.scala 29:58]
  wire  _T_5200 = ic_valid_ff & _T_196; // @[el2_ifu_mem_ctl.scala 740:64]
  wire  _T_5201 = ~perr_sel_invalidate; // @[el2_ifu_mem_ctl.scala 740:91]
  wire  _T_5202 = _T_5200 & _T_5201; // @[el2_ifu_mem_ctl.scala 740:89]
  wire  _T_5205 = _T_4472 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_5206 = perr_ic_index_ff == 6'h0; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_5208 = _T_5206 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_5210 = _T_5208 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_5211 = _T_5205 | _T_5210; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_5221 = _T_4476 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_5222 = perr_ic_index_ff == 6'h1; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_5224 = _T_5222 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_5226 = _T_5224 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_5227 = _T_5221 | _T_5226; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_5237 = _T_4480 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_5238 = perr_ic_index_ff == 6'h2; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_5240 = _T_5238 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_5242 = _T_5240 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_5243 = _T_5237 | _T_5242; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_5253 = _T_4484 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_5254 = perr_ic_index_ff == 6'h3; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_5256 = _T_5254 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_5258 = _T_5256 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_5259 = _T_5253 | _T_5258; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_5269 = _T_4488 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_5270 = perr_ic_index_ff == 6'h4; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_5272 = _T_5270 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_5274 = _T_5272 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_5275 = _T_5269 | _T_5274; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_5285 = _T_4492 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_5286 = perr_ic_index_ff == 6'h5; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_5288 = _T_5286 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_5290 = _T_5288 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_5291 = _T_5285 | _T_5290; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_5301 = _T_4496 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_5302 = perr_ic_index_ff == 6'h6; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_5304 = _T_5302 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_5306 = _T_5304 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_5307 = _T_5301 | _T_5306; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_5317 = _T_4500 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_5318 = perr_ic_index_ff == 6'h7; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_5320 = _T_5318 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_5322 = _T_5320 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_5323 = _T_5317 | _T_5322; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_5333 = _T_4504 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_5334 = perr_ic_index_ff == 6'h8; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_5336 = _T_5334 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_5338 = _T_5336 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_5339 = _T_5333 | _T_5338; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_5349 = _T_4508 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_5350 = perr_ic_index_ff == 6'h9; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_5352 = _T_5350 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_5354 = _T_5352 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_5355 = _T_5349 | _T_5354; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_5365 = _T_4512 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_5366 = perr_ic_index_ff == 6'ha; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_5368 = _T_5366 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_5370 = _T_5368 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_5371 = _T_5365 | _T_5370; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_5381 = _T_4516 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_5382 = perr_ic_index_ff == 6'hb; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_5384 = _T_5382 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_5386 = _T_5384 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_5387 = _T_5381 | _T_5386; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_5397 = _T_4520 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_5398 = perr_ic_index_ff == 6'hc; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_5400 = _T_5398 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_5402 = _T_5400 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_5403 = _T_5397 | _T_5402; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_5413 = _T_4524 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_5414 = perr_ic_index_ff == 6'hd; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_5416 = _T_5414 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_5418 = _T_5416 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_5419 = _T_5413 | _T_5418; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_5429 = _T_4528 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_5430 = perr_ic_index_ff == 6'he; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_5432 = _T_5430 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_5434 = _T_5432 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_5435 = _T_5429 | _T_5434; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_5445 = _T_4532 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_5446 = perr_ic_index_ff == 6'hf; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_5448 = _T_5446 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_5450 = _T_5448 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_5451 = _T_5445 | _T_5450; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_5461 = _T_4536 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_5462 = perr_ic_index_ff == 6'h10; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_5464 = _T_5462 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_5466 = _T_5464 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_5467 = _T_5461 | _T_5466; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_5477 = _T_4540 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_5478 = perr_ic_index_ff == 6'h11; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_5480 = _T_5478 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_5482 = _T_5480 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_5483 = _T_5477 | _T_5482; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_5493 = _T_4544 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_5494 = perr_ic_index_ff == 6'h12; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_5496 = _T_5494 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_5498 = _T_5496 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_5499 = _T_5493 | _T_5498; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_5509 = _T_4548 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_5510 = perr_ic_index_ff == 6'h13; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_5512 = _T_5510 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_5514 = _T_5512 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_5515 = _T_5509 | _T_5514; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_5525 = _T_4552 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_5526 = perr_ic_index_ff == 6'h14; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_5528 = _T_5526 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_5530 = _T_5528 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_5531 = _T_5525 | _T_5530; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_5541 = _T_4556 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_5542 = perr_ic_index_ff == 6'h15; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_5544 = _T_5542 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_5546 = _T_5544 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_5547 = _T_5541 | _T_5546; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_5557 = _T_4560 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_5558 = perr_ic_index_ff == 6'h16; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_5560 = _T_5558 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_5562 = _T_5560 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_5563 = _T_5557 | _T_5562; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_5573 = _T_4564 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_5574 = perr_ic_index_ff == 6'h17; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_5576 = _T_5574 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_5578 = _T_5576 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_5579 = _T_5573 | _T_5578; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_5589 = _T_4568 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_5590 = perr_ic_index_ff == 6'h18; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_5592 = _T_5590 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_5594 = _T_5592 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_5595 = _T_5589 | _T_5594; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_5605 = _T_4572 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_5606 = perr_ic_index_ff == 6'h19; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_5608 = _T_5606 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_5610 = _T_5608 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_5611 = _T_5605 | _T_5610; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_5621 = _T_4576 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_5622 = perr_ic_index_ff == 6'h1a; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_5624 = _T_5622 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_5626 = _T_5624 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_5627 = _T_5621 | _T_5626; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_5637 = _T_4580 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_5638 = perr_ic_index_ff == 6'h1b; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_5640 = _T_5638 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_5642 = _T_5640 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_5643 = _T_5637 | _T_5642; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_5653 = _T_4584 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_5654 = perr_ic_index_ff == 6'h1c; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_5656 = _T_5654 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_5658 = _T_5656 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_5659 = _T_5653 | _T_5658; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_5669 = _T_4588 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_5670 = perr_ic_index_ff == 6'h1d; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_5672 = _T_5670 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_5674 = _T_5672 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_5675 = _T_5669 | _T_5674; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_5685 = _T_4592 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_5686 = perr_ic_index_ff == 6'h1e; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_5688 = _T_5686 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_5690 = _T_5688 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_5691 = _T_5685 | _T_5690; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_5701 = _T_4596 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_5702 = perr_ic_index_ff == 6'h1f; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_5704 = _T_5702 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_5706 = _T_5704 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_5707 = _T_5701 | _T_5706; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_5717 = _T_4472 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_5720 = _T_5206 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_5722 = _T_5720 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_5723 = _T_5717 | _T_5722; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_5733 = _T_4476 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_5736 = _T_5222 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_5738 = _T_5736 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_5739 = _T_5733 | _T_5738; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_5749 = _T_4480 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_5752 = _T_5238 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_5754 = _T_5752 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_5755 = _T_5749 | _T_5754; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_5765 = _T_4484 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_5768 = _T_5254 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_5770 = _T_5768 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_5771 = _T_5765 | _T_5770; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_5781 = _T_4488 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_5784 = _T_5270 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_5786 = _T_5784 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_5787 = _T_5781 | _T_5786; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_5797 = _T_4492 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_5800 = _T_5286 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_5802 = _T_5800 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_5803 = _T_5797 | _T_5802; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_5813 = _T_4496 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_5816 = _T_5302 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_5818 = _T_5816 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_5819 = _T_5813 | _T_5818; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_5829 = _T_4500 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_5832 = _T_5318 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_5834 = _T_5832 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_5835 = _T_5829 | _T_5834; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_5845 = _T_4504 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_5848 = _T_5334 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_5850 = _T_5848 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_5851 = _T_5845 | _T_5850; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_5861 = _T_4508 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_5864 = _T_5350 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_5866 = _T_5864 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_5867 = _T_5861 | _T_5866; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_5877 = _T_4512 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_5880 = _T_5366 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_5882 = _T_5880 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_5883 = _T_5877 | _T_5882; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_5893 = _T_4516 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_5896 = _T_5382 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_5898 = _T_5896 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_5899 = _T_5893 | _T_5898; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_5909 = _T_4520 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_5912 = _T_5398 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_5914 = _T_5912 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_5915 = _T_5909 | _T_5914; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_5925 = _T_4524 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_5928 = _T_5414 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_5930 = _T_5928 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_5931 = _T_5925 | _T_5930; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_5941 = _T_4528 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_5944 = _T_5430 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_5946 = _T_5944 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_5947 = _T_5941 | _T_5946; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_5957 = _T_4532 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_5960 = _T_5446 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_5962 = _T_5960 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_5963 = _T_5957 | _T_5962; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_5973 = _T_4536 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_5976 = _T_5462 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_5978 = _T_5976 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_5979 = _T_5973 | _T_5978; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_5989 = _T_4540 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_5992 = _T_5478 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_5994 = _T_5992 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_5995 = _T_5989 | _T_5994; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_6005 = _T_4544 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_6008 = _T_5494 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_6010 = _T_6008 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_6011 = _T_6005 | _T_6010; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_6021 = _T_4548 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_6024 = _T_5510 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_6026 = _T_6024 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_6027 = _T_6021 | _T_6026; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_6037 = _T_4552 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_6040 = _T_5526 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_6042 = _T_6040 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_6043 = _T_6037 | _T_6042; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_6053 = _T_4556 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_6056 = _T_5542 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_6058 = _T_6056 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_6059 = _T_6053 | _T_6058; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_6069 = _T_4560 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_6072 = _T_5558 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_6074 = _T_6072 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_6075 = _T_6069 | _T_6074; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_6085 = _T_4564 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_6088 = _T_5574 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_6090 = _T_6088 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_6091 = _T_6085 | _T_6090; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_6101 = _T_4568 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_6104 = _T_5590 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_6106 = _T_6104 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_6107 = _T_6101 | _T_6106; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_6117 = _T_4572 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_6120 = _T_5606 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_6122 = _T_6120 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_6123 = _T_6117 | _T_6122; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_6133 = _T_4576 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_6136 = _T_5622 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_6138 = _T_6136 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_6139 = _T_6133 | _T_6138; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_6149 = _T_4580 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_6152 = _T_5638 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_6154 = _T_6152 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_6155 = _T_6149 | _T_6154; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_6165 = _T_4584 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_6168 = _T_5654 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_6170 = _T_6168 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_6171 = _T_6165 | _T_6170; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_6181 = _T_4588 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_6184 = _T_5670 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_6186 = _T_6184 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_6187 = _T_6181 | _T_6186; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_6197 = _T_4592 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_6200 = _T_5686 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_6202 = _T_6200 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_6203 = _T_6197 | _T_6202; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_6213 = _T_4596 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_6216 = _T_5702 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_6218 = _T_6216 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_6219 = _T_6213 | _T_6218; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_6229 = _T_4600 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_6230 = perr_ic_index_ff == 6'h20; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_6232 = _T_6230 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_6234 = _T_6232 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_6235 = _T_6229 | _T_6234; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_6245 = _T_4604 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_6246 = perr_ic_index_ff == 6'h21; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_6248 = _T_6246 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_6250 = _T_6248 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_6251 = _T_6245 | _T_6250; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_6261 = _T_4608 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_6262 = perr_ic_index_ff == 6'h22; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_6264 = _T_6262 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_6266 = _T_6264 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_6267 = _T_6261 | _T_6266; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_6277 = _T_4612 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_6278 = perr_ic_index_ff == 6'h23; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_6280 = _T_6278 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_6282 = _T_6280 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_6283 = _T_6277 | _T_6282; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_6293 = _T_4616 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_6294 = perr_ic_index_ff == 6'h24; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_6296 = _T_6294 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_6298 = _T_6296 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_6299 = _T_6293 | _T_6298; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_6309 = _T_4620 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_6310 = perr_ic_index_ff == 6'h25; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_6312 = _T_6310 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_6314 = _T_6312 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_6315 = _T_6309 | _T_6314; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_6325 = _T_4624 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_6326 = perr_ic_index_ff == 6'h26; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_6328 = _T_6326 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_6330 = _T_6328 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_6331 = _T_6325 | _T_6330; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_6341 = _T_4628 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_6342 = perr_ic_index_ff == 6'h27; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_6344 = _T_6342 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_6346 = _T_6344 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_6347 = _T_6341 | _T_6346; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_6357 = _T_4632 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_6358 = perr_ic_index_ff == 6'h28; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_6360 = _T_6358 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_6362 = _T_6360 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_6363 = _T_6357 | _T_6362; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_6373 = _T_4636 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_6374 = perr_ic_index_ff == 6'h29; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_6376 = _T_6374 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_6378 = _T_6376 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_6379 = _T_6373 | _T_6378; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_6389 = _T_4640 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_6390 = perr_ic_index_ff == 6'h2a; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_6392 = _T_6390 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_6394 = _T_6392 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_6395 = _T_6389 | _T_6394; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_6405 = _T_4644 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_6406 = perr_ic_index_ff == 6'h2b; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_6408 = _T_6406 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_6410 = _T_6408 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_6411 = _T_6405 | _T_6410; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_6421 = _T_4648 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_6422 = perr_ic_index_ff == 6'h2c; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_6424 = _T_6422 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_6426 = _T_6424 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_6427 = _T_6421 | _T_6426; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_6437 = _T_4652 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_6438 = perr_ic_index_ff == 6'h2d; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_6440 = _T_6438 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_6442 = _T_6440 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_6443 = _T_6437 | _T_6442; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_6453 = _T_4656 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_6454 = perr_ic_index_ff == 6'h2e; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_6456 = _T_6454 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_6458 = _T_6456 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_6459 = _T_6453 | _T_6458; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_6469 = _T_4660 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_6470 = perr_ic_index_ff == 6'h2f; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_6472 = _T_6470 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_6474 = _T_6472 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_6475 = _T_6469 | _T_6474; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_6485 = _T_4664 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_6486 = perr_ic_index_ff == 6'h30; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_6488 = _T_6486 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_6490 = _T_6488 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_6491 = _T_6485 | _T_6490; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_6501 = _T_4668 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_6502 = perr_ic_index_ff == 6'h31; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_6504 = _T_6502 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_6506 = _T_6504 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_6507 = _T_6501 | _T_6506; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_6517 = _T_4672 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_6518 = perr_ic_index_ff == 6'h32; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_6520 = _T_6518 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_6522 = _T_6520 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_6523 = _T_6517 | _T_6522; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_6533 = _T_4676 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_6534 = perr_ic_index_ff == 6'h33; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_6536 = _T_6534 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_6538 = _T_6536 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_6539 = _T_6533 | _T_6538; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_6549 = _T_4680 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_6550 = perr_ic_index_ff == 6'h34; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_6552 = _T_6550 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_6554 = _T_6552 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_6555 = _T_6549 | _T_6554; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_6565 = _T_4684 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_6566 = perr_ic_index_ff == 6'h35; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_6568 = _T_6566 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_6570 = _T_6568 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_6571 = _T_6565 | _T_6570; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_6581 = _T_4688 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_6582 = perr_ic_index_ff == 6'h36; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_6584 = _T_6582 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_6586 = _T_6584 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_6587 = _T_6581 | _T_6586; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_6597 = _T_4692 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_6598 = perr_ic_index_ff == 6'h37; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_6600 = _T_6598 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_6602 = _T_6600 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_6603 = _T_6597 | _T_6602; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_6613 = _T_4696 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_6614 = perr_ic_index_ff == 6'h38; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_6616 = _T_6614 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_6618 = _T_6616 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_6619 = _T_6613 | _T_6618; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_6629 = _T_4700 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_6630 = perr_ic_index_ff == 6'h39; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_6632 = _T_6630 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_6634 = _T_6632 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_6635 = _T_6629 | _T_6634; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_6645 = _T_4704 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_6646 = perr_ic_index_ff == 6'h3a; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_6648 = _T_6646 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_6650 = _T_6648 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_6651 = _T_6645 | _T_6650; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_6661 = _T_4708 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_6662 = perr_ic_index_ff == 6'h3b; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_6664 = _T_6662 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_6666 = _T_6664 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_6667 = _T_6661 | _T_6666; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_6677 = _T_4712 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_6678 = perr_ic_index_ff == 6'h3c; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_6680 = _T_6678 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_6682 = _T_6680 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_6683 = _T_6677 | _T_6682; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_6693 = _T_4716 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_6694 = perr_ic_index_ff == 6'h3d; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_6696 = _T_6694 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_6698 = _T_6696 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_6699 = _T_6693 | _T_6698; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_6709 = _T_4720 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_6710 = perr_ic_index_ff == 6'h3e; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_6712 = _T_6710 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_6714 = _T_6712 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_6715 = _T_6709 | _T_6714; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_6725 = _T_4724 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_6726 = perr_ic_index_ff == 6'h3f; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_6728 = _T_6726 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_6730 = _T_6728 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_6731 = _T_6725 | _T_6730; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_6741 = _T_4600 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_6744 = _T_6230 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_6746 = _T_6744 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_6747 = _T_6741 | _T_6746; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_6757 = _T_4604 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_6760 = _T_6246 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_6762 = _T_6760 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_6763 = _T_6757 | _T_6762; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_6773 = _T_4608 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_6776 = _T_6262 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_6778 = _T_6776 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_6779 = _T_6773 | _T_6778; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_6789 = _T_4612 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_6792 = _T_6278 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_6794 = _T_6792 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_6795 = _T_6789 | _T_6794; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_6805 = _T_4616 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_6808 = _T_6294 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_6810 = _T_6808 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_6811 = _T_6805 | _T_6810; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_6821 = _T_4620 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_6824 = _T_6310 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_6826 = _T_6824 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_6827 = _T_6821 | _T_6826; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_6837 = _T_4624 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_6840 = _T_6326 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_6842 = _T_6840 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_6843 = _T_6837 | _T_6842; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_6853 = _T_4628 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_6856 = _T_6342 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_6858 = _T_6856 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_6859 = _T_6853 | _T_6858; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_6869 = _T_4632 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_6872 = _T_6358 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_6874 = _T_6872 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_6875 = _T_6869 | _T_6874; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_6885 = _T_4636 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_6888 = _T_6374 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_6890 = _T_6888 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_6891 = _T_6885 | _T_6890; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_6901 = _T_4640 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_6904 = _T_6390 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_6906 = _T_6904 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_6907 = _T_6901 | _T_6906; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_6917 = _T_4644 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_6920 = _T_6406 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_6922 = _T_6920 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_6923 = _T_6917 | _T_6922; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_6933 = _T_4648 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_6936 = _T_6422 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_6938 = _T_6936 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_6939 = _T_6933 | _T_6938; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_6949 = _T_4652 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_6952 = _T_6438 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_6954 = _T_6952 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_6955 = _T_6949 | _T_6954; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_6965 = _T_4656 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_6968 = _T_6454 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_6970 = _T_6968 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_6971 = _T_6965 | _T_6970; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_6981 = _T_4660 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_6984 = _T_6470 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_6986 = _T_6984 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_6987 = _T_6981 | _T_6986; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_6997 = _T_4664 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_7000 = _T_6486 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_7002 = _T_7000 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_7003 = _T_6997 | _T_7002; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_7013 = _T_4668 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_7016 = _T_6502 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_7018 = _T_7016 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_7019 = _T_7013 | _T_7018; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_7029 = _T_4672 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_7032 = _T_6518 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_7034 = _T_7032 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_7035 = _T_7029 | _T_7034; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_7045 = _T_4676 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_7048 = _T_6534 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_7050 = _T_7048 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_7051 = _T_7045 | _T_7050; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_7061 = _T_4680 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_7064 = _T_6550 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_7066 = _T_7064 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_7067 = _T_7061 | _T_7066; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_7077 = _T_4684 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_7080 = _T_6566 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_7082 = _T_7080 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_7083 = _T_7077 | _T_7082; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_7093 = _T_4688 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_7096 = _T_6582 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_7098 = _T_7096 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_7099 = _T_7093 | _T_7098; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_7109 = _T_4692 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_7112 = _T_6598 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_7114 = _T_7112 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_7115 = _T_7109 | _T_7114; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_7125 = _T_4696 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_7128 = _T_6614 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_7130 = _T_7128 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_7131 = _T_7125 | _T_7130; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_7141 = _T_4700 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_7144 = _T_6630 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_7146 = _T_7144 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_7147 = _T_7141 | _T_7146; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_7157 = _T_4704 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_7160 = _T_6646 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_7162 = _T_7160 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_7163 = _T_7157 | _T_7162; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_7173 = _T_4708 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_7176 = _T_6662 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_7178 = _T_7176 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_7179 = _T_7173 | _T_7178; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_7189 = _T_4712 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_7192 = _T_6678 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_7194 = _T_7192 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_7195 = _T_7189 | _T_7194; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_7205 = _T_4716 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_7208 = _T_6694 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_7210 = _T_7208 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_7211 = _T_7205 | _T_7210; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_7221 = _T_4720 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_7224 = _T_6710 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_7226 = _T_7224 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_7227 = _T_7221 | _T_7226; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_7237 = _T_4724 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_7240 = _T_6726 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_7242 = _T_7240 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_7243 = _T_7237 | _T_7242; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_7253 = _T_4728 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire [6:0] _GEN_796 = {{1'd0}, perr_ic_index_ff}; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_7254 = _GEN_796 == 7'h40; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_7256 = _T_7254 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_7258 = _T_7256 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_7259 = _T_7253 | _T_7258; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_7269 = _T_4732 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_7270 = _GEN_796 == 7'h41; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_7272 = _T_7270 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_7274 = _T_7272 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_7275 = _T_7269 | _T_7274; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_7285 = _T_4736 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_7286 = _GEN_796 == 7'h42; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_7288 = _T_7286 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_7290 = _T_7288 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_7291 = _T_7285 | _T_7290; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_7301 = _T_4740 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_7302 = _GEN_796 == 7'h43; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_7304 = _T_7302 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_7306 = _T_7304 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_7307 = _T_7301 | _T_7306; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_7317 = _T_4744 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_7318 = _GEN_796 == 7'h44; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_7320 = _T_7318 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_7322 = _T_7320 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_7323 = _T_7317 | _T_7322; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_7333 = _T_4748 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_7334 = _GEN_796 == 7'h45; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_7336 = _T_7334 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_7338 = _T_7336 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_7339 = _T_7333 | _T_7338; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_7349 = _T_4752 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_7350 = _GEN_796 == 7'h46; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_7352 = _T_7350 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_7354 = _T_7352 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_7355 = _T_7349 | _T_7354; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_7365 = _T_4756 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_7366 = _GEN_796 == 7'h47; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_7368 = _T_7366 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_7370 = _T_7368 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_7371 = _T_7365 | _T_7370; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_7381 = _T_4760 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_7382 = _GEN_796 == 7'h48; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_7384 = _T_7382 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_7386 = _T_7384 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_7387 = _T_7381 | _T_7386; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_7397 = _T_4764 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_7398 = _GEN_796 == 7'h49; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_7400 = _T_7398 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_7402 = _T_7400 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_7403 = _T_7397 | _T_7402; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_7413 = _T_4768 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_7414 = _GEN_796 == 7'h4a; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_7416 = _T_7414 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_7418 = _T_7416 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_7419 = _T_7413 | _T_7418; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_7429 = _T_4772 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_7430 = _GEN_796 == 7'h4b; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_7432 = _T_7430 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_7434 = _T_7432 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_7435 = _T_7429 | _T_7434; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_7445 = _T_4776 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_7446 = _GEN_796 == 7'h4c; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_7448 = _T_7446 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_7450 = _T_7448 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_7451 = _T_7445 | _T_7450; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_7461 = _T_4780 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_7462 = _GEN_796 == 7'h4d; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_7464 = _T_7462 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_7466 = _T_7464 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_7467 = _T_7461 | _T_7466; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_7477 = _T_4784 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_7478 = _GEN_796 == 7'h4e; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_7480 = _T_7478 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_7482 = _T_7480 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_7483 = _T_7477 | _T_7482; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_7493 = _T_4788 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_7494 = _GEN_796 == 7'h4f; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_7496 = _T_7494 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_7498 = _T_7496 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_7499 = _T_7493 | _T_7498; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_7509 = _T_4792 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_7510 = _GEN_796 == 7'h50; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_7512 = _T_7510 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_7514 = _T_7512 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_7515 = _T_7509 | _T_7514; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_7525 = _T_4796 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_7526 = _GEN_796 == 7'h51; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_7528 = _T_7526 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_7530 = _T_7528 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_7531 = _T_7525 | _T_7530; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_7541 = _T_4800 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_7542 = _GEN_796 == 7'h52; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_7544 = _T_7542 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_7546 = _T_7544 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_7547 = _T_7541 | _T_7546; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_7557 = _T_4804 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_7558 = _GEN_796 == 7'h53; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_7560 = _T_7558 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_7562 = _T_7560 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_7563 = _T_7557 | _T_7562; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_7573 = _T_4808 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_7574 = _GEN_796 == 7'h54; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_7576 = _T_7574 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_7578 = _T_7576 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_7579 = _T_7573 | _T_7578; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_7589 = _T_4812 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_7590 = _GEN_796 == 7'h55; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_7592 = _T_7590 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_7594 = _T_7592 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_7595 = _T_7589 | _T_7594; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_7605 = _T_4816 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_7606 = _GEN_796 == 7'h56; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_7608 = _T_7606 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_7610 = _T_7608 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_7611 = _T_7605 | _T_7610; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_7621 = _T_4820 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_7622 = _GEN_796 == 7'h57; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_7624 = _T_7622 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_7626 = _T_7624 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_7627 = _T_7621 | _T_7626; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_7637 = _T_4824 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_7638 = _GEN_796 == 7'h58; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_7640 = _T_7638 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_7642 = _T_7640 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_7643 = _T_7637 | _T_7642; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_7653 = _T_4828 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_7654 = _GEN_796 == 7'h59; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_7656 = _T_7654 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_7658 = _T_7656 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_7659 = _T_7653 | _T_7658; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_7669 = _T_4832 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_7670 = _GEN_796 == 7'h5a; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_7672 = _T_7670 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_7674 = _T_7672 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_7675 = _T_7669 | _T_7674; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_7685 = _T_4836 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_7686 = _GEN_796 == 7'h5b; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_7688 = _T_7686 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_7690 = _T_7688 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_7691 = _T_7685 | _T_7690; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_7701 = _T_4840 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_7702 = _GEN_796 == 7'h5c; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_7704 = _T_7702 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_7706 = _T_7704 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_7707 = _T_7701 | _T_7706; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_7717 = _T_4844 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_7718 = _GEN_796 == 7'h5d; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_7720 = _T_7718 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_7722 = _T_7720 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_7723 = _T_7717 | _T_7722; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_7733 = _T_4848 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_7734 = _GEN_796 == 7'h5e; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_7736 = _T_7734 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_7738 = _T_7736 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_7739 = _T_7733 | _T_7738; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_7749 = _T_4852 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_7750 = _GEN_796 == 7'h5f; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_7752 = _T_7750 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_7754 = _T_7752 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_7755 = _T_7749 | _T_7754; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_7765 = _T_4728 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_7768 = _T_7254 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_7770 = _T_7768 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_7771 = _T_7765 | _T_7770; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_7781 = _T_4732 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_7784 = _T_7270 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_7786 = _T_7784 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_7787 = _T_7781 | _T_7786; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_7797 = _T_4736 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_7800 = _T_7286 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_7802 = _T_7800 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_7803 = _T_7797 | _T_7802; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_7813 = _T_4740 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_7816 = _T_7302 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_7818 = _T_7816 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_7819 = _T_7813 | _T_7818; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_7829 = _T_4744 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_7832 = _T_7318 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_7834 = _T_7832 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_7835 = _T_7829 | _T_7834; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_7845 = _T_4748 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_7848 = _T_7334 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_7850 = _T_7848 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_7851 = _T_7845 | _T_7850; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_7861 = _T_4752 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_7864 = _T_7350 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_7866 = _T_7864 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_7867 = _T_7861 | _T_7866; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_7877 = _T_4756 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_7880 = _T_7366 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_7882 = _T_7880 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_7883 = _T_7877 | _T_7882; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_7893 = _T_4760 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_7896 = _T_7382 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_7898 = _T_7896 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_7899 = _T_7893 | _T_7898; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_7909 = _T_4764 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_7912 = _T_7398 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_7914 = _T_7912 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_7915 = _T_7909 | _T_7914; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_7925 = _T_4768 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_7928 = _T_7414 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_7930 = _T_7928 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_7931 = _T_7925 | _T_7930; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_7941 = _T_4772 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_7944 = _T_7430 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_7946 = _T_7944 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_7947 = _T_7941 | _T_7946; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_7957 = _T_4776 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_7960 = _T_7446 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_7962 = _T_7960 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_7963 = _T_7957 | _T_7962; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_7973 = _T_4780 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_7976 = _T_7462 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_7978 = _T_7976 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_7979 = _T_7973 | _T_7978; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_7989 = _T_4784 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_7992 = _T_7478 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_7994 = _T_7992 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_7995 = _T_7989 | _T_7994; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_8005 = _T_4788 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_8008 = _T_7494 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_8010 = _T_8008 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_8011 = _T_8005 | _T_8010; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_8021 = _T_4792 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_8024 = _T_7510 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_8026 = _T_8024 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_8027 = _T_8021 | _T_8026; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_8037 = _T_4796 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_8040 = _T_7526 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_8042 = _T_8040 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_8043 = _T_8037 | _T_8042; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_8053 = _T_4800 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_8056 = _T_7542 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_8058 = _T_8056 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_8059 = _T_8053 | _T_8058; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_8069 = _T_4804 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_8072 = _T_7558 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_8074 = _T_8072 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_8075 = _T_8069 | _T_8074; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_8085 = _T_4808 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_8088 = _T_7574 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_8090 = _T_8088 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_8091 = _T_8085 | _T_8090; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_8101 = _T_4812 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_8104 = _T_7590 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_8106 = _T_8104 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_8107 = _T_8101 | _T_8106; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_8117 = _T_4816 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_8120 = _T_7606 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_8122 = _T_8120 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_8123 = _T_8117 | _T_8122; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_8133 = _T_4820 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_8136 = _T_7622 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_8138 = _T_8136 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_8139 = _T_8133 | _T_8138; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_8149 = _T_4824 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_8152 = _T_7638 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_8154 = _T_8152 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_8155 = _T_8149 | _T_8154; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_8165 = _T_4828 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_8168 = _T_7654 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_8170 = _T_8168 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_8171 = _T_8165 | _T_8170; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_8181 = _T_4832 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_8184 = _T_7670 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_8186 = _T_8184 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_8187 = _T_8181 | _T_8186; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_8197 = _T_4836 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_8200 = _T_7686 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_8202 = _T_8200 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_8203 = _T_8197 | _T_8202; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_8213 = _T_4840 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_8216 = _T_7702 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_8218 = _T_8216 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_8219 = _T_8213 | _T_8218; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_8229 = _T_4844 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_8232 = _T_7718 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_8234 = _T_8232 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_8235 = _T_8229 | _T_8234; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_8245 = _T_4848 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_8248 = _T_7734 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_8250 = _T_8248 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_8251 = _T_8245 | _T_8250; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_8261 = _T_4852 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_8264 = _T_7750 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_8266 = _T_8264 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_8267 = _T_8261 | _T_8266; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_8277 = _T_4856 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_8278 = _GEN_796 == 7'h60; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_8280 = _T_8278 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_8282 = _T_8280 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_8283 = _T_8277 | _T_8282; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_8293 = _T_4860 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_8294 = _GEN_796 == 7'h61; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_8296 = _T_8294 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_8298 = _T_8296 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_8299 = _T_8293 | _T_8298; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_8309 = _T_4864 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_8310 = _GEN_796 == 7'h62; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_8312 = _T_8310 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_8314 = _T_8312 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_8315 = _T_8309 | _T_8314; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_8325 = _T_4868 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_8326 = _GEN_796 == 7'h63; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_8328 = _T_8326 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_8330 = _T_8328 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_8331 = _T_8325 | _T_8330; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_8341 = _T_4872 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_8342 = _GEN_796 == 7'h64; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_8344 = _T_8342 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_8346 = _T_8344 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_8347 = _T_8341 | _T_8346; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_8357 = _T_4876 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_8358 = _GEN_796 == 7'h65; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_8360 = _T_8358 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_8362 = _T_8360 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_8363 = _T_8357 | _T_8362; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_8373 = _T_4880 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_8374 = _GEN_796 == 7'h66; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_8376 = _T_8374 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_8378 = _T_8376 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_8379 = _T_8373 | _T_8378; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_8389 = _T_4884 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_8390 = _GEN_796 == 7'h67; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_8392 = _T_8390 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_8394 = _T_8392 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_8395 = _T_8389 | _T_8394; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_8405 = _T_4888 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_8406 = _GEN_796 == 7'h68; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_8408 = _T_8406 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_8410 = _T_8408 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_8411 = _T_8405 | _T_8410; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_8421 = _T_4892 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_8422 = _GEN_796 == 7'h69; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_8424 = _T_8422 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_8426 = _T_8424 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_8427 = _T_8421 | _T_8426; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_8437 = _T_4896 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_8438 = _GEN_796 == 7'h6a; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_8440 = _T_8438 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_8442 = _T_8440 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_8443 = _T_8437 | _T_8442; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_8453 = _T_4900 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_8454 = _GEN_796 == 7'h6b; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_8456 = _T_8454 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_8458 = _T_8456 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_8459 = _T_8453 | _T_8458; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_8469 = _T_4904 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_8470 = _GEN_796 == 7'h6c; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_8472 = _T_8470 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_8474 = _T_8472 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_8475 = _T_8469 | _T_8474; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_8485 = _T_4908 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_8486 = _GEN_796 == 7'h6d; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_8488 = _T_8486 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_8490 = _T_8488 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_8491 = _T_8485 | _T_8490; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_8501 = _T_4912 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_8502 = _GEN_796 == 7'h6e; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_8504 = _T_8502 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_8506 = _T_8504 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_8507 = _T_8501 | _T_8506; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_8517 = _T_4916 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_8518 = _GEN_796 == 7'h6f; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_8520 = _T_8518 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_8522 = _T_8520 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_8523 = _T_8517 | _T_8522; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_8533 = _T_4920 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_8534 = _GEN_796 == 7'h70; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_8536 = _T_8534 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_8538 = _T_8536 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_8539 = _T_8533 | _T_8538; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_8549 = _T_4924 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_8550 = _GEN_796 == 7'h71; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_8552 = _T_8550 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_8554 = _T_8552 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_8555 = _T_8549 | _T_8554; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_8565 = _T_4928 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_8566 = _GEN_796 == 7'h72; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_8568 = _T_8566 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_8570 = _T_8568 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_8571 = _T_8565 | _T_8570; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_8581 = _T_4932 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_8582 = _GEN_796 == 7'h73; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_8584 = _T_8582 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_8586 = _T_8584 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_8587 = _T_8581 | _T_8586; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_8597 = _T_4936 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_8598 = _GEN_796 == 7'h74; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_8600 = _T_8598 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_8602 = _T_8600 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_8603 = _T_8597 | _T_8602; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_8613 = _T_4940 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_8614 = _GEN_796 == 7'h75; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_8616 = _T_8614 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_8618 = _T_8616 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_8619 = _T_8613 | _T_8618; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_8629 = _T_4944 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_8630 = _GEN_796 == 7'h76; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_8632 = _T_8630 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_8634 = _T_8632 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_8635 = _T_8629 | _T_8634; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_8645 = _T_4948 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_8646 = _GEN_796 == 7'h77; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_8648 = _T_8646 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_8650 = _T_8648 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_8651 = _T_8645 | _T_8650; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_8661 = _T_4952 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_8662 = _GEN_796 == 7'h78; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_8664 = _T_8662 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_8666 = _T_8664 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_8667 = _T_8661 | _T_8666; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_8677 = _T_4956 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_8678 = _GEN_796 == 7'h79; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_8680 = _T_8678 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_8682 = _T_8680 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_8683 = _T_8677 | _T_8682; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_8693 = _T_4960 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_8694 = _GEN_796 == 7'h7a; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_8696 = _T_8694 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_8698 = _T_8696 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_8699 = _T_8693 | _T_8698; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_8709 = _T_4964 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_8710 = _GEN_796 == 7'h7b; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_8712 = _T_8710 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_8714 = _T_8712 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_8715 = _T_8709 | _T_8714; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_8725 = _T_4968 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_8726 = _GEN_796 == 7'h7c; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_8728 = _T_8726 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_8730 = _T_8728 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_8731 = _T_8725 | _T_8730; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_8741 = _T_4972 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_8742 = _GEN_796 == 7'h7d; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_8744 = _T_8742 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_8746 = _T_8744 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_8747 = _T_8741 | _T_8746; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_8757 = _T_4976 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_8758 = _GEN_796 == 7'h7e; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_8760 = _T_8758 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_8762 = _T_8760 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_8763 = _T_8757 | _T_8762; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_8773 = _T_4980 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_8774 = _GEN_796 == 7'h7f; // @[el2_ifu_mem_ctl.scala 741:101]
  wire  _T_8776 = _T_8774 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_8778 = _T_8776 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_8779 = _T_8773 | _T_8778; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_8789 = _T_4856 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_8792 = _T_8278 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_8794 = _T_8792 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_8795 = _T_8789 | _T_8794; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_8805 = _T_4860 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_8808 = _T_8294 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_8810 = _T_8808 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_8811 = _T_8805 | _T_8810; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_8821 = _T_4864 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_8824 = _T_8310 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_8826 = _T_8824 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_8827 = _T_8821 | _T_8826; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_8837 = _T_4868 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_8840 = _T_8326 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_8842 = _T_8840 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_8843 = _T_8837 | _T_8842; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_8853 = _T_4872 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_8856 = _T_8342 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_8858 = _T_8856 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_8859 = _T_8853 | _T_8858; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_8869 = _T_4876 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_8872 = _T_8358 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_8874 = _T_8872 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_8875 = _T_8869 | _T_8874; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_8885 = _T_4880 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_8888 = _T_8374 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_8890 = _T_8888 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_8891 = _T_8885 | _T_8890; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_8901 = _T_4884 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_8904 = _T_8390 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_8906 = _T_8904 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_8907 = _T_8901 | _T_8906; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_8917 = _T_4888 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_8920 = _T_8406 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_8922 = _T_8920 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_8923 = _T_8917 | _T_8922; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_8933 = _T_4892 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_8936 = _T_8422 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_8938 = _T_8936 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_8939 = _T_8933 | _T_8938; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_8949 = _T_4896 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_8952 = _T_8438 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_8954 = _T_8952 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_8955 = _T_8949 | _T_8954; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_8965 = _T_4900 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_8968 = _T_8454 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_8970 = _T_8968 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_8971 = _T_8965 | _T_8970; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_8981 = _T_4904 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_8984 = _T_8470 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_8986 = _T_8984 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_8987 = _T_8981 | _T_8986; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_8997 = _T_4908 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_9000 = _T_8486 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_9002 = _T_9000 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_9003 = _T_8997 | _T_9002; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_9013 = _T_4912 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_9016 = _T_8502 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_9018 = _T_9016 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_9019 = _T_9013 | _T_9018; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_9029 = _T_4916 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_9032 = _T_8518 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_9034 = _T_9032 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_9035 = _T_9029 | _T_9034; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_9045 = _T_4920 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_9048 = _T_8534 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_9050 = _T_9048 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_9051 = _T_9045 | _T_9050; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_9061 = _T_4924 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_9064 = _T_8550 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_9066 = _T_9064 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_9067 = _T_9061 | _T_9066; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_9077 = _T_4928 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_9080 = _T_8566 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_9082 = _T_9080 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_9083 = _T_9077 | _T_9082; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_9093 = _T_4932 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_9096 = _T_8582 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_9098 = _T_9096 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_9099 = _T_9093 | _T_9098; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_9109 = _T_4936 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_9112 = _T_8598 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_9114 = _T_9112 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_9115 = _T_9109 | _T_9114; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_9125 = _T_4940 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_9128 = _T_8614 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_9130 = _T_9128 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_9131 = _T_9125 | _T_9130; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_9141 = _T_4944 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_9144 = _T_8630 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_9146 = _T_9144 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_9147 = _T_9141 | _T_9146; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_9157 = _T_4948 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_9160 = _T_8646 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_9162 = _T_9160 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_9163 = _T_9157 | _T_9162; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_9173 = _T_4952 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_9176 = _T_8662 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_9178 = _T_9176 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_9179 = _T_9173 | _T_9178; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_9189 = _T_4956 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_9192 = _T_8678 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_9194 = _T_9192 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_9195 = _T_9189 | _T_9194; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_9205 = _T_4960 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_9208 = _T_8694 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_9210 = _T_9208 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_9211 = _T_9205 | _T_9210; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_9221 = _T_4964 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_9224 = _T_8710 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_9226 = _T_9224 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_9227 = _T_9221 | _T_9226; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_9237 = _T_4968 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_9240 = _T_8726 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_9242 = _T_9240 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_9243 = _T_9237 | _T_9242; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_9253 = _T_4972 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_9256 = _T_8742 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_9258 = _T_9256 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_9259 = _T_9253 | _T_9258; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_9269 = _T_4976 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_9272 = _T_8758 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_9274 = _T_9272 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_9275 = _T_9269 | _T_9274; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_9285 = _T_4980 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:58]
  wire  _T_9288 = _T_8774 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 741:123]
  wire  _T_9290 = _T_9288 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 741:144]
  wire  _T_9291 = _T_9285 | _T_9290; // @[el2_ifu_mem_ctl.scala 741:80]
  wire  _T_10092 = ~fetch_uncacheable_ff; // @[el2_ifu_mem_ctl.scala 795:63]
  wire  _T_10093 = _T_10092 & ifc_fetch_req_f; // @[el2_ifu_mem_ctl.scala 795:85]
  wire [1:0] _T_10095 = _T_10093 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  reg  _T_10102; // @[el2_ifu_mem_ctl.scala 800:57]
  reg  _T_10103; // @[el2_ifu_mem_ctl.scala 801:56]
  reg  _T_10104; // @[el2_ifu_mem_ctl.scala 802:59]
  wire  _T_10105 = ~ifu_bus_arready_ff; // @[el2_ifu_mem_ctl.scala 803:80]
  wire  _T_10106 = ifu_bus_arvalid_ff & _T_10105; // @[el2_ifu_mem_ctl.scala 803:78]
  wire  _T_10107 = _T_10106 & miss_pending; // @[el2_ifu_mem_ctl.scala 803:100]
  reg  _T_10108; // @[el2_ifu_mem_ctl.scala 803:58]
  reg  _T_10109; // @[el2_ifu_mem_ctl.scala 804:58]
  wire  _T_10112 = io_dec_tlu_ic_diag_pkt_icache_dicawics[15:14] == 2'h3; // @[el2_ifu_mem_ctl.scala 811:71]
  wire  _T_10114 = io_dec_tlu_ic_diag_pkt_icache_dicawics[15:14] == 2'h2; // @[el2_ifu_mem_ctl.scala 811:124]
  wire  _T_10116 = io_dec_tlu_ic_diag_pkt_icache_dicawics[15:14] == 2'h1; // @[el2_ifu_mem_ctl.scala 812:50]
  wire  _T_10118 = io_dec_tlu_ic_diag_pkt_icache_dicawics[15:14] == 2'h0; // @[el2_ifu_mem_ctl.scala 812:103]
  wire [3:0] _T_10121 = {_T_10112,_T_10114,_T_10116,_T_10118}; // @[Cat.scala 29:58]
  wire  ic_debug_ict_array_sel_in = io_ic_debug_rd_en & io_ic_debug_tag_array; // @[el2_ifu_mem_ctl.scala 814:53]
  reg  _T_10132; // @[Reg.scala 27:20]
  assign io_ifu_miss_state_idle = miss_state == 3'h0; // @[el2_ifu_mem_ctl.scala 323:26]
  assign io_ifu_ic_mb_empty = _T_327 | _T_232; // @[el2_ifu_mem_ctl.scala 322:22]
  assign io_ic_dma_active = _T_11 | io_dec_tlu_flush_err_wb; // @[el2_ifu_mem_ctl.scala 187:20]
  assign io_ic_write_stall = write_ic_16_bytes & _T_3927; // @[el2_ifu_mem_ctl.scala 691:21]
  assign io_ifu_pmu_ic_miss = _T_10102; // @[el2_ifu_mem_ctl.scala 800:22]
  assign io_ifu_pmu_ic_hit = _T_10103; // @[el2_ifu_mem_ctl.scala 801:21]
  assign io_ifu_pmu_bus_error = _T_10104; // @[el2_ifu_mem_ctl.scala 802:24]
  assign io_ifu_pmu_bus_busy = _T_10108; // @[el2_ifu_mem_ctl.scala 803:23]
  assign io_ifu_pmu_bus_trxn = _T_10109; // @[el2_ifu_mem_ctl.scala 804:23]
  assign io_ifu_axi_awvalid = 1'h0; // @[el2_ifu_mem_ctl.scala 138:22]
  assign io_ifu_axi_awid = 3'h0; // @[el2_ifu_mem_ctl.scala 137:19]
  assign io_ifu_axi_awaddr = 32'h0; // @[el2_ifu_mem_ctl.scala 132:21]
  assign io_ifu_axi_awregion = 4'h0; // @[el2_ifu_mem_ctl.scala 136:23]
  assign io_ifu_axi_awlen = 8'h0; // @[el2_ifu_mem_ctl.scala 134:20]
  assign io_ifu_axi_awsize = 3'h0; // @[el2_ifu_mem_ctl.scala 145:21]
  assign io_ifu_axi_awburst = 2'h0; // @[el2_ifu_mem_ctl.scala 147:22]
  assign io_ifu_axi_awlock = 1'h0; // @[el2_ifu_mem_ctl.scala 142:21]
  assign io_ifu_axi_awcache = 4'h0; // @[el2_ifu_mem_ctl.scala 140:22]
  assign io_ifu_axi_awprot = 3'h0; // @[el2_ifu_mem_ctl.scala 133:21]
  assign io_ifu_axi_awqos = 4'h0; // @[el2_ifu_mem_ctl.scala 131:20]
  assign io_ifu_axi_wvalid = 1'h0; // @[el2_ifu_mem_ctl.scala 129:21]
  assign io_ifu_axi_wdata = 64'h0; // @[el2_ifu_mem_ctl.scala 130:20]
  assign io_ifu_axi_wstrb = 8'h0; // @[el2_ifu_mem_ctl.scala 139:20]
  assign io_ifu_axi_wlast = 1'h0; // @[el2_ifu_mem_ctl.scala 148:20]
  assign io_ifu_axi_bready = 1'h0; // @[el2_ifu_mem_ctl.scala 143:21]
  assign io_ifu_axi_arvalid = ifu_bus_cmd_valid; // @[el2_ifu_mem_ctl.scala 553:22]
  assign io_ifu_axi_arid = bus_rd_addr_count & _T_2521; // @[el2_ifu_mem_ctl.scala 554:19]
  assign io_ifu_axi_araddr = _T_2523 & _T_2525; // @[el2_ifu_mem_ctl.scala 555:21]
  assign io_ifu_axi_arregion = ifu_ic_req_addr_f[28:25]; // @[el2_ifu_mem_ctl.scala 558:23]
  assign io_ifu_axi_arlen = 8'h0; // @[el2_ifu_mem_ctl.scala 144:20]
  assign io_ifu_axi_arsize = 3'h3; // @[el2_ifu_mem_ctl.scala 556:21]
  assign io_ifu_axi_arburst = 2'h1; // @[el2_ifu_mem_ctl.scala 559:22]
  assign io_ifu_axi_arlock = 1'h0; // @[el2_ifu_mem_ctl.scala 135:21]
  assign io_ifu_axi_arcache = 4'hf; // @[el2_ifu_mem_ctl.scala 557:22]
  assign io_ifu_axi_arprot = 3'h0; // @[el2_ifu_mem_ctl.scala 146:21]
  assign io_ifu_axi_arqos = 4'h0; // @[el2_ifu_mem_ctl.scala 141:20]
  assign io_ifu_axi_rready = 1'h1; // @[el2_ifu_mem_ctl.scala 560:21]
  assign io_iccm_dma_ecc_error = |iccm_double_ecc_error; // @[el2_ifu_mem_ctl.scala 650:25]
  assign io_iccm_dma_rvalid = iccm_dma_rvalid; // @[el2_ifu_mem_ctl.scala 648:22]
  assign io_iccm_dma_rdata = iccm_dma_rdata; // @[el2_ifu_mem_ctl.scala 652:21]
  assign io_iccm_dma_rtag = iccm_dma_rtag; // @[el2_ifu_mem_ctl.scala 643:20]
  assign io_iccm_ready = _T_2624 & _T_2618; // @[el2_ifu_mem_ctl.scala 623:17]
  assign io_ic_rw_addr = _T_341 | _T_342; // @[el2_ifu_mem_ctl.scala 332:17]
  assign io_ic_wr_en = 2'h0; // @[el2_ifu_mem_ctl.scala 690:15]
  assign io_ic_rd_en = _T_3905 | _T_3910; // @[el2_ifu_mem_ctl.scala 681:15]
  assign io_ic_wr_data_0 = ic_wr_16bytes_data[70:0]; // @[el2_ifu_mem_ctl.scala 339:17]
  assign io_ic_wr_data_1 = ic_wr_16bytes_data[141:71]; // @[el2_ifu_mem_ctl.scala 339:17]
  assign io_ic_debug_wr_data = io_dec_tlu_ic_diag_pkt_icache_wrdata; // @[el2_ifu_mem_ctl.scala 340:23]
  assign io_ifu_ic_debug_rd_data = _T_1212; // @[el2_ifu_mem_ctl.scala 348:27]
  assign io_ic_debug_addr = io_dec_tlu_ic_diag_pkt_icache_dicawics[9:0]; // @[el2_ifu_mem_ctl.scala 807:20]
  assign io_ic_debug_rd_en = io_dec_tlu_ic_diag_pkt_icache_rd_valid; // @[el2_ifu_mem_ctl.scala 809:21]
  assign io_ic_debug_wr_en = io_dec_tlu_ic_diag_pkt_icache_wr_valid; // @[el2_ifu_mem_ctl.scala 810:21]
  assign io_ic_debug_tag_array = io_dec_tlu_ic_diag_pkt_icache_dicawics[16]; // @[el2_ifu_mem_ctl.scala 808:25]
  assign io_ic_debug_way = _T_10121[1:0]; // @[el2_ifu_mem_ctl.scala 811:19]
  assign io_ic_tag_valid = ic_tag_valid_unq & _T_10095; // @[el2_ifu_mem_ctl.scala 795:19]
  assign io_iccm_rw_addr = _T_3059[14:0]; // @[el2_ifu_mem_ctl.scala 654:19]
  assign io_iccm_wren = _T_2628 | iccm_correct_ecc; // @[el2_ifu_mem_ctl.scala 625:16]
  assign io_iccm_rden = _T_2632 | _T_2633; // @[el2_ifu_mem_ctl.scala 626:16]
  assign io_iccm_wr_data = _T_3034 ? _T_3035 : _T_3042; // @[el2_ifu_mem_ctl.scala 631:19]
  assign io_iccm_wr_size = _T_2638 & io_dma_mem_sz; // @[el2_ifu_mem_ctl.scala 628:19]
  assign io_ic_hit_f = _T_264 | _T_265; // @[el2_ifu_mem_ctl.scala 284:15]
  assign io_ic_access_fault_f = _T_2406 & _T_318; // @[el2_ifu_mem_ctl.scala 379:24]
  assign io_ic_access_fault_type_f = io_iccm_rd_ecc_double_err ? 2'h1 : _T_1276; // @[el2_ifu_mem_ctl.scala 380:29]
  assign io_iccm_rd_ecc_single_err = _T_3850 & ifc_fetch_req_f; // @[el2_ifu_mem_ctl.scala 667:29]
  assign io_iccm_rd_ecc_double_err = iccm_dma_ecc_error_in & ifc_iccm_access_f; // @[el2_ifu_mem_ctl.scala 668:29]
  assign io_ic_error_start = _T_1200 | ic_rd_parity_final_err; // @[el2_ifu_mem_ctl.scala 342:21]
  assign io_ifu_async_error_start = io_iccm_rd_ecc_single_err | io_ic_error_start; // @[el2_ifu_mem_ctl.scala 186:28]
  assign io_iccm_dma_sb_error = _T_3 & dma_iccm_req_f; // @[el2_ifu_mem_ctl.scala 185:24]
  assign io_ic_fetch_val_f = {1'h0,fetch_req_f_qual}; // @[el2_ifu_mem_ctl.scala 384:21]
  assign io_ic_data_f = io_ic_rd_data[31:0]; // @[el2_ifu_mem_ctl.scala 376:16]
  assign io_ic_premux_data = ic_premux_data[63:0]; // @[el2_ifu_mem_ctl.scala 373:21]
  assign io_ic_sel_premux_data = fetch_req_iccm_f | sel_byp_data; // @[el2_ifu_mem_ctl.scala 374:25]
  assign io_ifu_ic_debug_rd_data_valid = _T_10132; // @[el2_ifu_mem_ctl.scala 818:33]
  assign io_iccm_buf_correct_ecc = iccm_correct_ecc & _T_2411; // @[el2_ifu_mem_ctl.scala 472:27]
  assign io_iccm_correction_state = _T_2439 ? 1'h0 : _GEN_59; // @[el2_ifu_mem_ctl.scala 507:28 el2_ifu_mem_ctl.scala 520:32 el2_ifu_mem_ctl.scala 527:32 el2_ifu_mem_ctl.scala 534:32]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  flush_final_f = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  ifc_fetch_req_f_raw = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  miss_state = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  scnd_miss_req_q = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  ifu_fetch_addr_int_f = _RAND_4[30:0];
  _RAND_5 = {1{`RANDOM}};
  ifc_iccm_access_f = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  iccm_dma_rvalid_in = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  dma_iccm_req_f = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  perr_state = _RAND_8[2:0];
  _RAND_9 = {1{`RANDOM}};
  err_stop_state = _RAND_9[1:0];
  _RAND_10 = {1{`RANDOM}};
  reset_all_tags = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  ifc_region_acc_fault_final_f = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  ifu_bus_rvalid_unq_ff = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  bus_ifu_bus_clk_en_ff = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  uncacheable_miss_ff = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  bus_data_beat_count = _RAND_15[2:0];
  _RAND_16 = {1{`RANDOM}};
  ic_miss_buff_data_valid = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  imb_ff = _RAND_17[30:0];
  _RAND_18 = {1{`RANDOM}};
  last_data_recieved_ff = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  sel_mb_addr_ff = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  way_status_mb_scnd_ff = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  _T_5115 = _RAND_21[6:0];
  _RAND_22 = {1{`RANDOM}};
  _T_4471 = _RAND_22[2:0];
  _RAND_23 = {1{`RANDOM}};
  _T_4467 = _RAND_23[2:0];
  _RAND_24 = {1{`RANDOM}};
  _T_4463 = _RAND_24[2:0];
  _RAND_25 = {1{`RANDOM}};
  _T_4459 = _RAND_25[2:0];
  _RAND_26 = {1{`RANDOM}};
  _T_4455 = _RAND_26[2:0];
  _RAND_27 = {1{`RANDOM}};
  _T_4451 = _RAND_27[2:0];
  _RAND_28 = {1{`RANDOM}};
  _T_4447 = _RAND_28[2:0];
  _RAND_29 = {1{`RANDOM}};
  _T_4443 = _RAND_29[2:0];
  _RAND_30 = {1{`RANDOM}};
  _T_4439 = _RAND_30[2:0];
  _RAND_31 = {1{`RANDOM}};
  _T_4435 = _RAND_31[2:0];
  _RAND_32 = {1{`RANDOM}};
  _T_4431 = _RAND_32[2:0];
  _RAND_33 = {1{`RANDOM}};
  _T_4427 = _RAND_33[2:0];
  _RAND_34 = {1{`RANDOM}};
  _T_4423 = _RAND_34[2:0];
  _RAND_35 = {1{`RANDOM}};
  _T_4419 = _RAND_35[2:0];
  _RAND_36 = {1{`RANDOM}};
  _T_4415 = _RAND_36[2:0];
  _RAND_37 = {1{`RANDOM}};
  _T_4411 = _RAND_37[2:0];
  _RAND_38 = {1{`RANDOM}};
  _T_4407 = _RAND_38[2:0];
  _RAND_39 = {1{`RANDOM}};
  _T_4403 = _RAND_39[2:0];
  _RAND_40 = {1{`RANDOM}};
  _T_4399 = _RAND_40[2:0];
  _RAND_41 = {1{`RANDOM}};
  _T_4395 = _RAND_41[2:0];
  _RAND_42 = {1{`RANDOM}};
  _T_4391 = _RAND_42[2:0];
  _RAND_43 = {1{`RANDOM}};
  _T_4387 = _RAND_43[2:0];
  _RAND_44 = {1{`RANDOM}};
  _T_4383 = _RAND_44[2:0];
  _RAND_45 = {1{`RANDOM}};
  _T_4379 = _RAND_45[2:0];
  _RAND_46 = {1{`RANDOM}};
  _T_4375 = _RAND_46[2:0];
  _RAND_47 = {1{`RANDOM}};
  _T_4371 = _RAND_47[2:0];
  _RAND_48 = {1{`RANDOM}};
  _T_4367 = _RAND_48[2:0];
  _RAND_49 = {1{`RANDOM}};
  _T_4363 = _RAND_49[2:0];
  _RAND_50 = {1{`RANDOM}};
  _T_4359 = _RAND_50[2:0];
  _RAND_51 = {1{`RANDOM}};
  _T_4355 = _RAND_51[2:0];
  _RAND_52 = {1{`RANDOM}};
  _T_4351 = _RAND_52[2:0];
  _RAND_53 = {1{`RANDOM}};
  _T_4347 = _RAND_53[2:0];
  _RAND_54 = {1{`RANDOM}};
  _T_4343 = _RAND_54[2:0];
  _RAND_55 = {1{`RANDOM}};
  _T_4339 = _RAND_55[2:0];
  _RAND_56 = {1{`RANDOM}};
  _T_4335 = _RAND_56[2:0];
  _RAND_57 = {1{`RANDOM}};
  _T_4331 = _RAND_57[2:0];
  _RAND_58 = {1{`RANDOM}};
  _T_4327 = _RAND_58[2:0];
  _RAND_59 = {1{`RANDOM}};
  _T_4323 = _RAND_59[2:0];
  _RAND_60 = {1{`RANDOM}};
  _T_4319 = _RAND_60[2:0];
  _RAND_61 = {1{`RANDOM}};
  _T_4315 = _RAND_61[2:0];
  _RAND_62 = {1{`RANDOM}};
  _T_4311 = _RAND_62[2:0];
  _RAND_63 = {1{`RANDOM}};
  _T_4307 = _RAND_63[2:0];
  _RAND_64 = {1{`RANDOM}};
  _T_4303 = _RAND_64[2:0];
  _RAND_65 = {1{`RANDOM}};
  _T_4299 = _RAND_65[2:0];
  _RAND_66 = {1{`RANDOM}};
  _T_4295 = _RAND_66[2:0];
  _RAND_67 = {1{`RANDOM}};
  _T_4291 = _RAND_67[2:0];
  _RAND_68 = {1{`RANDOM}};
  _T_4287 = _RAND_68[2:0];
  _RAND_69 = {1{`RANDOM}};
  _T_4283 = _RAND_69[2:0];
  _RAND_70 = {1{`RANDOM}};
  _T_4279 = _RAND_70[2:0];
  _RAND_71 = {1{`RANDOM}};
  _T_4275 = _RAND_71[2:0];
  _RAND_72 = {1{`RANDOM}};
  _T_4271 = _RAND_72[2:0];
  _RAND_73 = {1{`RANDOM}};
  _T_4267 = _RAND_73[2:0];
  _RAND_74 = {1{`RANDOM}};
  _T_4263 = _RAND_74[2:0];
  _RAND_75 = {1{`RANDOM}};
  _T_4259 = _RAND_75[2:0];
  _RAND_76 = {1{`RANDOM}};
  _T_4255 = _RAND_76[2:0];
  _RAND_77 = {1{`RANDOM}};
  _T_4251 = _RAND_77[2:0];
  _RAND_78 = {1{`RANDOM}};
  _T_4247 = _RAND_78[2:0];
  _RAND_79 = {1{`RANDOM}};
  _T_4243 = _RAND_79[2:0];
  _RAND_80 = {1{`RANDOM}};
  _T_4239 = _RAND_80[2:0];
  _RAND_81 = {1{`RANDOM}};
  _T_4235 = _RAND_81[2:0];
  _RAND_82 = {1{`RANDOM}};
  _T_4231 = _RAND_82[2:0];
  _RAND_83 = {1{`RANDOM}};
  _T_4227 = _RAND_83[2:0];
  _RAND_84 = {1{`RANDOM}};
  _T_4223 = _RAND_84[2:0];
  _RAND_85 = {1{`RANDOM}};
  _T_4219 = _RAND_85[2:0];
  _RAND_86 = {1{`RANDOM}};
  _T_4215 = _RAND_86[2:0];
  _RAND_87 = {1{`RANDOM}};
  _T_4211 = _RAND_87[2:0];
  _RAND_88 = {1{`RANDOM}};
  _T_4207 = _RAND_88[2:0];
  _RAND_89 = {1{`RANDOM}};
  _T_4203 = _RAND_89[2:0];
  _RAND_90 = {1{`RANDOM}};
  _T_4199 = _RAND_90[2:0];
  _RAND_91 = {1{`RANDOM}};
  _T_4195 = _RAND_91[2:0];
  _RAND_92 = {1{`RANDOM}};
  _T_4191 = _RAND_92[2:0];
  _RAND_93 = {1{`RANDOM}};
  _T_4187 = _RAND_93[2:0];
  _RAND_94 = {1{`RANDOM}};
  _T_4183 = _RAND_94[2:0];
  _RAND_95 = {1{`RANDOM}};
  _T_4179 = _RAND_95[2:0];
  _RAND_96 = {1{`RANDOM}};
  _T_4175 = _RAND_96[2:0];
  _RAND_97 = {1{`RANDOM}};
  _T_4171 = _RAND_97[2:0];
  _RAND_98 = {1{`RANDOM}};
  _T_4167 = _RAND_98[2:0];
  _RAND_99 = {1{`RANDOM}};
  _T_4163 = _RAND_99[2:0];
  _RAND_100 = {1{`RANDOM}};
  _T_4159 = _RAND_100[2:0];
  _RAND_101 = {1{`RANDOM}};
  _T_4155 = _RAND_101[2:0];
  _RAND_102 = {1{`RANDOM}};
  _T_4151 = _RAND_102[2:0];
  _RAND_103 = {1{`RANDOM}};
  _T_4147 = _RAND_103[2:0];
  _RAND_104 = {1{`RANDOM}};
  _T_4143 = _RAND_104[2:0];
  _RAND_105 = {1{`RANDOM}};
  _T_4139 = _RAND_105[2:0];
  _RAND_106 = {1{`RANDOM}};
  _T_4135 = _RAND_106[2:0];
  _RAND_107 = {1{`RANDOM}};
  _T_4131 = _RAND_107[2:0];
  _RAND_108 = {1{`RANDOM}};
  _T_4127 = _RAND_108[2:0];
  _RAND_109 = {1{`RANDOM}};
  _T_4123 = _RAND_109[2:0];
  _RAND_110 = {1{`RANDOM}};
  _T_4119 = _RAND_110[2:0];
  _RAND_111 = {1{`RANDOM}};
  _T_4115 = _RAND_111[2:0];
  _RAND_112 = {1{`RANDOM}};
  _T_4111 = _RAND_112[2:0];
  _RAND_113 = {1{`RANDOM}};
  _T_4107 = _RAND_113[2:0];
  _RAND_114 = {1{`RANDOM}};
  _T_4103 = _RAND_114[2:0];
  _RAND_115 = {1{`RANDOM}};
  _T_4099 = _RAND_115[2:0];
  _RAND_116 = {1{`RANDOM}};
  _T_4095 = _RAND_116[2:0];
  _RAND_117 = {1{`RANDOM}};
  _T_4091 = _RAND_117[2:0];
  _RAND_118 = {1{`RANDOM}};
  _T_4087 = _RAND_118[2:0];
  _RAND_119 = {1{`RANDOM}};
  _T_4083 = _RAND_119[2:0];
  _RAND_120 = {1{`RANDOM}};
  _T_4079 = _RAND_120[2:0];
  _RAND_121 = {1{`RANDOM}};
  _T_4075 = _RAND_121[2:0];
  _RAND_122 = {1{`RANDOM}};
  _T_4071 = _RAND_122[2:0];
  _RAND_123 = {1{`RANDOM}};
  _T_4067 = _RAND_123[2:0];
  _RAND_124 = {1{`RANDOM}};
  _T_4063 = _RAND_124[2:0];
  _RAND_125 = {1{`RANDOM}};
  _T_4059 = _RAND_125[2:0];
  _RAND_126 = {1{`RANDOM}};
  _T_4055 = _RAND_126[2:0];
  _RAND_127 = {1{`RANDOM}};
  _T_4051 = _RAND_127[2:0];
  _RAND_128 = {1{`RANDOM}};
  _T_4047 = _RAND_128[2:0];
  _RAND_129 = {1{`RANDOM}};
  _T_4043 = _RAND_129[2:0];
  _RAND_130 = {1{`RANDOM}};
  _T_4039 = _RAND_130[2:0];
  _RAND_131 = {1{`RANDOM}};
  _T_4035 = _RAND_131[2:0];
  _RAND_132 = {1{`RANDOM}};
  _T_4031 = _RAND_132[2:0];
  _RAND_133 = {1{`RANDOM}};
  _T_4027 = _RAND_133[2:0];
  _RAND_134 = {1{`RANDOM}};
  _T_4023 = _RAND_134[2:0];
  _RAND_135 = {1{`RANDOM}};
  _T_4019 = _RAND_135[2:0];
  _RAND_136 = {1{`RANDOM}};
  _T_4015 = _RAND_136[2:0];
  _RAND_137 = {1{`RANDOM}};
  _T_4011 = _RAND_137[2:0];
  _RAND_138 = {1{`RANDOM}};
  _T_4007 = _RAND_138[2:0];
  _RAND_139 = {1{`RANDOM}};
  _T_4003 = _RAND_139[2:0];
  _RAND_140 = {1{`RANDOM}};
  _T_3999 = _RAND_140[2:0];
  _RAND_141 = {1{`RANDOM}};
  _T_3995 = _RAND_141[2:0];
  _RAND_142 = {1{`RANDOM}};
  _T_3991 = _RAND_142[2:0];
  _RAND_143 = {1{`RANDOM}};
  _T_3987 = _RAND_143[2:0];
  _RAND_144 = {1{`RANDOM}};
  _T_3983 = _RAND_144[2:0];
  _RAND_145 = {1{`RANDOM}};
  _T_3979 = _RAND_145[2:0];
  _RAND_146 = {1{`RANDOM}};
  _T_3975 = _RAND_146[2:0];
  _RAND_147 = {1{`RANDOM}};
  _T_3971 = _RAND_147[2:0];
  _RAND_148 = {1{`RANDOM}};
  _T_3967 = _RAND_148[2:0];
  _RAND_149 = {1{`RANDOM}};
  _T_3963 = _RAND_149[2:0];
  _RAND_150 = {1{`RANDOM}};
  uncacheable_miss_scnd_ff = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  imb_scnd_ff = _RAND_151[30:0];
  _RAND_152 = {1{`RANDOM}};
  ifu_bus_rid_ff = _RAND_152[2:0];
  _RAND_153 = {1{`RANDOM}};
  ifu_bus_rresp_ff = _RAND_153[1:0];
  _RAND_154 = {1{`RANDOM}};
  ifu_wr_data_comb_err_ff = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  way_status_mb_ff = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  tagv_mb_ff = _RAND_156[1:0];
  _RAND_157 = {1{`RANDOM}};
  reset_ic_ff = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  fetch_uncacheable_ff = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  miss_addr = _RAND_159[25:0];
  _RAND_160 = {1{`RANDOM}};
  ifc_region_acc_fault_f = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  bus_rd_addr_count = _RAND_161[2:0];
  _RAND_162 = {1{`RANDOM}};
  ic_act_miss_f_delayed = _RAND_162[0:0];
  _RAND_163 = {2{`RANDOM}};
  ifu_bus_rdata_ff = _RAND_163[63:0];
  _RAND_164 = {2{`RANDOM}};
  _T_1296 = _RAND_164[63:0];
  _RAND_165 = {2{`RANDOM}};
  _T_1298 = _RAND_165[63:0];
  _RAND_166 = {2{`RANDOM}};
  _T_1300 = _RAND_166[63:0];
  _RAND_167 = {2{`RANDOM}};
  _T_1302 = _RAND_167[63:0];
  _RAND_168 = {2{`RANDOM}};
  _T_1304 = _RAND_168[63:0];
  _RAND_169 = {2{`RANDOM}};
  _T_1306 = _RAND_169[63:0];
  _RAND_170 = {2{`RANDOM}};
  _T_1308 = _RAND_170[63:0];
  _RAND_171 = {2{`RANDOM}};
  _T_1310 = _RAND_171[63:0];
  _RAND_172 = {2{`RANDOM}};
  _T_1312 = _RAND_172[63:0];
  _RAND_173 = {2{`RANDOM}};
  _T_1314 = _RAND_173[63:0];
  _RAND_174 = {2{`RANDOM}};
  _T_1316 = _RAND_174[63:0];
  _RAND_175 = {2{`RANDOM}};
  _T_1318 = _RAND_175[63:0];
  _RAND_176 = {2{`RANDOM}};
  _T_1320 = _RAND_176[63:0];
  _RAND_177 = {2{`RANDOM}};
  _T_1322 = _RAND_177[63:0];
  _RAND_178 = {2{`RANDOM}};
  _T_1324 = _RAND_178[63:0];
  _RAND_179 = {2{`RANDOM}};
  _T_1326 = _RAND_179[63:0];
  _RAND_180 = {1{`RANDOM}};
  ic_crit_wd_rdy_new_ff = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  ic_miss_buff_data_error = _RAND_181[7:0];
  _RAND_182 = {1{`RANDOM}};
  ic_debug_ict_array_sel_ff = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  ic_tag_valid_out_1_0 = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  ic_tag_valid_out_1_1 = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  ic_tag_valid_out_1_2 = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  ic_tag_valid_out_1_3 = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  ic_tag_valid_out_1_4 = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  ic_tag_valid_out_1_5 = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  ic_tag_valid_out_1_6 = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  ic_tag_valid_out_1_7 = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  ic_tag_valid_out_1_8 = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  ic_tag_valid_out_1_9 = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  ic_tag_valid_out_1_10 = _RAND_193[0:0];
  _RAND_194 = {1{`RANDOM}};
  ic_tag_valid_out_1_11 = _RAND_194[0:0];
  _RAND_195 = {1{`RANDOM}};
  ic_tag_valid_out_1_12 = _RAND_195[0:0];
  _RAND_196 = {1{`RANDOM}};
  ic_tag_valid_out_1_13 = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  ic_tag_valid_out_1_14 = _RAND_197[0:0];
  _RAND_198 = {1{`RANDOM}};
  ic_tag_valid_out_1_15 = _RAND_198[0:0];
  _RAND_199 = {1{`RANDOM}};
  ic_tag_valid_out_1_16 = _RAND_199[0:0];
  _RAND_200 = {1{`RANDOM}};
  ic_tag_valid_out_1_17 = _RAND_200[0:0];
  _RAND_201 = {1{`RANDOM}};
  ic_tag_valid_out_1_18 = _RAND_201[0:0];
  _RAND_202 = {1{`RANDOM}};
  ic_tag_valid_out_1_19 = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  ic_tag_valid_out_1_20 = _RAND_203[0:0];
  _RAND_204 = {1{`RANDOM}};
  ic_tag_valid_out_1_21 = _RAND_204[0:0];
  _RAND_205 = {1{`RANDOM}};
  ic_tag_valid_out_1_22 = _RAND_205[0:0];
  _RAND_206 = {1{`RANDOM}};
  ic_tag_valid_out_1_23 = _RAND_206[0:0];
  _RAND_207 = {1{`RANDOM}};
  ic_tag_valid_out_1_24 = _RAND_207[0:0];
  _RAND_208 = {1{`RANDOM}};
  ic_tag_valid_out_1_25 = _RAND_208[0:0];
  _RAND_209 = {1{`RANDOM}};
  ic_tag_valid_out_1_26 = _RAND_209[0:0];
  _RAND_210 = {1{`RANDOM}};
  ic_tag_valid_out_1_27 = _RAND_210[0:0];
  _RAND_211 = {1{`RANDOM}};
  ic_tag_valid_out_1_28 = _RAND_211[0:0];
  _RAND_212 = {1{`RANDOM}};
  ic_tag_valid_out_1_29 = _RAND_212[0:0];
  _RAND_213 = {1{`RANDOM}};
  ic_tag_valid_out_1_30 = _RAND_213[0:0];
  _RAND_214 = {1{`RANDOM}};
  ic_tag_valid_out_1_31 = _RAND_214[0:0];
  _RAND_215 = {1{`RANDOM}};
  ic_tag_valid_out_1_32 = _RAND_215[0:0];
  _RAND_216 = {1{`RANDOM}};
  ic_tag_valid_out_1_33 = _RAND_216[0:0];
  _RAND_217 = {1{`RANDOM}};
  ic_tag_valid_out_1_34 = _RAND_217[0:0];
  _RAND_218 = {1{`RANDOM}};
  ic_tag_valid_out_1_35 = _RAND_218[0:0];
  _RAND_219 = {1{`RANDOM}};
  ic_tag_valid_out_1_36 = _RAND_219[0:0];
  _RAND_220 = {1{`RANDOM}};
  ic_tag_valid_out_1_37 = _RAND_220[0:0];
  _RAND_221 = {1{`RANDOM}};
  ic_tag_valid_out_1_38 = _RAND_221[0:0];
  _RAND_222 = {1{`RANDOM}};
  ic_tag_valid_out_1_39 = _RAND_222[0:0];
  _RAND_223 = {1{`RANDOM}};
  ic_tag_valid_out_1_40 = _RAND_223[0:0];
  _RAND_224 = {1{`RANDOM}};
  ic_tag_valid_out_1_41 = _RAND_224[0:0];
  _RAND_225 = {1{`RANDOM}};
  ic_tag_valid_out_1_42 = _RAND_225[0:0];
  _RAND_226 = {1{`RANDOM}};
  ic_tag_valid_out_1_43 = _RAND_226[0:0];
  _RAND_227 = {1{`RANDOM}};
  ic_tag_valid_out_1_44 = _RAND_227[0:0];
  _RAND_228 = {1{`RANDOM}};
  ic_tag_valid_out_1_45 = _RAND_228[0:0];
  _RAND_229 = {1{`RANDOM}};
  ic_tag_valid_out_1_46 = _RAND_229[0:0];
  _RAND_230 = {1{`RANDOM}};
  ic_tag_valid_out_1_47 = _RAND_230[0:0];
  _RAND_231 = {1{`RANDOM}};
  ic_tag_valid_out_1_48 = _RAND_231[0:0];
  _RAND_232 = {1{`RANDOM}};
  ic_tag_valid_out_1_49 = _RAND_232[0:0];
  _RAND_233 = {1{`RANDOM}};
  ic_tag_valid_out_1_50 = _RAND_233[0:0];
  _RAND_234 = {1{`RANDOM}};
  ic_tag_valid_out_1_51 = _RAND_234[0:0];
  _RAND_235 = {1{`RANDOM}};
  ic_tag_valid_out_1_52 = _RAND_235[0:0];
  _RAND_236 = {1{`RANDOM}};
  ic_tag_valid_out_1_53 = _RAND_236[0:0];
  _RAND_237 = {1{`RANDOM}};
  ic_tag_valid_out_1_54 = _RAND_237[0:0];
  _RAND_238 = {1{`RANDOM}};
  ic_tag_valid_out_1_55 = _RAND_238[0:0];
  _RAND_239 = {1{`RANDOM}};
  ic_tag_valid_out_1_56 = _RAND_239[0:0];
  _RAND_240 = {1{`RANDOM}};
  ic_tag_valid_out_1_57 = _RAND_240[0:0];
  _RAND_241 = {1{`RANDOM}};
  ic_tag_valid_out_1_58 = _RAND_241[0:0];
  _RAND_242 = {1{`RANDOM}};
  ic_tag_valid_out_1_59 = _RAND_242[0:0];
  _RAND_243 = {1{`RANDOM}};
  ic_tag_valid_out_1_60 = _RAND_243[0:0];
  _RAND_244 = {1{`RANDOM}};
  ic_tag_valid_out_1_61 = _RAND_244[0:0];
  _RAND_245 = {1{`RANDOM}};
  ic_tag_valid_out_1_62 = _RAND_245[0:0];
  _RAND_246 = {1{`RANDOM}};
  ic_tag_valid_out_1_63 = _RAND_246[0:0];
  _RAND_247 = {1{`RANDOM}};
  ic_tag_valid_out_1_64 = _RAND_247[0:0];
  _RAND_248 = {1{`RANDOM}};
  ic_tag_valid_out_1_65 = _RAND_248[0:0];
  _RAND_249 = {1{`RANDOM}};
  ic_tag_valid_out_1_66 = _RAND_249[0:0];
  _RAND_250 = {1{`RANDOM}};
  ic_tag_valid_out_1_67 = _RAND_250[0:0];
  _RAND_251 = {1{`RANDOM}};
  ic_tag_valid_out_1_68 = _RAND_251[0:0];
  _RAND_252 = {1{`RANDOM}};
  ic_tag_valid_out_1_69 = _RAND_252[0:0];
  _RAND_253 = {1{`RANDOM}};
  ic_tag_valid_out_1_70 = _RAND_253[0:0];
  _RAND_254 = {1{`RANDOM}};
  ic_tag_valid_out_1_71 = _RAND_254[0:0];
  _RAND_255 = {1{`RANDOM}};
  ic_tag_valid_out_1_72 = _RAND_255[0:0];
  _RAND_256 = {1{`RANDOM}};
  ic_tag_valid_out_1_73 = _RAND_256[0:0];
  _RAND_257 = {1{`RANDOM}};
  ic_tag_valid_out_1_74 = _RAND_257[0:0];
  _RAND_258 = {1{`RANDOM}};
  ic_tag_valid_out_1_75 = _RAND_258[0:0];
  _RAND_259 = {1{`RANDOM}};
  ic_tag_valid_out_1_76 = _RAND_259[0:0];
  _RAND_260 = {1{`RANDOM}};
  ic_tag_valid_out_1_77 = _RAND_260[0:0];
  _RAND_261 = {1{`RANDOM}};
  ic_tag_valid_out_1_78 = _RAND_261[0:0];
  _RAND_262 = {1{`RANDOM}};
  ic_tag_valid_out_1_79 = _RAND_262[0:0];
  _RAND_263 = {1{`RANDOM}};
  ic_tag_valid_out_1_80 = _RAND_263[0:0];
  _RAND_264 = {1{`RANDOM}};
  ic_tag_valid_out_1_81 = _RAND_264[0:0];
  _RAND_265 = {1{`RANDOM}};
  ic_tag_valid_out_1_82 = _RAND_265[0:0];
  _RAND_266 = {1{`RANDOM}};
  ic_tag_valid_out_1_83 = _RAND_266[0:0];
  _RAND_267 = {1{`RANDOM}};
  ic_tag_valid_out_1_84 = _RAND_267[0:0];
  _RAND_268 = {1{`RANDOM}};
  ic_tag_valid_out_1_85 = _RAND_268[0:0];
  _RAND_269 = {1{`RANDOM}};
  ic_tag_valid_out_1_86 = _RAND_269[0:0];
  _RAND_270 = {1{`RANDOM}};
  ic_tag_valid_out_1_87 = _RAND_270[0:0];
  _RAND_271 = {1{`RANDOM}};
  ic_tag_valid_out_1_88 = _RAND_271[0:0];
  _RAND_272 = {1{`RANDOM}};
  ic_tag_valid_out_1_89 = _RAND_272[0:0];
  _RAND_273 = {1{`RANDOM}};
  ic_tag_valid_out_1_90 = _RAND_273[0:0];
  _RAND_274 = {1{`RANDOM}};
  ic_tag_valid_out_1_91 = _RAND_274[0:0];
  _RAND_275 = {1{`RANDOM}};
  ic_tag_valid_out_1_92 = _RAND_275[0:0];
  _RAND_276 = {1{`RANDOM}};
  ic_tag_valid_out_1_93 = _RAND_276[0:0];
  _RAND_277 = {1{`RANDOM}};
  ic_tag_valid_out_1_94 = _RAND_277[0:0];
  _RAND_278 = {1{`RANDOM}};
  ic_tag_valid_out_1_95 = _RAND_278[0:0];
  _RAND_279 = {1{`RANDOM}};
  ic_tag_valid_out_1_96 = _RAND_279[0:0];
  _RAND_280 = {1{`RANDOM}};
  ic_tag_valid_out_1_97 = _RAND_280[0:0];
  _RAND_281 = {1{`RANDOM}};
  ic_tag_valid_out_1_98 = _RAND_281[0:0];
  _RAND_282 = {1{`RANDOM}};
  ic_tag_valid_out_1_99 = _RAND_282[0:0];
  _RAND_283 = {1{`RANDOM}};
  ic_tag_valid_out_1_100 = _RAND_283[0:0];
  _RAND_284 = {1{`RANDOM}};
  ic_tag_valid_out_1_101 = _RAND_284[0:0];
  _RAND_285 = {1{`RANDOM}};
  ic_tag_valid_out_1_102 = _RAND_285[0:0];
  _RAND_286 = {1{`RANDOM}};
  ic_tag_valid_out_1_103 = _RAND_286[0:0];
  _RAND_287 = {1{`RANDOM}};
  ic_tag_valid_out_1_104 = _RAND_287[0:0];
  _RAND_288 = {1{`RANDOM}};
  ic_tag_valid_out_1_105 = _RAND_288[0:0];
  _RAND_289 = {1{`RANDOM}};
  ic_tag_valid_out_1_106 = _RAND_289[0:0];
  _RAND_290 = {1{`RANDOM}};
  ic_tag_valid_out_1_107 = _RAND_290[0:0];
  _RAND_291 = {1{`RANDOM}};
  ic_tag_valid_out_1_108 = _RAND_291[0:0];
  _RAND_292 = {1{`RANDOM}};
  ic_tag_valid_out_1_109 = _RAND_292[0:0];
  _RAND_293 = {1{`RANDOM}};
  ic_tag_valid_out_1_110 = _RAND_293[0:0];
  _RAND_294 = {1{`RANDOM}};
  ic_tag_valid_out_1_111 = _RAND_294[0:0];
  _RAND_295 = {1{`RANDOM}};
  ic_tag_valid_out_1_112 = _RAND_295[0:0];
  _RAND_296 = {1{`RANDOM}};
  ic_tag_valid_out_1_113 = _RAND_296[0:0];
  _RAND_297 = {1{`RANDOM}};
  ic_tag_valid_out_1_114 = _RAND_297[0:0];
  _RAND_298 = {1{`RANDOM}};
  ic_tag_valid_out_1_115 = _RAND_298[0:0];
  _RAND_299 = {1{`RANDOM}};
  ic_tag_valid_out_1_116 = _RAND_299[0:0];
  _RAND_300 = {1{`RANDOM}};
  ic_tag_valid_out_1_117 = _RAND_300[0:0];
  _RAND_301 = {1{`RANDOM}};
  ic_tag_valid_out_1_118 = _RAND_301[0:0];
  _RAND_302 = {1{`RANDOM}};
  ic_tag_valid_out_1_119 = _RAND_302[0:0];
  _RAND_303 = {1{`RANDOM}};
  ic_tag_valid_out_1_120 = _RAND_303[0:0];
  _RAND_304 = {1{`RANDOM}};
  ic_tag_valid_out_1_121 = _RAND_304[0:0];
  _RAND_305 = {1{`RANDOM}};
  ic_tag_valid_out_1_122 = _RAND_305[0:0];
  _RAND_306 = {1{`RANDOM}};
  ic_tag_valid_out_1_123 = _RAND_306[0:0];
  _RAND_307 = {1{`RANDOM}};
  ic_tag_valid_out_1_124 = _RAND_307[0:0];
  _RAND_308 = {1{`RANDOM}};
  ic_tag_valid_out_1_125 = _RAND_308[0:0];
  _RAND_309 = {1{`RANDOM}};
  ic_tag_valid_out_1_126 = _RAND_309[0:0];
  _RAND_310 = {1{`RANDOM}};
  ic_tag_valid_out_1_127 = _RAND_310[0:0];
  _RAND_311 = {1{`RANDOM}};
  ic_tag_valid_out_0_0 = _RAND_311[0:0];
  _RAND_312 = {1{`RANDOM}};
  ic_tag_valid_out_0_1 = _RAND_312[0:0];
  _RAND_313 = {1{`RANDOM}};
  ic_tag_valid_out_0_2 = _RAND_313[0:0];
  _RAND_314 = {1{`RANDOM}};
  ic_tag_valid_out_0_3 = _RAND_314[0:0];
  _RAND_315 = {1{`RANDOM}};
  ic_tag_valid_out_0_4 = _RAND_315[0:0];
  _RAND_316 = {1{`RANDOM}};
  ic_tag_valid_out_0_5 = _RAND_316[0:0];
  _RAND_317 = {1{`RANDOM}};
  ic_tag_valid_out_0_6 = _RAND_317[0:0];
  _RAND_318 = {1{`RANDOM}};
  ic_tag_valid_out_0_7 = _RAND_318[0:0];
  _RAND_319 = {1{`RANDOM}};
  ic_tag_valid_out_0_8 = _RAND_319[0:0];
  _RAND_320 = {1{`RANDOM}};
  ic_tag_valid_out_0_9 = _RAND_320[0:0];
  _RAND_321 = {1{`RANDOM}};
  ic_tag_valid_out_0_10 = _RAND_321[0:0];
  _RAND_322 = {1{`RANDOM}};
  ic_tag_valid_out_0_11 = _RAND_322[0:0];
  _RAND_323 = {1{`RANDOM}};
  ic_tag_valid_out_0_12 = _RAND_323[0:0];
  _RAND_324 = {1{`RANDOM}};
  ic_tag_valid_out_0_13 = _RAND_324[0:0];
  _RAND_325 = {1{`RANDOM}};
  ic_tag_valid_out_0_14 = _RAND_325[0:0];
  _RAND_326 = {1{`RANDOM}};
  ic_tag_valid_out_0_15 = _RAND_326[0:0];
  _RAND_327 = {1{`RANDOM}};
  ic_tag_valid_out_0_16 = _RAND_327[0:0];
  _RAND_328 = {1{`RANDOM}};
  ic_tag_valid_out_0_17 = _RAND_328[0:0];
  _RAND_329 = {1{`RANDOM}};
  ic_tag_valid_out_0_18 = _RAND_329[0:0];
  _RAND_330 = {1{`RANDOM}};
  ic_tag_valid_out_0_19 = _RAND_330[0:0];
  _RAND_331 = {1{`RANDOM}};
  ic_tag_valid_out_0_20 = _RAND_331[0:0];
  _RAND_332 = {1{`RANDOM}};
  ic_tag_valid_out_0_21 = _RAND_332[0:0];
  _RAND_333 = {1{`RANDOM}};
  ic_tag_valid_out_0_22 = _RAND_333[0:0];
  _RAND_334 = {1{`RANDOM}};
  ic_tag_valid_out_0_23 = _RAND_334[0:0];
  _RAND_335 = {1{`RANDOM}};
  ic_tag_valid_out_0_24 = _RAND_335[0:0];
  _RAND_336 = {1{`RANDOM}};
  ic_tag_valid_out_0_25 = _RAND_336[0:0];
  _RAND_337 = {1{`RANDOM}};
  ic_tag_valid_out_0_26 = _RAND_337[0:0];
  _RAND_338 = {1{`RANDOM}};
  ic_tag_valid_out_0_27 = _RAND_338[0:0];
  _RAND_339 = {1{`RANDOM}};
  ic_tag_valid_out_0_28 = _RAND_339[0:0];
  _RAND_340 = {1{`RANDOM}};
  ic_tag_valid_out_0_29 = _RAND_340[0:0];
  _RAND_341 = {1{`RANDOM}};
  ic_tag_valid_out_0_30 = _RAND_341[0:0];
  _RAND_342 = {1{`RANDOM}};
  ic_tag_valid_out_0_31 = _RAND_342[0:0];
  _RAND_343 = {1{`RANDOM}};
  ic_tag_valid_out_0_32 = _RAND_343[0:0];
  _RAND_344 = {1{`RANDOM}};
  ic_tag_valid_out_0_33 = _RAND_344[0:0];
  _RAND_345 = {1{`RANDOM}};
  ic_tag_valid_out_0_34 = _RAND_345[0:0];
  _RAND_346 = {1{`RANDOM}};
  ic_tag_valid_out_0_35 = _RAND_346[0:0];
  _RAND_347 = {1{`RANDOM}};
  ic_tag_valid_out_0_36 = _RAND_347[0:0];
  _RAND_348 = {1{`RANDOM}};
  ic_tag_valid_out_0_37 = _RAND_348[0:0];
  _RAND_349 = {1{`RANDOM}};
  ic_tag_valid_out_0_38 = _RAND_349[0:0];
  _RAND_350 = {1{`RANDOM}};
  ic_tag_valid_out_0_39 = _RAND_350[0:0];
  _RAND_351 = {1{`RANDOM}};
  ic_tag_valid_out_0_40 = _RAND_351[0:0];
  _RAND_352 = {1{`RANDOM}};
  ic_tag_valid_out_0_41 = _RAND_352[0:0];
  _RAND_353 = {1{`RANDOM}};
  ic_tag_valid_out_0_42 = _RAND_353[0:0];
  _RAND_354 = {1{`RANDOM}};
  ic_tag_valid_out_0_43 = _RAND_354[0:0];
  _RAND_355 = {1{`RANDOM}};
  ic_tag_valid_out_0_44 = _RAND_355[0:0];
  _RAND_356 = {1{`RANDOM}};
  ic_tag_valid_out_0_45 = _RAND_356[0:0];
  _RAND_357 = {1{`RANDOM}};
  ic_tag_valid_out_0_46 = _RAND_357[0:0];
  _RAND_358 = {1{`RANDOM}};
  ic_tag_valid_out_0_47 = _RAND_358[0:0];
  _RAND_359 = {1{`RANDOM}};
  ic_tag_valid_out_0_48 = _RAND_359[0:0];
  _RAND_360 = {1{`RANDOM}};
  ic_tag_valid_out_0_49 = _RAND_360[0:0];
  _RAND_361 = {1{`RANDOM}};
  ic_tag_valid_out_0_50 = _RAND_361[0:0];
  _RAND_362 = {1{`RANDOM}};
  ic_tag_valid_out_0_51 = _RAND_362[0:0];
  _RAND_363 = {1{`RANDOM}};
  ic_tag_valid_out_0_52 = _RAND_363[0:0];
  _RAND_364 = {1{`RANDOM}};
  ic_tag_valid_out_0_53 = _RAND_364[0:0];
  _RAND_365 = {1{`RANDOM}};
  ic_tag_valid_out_0_54 = _RAND_365[0:0];
  _RAND_366 = {1{`RANDOM}};
  ic_tag_valid_out_0_55 = _RAND_366[0:0];
  _RAND_367 = {1{`RANDOM}};
  ic_tag_valid_out_0_56 = _RAND_367[0:0];
  _RAND_368 = {1{`RANDOM}};
  ic_tag_valid_out_0_57 = _RAND_368[0:0];
  _RAND_369 = {1{`RANDOM}};
  ic_tag_valid_out_0_58 = _RAND_369[0:0];
  _RAND_370 = {1{`RANDOM}};
  ic_tag_valid_out_0_59 = _RAND_370[0:0];
  _RAND_371 = {1{`RANDOM}};
  ic_tag_valid_out_0_60 = _RAND_371[0:0];
  _RAND_372 = {1{`RANDOM}};
  ic_tag_valid_out_0_61 = _RAND_372[0:0];
  _RAND_373 = {1{`RANDOM}};
  ic_tag_valid_out_0_62 = _RAND_373[0:0];
  _RAND_374 = {1{`RANDOM}};
  ic_tag_valid_out_0_63 = _RAND_374[0:0];
  _RAND_375 = {1{`RANDOM}};
  ic_tag_valid_out_0_64 = _RAND_375[0:0];
  _RAND_376 = {1{`RANDOM}};
  ic_tag_valid_out_0_65 = _RAND_376[0:0];
  _RAND_377 = {1{`RANDOM}};
  ic_tag_valid_out_0_66 = _RAND_377[0:0];
  _RAND_378 = {1{`RANDOM}};
  ic_tag_valid_out_0_67 = _RAND_378[0:0];
  _RAND_379 = {1{`RANDOM}};
  ic_tag_valid_out_0_68 = _RAND_379[0:0];
  _RAND_380 = {1{`RANDOM}};
  ic_tag_valid_out_0_69 = _RAND_380[0:0];
  _RAND_381 = {1{`RANDOM}};
  ic_tag_valid_out_0_70 = _RAND_381[0:0];
  _RAND_382 = {1{`RANDOM}};
  ic_tag_valid_out_0_71 = _RAND_382[0:0];
  _RAND_383 = {1{`RANDOM}};
  ic_tag_valid_out_0_72 = _RAND_383[0:0];
  _RAND_384 = {1{`RANDOM}};
  ic_tag_valid_out_0_73 = _RAND_384[0:0];
  _RAND_385 = {1{`RANDOM}};
  ic_tag_valid_out_0_74 = _RAND_385[0:0];
  _RAND_386 = {1{`RANDOM}};
  ic_tag_valid_out_0_75 = _RAND_386[0:0];
  _RAND_387 = {1{`RANDOM}};
  ic_tag_valid_out_0_76 = _RAND_387[0:0];
  _RAND_388 = {1{`RANDOM}};
  ic_tag_valid_out_0_77 = _RAND_388[0:0];
  _RAND_389 = {1{`RANDOM}};
  ic_tag_valid_out_0_78 = _RAND_389[0:0];
  _RAND_390 = {1{`RANDOM}};
  ic_tag_valid_out_0_79 = _RAND_390[0:0];
  _RAND_391 = {1{`RANDOM}};
  ic_tag_valid_out_0_80 = _RAND_391[0:0];
  _RAND_392 = {1{`RANDOM}};
  ic_tag_valid_out_0_81 = _RAND_392[0:0];
  _RAND_393 = {1{`RANDOM}};
  ic_tag_valid_out_0_82 = _RAND_393[0:0];
  _RAND_394 = {1{`RANDOM}};
  ic_tag_valid_out_0_83 = _RAND_394[0:0];
  _RAND_395 = {1{`RANDOM}};
  ic_tag_valid_out_0_84 = _RAND_395[0:0];
  _RAND_396 = {1{`RANDOM}};
  ic_tag_valid_out_0_85 = _RAND_396[0:0];
  _RAND_397 = {1{`RANDOM}};
  ic_tag_valid_out_0_86 = _RAND_397[0:0];
  _RAND_398 = {1{`RANDOM}};
  ic_tag_valid_out_0_87 = _RAND_398[0:0];
  _RAND_399 = {1{`RANDOM}};
  ic_tag_valid_out_0_88 = _RAND_399[0:0];
  _RAND_400 = {1{`RANDOM}};
  ic_tag_valid_out_0_89 = _RAND_400[0:0];
  _RAND_401 = {1{`RANDOM}};
  ic_tag_valid_out_0_90 = _RAND_401[0:0];
  _RAND_402 = {1{`RANDOM}};
  ic_tag_valid_out_0_91 = _RAND_402[0:0];
  _RAND_403 = {1{`RANDOM}};
  ic_tag_valid_out_0_92 = _RAND_403[0:0];
  _RAND_404 = {1{`RANDOM}};
  ic_tag_valid_out_0_93 = _RAND_404[0:0];
  _RAND_405 = {1{`RANDOM}};
  ic_tag_valid_out_0_94 = _RAND_405[0:0];
  _RAND_406 = {1{`RANDOM}};
  ic_tag_valid_out_0_95 = _RAND_406[0:0];
  _RAND_407 = {1{`RANDOM}};
  ic_tag_valid_out_0_96 = _RAND_407[0:0];
  _RAND_408 = {1{`RANDOM}};
  ic_tag_valid_out_0_97 = _RAND_408[0:0];
  _RAND_409 = {1{`RANDOM}};
  ic_tag_valid_out_0_98 = _RAND_409[0:0];
  _RAND_410 = {1{`RANDOM}};
  ic_tag_valid_out_0_99 = _RAND_410[0:0];
  _RAND_411 = {1{`RANDOM}};
  ic_tag_valid_out_0_100 = _RAND_411[0:0];
  _RAND_412 = {1{`RANDOM}};
  ic_tag_valid_out_0_101 = _RAND_412[0:0];
  _RAND_413 = {1{`RANDOM}};
  ic_tag_valid_out_0_102 = _RAND_413[0:0];
  _RAND_414 = {1{`RANDOM}};
  ic_tag_valid_out_0_103 = _RAND_414[0:0];
  _RAND_415 = {1{`RANDOM}};
  ic_tag_valid_out_0_104 = _RAND_415[0:0];
  _RAND_416 = {1{`RANDOM}};
  ic_tag_valid_out_0_105 = _RAND_416[0:0];
  _RAND_417 = {1{`RANDOM}};
  ic_tag_valid_out_0_106 = _RAND_417[0:0];
  _RAND_418 = {1{`RANDOM}};
  ic_tag_valid_out_0_107 = _RAND_418[0:0];
  _RAND_419 = {1{`RANDOM}};
  ic_tag_valid_out_0_108 = _RAND_419[0:0];
  _RAND_420 = {1{`RANDOM}};
  ic_tag_valid_out_0_109 = _RAND_420[0:0];
  _RAND_421 = {1{`RANDOM}};
  ic_tag_valid_out_0_110 = _RAND_421[0:0];
  _RAND_422 = {1{`RANDOM}};
  ic_tag_valid_out_0_111 = _RAND_422[0:0];
  _RAND_423 = {1{`RANDOM}};
  ic_tag_valid_out_0_112 = _RAND_423[0:0];
  _RAND_424 = {1{`RANDOM}};
  ic_tag_valid_out_0_113 = _RAND_424[0:0];
  _RAND_425 = {1{`RANDOM}};
  ic_tag_valid_out_0_114 = _RAND_425[0:0];
  _RAND_426 = {1{`RANDOM}};
  ic_tag_valid_out_0_115 = _RAND_426[0:0];
  _RAND_427 = {1{`RANDOM}};
  ic_tag_valid_out_0_116 = _RAND_427[0:0];
  _RAND_428 = {1{`RANDOM}};
  ic_tag_valid_out_0_117 = _RAND_428[0:0];
  _RAND_429 = {1{`RANDOM}};
  ic_tag_valid_out_0_118 = _RAND_429[0:0];
  _RAND_430 = {1{`RANDOM}};
  ic_tag_valid_out_0_119 = _RAND_430[0:0];
  _RAND_431 = {1{`RANDOM}};
  ic_tag_valid_out_0_120 = _RAND_431[0:0];
  _RAND_432 = {1{`RANDOM}};
  ic_tag_valid_out_0_121 = _RAND_432[0:0];
  _RAND_433 = {1{`RANDOM}};
  ic_tag_valid_out_0_122 = _RAND_433[0:0];
  _RAND_434 = {1{`RANDOM}};
  ic_tag_valid_out_0_123 = _RAND_434[0:0];
  _RAND_435 = {1{`RANDOM}};
  ic_tag_valid_out_0_124 = _RAND_435[0:0];
  _RAND_436 = {1{`RANDOM}};
  ic_tag_valid_out_0_125 = _RAND_436[0:0];
  _RAND_437 = {1{`RANDOM}};
  ic_tag_valid_out_0_126 = _RAND_437[0:0];
  _RAND_438 = {1{`RANDOM}};
  ic_tag_valid_out_0_127 = _RAND_438[0:0];
  _RAND_439 = {1{`RANDOM}};
  ic_debug_way_ff = _RAND_439[1:0];
  _RAND_440 = {1{`RANDOM}};
  ic_debug_rd_en_ff = _RAND_440[0:0];
  _RAND_441 = {3{`RANDOM}};
  _T_1212 = _RAND_441[70:0];
  _RAND_442 = {1{`RANDOM}};
  perr_ic_index_ff = _RAND_442[5:0];
  _RAND_443 = {1{`RANDOM}};
  dma_sb_err_state_ff = _RAND_443[0:0];
  _RAND_444 = {1{`RANDOM}};
  ifu_bus_cmd_valid = _RAND_444[0:0];
  _RAND_445 = {1{`RANDOM}};
  bus_cmd_beat_count = _RAND_445[2:0];
  _RAND_446 = {1{`RANDOM}};
  ifu_bus_arready_unq_ff = _RAND_446[0:0];
  _RAND_447 = {1{`RANDOM}};
  ifu_bus_arvalid_ff = _RAND_447[0:0];
  _RAND_448 = {1{`RANDOM}};
  ifc_dma_access_ok_prev = _RAND_448[0:0];
  _RAND_449 = {2{`RANDOM}};
  iccm_ecc_corr_data_ff = _RAND_449[38:0];
  _RAND_450 = {1{`RANDOM}};
  dma_mem_addr_ff = _RAND_450[1:0];
  _RAND_451 = {1{`RANDOM}};
  dma_mem_tag_ff = _RAND_451[2:0];
  _RAND_452 = {1{`RANDOM}};
  iccm_dma_rtag = _RAND_452[2:0];
  _RAND_453 = {1{`RANDOM}};
  iccm_dma_rvalid = _RAND_453[0:0];
  _RAND_454 = {2{`RANDOM}};
  iccm_dma_rdata = _RAND_454[63:0];
  _RAND_455 = {1{`RANDOM}};
  iccm_ecc_corr_index_ff = _RAND_455[13:0];
  _RAND_456 = {1{`RANDOM}};
  iccm_rd_ecc_single_err_ff = _RAND_456[0:0];
  _RAND_457 = {1{`RANDOM}};
  iccm_rw_addr_f = _RAND_457[13:0];
  _RAND_458 = {1{`RANDOM}};
  ifu_status_wr_addr_ff = _RAND_458[6:0];
  _RAND_459 = {1{`RANDOM}};
  way_status_wr_en_ff = _RAND_459[0:0];
  _RAND_460 = {1{`RANDOM}};
  way_status_new_ff = _RAND_460[2:0];
  _RAND_461 = {1{`RANDOM}};
  ifu_tag_wren_ff = _RAND_461[1:0];
  _RAND_462 = {1{`RANDOM}};
  ic_valid_ff = _RAND_462[0:0];
  _RAND_463 = {1{`RANDOM}};
  _T_10102 = _RAND_463[0:0];
  _RAND_464 = {1{`RANDOM}};
  _T_10103 = _RAND_464[0:0];
  _RAND_465 = {1{`RANDOM}};
  _T_10104 = _RAND_465[0:0];
  _RAND_466 = {1{`RANDOM}};
  _T_10108 = _RAND_466[0:0];
  _RAND_467 = {1{`RANDOM}};
  _T_10109 = _RAND_467[0:0];
  _RAND_468 = {1{`RANDOM}};
  _T_10132 = _RAND_468[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      flush_final_f <= 1'h0;
    end else begin
      flush_final_f <= io_exu_flush_final;
    end
    if (reset) begin
      ifc_fetch_req_f_raw <= 1'h0;
    end else begin
      ifc_fetch_req_f_raw <= ifc_fetch_req_qual_bf;
    end
    if (reset) begin
      miss_state <= 3'h0;
    end else if (miss_state_en) begin
      if (_T_25) begin
        if (_T_27) begin
          miss_state <= 3'h1;
        end else begin
          miss_state <= 3'h2;
        end
      end else if (_T_32) begin
        if (_T_37) begin
          miss_state <= 3'h0;
        end else if (_T_41) begin
          miss_state <= 3'h3;
        end else if (_T_48) begin
          miss_state <= 3'h4;
        end else if (_T_52) begin
          miss_state <= 3'h0;
        end else if (_T_62) begin
          miss_state <= 3'h6;
        end else if (_T_72) begin
          miss_state <= 3'h6;
        end else if (_T_80) begin
          miss_state <= 3'h0;
        end else if (_T_85) begin
          miss_state <= 3'h2;
        end else begin
          miss_state <= 3'h0;
        end
      end else if (_T_103) begin
        miss_state <= 3'h0;
      end else if (_T_107) begin
        if (_T_114) begin
          miss_state <= 3'h2;
        end else begin
          miss_state <= 3'h0;
        end
      end else if (_T_122) begin
        if (_T_127) begin
          miss_state <= 3'h2;
        end else begin
          miss_state <= 3'h0;
        end
      end else if (_T_133) begin
        if (_T_138) begin
          miss_state <= 3'h5;
        end else if (_T_144) begin
          miss_state <= 3'h7;
        end else begin
          miss_state <= 3'h0;
        end
      end else if (_T_152) begin
        if (io_dec_tlu_force_halt) begin
          miss_state <= 3'h0;
        end else if (io_exu_flush_final) begin
          if (_T_33) begin
            miss_state <= 3'h0;
          end else begin
            miss_state <= 3'h2;
          end
        end else begin
          miss_state <= 3'h1;
        end
      end else if (_T_161) begin
        if (io_dec_tlu_force_halt) begin
          miss_state <= 3'h0;
        end else if (io_exu_flush_final) begin
          if (_T_33) begin
            miss_state <= 3'h0;
          end else begin
            miss_state <= 3'h2;
          end
        end else begin
          miss_state <= 3'h0;
        end
      end else begin
        miss_state <= 3'h0;
      end
    end
    if (reset) begin
      ifu_fetch_addr_int_f <= 31'h0;
    end else begin
      ifu_fetch_addr_int_f <= io_ifc_fetch_addr_bf;
    end
    if (reset) begin
      ifc_iccm_access_f <= 1'h0;
    end else begin
      ifc_iccm_access_f <= io_ifc_iccm_access_bf;
    end
    if (reset) begin
      ifc_region_acc_fault_final_f <= 1'h0;
    end else begin
      ifc_region_acc_fault_final_f <= io_ifc_region_acc_fault_bf;
    end
    if (reset) begin
      ifu_bus_rvalid_unq_ff <= 1'h0;
    end else if (io_ifu_bus_clk_en) begin
      ifu_bus_rvalid_unq_ff <= io_ifu_axi_rvalid;
    end
    if (reset) begin
      uncacheable_miss_ff <= 1'h0;
    end else if (scnd_miss_req) begin
      uncacheable_miss_ff <= uncacheable_miss_scnd_ff;
    end else if (!(sel_hold_imb)) begin
      uncacheable_miss_ff <= io_ifc_fetch_uncacheable_bf;
    end
    if (scnd_miss_req) begin
      imb_ff <= imb_scnd_ff;
    end else if (!(sel_hold_imb)) begin
      imb_ff <= io_ifc_fetch_addr_bf;
    end
    if (reset) begin
      way_status_mb_scnd_ff <= 1'h0;
    end else if (!(_T_17)) begin
      way_status_mb_scnd_ff <= way_status;
    end
    if (reset) begin
      _T_4471 <= 3'h0;
    end else if (_T_4470) begin
      _T_4471 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4467 <= 3'h0;
    end else if (_T_4466) begin
      _T_4467 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4463 <= 3'h0;
    end else if (_T_4462) begin
      _T_4463 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4459 <= 3'h0;
    end else if (_T_4458) begin
      _T_4459 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4455 <= 3'h0;
    end else if (_T_4454) begin
      _T_4455 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4451 <= 3'h0;
    end else if (_T_4450) begin
      _T_4451 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4447 <= 3'h0;
    end else if (_T_4446) begin
      _T_4447 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4443 <= 3'h0;
    end else if (_T_4442) begin
      _T_4443 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4439 <= 3'h0;
    end else if (_T_4438) begin
      _T_4439 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4435 <= 3'h0;
    end else if (_T_4434) begin
      _T_4435 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4431 <= 3'h0;
    end else if (_T_4430) begin
      _T_4431 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4427 <= 3'h0;
    end else if (_T_4426) begin
      _T_4427 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4423 <= 3'h0;
    end else if (_T_4422) begin
      _T_4423 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4419 <= 3'h0;
    end else if (_T_4418) begin
      _T_4419 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4415 <= 3'h0;
    end else if (_T_4414) begin
      _T_4415 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4411 <= 3'h0;
    end else if (_T_4410) begin
      _T_4411 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4407 <= 3'h0;
    end else if (_T_4406) begin
      _T_4407 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4403 <= 3'h0;
    end else if (_T_4402) begin
      _T_4403 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4399 <= 3'h0;
    end else if (_T_4398) begin
      _T_4399 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4395 <= 3'h0;
    end else if (_T_4394) begin
      _T_4395 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4391 <= 3'h0;
    end else if (_T_4390) begin
      _T_4391 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4387 <= 3'h0;
    end else if (_T_4386) begin
      _T_4387 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4383 <= 3'h0;
    end else if (_T_4382) begin
      _T_4383 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4379 <= 3'h0;
    end else if (_T_4378) begin
      _T_4379 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4375 <= 3'h0;
    end else if (_T_4374) begin
      _T_4375 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4371 <= 3'h0;
    end else if (_T_4370) begin
      _T_4371 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4367 <= 3'h0;
    end else if (_T_4366) begin
      _T_4367 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4363 <= 3'h0;
    end else if (_T_4362) begin
      _T_4363 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4359 <= 3'h0;
    end else if (_T_4358) begin
      _T_4359 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4355 <= 3'h0;
    end else if (_T_4354) begin
      _T_4355 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4351 <= 3'h0;
    end else if (_T_4350) begin
      _T_4351 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4347 <= 3'h0;
    end else if (_T_4346) begin
      _T_4347 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4343 <= 3'h0;
    end else if (_T_4342) begin
      _T_4343 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4339 <= 3'h0;
    end else if (_T_4338) begin
      _T_4339 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4335 <= 3'h0;
    end else if (_T_4334) begin
      _T_4335 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4331 <= 3'h0;
    end else if (_T_4330) begin
      _T_4331 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4327 <= 3'h0;
    end else if (_T_4326) begin
      _T_4327 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4323 <= 3'h0;
    end else if (_T_4322) begin
      _T_4323 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4319 <= 3'h0;
    end else if (_T_4318) begin
      _T_4319 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4315 <= 3'h0;
    end else if (_T_4314) begin
      _T_4315 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4311 <= 3'h0;
    end else if (_T_4310) begin
      _T_4311 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4307 <= 3'h0;
    end else if (_T_4306) begin
      _T_4307 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4303 <= 3'h0;
    end else if (_T_4302) begin
      _T_4303 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4299 <= 3'h0;
    end else if (_T_4298) begin
      _T_4299 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4295 <= 3'h0;
    end else if (_T_4294) begin
      _T_4295 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4291 <= 3'h0;
    end else if (_T_4290) begin
      _T_4291 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4287 <= 3'h0;
    end else if (_T_4286) begin
      _T_4287 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4283 <= 3'h0;
    end else if (_T_4282) begin
      _T_4283 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4279 <= 3'h0;
    end else if (_T_4278) begin
      _T_4279 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4275 <= 3'h0;
    end else if (_T_4274) begin
      _T_4275 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4271 <= 3'h0;
    end else if (_T_4270) begin
      _T_4271 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4267 <= 3'h0;
    end else if (_T_4266) begin
      _T_4267 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4263 <= 3'h0;
    end else if (_T_4262) begin
      _T_4263 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4259 <= 3'h0;
    end else if (_T_4258) begin
      _T_4259 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4255 <= 3'h0;
    end else if (_T_4254) begin
      _T_4255 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4251 <= 3'h0;
    end else if (_T_4250) begin
      _T_4251 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4247 <= 3'h0;
    end else if (_T_4246) begin
      _T_4247 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4243 <= 3'h0;
    end else if (_T_4242) begin
      _T_4243 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4239 <= 3'h0;
    end else if (_T_4238) begin
      _T_4239 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4235 <= 3'h0;
    end else if (_T_4234) begin
      _T_4235 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4231 <= 3'h0;
    end else if (_T_4230) begin
      _T_4231 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4227 <= 3'h0;
    end else if (_T_4226) begin
      _T_4227 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4223 <= 3'h0;
    end else if (_T_4222) begin
      _T_4223 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4219 <= 3'h0;
    end else if (_T_4218) begin
      _T_4219 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4215 <= 3'h0;
    end else if (_T_4214) begin
      _T_4215 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4211 <= 3'h0;
    end else if (_T_4210) begin
      _T_4211 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4207 <= 3'h0;
    end else if (_T_4206) begin
      _T_4207 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4203 <= 3'h0;
    end else if (_T_4202) begin
      _T_4203 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4199 <= 3'h0;
    end else if (_T_4198) begin
      _T_4199 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4195 <= 3'h0;
    end else if (_T_4194) begin
      _T_4195 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4191 <= 3'h0;
    end else if (_T_4190) begin
      _T_4191 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4187 <= 3'h0;
    end else if (_T_4186) begin
      _T_4187 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4183 <= 3'h0;
    end else if (_T_4182) begin
      _T_4183 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4179 <= 3'h0;
    end else if (_T_4178) begin
      _T_4179 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4175 <= 3'h0;
    end else if (_T_4174) begin
      _T_4175 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4171 <= 3'h0;
    end else if (_T_4170) begin
      _T_4171 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4167 <= 3'h0;
    end else if (_T_4166) begin
      _T_4167 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4163 <= 3'h0;
    end else if (_T_4162) begin
      _T_4163 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4159 <= 3'h0;
    end else if (_T_4158) begin
      _T_4159 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4155 <= 3'h0;
    end else if (_T_4154) begin
      _T_4155 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4151 <= 3'h0;
    end else if (_T_4150) begin
      _T_4151 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4147 <= 3'h0;
    end else if (_T_4146) begin
      _T_4147 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4143 <= 3'h0;
    end else if (_T_4142) begin
      _T_4143 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4139 <= 3'h0;
    end else if (_T_4138) begin
      _T_4139 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4135 <= 3'h0;
    end else if (_T_4134) begin
      _T_4135 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4131 <= 3'h0;
    end else if (_T_4130) begin
      _T_4131 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4127 <= 3'h0;
    end else if (_T_4126) begin
      _T_4127 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4123 <= 3'h0;
    end else if (_T_4122) begin
      _T_4123 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4119 <= 3'h0;
    end else if (_T_4118) begin
      _T_4119 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4115 <= 3'h0;
    end else if (_T_4114) begin
      _T_4115 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4111 <= 3'h0;
    end else if (_T_4110) begin
      _T_4111 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4107 <= 3'h0;
    end else if (_T_4106) begin
      _T_4107 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4103 <= 3'h0;
    end else if (_T_4102) begin
      _T_4103 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4099 <= 3'h0;
    end else if (_T_4098) begin
      _T_4099 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4095 <= 3'h0;
    end else if (_T_4094) begin
      _T_4095 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4091 <= 3'h0;
    end else if (_T_4090) begin
      _T_4091 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4087 <= 3'h0;
    end else if (_T_4086) begin
      _T_4087 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4083 <= 3'h0;
    end else if (_T_4082) begin
      _T_4083 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4079 <= 3'h0;
    end else if (_T_4078) begin
      _T_4079 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4075 <= 3'h0;
    end else if (_T_4074) begin
      _T_4075 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4071 <= 3'h0;
    end else if (_T_4070) begin
      _T_4071 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4067 <= 3'h0;
    end else if (_T_4066) begin
      _T_4067 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4063 <= 3'h0;
    end else if (_T_4062) begin
      _T_4063 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4059 <= 3'h0;
    end else if (_T_4058) begin
      _T_4059 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4055 <= 3'h0;
    end else if (_T_4054) begin
      _T_4055 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4051 <= 3'h0;
    end else if (_T_4050) begin
      _T_4051 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4047 <= 3'h0;
    end else if (_T_4046) begin
      _T_4047 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4043 <= 3'h0;
    end else if (_T_4042) begin
      _T_4043 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4039 <= 3'h0;
    end else if (_T_4038) begin
      _T_4039 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4035 <= 3'h0;
    end else if (_T_4034) begin
      _T_4035 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4031 <= 3'h0;
    end else if (_T_4030) begin
      _T_4031 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4027 <= 3'h0;
    end else if (_T_4026) begin
      _T_4027 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4023 <= 3'h0;
    end else if (_T_4022) begin
      _T_4023 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4019 <= 3'h0;
    end else if (_T_4018) begin
      _T_4019 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4015 <= 3'h0;
    end else if (_T_4014) begin
      _T_4015 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4011 <= 3'h0;
    end else if (_T_4010) begin
      _T_4011 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4007 <= 3'h0;
    end else if (_T_4006) begin
      _T_4007 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4003 <= 3'h0;
    end else if (_T_4002) begin
      _T_4003 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3999 <= 3'h0;
    end else if (_T_3998) begin
      _T_3999 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3995 <= 3'h0;
    end else if (_T_3994) begin
      _T_3995 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3991 <= 3'h0;
    end else if (_T_3990) begin
      _T_3991 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3987 <= 3'h0;
    end else if (_T_3986) begin
      _T_3987 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3983 <= 3'h0;
    end else if (_T_3982) begin
      _T_3983 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3979 <= 3'h0;
    end else if (_T_3978) begin
      _T_3979 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3975 <= 3'h0;
    end else if (_T_3974) begin
      _T_3975 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3971 <= 3'h0;
    end else if (_T_3970) begin
      _T_3971 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3967 <= 3'h0;
    end else if (_T_3966) begin
      _T_3967 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3963 <= 3'h0;
    end else if (_T_3962) begin
      _T_3963 <= way_status_new_ff;
    end
    if (reset) begin
      uncacheable_miss_scnd_ff <= 1'h0;
    end else if (!(sel_hold_imb_scnd)) begin
      uncacheable_miss_scnd_ff <= io_ifc_fetch_uncacheable_bf;
    end
    if (reset) begin
      imb_scnd_ff <= 31'h0;
    end else if (!(sel_hold_imb_scnd)) begin
      imb_scnd_ff <= io_ifc_fetch_addr_bf;
    end
    if (reset) begin
      ifu_bus_rid_ff <= 3'h0;
    end else if (io_ifu_bus_clk_en) begin
      ifu_bus_rid_ff <= io_ifu_axi_rid;
    end
    if (reset) begin
      ifu_bus_rresp_ff <= 2'h0;
    end else if (io_ifu_bus_clk_en) begin
      ifu_bus_rresp_ff <= io_ifu_axi_rresp;
    end
    if (reset) begin
      way_status_mb_ff <= 1'h0;
    end else if (_T_279) begin
      way_status_mb_ff <= way_status_mb_scnd_ff;
    end else if (_T_281) begin
      way_status_mb_ff <= replace_way_mb_any_0;
    end else if (!(miss_pending)) begin
      way_status_mb_ff <= way_status;
    end
    if (reset) begin
      tagv_mb_ff <= 2'h0;
    end else if (scnd_miss_req) begin
      tagv_mb_ff <= _T_290;
    end else if (!(miss_pending)) begin
      tagv_mb_ff <= 2'h0;
    end
    reset_ic_ff <= _T_299 & _T_300;
    if (reset) begin
      fetch_uncacheable_ff <= 1'h0;
    end else begin
      fetch_uncacheable_ff <= io_ifc_fetch_uncacheable_bf;
    end
    if (reset) begin
      miss_addr <= 26'h0;
    end else if (_T_232) begin
      miss_addr <= imb_ff[30:5];
    end else if (scnd_miss_req_q) begin
      miss_addr <= imb_scnd_ff[30:5];
    end
    if (reset) begin
      ifc_region_acc_fault_f <= 1'h0;
    end else begin
      ifc_region_acc_fault_f <= io_ifc_region_acc_fault_bf;
    end
    if (reset) begin
      bus_rd_addr_count <= 3'h0;
    end else if (_T_2564) begin
      if (_T_232) begin
        bus_rd_addr_count <= imb_ff[4:2];
      end else if (scnd_miss_req_q) begin
        bus_rd_addr_count <= imb_scnd_ff[4:2];
      end else if (bus_cmd_sent) begin
        bus_rd_addr_count <= _T_2560;
      end
    end
    if (reset) begin
      ifu_bus_rdata_ff <= 64'h0;
    end else if (io_ifu_bus_clk_en) begin
      ifu_bus_rdata_ff <= io_ifu_axi_rdata;
    end
    if (reset) begin
      _T_1296 <= 64'h0;
    end else if (write_fill_data_0) begin
      _T_1296 <= io_ifu_axi_rdata;
    end
    if (reset) begin
      _T_1298 <= 64'h0;
    end else if (write_fill_data_0) begin
      _T_1298 <= io_ifu_axi_rdata;
    end
    if (reset) begin
      _T_1300 <= 64'h0;
    end else if (write_fill_data_1) begin
      _T_1300 <= io_ifu_axi_rdata;
    end
    if (reset) begin
      _T_1302 <= 64'h0;
    end else if (write_fill_data_1) begin
      _T_1302 <= io_ifu_axi_rdata;
    end
    if (reset) begin
      _T_1304 <= 64'h0;
    end else if (write_fill_data_2) begin
      _T_1304 <= io_ifu_axi_rdata;
    end
    if (reset) begin
      _T_1306 <= 64'h0;
    end else if (write_fill_data_2) begin
      _T_1306 <= io_ifu_axi_rdata;
    end
    if (reset) begin
      _T_1308 <= 64'h0;
    end else if (write_fill_data_3) begin
      _T_1308 <= io_ifu_axi_rdata;
    end
    if (reset) begin
      _T_1310 <= 64'h0;
    end else if (write_fill_data_3) begin
      _T_1310 <= io_ifu_axi_rdata;
    end
    if (reset) begin
      _T_1312 <= 64'h0;
    end else if (write_fill_data_4) begin
      _T_1312 <= io_ifu_axi_rdata;
    end
    if (reset) begin
      _T_1314 <= 64'h0;
    end else if (write_fill_data_4) begin
      _T_1314 <= io_ifu_axi_rdata;
    end
    if (reset) begin
      _T_1316 <= 64'h0;
    end else if (write_fill_data_5) begin
      _T_1316 <= io_ifu_axi_rdata;
    end
    if (reset) begin
      _T_1318 <= 64'h0;
    end else if (write_fill_data_5) begin
      _T_1318 <= io_ifu_axi_rdata;
    end
    if (reset) begin
      _T_1320 <= 64'h0;
    end else if (write_fill_data_6) begin
      _T_1320 <= io_ifu_axi_rdata;
    end
    if (reset) begin
      _T_1322 <= 64'h0;
    end else if (write_fill_data_6) begin
      _T_1322 <= io_ifu_axi_rdata;
    end
    if (reset) begin
      _T_1324 <= 64'h0;
    end else if (write_fill_data_7) begin
      _T_1324 <= io_ifu_axi_rdata;
    end
    if (reset) begin
      _T_1326 <= 64'h0;
    end else if (write_fill_data_7) begin
      _T_1326 <= io_ifu_axi_rdata;
    end
    if (reset) begin
      ic_debug_ict_array_sel_ff <= 1'h0;
    end else if (debug_c1_clken) begin
      ic_debug_ict_array_sel_ff <= ic_debug_ict_array_sel_in;
    end
    if (reset) begin
      ic_tag_valid_out_1_0 <= 1'h0;
    end else if (_T_5723) begin
      ic_tag_valid_out_1_0 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_1 <= 1'h0;
    end else if (_T_5739) begin
      ic_tag_valid_out_1_1 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_2 <= 1'h0;
    end else if (_T_5755) begin
      ic_tag_valid_out_1_2 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_3 <= 1'h0;
    end else if (_T_5771) begin
      ic_tag_valid_out_1_3 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_4 <= 1'h0;
    end else if (_T_5787) begin
      ic_tag_valid_out_1_4 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_5 <= 1'h0;
    end else if (_T_5803) begin
      ic_tag_valid_out_1_5 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_6 <= 1'h0;
    end else if (_T_5819) begin
      ic_tag_valid_out_1_6 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_7 <= 1'h0;
    end else if (_T_5835) begin
      ic_tag_valid_out_1_7 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_8 <= 1'h0;
    end else if (_T_5851) begin
      ic_tag_valid_out_1_8 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_9 <= 1'h0;
    end else if (_T_5867) begin
      ic_tag_valid_out_1_9 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_10 <= 1'h0;
    end else if (_T_5883) begin
      ic_tag_valid_out_1_10 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_11 <= 1'h0;
    end else if (_T_5899) begin
      ic_tag_valid_out_1_11 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_12 <= 1'h0;
    end else if (_T_5915) begin
      ic_tag_valid_out_1_12 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_13 <= 1'h0;
    end else if (_T_5931) begin
      ic_tag_valid_out_1_13 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_14 <= 1'h0;
    end else if (_T_5947) begin
      ic_tag_valid_out_1_14 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_15 <= 1'h0;
    end else if (_T_5963) begin
      ic_tag_valid_out_1_15 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_16 <= 1'h0;
    end else if (_T_5979) begin
      ic_tag_valid_out_1_16 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_17 <= 1'h0;
    end else if (_T_5995) begin
      ic_tag_valid_out_1_17 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_18 <= 1'h0;
    end else if (_T_6011) begin
      ic_tag_valid_out_1_18 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_19 <= 1'h0;
    end else if (_T_6027) begin
      ic_tag_valid_out_1_19 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_20 <= 1'h0;
    end else if (_T_6043) begin
      ic_tag_valid_out_1_20 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_21 <= 1'h0;
    end else if (_T_6059) begin
      ic_tag_valid_out_1_21 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_22 <= 1'h0;
    end else if (_T_6075) begin
      ic_tag_valid_out_1_22 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_23 <= 1'h0;
    end else if (_T_6091) begin
      ic_tag_valid_out_1_23 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_24 <= 1'h0;
    end else if (_T_6107) begin
      ic_tag_valid_out_1_24 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_25 <= 1'h0;
    end else if (_T_6123) begin
      ic_tag_valid_out_1_25 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_26 <= 1'h0;
    end else if (_T_6139) begin
      ic_tag_valid_out_1_26 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_27 <= 1'h0;
    end else if (_T_6155) begin
      ic_tag_valid_out_1_27 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_28 <= 1'h0;
    end else if (_T_6171) begin
      ic_tag_valid_out_1_28 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_29 <= 1'h0;
    end else if (_T_6187) begin
      ic_tag_valid_out_1_29 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_30 <= 1'h0;
    end else if (_T_6203) begin
      ic_tag_valid_out_1_30 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_31 <= 1'h0;
    end else if (_T_6219) begin
      ic_tag_valid_out_1_31 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_32 <= 1'h0;
    end else if (_T_6747) begin
      ic_tag_valid_out_1_32 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_33 <= 1'h0;
    end else if (_T_6763) begin
      ic_tag_valid_out_1_33 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_34 <= 1'h0;
    end else if (_T_6779) begin
      ic_tag_valid_out_1_34 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_35 <= 1'h0;
    end else if (_T_6795) begin
      ic_tag_valid_out_1_35 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_36 <= 1'h0;
    end else if (_T_6811) begin
      ic_tag_valid_out_1_36 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_37 <= 1'h0;
    end else if (_T_6827) begin
      ic_tag_valid_out_1_37 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_38 <= 1'h0;
    end else if (_T_6843) begin
      ic_tag_valid_out_1_38 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_39 <= 1'h0;
    end else if (_T_6859) begin
      ic_tag_valid_out_1_39 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_40 <= 1'h0;
    end else if (_T_6875) begin
      ic_tag_valid_out_1_40 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_41 <= 1'h0;
    end else if (_T_6891) begin
      ic_tag_valid_out_1_41 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_42 <= 1'h0;
    end else if (_T_6907) begin
      ic_tag_valid_out_1_42 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_43 <= 1'h0;
    end else if (_T_6923) begin
      ic_tag_valid_out_1_43 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_44 <= 1'h0;
    end else if (_T_6939) begin
      ic_tag_valid_out_1_44 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_45 <= 1'h0;
    end else if (_T_6955) begin
      ic_tag_valid_out_1_45 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_46 <= 1'h0;
    end else if (_T_6971) begin
      ic_tag_valid_out_1_46 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_47 <= 1'h0;
    end else if (_T_6987) begin
      ic_tag_valid_out_1_47 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_48 <= 1'h0;
    end else if (_T_7003) begin
      ic_tag_valid_out_1_48 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_49 <= 1'h0;
    end else if (_T_7019) begin
      ic_tag_valid_out_1_49 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_50 <= 1'h0;
    end else if (_T_7035) begin
      ic_tag_valid_out_1_50 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_51 <= 1'h0;
    end else if (_T_7051) begin
      ic_tag_valid_out_1_51 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_52 <= 1'h0;
    end else if (_T_7067) begin
      ic_tag_valid_out_1_52 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_53 <= 1'h0;
    end else if (_T_7083) begin
      ic_tag_valid_out_1_53 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_54 <= 1'h0;
    end else if (_T_7099) begin
      ic_tag_valid_out_1_54 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_55 <= 1'h0;
    end else if (_T_7115) begin
      ic_tag_valid_out_1_55 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_56 <= 1'h0;
    end else if (_T_7131) begin
      ic_tag_valid_out_1_56 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_57 <= 1'h0;
    end else if (_T_7147) begin
      ic_tag_valid_out_1_57 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_58 <= 1'h0;
    end else if (_T_7163) begin
      ic_tag_valid_out_1_58 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_59 <= 1'h0;
    end else if (_T_7179) begin
      ic_tag_valid_out_1_59 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_60 <= 1'h0;
    end else if (_T_7195) begin
      ic_tag_valid_out_1_60 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_61 <= 1'h0;
    end else if (_T_7211) begin
      ic_tag_valid_out_1_61 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_62 <= 1'h0;
    end else if (_T_7227) begin
      ic_tag_valid_out_1_62 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_63 <= 1'h0;
    end else if (_T_7243) begin
      ic_tag_valid_out_1_63 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_64 <= 1'h0;
    end else if (_T_7771) begin
      ic_tag_valid_out_1_64 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_65 <= 1'h0;
    end else if (_T_7787) begin
      ic_tag_valid_out_1_65 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_66 <= 1'h0;
    end else if (_T_7803) begin
      ic_tag_valid_out_1_66 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_67 <= 1'h0;
    end else if (_T_7819) begin
      ic_tag_valid_out_1_67 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_68 <= 1'h0;
    end else if (_T_7835) begin
      ic_tag_valid_out_1_68 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_69 <= 1'h0;
    end else if (_T_7851) begin
      ic_tag_valid_out_1_69 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_70 <= 1'h0;
    end else if (_T_7867) begin
      ic_tag_valid_out_1_70 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_71 <= 1'h0;
    end else if (_T_7883) begin
      ic_tag_valid_out_1_71 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_72 <= 1'h0;
    end else if (_T_7899) begin
      ic_tag_valid_out_1_72 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_73 <= 1'h0;
    end else if (_T_7915) begin
      ic_tag_valid_out_1_73 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_74 <= 1'h0;
    end else if (_T_7931) begin
      ic_tag_valid_out_1_74 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_75 <= 1'h0;
    end else if (_T_7947) begin
      ic_tag_valid_out_1_75 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_76 <= 1'h0;
    end else if (_T_7963) begin
      ic_tag_valid_out_1_76 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_77 <= 1'h0;
    end else if (_T_7979) begin
      ic_tag_valid_out_1_77 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_78 <= 1'h0;
    end else if (_T_7995) begin
      ic_tag_valid_out_1_78 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_79 <= 1'h0;
    end else if (_T_8011) begin
      ic_tag_valid_out_1_79 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_80 <= 1'h0;
    end else if (_T_8027) begin
      ic_tag_valid_out_1_80 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_81 <= 1'h0;
    end else if (_T_8043) begin
      ic_tag_valid_out_1_81 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_82 <= 1'h0;
    end else if (_T_8059) begin
      ic_tag_valid_out_1_82 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_83 <= 1'h0;
    end else if (_T_8075) begin
      ic_tag_valid_out_1_83 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_84 <= 1'h0;
    end else if (_T_8091) begin
      ic_tag_valid_out_1_84 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_85 <= 1'h0;
    end else if (_T_8107) begin
      ic_tag_valid_out_1_85 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_86 <= 1'h0;
    end else if (_T_8123) begin
      ic_tag_valid_out_1_86 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_87 <= 1'h0;
    end else if (_T_8139) begin
      ic_tag_valid_out_1_87 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_88 <= 1'h0;
    end else if (_T_8155) begin
      ic_tag_valid_out_1_88 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_89 <= 1'h0;
    end else if (_T_8171) begin
      ic_tag_valid_out_1_89 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_90 <= 1'h0;
    end else if (_T_8187) begin
      ic_tag_valid_out_1_90 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_91 <= 1'h0;
    end else if (_T_8203) begin
      ic_tag_valid_out_1_91 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_92 <= 1'h0;
    end else if (_T_8219) begin
      ic_tag_valid_out_1_92 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_93 <= 1'h0;
    end else if (_T_8235) begin
      ic_tag_valid_out_1_93 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_94 <= 1'h0;
    end else if (_T_8251) begin
      ic_tag_valid_out_1_94 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_95 <= 1'h0;
    end else if (_T_8267) begin
      ic_tag_valid_out_1_95 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_96 <= 1'h0;
    end else if (_T_8795) begin
      ic_tag_valid_out_1_96 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_97 <= 1'h0;
    end else if (_T_8811) begin
      ic_tag_valid_out_1_97 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_98 <= 1'h0;
    end else if (_T_8827) begin
      ic_tag_valid_out_1_98 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_99 <= 1'h0;
    end else if (_T_8843) begin
      ic_tag_valid_out_1_99 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_100 <= 1'h0;
    end else if (_T_8859) begin
      ic_tag_valid_out_1_100 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_101 <= 1'h0;
    end else if (_T_8875) begin
      ic_tag_valid_out_1_101 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_102 <= 1'h0;
    end else if (_T_8891) begin
      ic_tag_valid_out_1_102 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_103 <= 1'h0;
    end else if (_T_8907) begin
      ic_tag_valid_out_1_103 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_104 <= 1'h0;
    end else if (_T_8923) begin
      ic_tag_valid_out_1_104 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_105 <= 1'h0;
    end else if (_T_8939) begin
      ic_tag_valid_out_1_105 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_106 <= 1'h0;
    end else if (_T_8955) begin
      ic_tag_valid_out_1_106 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_107 <= 1'h0;
    end else if (_T_8971) begin
      ic_tag_valid_out_1_107 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_108 <= 1'h0;
    end else if (_T_8987) begin
      ic_tag_valid_out_1_108 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_109 <= 1'h0;
    end else if (_T_9003) begin
      ic_tag_valid_out_1_109 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_110 <= 1'h0;
    end else if (_T_9019) begin
      ic_tag_valid_out_1_110 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_111 <= 1'h0;
    end else if (_T_9035) begin
      ic_tag_valid_out_1_111 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_112 <= 1'h0;
    end else if (_T_9051) begin
      ic_tag_valid_out_1_112 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_113 <= 1'h0;
    end else if (_T_9067) begin
      ic_tag_valid_out_1_113 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_114 <= 1'h0;
    end else if (_T_9083) begin
      ic_tag_valid_out_1_114 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_115 <= 1'h0;
    end else if (_T_9099) begin
      ic_tag_valid_out_1_115 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_116 <= 1'h0;
    end else if (_T_9115) begin
      ic_tag_valid_out_1_116 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_117 <= 1'h0;
    end else if (_T_9131) begin
      ic_tag_valid_out_1_117 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_118 <= 1'h0;
    end else if (_T_9147) begin
      ic_tag_valid_out_1_118 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_119 <= 1'h0;
    end else if (_T_9163) begin
      ic_tag_valid_out_1_119 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_120 <= 1'h0;
    end else if (_T_9179) begin
      ic_tag_valid_out_1_120 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_121 <= 1'h0;
    end else if (_T_9195) begin
      ic_tag_valid_out_1_121 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_122 <= 1'h0;
    end else if (_T_9211) begin
      ic_tag_valid_out_1_122 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_123 <= 1'h0;
    end else if (_T_9227) begin
      ic_tag_valid_out_1_123 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_124 <= 1'h0;
    end else if (_T_9243) begin
      ic_tag_valid_out_1_124 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_125 <= 1'h0;
    end else if (_T_9259) begin
      ic_tag_valid_out_1_125 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_126 <= 1'h0;
    end else if (_T_9275) begin
      ic_tag_valid_out_1_126 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_1_127 <= 1'h0;
    end else if (_T_9291) begin
      ic_tag_valid_out_1_127 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_0 <= 1'h0;
    end else if (_T_5211) begin
      ic_tag_valid_out_0_0 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_1 <= 1'h0;
    end else if (_T_5227) begin
      ic_tag_valid_out_0_1 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_2 <= 1'h0;
    end else if (_T_5243) begin
      ic_tag_valid_out_0_2 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_3 <= 1'h0;
    end else if (_T_5259) begin
      ic_tag_valid_out_0_3 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_4 <= 1'h0;
    end else if (_T_5275) begin
      ic_tag_valid_out_0_4 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_5 <= 1'h0;
    end else if (_T_5291) begin
      ic_tag_valid_out_0_5 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_6 <= 1'h0;
    end else if (_T_5307) begin
      ic_tag_valid_out_0_6 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_7 <= 1'h0;
    end else if (_T_5323) begin
      ic_tag_valid_out_0_7 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_8 <= 1'h0;
    end else if (_T_5339) begin
      ic_tag_valid_out_0_8 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_9 <= 1'h0;
    end else if (_T_5355) begin
      ic_tag_valid_out_0_9 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_10 <= 1'h0;
    end else if (_T_5371) begin
      ic_tag_valid_out_0_10 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_11 <= 1'h0;
    end else if (_T_5387) begin
      ic_tag_valid_out_0_11 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_12 <= 1'h0;
    end else if (_T_5403) begin
      ic_tag_valid_out_0_12 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_13 <= 1'h0;
    end else if (_T_5419) begin
      ic_tag_valid_out_0_13 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_14 <= 1'h0;
    end else if (_T_5435) begin
      ic_tag_valid_out_0_14 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_15 <= 1'h0;
    end else if (_T_5451) begin
      ic_tag_valid_out_0_15 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_16 <= 1'h0;
    end else if (_T_5467) begin
      ic_tag_valid_out_0_16 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_17 <= 1'h0;
    end else if (_T_5483) begin
      ic_tag_valid_out_0_17 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_18 <= 1'h0;
    end else if (_T_5499) begin
      ic_tag_valid_out_0_18 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_19 <= 1'h0;
    end else if (_T_5515) begin
      ic_tag_valid_out_0_19 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_20 <= 1'h0;
    end else if (_T_5531) begin
      ic_tag_valid_out_0_20 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_21 <= 1'h0;
    end else if (_T_5547) begin
      ic_tag_valid_out_0_21 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_22 <= 1'h0;
    end else if (_T_5563) begin
      ic_tag_valid_out_0_22 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_23 <= 1'h0;
    end else if (_T_5579) begin
      ic_tag_valid_out_0_23 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_24 <= 1'h0;
    end else if (_T_5595) begin
      ic_tag_valid_out_0_24 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_25 <= 1'h0;
    end else if (_T_5611) begin
      ic_tag_valid_out_0_25 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_26 <= 1'h0;
    end else if (_T_5627) begin
      ic_tag_valid_out_0_26 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_27 <= 1'h0;
    end else if (_T_5643) begin
      ic_tag_valid_out_0_27 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_28 <= 1'h0;
    end else if (_T_5659) begin
      ic_tag_valid_out_0_28 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_29 <= 1'h0;
    end else if (_T_5675) begin
      ic_tag_valid_out_0_29 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_30 <= 1'h0;
    end else if (_T_5691) begin
      ic_tag_valid_out_0_30 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_31 <= 1'h0;
    end else if (_T_5707) begin
      ic_tag_valid_out_0_31 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_32 <= 1'h0;
    end else if (_T_6235) begin
      ic_tag_valid_out_0_32 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_33 <= 1'h0;
    end else if (_T_6251) begin
      ic_tag_valid_out_0_33 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_34 <= 1'h0;
    end else if (_T_6267) begin
      ic_tag_valid_out_0_34 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_35 <= 1'h0;
    end else if (_T_6283) begin
      ic_tag_valid_out_0_35 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_36 <= 1'h0;
    end else if (_T_6299) begin
      ic_tag_valid_out_0_36 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_37 <= 1'h0;
    end else if (_T_6315) begin
      ic_tag_valid_out_0_37 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_38 <= 1'h0;
    end else if (_T_6331) begin
      ic_tag_valid_out_0_38 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_39 <= 1'h0;
    end else if (_T_6347) begin
      ic_tag_valid_out_0_39 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_40 <= 1'h0;
    end else if (_T_6363) begin
      ic_tag_valid_out_0_40 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_41 <= 1'h0;
    end else if (_T_6379) begin
      ic_tag_valid_out_0_41 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_42 <= 1'h0;
    end else if (_T_6395) begin
      ic_tag_valid_out_0_42 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_43 <= 1'h0;
    end else if (_T_6411) begin
      ic_tag_valid_out_0_43 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_44 <= 1'h0;
    end else if (_T_6427) begin
      ic_tag_valid_out_0_44 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_45 <= 1'h0;
    end else if (_T_6443) begin
      ic_tag_valid_out_0_45 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_46 <= 1'h0;
    end else if (_T_6459) begin
      ic_tag_valid_out_0_46 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_47 <= 1'h0;
    end else if (_T_6475) begin
      ic_tag_valid_out_0_47 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_48 <= 1'h0;
    end else if (_T_6491) begin
      ic_tag_valid_out_0_48 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_49 <= 1'h0;
    end else if (_T_6507) begin
      ic_tag_valid_out_0_49 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_50 <= 1'h0;
    end else if (_T_6523) begin
      ic_tag_valid_out_0_50 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_51 <= 1'h0;
    end else if (_T_6539) begin
      ic_tag_valid_out_0_51 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_52 <= 1'h0;
    end else if (_T_6555) begin
      ic_tag_valid_out_0_52 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_53 <= 1'h0;
    end else if (_T_6571) begin
      ic_tag_valid_out_0_53 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_54 <= 1'h0;
    end else if (_T_6587) begin
      ic_tag_valid_out_0_54 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_55 <= 1'h0;
    end else if (_T_6603) begin
      ic_tag_valid_out_0_55 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_56 <= 1'h0;
    end else if (_T_6619) begin
      ic_tag_valid_out_0_56 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_57 <= 1'h0;
    end else if (_T_6635) begin
      ic_tag_valid_out_0_57 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_58 <= 1'h0;
    end else if (_T_6651) begin
      ic_tag_valid_out_0_58 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_59 <= 1'h0;
    end else if (_T_6667) begin
      ic_tag_valid_out_0_59 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_60 <= 1'h0;
    end else if (_T_6683) begin
      ic_tag_valid_out_0_60 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_61 <= 1'h0;
    end else if (_T_6699) begin
      ic_tag_valid_out_0_61 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_62 <= 1'h0;
    end else if (_T_6715) begin
      ic_tag_valid_out_0_62 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_63 <= 1'h0;
    end else if (_T_6731) begin
      ic_tag_valid_out_0_63 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_64 <= 1'h0;
    end else if (_T_7259) begin
      ic_tag_valid_out_0_64 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_65 <= 1'h0;
    end else if (_T_7275) begin
      ic_tag_valid_out_0_65 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_66 <= 1'h0;
    end else if (_T_7291) begin
      ic_tag_valid_out_0_66 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_67 <= 1'h0;
    end else if (_T_7307) begin
      ic_tag_valid_out_0_67 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_68 <= 1'h0;
    end else if (_T_7323) begin
      ic_tag_valid_out_0_68 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_69 <= 1'h0;
    end else if (_T_7339) begin
      ic_tag_valid_out_0_69 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_70 <= 1'h0;
    end else if (_T_7355) begin
      ic_tag_valid_out_0_70 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_71 <= 1'h0;
    end else if (_T_7371) begin
      ic_tag_valid_out_0_71 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_72 <= 1'h0;
    end else if (_T_7387) begin
      ic_tag_valid_out_0_72 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_73 <= 1'h0;
    end else if (_T_7403) begin
      ic_tag_valid_out_0_73 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_74 <= 1'h0;
    end else if (_T_7419) begin
      ic_tag_valid_out_0_74 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_75 <= 1'h0;
    end else if (_T_7435) begin
      ic_tag_valid_out_0_75 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_76 <= 1'h0;
    end else if (_T_7451) begin
      ic_tag_valid_out_0_76 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_77 <= 1'h0;
    end else if (_T_7467) begin
      ic_tag_valid_out_0_77 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_78 <= 1'h0;
    end else if (_T_7483) begin
      ic_tag_valid_out_0_78 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_79 <= 1'h0;
    end else if (_T_7499) begin
      ic_tag_valid_out_0_79 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_80 <= 1'h0;
    end else if (_T_7515) begin
      ic_tag_valid_out_0_80 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_81 <= 1'h0;
    end else if (_T_7531) begin
      ic_tag_valid_out_0_81 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_82 <= 1'h0;
    end else if (_T_7547) begin
      ic_tag_valid_out_0_82 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_83 <= 1'h0;
    end else if (_T_7563) begin
      ic_tag_valid_out_0_83 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_84 <= 1'h0;
    end else if (_T_7579) begin
      ic_tag_valid_out_0_84 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_85 <= 1'h0;
    end else if (_T_7595) begin
      ic_tag_valid_out_0_85 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_86 <= 1'h0;
    end else if (_T_7611) begin
      ic_tag_valid_out_0_86 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_87 <= 1'h0;
    end else if (_T_7627) begin
      ic_tag_valid_out_0_87 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_88 <= 1'h0;
    end else if (_T_7643) begin
      ic_tag_valid_out_0_88 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_89 <= 1'h0;
    end else if (_T_7659) begin
      ic_tag_valid_out_0_89 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_90 <= 1'h0;
    end else if (_T_7675) begin
      ic_tag_valid_out_0_90 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_91 <= 1'h0;
    end else if (_T_7691) begin
      ic_tag_valid_out_0_91 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_92 <= 1'h0;
    end else if (_T_7707) begin
      ic_tag_valid_out_0_92 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_93 <= 1'h0;
    end else if (_T_7723) begin
      ic_tag_valid_out_0_93 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_94 <= 1'h0;
    end else if (_T_7739) begin
      ic_tag_valid_out_0_94 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_95 <= 1'h0;
    end else if (_T_7755) begin
      ic_tag_valid_out_0_95 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_96 <= 1'h0;
    end else if (_T_8283) begin
      ic_tag_valid_out_0_96 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_97 <= 1'h0;
    end else if (_T_8299) begin
      ic_tag_valid_out_0_97 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_98 <= 1'h0;
    end else if (_T_8315) begin
      ic_tag_valid_out_0_98 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_99 <= 1'h0;
    end else if (_T_8331) begin
      ic_tag_valid_out_0_99 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_100 <= 1'h0;
    end else if (_T_8347) begin
      ic_tag_valid_out_0_100 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_101 <= 1'h0;
    end else if (_T_8363) begin
      ic_tag_valid_out_0_101 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_102 <= 1'h0;
    end else if (_T_8379) begin
      ic_tag_valid_out_0_102 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_103 <= 1'h0;
    end else if (_T_8395) begin
      ic_tag_valid_out_0_103 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_104 <= 1'h0;
    end else if (_T_8411) begin
      ic_tag_valid_out_0_104 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_105 <= 1'h0;
    end else if (_T_8427) begin
      ic_tag_valid_out_0_105 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_106 <= 1'h0;
    end else if (_T_8443) begin
      ic_tag_valid_out_0_106 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_107 <= 1'h0;
    end else if (_T_8459) begin
      ic_tag_valid_out_0_107 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_108 <= 1'h0;
    end else if (_T_8475) begin
      ic_tag_valid_out_0_108 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_109 <= 1'h0;
    end else if (_T_8491) begin
      ic_tag_valid_out_0_109 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_110 <= 1'h0;
    end else if (_T_8507) begin
      ic_tag_valid_out_0_110 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_111 <= 1'h0;
    end else if (_T_8523) begin
      ic_tag_valid_out_0_111 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_112 <= 1'h0;
    end else if (_T_8539) begin
      ic_tag_valid_out_0_112 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_113 <= 1'h0;
    end else if (_T_8555) begin
      ic_tag_valid_out_0_113 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_114 <= 1'h0;
    end else if (_T_8571) begin
      ic_tag_valid_out_0_114 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_115 <= 1'h0;
    end else if (_T_8587) begin
      ic_tag_valid_out_0_115 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_116 <= 1'h0;
    end else if (_T_8603) begin
      ic_tag_valid_out_0_116 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_117 <= 1'h0;
    end else if (_T_8619) begin
      ic_tag_valid_out_0_117 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_118 <= 1'h0;
    end else if (_T_8635) begin
      ic_tag_valid_out_0_118 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_119 <= 1'h0;
    end else if (_T_8651) begin
      ic_tag_valid_out_0_119 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_120 <= 1'h0;
    end else if (_T_8667) begin
      ic_tag_valid_out_0_120 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_121 <= 1'h0;
    end else if (_T_8683) begin
      ic_tag_valid_out_0_121 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_122 <= 1'h0;
    end else if (_T_8699) begin
      ic_tag_valid_out_0_122 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_123 <= 1'h0;
    end else if (_T_8715) begin
      ic_tag_valid_out_0_123 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_124 <= 1'h0;
    end else if (_T_8731) begin
      ic_tag_valid_out_0_124 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_125 <= 1'h0;
    end else if (_T_8747) begin
      ic_tag_valid_out_0_125 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_126 <= 1'h0;
    end else if (_T_8763) begin
      ic_tag_valid_out_0_126 <= _T_5202;
    end
    if (reset) begin
      ic_tag_valid_out_0_127 <= 1'h0;
    end else if (_T_8779) begin
      ic_tag_valid_out_0_127 <= _T_5202;
    end
    if (reset) begin
      ic_debug_way_ff <= 2'h0;
    end else if (debug_c1_clken) begin
      ic_debug_way_ff <= io_ic_debug_way;
    end
    if (reset) begin
      _T_1212 <= 71'h0;
    end else if (ic_debug_ict_array_sel_ff) begin
      _T_1212 <= {{5'd0}, _T_1211};
    end else begin
      _T_1212 <= io_ic_debug_rd_data;
    end
    if (reset) begin
      ifu_bus_cmd_valid <= 1'h0;
    end else if (_T_2513) begin
      ifu_bus_cmd_valid <= ifc_bus_ic_req_ff_in;
    end
    if (reset) begin
      bus_cmd_beat_count <= 3'h0;
    end else if (_T_2588) begin
      bus_cmd_beat_count <= bus_new_cmd_beat_count;
    end
    if (reset) begin
      ifu_bus_arready_unq_ff <= 1'h0;
    end else if (io_ifu_bus_clk_en) begin
      ifu_bus_arready_unq_ff <= io_ifu_axi_arready;
    end
    if (reset) begin
      ifu_bus_arvalid_ff <= 1'h0;
    end else if (io_ifu_bus_clk_en) begin
      ifu_bus_arvalid_ff <= io_ifu_axi_arvalid;
    end
  end
  always @(posedge io_free_clk) begin
    if (reset) begin
      scnd_miss_req_q <= 1'h0;
    end else begin
      scnd_miss_req_q <= scnd_miss_req_in;
    end
    if (reset) begin
      iccm_dma_rvalid_in <= 1'h0;
    end else begin
      iccm_dma_rvalid_in <= _T_2632;
    end
    if (reset) begin
      dma_iccm_req_f <= 1'h0;
    end else begin
      dma_iccm_req_f <= io_dma_iccm_req;
    end
    if (reset) begin
      perr_state <= 3'h0;
    end else if (perr_state_en) begin
      if (_T_2414) begin
        if (io_iccm_dma_sb_error) begin
          perr_state <= 3'h4;
        end else if (_T_2416) begin
          perr_state <= 3'h1;
        end else begin
          perr_state <= 3'h2;
        end
      end else if (_T_2426) begin
        perr_state <= 3'h0;
      end else if (_T_2429) begin
        if (_T_2431) begin
          perr_state <= 3'h0;
        end else begin
          perr_state <= 3'h3;
        end
      end else if (_T_2435) begin
        if (io_dec_tlu_force_halt) begin
          perr_state <= 3'h0;
        end else begin
          perr_state <= 3'h3;
        end
      end else begin
        perr_state <= 3'h0;
      end
    end
    if (reset) begin
      err_stop_state <= 2'h0;
    end else if (err_stop_state_en) begin
      if (_T_2439) begin
        err_stop_state <= 2'h1;
      end else if (_T_2444) begin
        if (_T_2446) begin
          err_stop_state <= 2'h0;
        end else if (_T_2467) begin
          err_stop_state <= 2'h3;
        end else if (io_ifu_fetch_val[0]) begin
          err_stop_state <= 2'h2;
        end else begin
          err_stop_state <= 2'h1;
        end
      end else if (_T_2471) begin
        if (_T_2446) begin
          err_stop_state <= 2'h0;
        end else if (io_ifu_fetch_val[0]) begin
          err_stop_state <= 2'h3;
        end else begin
          err_stop_state <= 2'h2;
        end
      end else if (_T_2488) begin
        if (_T_2492) begin
          err_stop_state <= 2'h0;
        end else if (io_dec_tlu_flush_err_wb) begin
          err_stop_state <= 2'h1;
        end else begin
          err_stop_state <= 2'h3;
        end
      end else begin
        err_stop_state <= 2'h0;
      end
    end
    if (reset) begin
      bus_ifu_bus_clk_en_ff <= 1'h0;
    end else begin
      bus_ifu_bus_clk_en_ff <= io_ifu_bus_clk_en;
    end
    if (reset) begin
      bus_data_beat_count <= 3'h0;
    end else begin
      bus_data_beat_count <= bus_new_data_beat_count;
    end
    if (reset) begin
      ic_miss_buff_data_valid <= 8'h0;
    end else begin
      ic_miss_buff_data_valid <= _T_1357;
    end
    if (reset) begin
      last_data_recieved_ff <= 1'h0;
    end else begin
      last_data_recieved_ff <= last_data_recieved_in;
    end
    if (reset) begin
      sel_mb_addr_ff <= 1'h0;
    end else begin
      sel_mb_addr_ff <= sel_mb_addr;
    end
    if (reset) begin
      _T_5115 <= 7'h0;
    end else if (_T_3936) begin
      _T_5115 <= io_ic_debug_addr[9:3];
    end else begin
      _T_5115 <= ifu_ic_rw_int_addr[11:5];
    end
    if (reset) begin
      ifu_wr_data_comb_err_ff <= 1'h0;
    end else begin
      ifu_wr_data_comb_err_ff <= ifu_wr_cumulative_err;
    end
    if (reset) begin
      ic_act_miss_f_delayed <= 1'h0;
    end else begin
      ic_act_miss_f_delayed <= ic_act_miss_f;
    end
    if (reset) begin
      ic_crit_wd_rdy_new_ff <= 1'h0;
    end else begin
      ic_crit_wd_rdy_new_ff <= ic_crit_wd_rdy_new_in;
    end
    if (reset) begin
      ic_miss_buff_data_error <= 8'h0;
    end else begin
      ic_miss_buff_data_error <= _T_1397;
    end
    if (reset) begin
      ic_debug_rd_en_ff <= 1'h0;
    end else begin
      ic_debug_rd_en_ff <= io_ic_debug_rd_en;
    end
    if (reset) begin
      ifc_dma_access_ok_prev <= 1'h0;
    end else begin
      ifc_dma_access_ok_prev <= ifc_dma_access_ok_d;
    end
    if (reset) begin
      iccm_ecc_corr_data_ff <= 39'h0;
    end else if (iccm_ecc_write_status) begin
      iccm_ecc_corr_data_ff <= _T_3871;
    end
    if (reset) begin
      dma_mem_addr_ff <= 2'h0;
    end else begin
      dma_mem_addr_ff <= io_dma_mem_addr[3:2];
    end
    if (reset) begin
      dma_mem_tag_ff <= 3'h0;
    end else begin
      dma_mem_tag_ff <= io_dma_mem_tag;
    end
    if (reset) begin
      iccm_dma_rtag <= 3'h0;
    end else begin
      iccm_dma_rtag <= dma_mem_tag_ff;
    end
    if (reset) begin
      iccm_dma_rvalid <= 1'h0;
    end else begin
      iccm_dma_rvalid <= iccm_dma_rvalid_in;
    end
    if (reset) begin
      iccm_dma_rdata <= 64'h0;
    end else if (iccm_dma_ecc_error_in) begin
      iccm_dma_rdata <= _T_3046;
    end else begin
      iccm_dma_rdata <= _T_3047;
    end
    if (reset) begin
      iccm_ecc_corr_index_ff <= 14'h0;
    end else if (iccm_ecc_write_status) begin
      if (iccm_single_ecc_error[0]) begin
        iccm_ecc_corr_index_ff <= iccm_rw_addr_f;
      end else begin
        iccm_ecc_corr_index_ff <= _T_3867;
      end
    end
    if (reset) begin
      iccm_rd_ecc_single_err_ff <= 1'h0;
    end else begin
      iccm_rd_ecc_single_err_ff <= iccm_rd_ecc_single_err_hold_in;
    end
    if (reset) begin
      iccm_rw_addr_f <= 14'h0;
    end else begin
      iccm_rw_addr_f <= io_iccm_rw_addr[14:1];
    end
    if (reset) begin
      ifu_status_wr_addr_ff <= 7'h0;
    end else if (_T_3936) begin
      ifu_status_wr_addr_ff <= io_ic_debug_addr[9:3];
    end else begin
      ifu_status_wr_addr_ff <= ifu_status_wr_addr[11:5];
    end
    if (reset) begin
      way_status_wr_en_ff <= 1'h0;
    end else begin
      way_status_wr_en_ff <= way_status_wr_en_w_debug;
    end
    if (reset) begin
      way_status_new_ff <= 3'h0;
    end else if (_T_3939) begin
      way_status_new_ff <= _T_3943;
    end else begin
      way_status_new_ff <= {{2'd0}, way_status_new};
    end
    if (reset) begin
      ifu_tag_wren_ff <= 2'h0;
    end else begin
      ifu_tag_wren_ff <= ifu_tag_wren_w_debug;
    end
    if (reset) begin
      ic_valid_ff <= 1'h0;
    end else if (_T_3939) begin
      ic_valid_ff <= io_ic_debug_wr_data[0];
    end else begin
      ic_valid_ff <= ic_valid;
    end
    if (reset) begin
      _T_10132 <= 1'h0;
    end else if (ic_debug_rd_en_ff) begin
      _T_10132 <= ic_debug_rd_en_ff;
    end
  end
  always @(posedge io_active_clk) begin
    if (reset) begin
      reset_all_tags <= 1'h0;
    end else begin
      reset_all_tags <= io_dec_tlu_fence_i_wb;
    end
    if (reset) begin
      perr_ic_index_ff <= 6'h0;
    end else if (perr_sb_write_status) begin
      perr_ic_index_ff <= ifu_ic_rw_int_addr_ff;
    end
    if (reset) begin
      dma_sb_err_state_ff <= 1'h0;
    end else begin
      dma_sb_err_state_ff <= _T_7;
    end
    if (reset) begin
      _T_10102 <= 1'h0;
    end else begin
      _T_10102 <= ic_act_miss_f;
    end
    if (reset) begin
      _T_10103 <= 1'h0;
    end else begin
      _T_10103 <= ic_act_hit_f;
    end
    if (reset) begin
      _T_10104 <= 1'h0;
    end else begin
      _T_10104 <= ifc_bus_acc_fault_f;
    end
    if (reset) begin
      _T_10108 <= 1'h0;
    end else begin
      _T_10108 <= _T_10107;
    end
    if (reset) begin
      _T_10109 <= 1'h0;
    end else begin
      _T_10109 <= bus_cmd_sent;
    end
  end
endmodule
