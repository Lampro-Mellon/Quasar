module rvclkhdr(
  output  io_l1clk,
  input   io_clk,
  input   io_en,
  input   io_scan_mode
);
  wire  clkhdr_Q; // @[lib.scala 334:26]
  wire  clkhdr_CK; // @[lib.scala 334:26]
  wire  clkhdr_EN; // @[lib.scala 334:26]
  wire  clkhdr_SE; // @[lib.scala 334:26]
  gated_latch clkhdr ( // @[lib.scala 334:26]
    .Q(clkhdr_Q),
    .CK(clkhdr_CK),
    .EN(clkhdr_EN),
    .SE(clkhdr_SE)
  );
  assign io_l1clk = clkhdr_Q; // @[lib.scala 335:14]
  assign clkhdr_CK = io_clk; // @[lib.scala 336:18]
  assign clkhdr_EN = io_en; // @[lib.scala 337:18]
  assign clkhdr_SE = io_scan_mode; // @[lib.scala 338:18]
endmodule
module ifu_mem_ctl(
  input         clock,
  input         reset,
  input         io_free_clk,
  input         io_active_clk,
  input         io_exu_flush_final,
  input         io_dec_mem_ctrl_dec_tlu_flush_err_wb,
  input         io_dec_mem_ctrl_dec_tlu_i0_commit_cmt,
  input         io_dec_mem_ctrl_dec_tlu_force_halt,
  input         io_dec_mem_ctrl_dec_tlu_fence_i_wb,
  input  [70:0] io_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_wrdata,
  input  [16:0] io_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_dicawics,
  input         io_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_rd_valid,
  input         io_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_wr_valid,
  input         io_dec_mem_ctrl_dec_tlu_core_ecc_disable,
  output        io_dec_mem_ctrl_ifu_pmu_ic_miss,
  output        io_dec_mem_ctrl_ifu_pmu_ic_hit,
  output        io_dec_mem_ctrl_ifu_pmu_bus_error,
  output        io_dec_mem_ctrl_ifu_pmu_bus_busy,
  output        io_dec_mem_ctrl_ifu_pmu_bus_trxn,
  output        io_dec_mem_ctrl_ifu_ic_error_start,
  output        io_dec_mem_ctrl_ifu_iccm_rd_ecc_single_err,
  output [70:0] io_dec_mem_ctrl_ifu_ic_debug_rd_data,
  output        io_dec_mem_ctrl_ifu_ic_debug_rd_data_valid,
  output        io_dec_mem_ctrl_ifu_miss_state_idle,
  input  [30:0] io_ifc_fetch_addr_bf,
  input         io_ifc_fetch_uncacheable_bf,
  input         io_ifc_fetch_req_bf,
  input         io_ifc_fetch_req_bf_raw,
  input         io_ifc_iccm_access_bf,
  input         io_ifc_region_acc_fault_bf,
  input         io_ifc_dma_access_ok,
  input         io_ifu_bp_hit_taken_f,
  input         io_ifu_bp_inst_mask_f,
  input         io_ifu_axi_ar_ready,
  output        io_ifu_axi_ar_valid,
  output [2:0]  io_ifu_axi_ar_bits_id,
  output [31:0] io_ifu_axi_ar_bits_addr,
  output [3:0]  io_ifu_axi_ar_bits_region,
  output        io_ifu_axi_r_ready,
  input         io_ifu_axi_r_valid,
  input  [2:0]  io_ifu_axi_r_bits_id,
  input  [63:0] io_ifu_axi_r_bits_data,
  input  [1:0]  io_ifu_axi_r_bits_resp,
  input         io_ifu_bus_clk_en,
  input         io_dma_mem_ctl_dma_iccm_req,
  input  [31:0] io_dma_mem_ctl_dma_mem_addr,
  input  [2:0]  io_dma_mem_ctl_dma_mem_sz,
  input         io_dma_mem_ctl_dma_mem_write,
  input  [63:0] io_dma_mem_ctl_dma_mem_wdata,
  input  [2:0]  io_dma_mem_ctl_dma_mem_tag,
  output [14:0] io_iccm_rw_addr,
  output        io_iccm_buf_correct_ecc,
  output        io_iccm_correction_state,
  output        io_iccm_wren,
  output        io_iccm_rden,
  output [2:0]  io_iccm_wr_size,
  output [77:0] io_iccm_wr_data,
  input  [63:0] io_iccm_rd_data,
  input  [77:0] io_iccm_rd_data_ecc,
  output [30:0] io_ic_rw_addr,
  output [1:0]  io_ic_tag_valid,
  output [1:0]  io_ic_wr_en,
  output        io_ic_rd_en,
  output [70:0] io_ic_wr_data_0,
  output [70:0] io_ic_wr_data_1,
  output [70:0] io_ic_debug_wr_data,
  output [9:0]  io_ic_debug_addr,
  input  [63:0] io_ic_rd_data,
  input  [70:0] io_ic_debug_rd_data,
  input  [25:0] io_ic_tag_debug_rd_data,
  input  [1:0]  io_ic_eccerr,
  input  [1:0]  io_ic_rd_hit,
  input         io_ic_tag_perr,
  output        io_ic_debug_rd_en,
  output        io_ic_debug_wr_en,
  output        io_ic_debug_tag_array,
  output [1:0]  io_ic_debug_way,
  output [63:0] io_ic_premux_data,
  output        io_ic_sel_premux_data,
  input  [1:0]  io_ifu_fetch_val,
  output        io_ifu_ic_mb_empty,
  output        io_ic_dma_active,
  output        io_ic_write_stall,
  output        io_iccm_dma_ecc_error,
  output        io_iccm_dma_rvalid,
  output [63:0] io_iccm_dma_rdata,
  output [2:0]  io_iccm_dma_rtag,
  output        io_iccm_ready,
  input         io_dec_tlu_flush_lower_wb,
  output        io_iccm_rd_ecc_double_err,
  output        io_iccm_dma_sb_error,
  output        io_ic_hit_f,
  output        io_ic_access_fault_f,
  output [1:0]  io_ic_access_fault_type_f,
  output        io_ifu_async_error_start,
  output [1:0]  io_ic_fetch_val_f,
  output [31:0] io_ic_data_f,
  input         io_scan_mode
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [63:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [95:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [63:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [63:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
`endif // RANDOMIZE_REG_INIT
  wire  rvclkhdr_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_1_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_1_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_1_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_1_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_2_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_2_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_2_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_2_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_3_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_3_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_3_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_3_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_4_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_4_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_4_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_4_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_5_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_5_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_5_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_5_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_6_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_6_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_6_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_6_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_7_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_7_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_7_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_7_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_8_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_8_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_8_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_8_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_9_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_9_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_9_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_9_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_10_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_10_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_10_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_10_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_11_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_11_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_11_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_11_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_12_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_12_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_12_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_12_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_13_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_13_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_13_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_13_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_14_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_14_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_14_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_14_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_15_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_15_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_15_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_15_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_16_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_16_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_16_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_16_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_17_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_17_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_17_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_17_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_18_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_18_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_18_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_18_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_19_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_19_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_19_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_19_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_20_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_20_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_20_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_20_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_21_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_21_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_21_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_21_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_22_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_22_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_22_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_22_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_23_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_23_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_23_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_23_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_24_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_24_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_24_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_24_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_25_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_25_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_25_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_25_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_26_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_26_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_26_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_26_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_27_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_27_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_27_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_27_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_28_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_28_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_28_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_28_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_29_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_29_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_29_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_29_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_30_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_30_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_30_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_30_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_31_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_31_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_31_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_31_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_32_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_32_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_32_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_32_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_33_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_33_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_33_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_33_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_34_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_34_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_34_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_34_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_35_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_35_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_35_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_35_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_36_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_36_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_36_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_36_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_37_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_37_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_37_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_37_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_38_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_38_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_38_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_38_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_39_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_39_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_39_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_39_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_40_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_40_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_40_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_40_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_41_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_41_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_41_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_41_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_42_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_42_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_42_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_42_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_43_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_43_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_43_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_43_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_44_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_44_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_44_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_44_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_45_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_45_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_45_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_45_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_46_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_46_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_46_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_46_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_47_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_47_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_47_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_47_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_48_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_48_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_48_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_48_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_49_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_49_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_49_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_49_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_50_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_50_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_50_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_50_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_51_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_51_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_51_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_51_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_52_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_52_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_52_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_52_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_53_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_53_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_53_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_53_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_54_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_54_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_54_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_54_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_55_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_55_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_55_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_55_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_56_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_56_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_56_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_56_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_57_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_57_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_57_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_57_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_58_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_58_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_58_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_58_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_59_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_59_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_59_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_59_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_60_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_60_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_60_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_60_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_61_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_61_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_61_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_61_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_62_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_62_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_62_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_62_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_63_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_63_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_63_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_63_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_64_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_64_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_64_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_64_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_65_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_65_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_65_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_65_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_66_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_66_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_66_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_66_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_67_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_67_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_67_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_67_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_68_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_68_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_68_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_68_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_69_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_69_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_69_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_69_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_70_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_70_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_70_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_70_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_71_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_71_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_71_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_71_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_72_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_72_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_72_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_72_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_73_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_73_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_73_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_73_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_74_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_74_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_74_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_74_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_75_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_75_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_75_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_75_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_76_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_76_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_76_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_76_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_77_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_77_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_77_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_77_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_78_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_78_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_78_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_78_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_79_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_79_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_79_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_79_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_80_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_80_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_80_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_80_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_81_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_81_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_81_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_81_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_82_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_82_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_82_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_82_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_83_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_83_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_83_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_83_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_84_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_84_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_84_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_84_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_85_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_85_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_85_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_85_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_86_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_86_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_86_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_86_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_87_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_87_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_87_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_87_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_88_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_88_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_88_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_88_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_89_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_89_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_89_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_89_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_90_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_90_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_90_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_90_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_91_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_91_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_91_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_91_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_92_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_92_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_92_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_92_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_93_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_93_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_93_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_93_io_scan_mode; // @[lib.scala 343:22]
  reg  flush_final_f; // @[ifu_mem_ctl.scala 90:53]
  reg  ifc_fetch_req_f_raw; // @[ifu_mem_ctl.scala 227:61]
  wire  _T_319 = ~io_exu_flush_final; // @[ifu_mem_ctl.scala 228:44]
  wire  ifc_fetch_req_f = ifc_fetch_req_f_raw & _T_319; // @[ifu_mem_ctl.scala 228:42]
  wire  _T = io_ifc_fetch_req_bf_raw | ifc_fetch_req_f; // @[ifu_mem_ctl.scala 91:53]
  reg [2:0] miss_state; // @[Reg.scala 27:20]
  wire  miss_pending = miss_state != 3'h0; // @[ifu_mem_ctl.scala 159:30]
  wire  _T_1 = _T | miss_pending; // @[ifu_mem_ctl.scala 91:71]
  wire  _T_2 = _T_1 | io_exu_flush_final; // @[ifu_mem_ctl.scala 91:86]
  reg  scnd_miss_req_q; // @[ifu_mem_ctl.scala 464:52]
  wire  scnd_miss_req = scnd_miss_req_q & _T_319; // @[ifu_mem_ctl.scala 466:36]
  wire  debug_c1_clken = io_ic_debug_rd_en | io_ic_debug_wr_en; // @[ifu_mem_ctl.scala 92:42]
  wire [3:0] ic_fetch_val_int_f = {2'h0,io_ic_fetch_val_f}; // @[Cat.scala 29:58]
  reg [30:0] ifu_fetch_addr_int_f; // @[ifu_mem_ctl.scala 214:63]
  wire [4:0] _GEN_435 = {{1'd0}, ic_fetch_val_int_f}; // @[ifu_mem_ctl.scala 602:53]
  wire [4:0] ic_fetch_val_shift_right = _GEN_435 << ifu_fetch_addr_int_f[0]; // @[ifu_mem_ctl.scala 602:53]
  wire  _T_3129 = |ic_fetch_val_shift_right[3:2]; // @[ifu_mem_ctl.scala 605:91]
  wire  _T_3131 = _T_3129 & _T_319; // @[ifu_mem_ctl.scala 605:95]
  reg  ifc_iccm_access_f; // @[ifu_mem_ctl.scala 229:60]
  wire  fetch_req_iccm_f = ifc_fetch_req_f & ifc_iccm_access_f; // @[ifu_mem_ctl.scala 181:46]
  wire  _T_3132 = _T_3131 & fetch_req_iccm_f; // @[ifu_mem_ctl.scala 605:117]
  reg  iccm_dma_rvalid_in; // @[ifu_mem_ctl.scala 591:59]
  wire  _T_3133 = _T_3132 | iccm_dma_rvalid_in; // @[ifu_mem_ctl.scala 605:134]
  wire  _T_3134 = ~io_dec_mem_ctrl_dec_tlu_core_ecc_disable; // @[ifu_mem_ctl.scala 605:158]
  wire  _T_3135 = _T_3133 & _T_3134; // @[ifu_mem_ctl.scala 605:156]
  wire  _T_3121 = |ic_fetch_val_shift_right[1:0]; // @[ifu_mem_ctl.scala 605:91]
  wire  _T_3123 = _T_3121 & _T_319; // @[ifu_mem_ctl.scala 605:95]
  wire  _T_3124 = _T_3123 & fetch_req_iccm_f; // @[ifu_mem_ctl.scala 605:117]
  wire  _T_3125 = _T_3124 | iccm_dma_rvalid_in; // @[ifu_mem_ctl.scala 605:134]
  wire  _T_3127 = _T_3125 & _T_3134; // @[ifu_mem_ctl.scala 605:156]
  wire [1:0] iccm_ecc_word_enable = {_T_3135,_T_3127}; // @[Cat.scala 29:58]
  wire  _T_3620 = ^io_iccm_rd_data_ecc[70:39]; // @[lib.scala 193:30]
  wire  _T_3621 = ^io_iccm_rd_data_ecc[77:71]; // @[lib.scala 193:44]
  wire  _T_3622 = _T_3620 ^ _T_3621; // @[lib.scala 193:35]
  wire [5:0] _T_3630 = {io_iccm_rd_data_ecc[70],io_iccm_rd_data_ecc[69],io_iccm_rd_data_ecc[68],io_iccm_rd_data_ecc[67],io_iccm_rd_data_ecc[66],io_iccm_rd_data_ecc[65]}; // @[lib.scala 193:76]
  wire  _T_3631 = ^_T_3630; // @[lib.scala 193:83]
  wire  _T_3632 = io_iccm_rd_data_ecc[76] ^ _T_3631; // @[lib.scala 193:71]
  wire [6:0] _T_3639 = {io_iccm_rd_data_ecc[56],io_iccm_rd_data_ecc[55],io_iccm_rd_data_ecc[54],io_iccm_rd_data_ecc[53],io_iccm_rd_data_ecc[52],io_iccm_rd_data_ecc[51],io_iccm_rd_data_ecc[50]}; // @[lib.scala 193:103]
  wire [14:0] _T_3647 = {io_iccm_rd_data_ecc[64],io_iccm_rd_data_ecc[63],io_iccm_rd_data_ecc[62],io_iccm_rd_data_ecc[61],io_iccm_rd_data_ecc[60],io_iccm_rd_data_ecc[59],io_iccm_rd_data_ecc[58],io_iccm_rd_data_ecc[57],_T_3639}; // @[lib.scala 193:103]
  wire  _T_3648 = ^_T_3647; // @[lib.scala 193:110]
  wire  _T_3649 = io_iccm_rd_data_ecc[75] ^ _T_3648; // @[lib.scala 193:98]
  wire [6:0] _T_3656 = {io_iccm_rd_data_ecc[49],io_iccm_rd_data_ecc[48],io_iccm_rd_data_ecc[47],io_iccm_rd_data_ecc[46],io_iccm_rd_data_ecc[45],io_iccm_rd_data_ecc[44],io_iccm_rd_data_ecc[43]}; // @[lib.scala 193:130]
  wire [14:0] _T_3664 = {io_iccm_rd_data_ecc[64],io_iccm_rd_data_ecc[63],io_iccm_rd_data_ecc[62],io_iccm_rd_data_ecc[61],io_iccm_rd_data_ecc[60],io_iccm_rd_data_ecc[59],io_iccm_rd_data_ecc[58],io_iccm_rd_data_ecc[57],_T_3656}; // @[lib.scala 193:130]
  wire  _T_3665 = ^_T_3664; // @[lib.scala 193:137]
  wire  _T_3666 = io_iccm_rd_data_ecc[74] ^ _T_3665; // @[lib.scala 193:125]
  wire [8:0] _T_3675 = {io_iccm_rd_data_ecc[54],io_iccm_rd_data_ecc[53],io_iccm_rd_data_ecc[49],io_iccm_rd_data_ecc[48],io_iccm_rd_data_ecc[47],io_iccm_rd_data_ecc[46],io_iccm_rd_data_ecc[42],io_iccm_rd_data_ecc[41],io_iccm_rd_data_ecc[40]}; // @[lib.scala 193:157]
  wire [17:0] _T_3684 = {io_iccm_rd_data_ecc[70],io_iccm_rd_data_ecc[69],io_iccm_rd_data_ecc[68],io_iccm_rd_data_ecc[64],io_iccm_rd_data_ecc[63],io_iccm_rd_data_ecc[62],io_iccm_rd_data_ecc[61],io_iccm_rd_data_ecc[56],io_iccm_rd_data_ecc[55],_T_3675}; // @[lib.scala 193:157]
  wire  _T_3685 = ^_T_3684; // @[lib.scala 193:164]
  wire  _T_3686 = io_iccm_rd_data_ecc[73] ^ _T_3685; // @[lib.scala 193:152]
  wire [8:0] _T_3695 = {io_iccm_rd_data_ecc[52],io_iccm_rd_data_ecc[51],io_iccm_rd_data_ecc[49],io_iccm_rd_data_ecc[48],io_iccm_rd_data_ecc[45],io_iccm_rd_data_ecc[44],io_iccm_rd_data_ecc[42],io_iccm_rd_data_ecc[41],io_iccm_rd_data_ecc[39]}; // @[lib.scala 193:184]
  wire [17:0] _T_3704 = {io_iccm_rd_data_ecc[70],io_iccm_rd_data_ecc[67],io_iccm_rd_data_ecc[66],io_iccm_rd_data_ecc[64],io_iccm_rd_data_ecc[63],io_iccm_rd_data_ecc[60],io_iccm_rd_data_ecc[59],io_iccm_rd_data_ecc[56],io_iccm_rd_data_ecc[55],_T_3695}; // @[lib.scala 193:184]
  wire  _T_3705 = ^_T_3704; // @[lib.scala 193:191]
  wire  _T_3706 = io_iccm_rd_data_ecc[72] ^ _T_3705; // @[lib.scala 193:179]
  wire [8:0] _T_3715 = {io_iccm_rd_data_ecc[52],io_iccm_rd_data_ecc[50],io_iccm_rd_data_ecc[49],io_iccm_rd_data_ecc[47],io_iccm_rd_data_ecc[45],io_iccm_rd_data_ecc[43],io_iccm_rd_data_ecc[42],io_iccm_rd_data_ecc[40],io_iccm_rd_data_ecc[39]}; // @[lib.scala 193:211]
  wire [17:0] _T_3724 = {io_iccm_rd_data_ecc[69],io_iccm_rd_data_ecc[67],io_iccm_rd_data_ecc[65],io_iccm_rd_data_ecc[64],io_iccm_rd_data_ecc[62],io_iccm_rd_data_ecc[60],io_iccm_rd_data_ecc[58],io_iccm_rd_data_ecc[56],io_iccm_rd_data_ecc[54],_T_3715}; // @[lib.scala 193:211]
  wire  _T_3725 = ^_T_3724; // @[lib.scala 193:218]
  wire  _T_3726 = io_iccm_rd_data_ecc[71] ^ _T_3725; // @[lib.scala 193:206]
  wire [6:0] _T_3732 = {_T_3622,_T_3632,_T_3649,_T_3666,_T_3686,_T_3706,_T_3726}; // @[Cat.scala 29:58]
  wire  _T_3733 = _T_3732 != 7'h0; // @[lib.scala 194:44]
  wire  _T_3734 = iccm_ecc_word_enable[1] & _T_3733; // @[lib.scala 194:32]
  wire  _T_3736 = _T_3734 & _T_3732[6]; // @[lib.scala 194:53]
  wire  _T_3235 = ^io_iccm_rd_data_ecc[31:0]; // @[lib.scala 193:30]
  wire  _T_3236 = ^io_iccm_rd_data_ecc[38:32]; // @[lib.scala 193:44]
  wire  _T_3237 = _T_3235 ^ _T_3236; // @[lib.scala 193:35]
  wire [5:0] _T_3245 = {io_iccm_rd_data_ecc[31],io_iccm_rd_data_ecc[30],io_iccm_rd_data_ecc[29],io_iccm_rd_data_ecc[28],io_iccm_rd_data_ecc[27],io_iccm_rd_data_ecc[26]}; // @[lib.scala 193:76]
  wire  _T_3246 = ^_T_3245; // @[lib.scala 193:83]
  wire  _T_3247 = io_iccm_rd_data_ecc[37] ^ _T_3246; // @[lib.scala 193:71]
  wire [6:0] _T_3254 = {io_iccm_rd_data_ecc[17],io_iccm_rd_data_ecc[16],io_iccm_rd_data_ecc[15],io_iccm_rd_data_ecc[14],io_iccm_rd_data_ecc[13],io_iccm_rd_data_ecc[12],io_iccm_rd_data_ecc[11]}; // @[lib.scala 193:103]
  wire [14:0] _T_3262 = {io_iccm_rd_data_ecc[25],io_iccm_rd_data_ecc[24],io_iccm_rd_data_ecc[23],io_iccm_rd_data_ecc[22],io_iccm_rd_data_ecc[21],io_iccm_rd_data_ecc[20],io_iccm_rd_data_ecc[19],io_iccm_rd_data_ecc[18],_T_3254}; // @[lib.scala 193:103]
  wire  _T_3263 = ^_T_3262; // @[lib.scala 193:110]
  wire  _T_3264 = io_iccm_rd_data_ecc[36] ^ _T_3263; // @[lib.scala 193:98]
  wire [6:0] _T_3271 = {io_iccm_rd_data_ecc[10],io_iccm_rd_data_ecc[9],io_iccm_rd_data_ecc[8],io_iccm_rd_data_ecc[7],io_iccm_rd_data_ecc[6],io_iccm_rd_data_ecc[5],io_iccm_rd_data_ecc[4]}; // @[lib.scala 193:130]
  wire [14:0] _T_3279 = {io_iccm_rd_data_ecc[25],io_iccm_rd_data_ecc[24],io_iccm_rd_data_ecc[23],io_iccm_rd_data_ecc[22],io_iccm_rd_data_ecc[21],io_iccm_rd_data_ecc[20],io_iccm_rd_data_ecc[19],io_iccm_rd_data_ecc[18],_T_3271}; // @[lib.scala 193:130]
  wire  _T_3280 = ^_T_3279; // @[lib.scala 193:137]
  wire  _T_3281 = io_iccm_rd_data_ecc[35] ^ _T_3280; // @[lib.scala 193:125]
  wire [8:0] _T_3290 = {io_iccm_rd_data_ecc[15],io_iccm_rd_data_ecc[14],io_iccm_rd_data_ecc[10],io_iccm_rd_data_ecc[9],io_iccm_rd_data_ecc[8],io_iccm_rd_data_ecc[7],io_iccm_rd_data_ecc[3],io_iccm_rd_data_ecc[2],io_iccm_rd_data_ecc[1]}; // @[lib.scala 193:157]
  wire [17:0] _T_3299 = {io_iccm_rd_data_ecc[31],io_iccm_rd_data_ecc[30],io_iccm_rd_data_ecc[29],io_iccm_rd_data_ecc[25],io_iccm_rd_data_ecc[24],io_iccm_rd_data_ecc[23],io_iccm_rd_data_ecc[22],io_iccm_rd_data_ecc[17],io_iccm_rd_data_ecc[16],_T_3290}; // @[lib.scala 193:157]
  wire  _T_3300 = ^_T_3299; // @[lib.scala 193:164]
  wire  _T_3301 = io_iccm_rd_data_ecc[34] ^ _T_3300; // @[lib.scala 193:152]
  wire [8:0] _T_3310 = {io_iccm_rd_data_ecc[13],io_iccm_rd_data_ecc[12],io_iccm_rd_data_ecc[10],io_iccm_rd_data_ecc[9],io_iccm_rd_data_ecc[6],io_iccm_rd_data_ecc[5],io_iccm_rd_data_ecc[3],io_iccm_rd_data_ecc[2],io_iccm_rd_data_ecc[0]}; // @[lib.scala 193:184]
  wire [17:0] _T_3319 = {io_iccm_rd_data_ecc[31],io_iccm_rd_data_ecc[28],io_iccm_rd_data_ecc[27],io_iccm_rd_data_ecc[25],io_iccm_rd_data_ecc[24],io_iccm_rd_data_ecc[21],io_iccm_rd_data_ecc[20],io_iccm_rd_data_ecc[17],io_iccm_rd_data_ecc[16],_T_3310}; // @[lib.scala 193:184]
  wire  _T_3320 = ^_T_3319; // @[lib.scala 193:191]
  wire  _T_3321 = io_iccm_rd_data_ecc[33] ^ _T_3320; // @[lib.scala 193:179]
  wire [8:0] _T_3330 = {io_iccm_rd_data_ecc[13],io_iccm_rd_data_ecc[11],io_iccm_rd_data_ecc[10],io_iccm_rd_data_ecc[8],io_iccm_rd_data_ecc[6],io_iccm_rd_data_ecc[4],io_iccm_rd_data_ecc[3],io_iccm_rd_data_ecc[1],io_iccm_rd_data_ecc[0]}; // @[lib.scala 193:211]
  wire [17:0] _T_3339 = {io_iccm_rd_data_ecc[30],io_iccm_rd_data_ecc[28],io_iccm_rd_data_ecc[26],io_iccm_rd_data_ecc[25],io_iccm_rd_data_ecc[23],io_iccm_rd_data_ecc[21],io_iccm_rd_data_ecc[19],io_iccm_rd_data_ecc[17],io_iccm_rd_data_ecc[15],_T_3330}; // @[lib.scala 193:211]
  wire  _T_3340 = ^_T_3339; // @[lib.scala 193:218]
  wire  _T_3341 = io_iccm_rd_data_ecc[32] ^ _T_3340; // @[lib.scala 193:206]
  wire [6:0] _T_3347 = {_T_3237,_T_3247,_T_3264,_T_3281,_T_3301,_T_3321,_T_3341}; // @[Cat.scala 29:58]
  wire  _T_3348 = _T_3347 != 7'h0; // @[lib.scala 194:44]
  wire  _T_3349 = iccm_ecc_word_enable[0] & _T_3348; // @[lib.scala 194:32]
  wire  _T_3351 = _T_3349 & _T_3347[6]; // @[lib.scala 194:53]
  wire [1:0] iccm_single_ecc_error = {_T_3736,_T_3351}; // @[Cat.scala 29:58]
  wire  _T_3 = |iccm_single_ecc_error; // @[ifu_mem_ctl.scala 95:52]
  reg  dma_iccm_req_f; // @[ifu_mem_ctl.scala 568:51]
  wire  _T_6 = io_dec_mem_ctrl_ifu_iccm_rd_ecc_single_err | io_dec_mem_ctrl_ifu_ic_error_start; // @[ifu_mem_ctl.scala 96:74]
  reg [2:0] perr_state; // @[Reg.scala 27:20]
  wire  _T_7 = perr_state == 3'h4; // @[ifu_mem_ctl.scala 97:54]
  wire  iccm_correct_ecc = perr_state == 3'h3; // @[ifu_mem_ctl.scala 392:34]
  wire  _T_8 = iccm_correct_ecc | _T_7; // @[ifu_mem_ctl.scala 97:40]
  reg [1:0] err_stop_state; // @[Reg.scala 27:20]
  wire  _T_9 = err_stop_state == 2'h3; // @[ifu_mem_ctl.scala 97:90]
  wire  _T_10 = _T_8 | _T_9; // @[ifu_mem_ctl.scala 97:72]
  wire  _T_2526 = 2'h0 == err_stop_state; // @[Conditional.scala 37:30]
  wire  _T_2531 = 2'h1 == err_stop_state; // @[Conditional.scala 37:30]
  wire  _T_2551 = io_ifu_fetch_val == 2'h3; // @[ifu_mem_ctl.scala 441:48]
  wire  two_byte_instr = io_ic_data_f[1:0] != 2'h3; // @[ifu_mem_ctl.scala 306:42]
  wire  _T_2553 = io_ifu_fetch_val[0] & two_byte_instr; // @[ifu_mem_ctl.scala 441:79]
  wire  _T_2554 = _T_2551 | _T_2553; // @[ifu_mem_ctl.scala 441:56]
  wire  _T_2555 = io_exu_flush_final | io_dec_mem_ctrl_dec_tlu_i0_commit_cmt; // @[ifu_mem_ctl.scala 441:122]
  wire  _T_2556 = ~_T_2555; // @[ifu_mem_ctl.scala 441:101]
  wire  _T_2557 = _T_2554 & _T_2556; // @[ifu_mem_ctl.scala 441:99]
  wire  _T_2558 = 2'h2 == err_stop_state; // @[Conditional.scala 37:30]
  wire  _T_2572 = io_ifu_fetch_val[0] & _T_319; // @[ifu_mem_ctl.scala 448:45]
  wire  _T_2573 = ~io_dec_mem_ctrl_dec_tlu_i0_commit_cmt; // @[ifu_mem_ctl.scala 448:69]
  wire  _T_2574 = _T_2572 & _T_2573; // @[ifu_mem_ctl.scala 448:67]
  wire  _T_2575 = 2'h3 == err_stop_state; // @[Conditional.scala 37:30]
  wire  _GEN_37 = _T_2558 ? _T_2574 : _T_2575; // @[Conditional.scala 39:67]
  wire  _GEN_41 = _T_2531 ? _T_2557 : _GEN_37; // @[Conditional.scala 39:67]
  wire  err_stop_fetch = _T_2526 ? 1'h0 : _GEN_41; // @[Conditional.scala 40:58]
  wire  _T_11 = _T_10 | err_stop_fetch; // @[ifu_mem_ctl.scala 97:112]
  wire  _T_13 = io_ifu_axi_r_valid & io_ifu_bus_clk_en; // @[ifu_mem_ctl.scala 99:44]
  wire  _T_14 = _T_13 & io_ifu_axi_r_ready; // @[ifu_mem_ctl.scala 99:65]
  wire  _T_227 = |io_ic_rd_hit; // @[ifu_mem_ctl.scala 189:37]
  wire  _T_228 = ~_T_227; // @[ifu_mem_ctl.scala 189:23]
  reg  reset_all_tags; // @[ifu_mem_ctl.scala 637:53]
  wire  _T_229 = _T_228 | reset_all_tags; // @[ifu_mem_ctl.scala 189:41]
  wire  _T_207 = ~ifc_iccm_access_f; // @[ifu_mem_ctl.scala 180:48]
  wire  _T_208 = ifc_fetch_req_f & _T_207; // @[ifu_mem_ctl.scala 180:46]
  reg  ifc_region_acc_fault_final_f; // @[ifu_mem_ctl.scala 231:71]
  wire  _T_209 = ~ifc_region_acc_fault_final_f; // @[ifu_mem_ctl.scala 180:69]
  wire  fetch_req_icache_f = _T_208 & _T_209; // @[ifu_mem_ctl.scala 180:67]
  wire  _T_230 = _T_229 & fetch_req_icache_f; // @[ifu_mem_ctl.scala 189:59]
  wire  _T_231 = ~miss_pending; // @[ifu_mem_ctl.scala 189:82]
  wire  _T_232 = _T_230 & _T_231; // @[ifu_mem_ctl.scala 189:80]
  wire  _T_233 = _T_232 | scnd_miss_req; // @[ifu_mem_ctl.scala 189:97]
  wire  ic_act_miss_f = _T_233 & _T_209; // @[ifu_mem_ctl.scala 189:114]
  reg  ifu_bus_rvalid_unq_ff; // @[ifu_mem_ctl.scala 510:56]
  reg  bus_ifu_bus_clk_en_ff; // @[ifu_mem_ctl.scala 463:61]
  wire  ifu_bus_rvalid_ff = ifu_bus_rvalid_unq_ff & bus_ifu_bus_clk_en_ff; // @[ifu_mem_ctl.scala 524:49]
  wire  bus_ifu_wr_en_ff = ifu_bus_rvalid_ff & miss_pending; // @[ifu_mem_ctl.scala 552:41]
  reg  uncacheable_miss_ff; // @[ifu_mem_ctl.scala 216:62]
  reg [2:0] bus_data_beat_count; // @[ifu_mem_ctl.scala 533:56]
  wire  _T_2672 = bus_data_beat_count == 3'h1; // @[ifu_mem_ctl.scala 550:69]
  wire  _T_2673 = &bus_data_beat_count; // @[ifu_mem_ctl.scala 550:101]
  wire  bus_last_data_beat = uncacheable_miss_ff ? _T_2672 : _T_2673; // @[ifu_mem_ctl.scala 550:28]
  wire  _T_2624 = bus_ifu_wr_en_ff & bus_last_data_beat; // @[ifu_mem_ctl.scala 529:68]
  wire  _T_2625 = ic_act_miss_f | _T_2624; // @[ifu_mem_ctl.scala 529:48]
  wire  bus_reset_data_beat_cnt = _T_2625 | io_dec_mem_ctrl_dec_tlu_force_halt; // @[ifu_mem_ctl.scala 529:91]
  wire  _T_2621 = ~bus_last_data_beat; // @[ifu_mem_ctl.scala 528:50]
  wire  _T_2622 = bus_ifu_wr_en_ff & _T_2621; // @[ifu_mem_ctl.scala 528:48]
  wire  _T_2623 = ~io_dec_mem_ctrl_dec_tlu_force_halt; // @[ifu_mem_ctl.scala 528:72]
  wire  bus_inc_data_beat_cnt = _T_2622 & _T_2623; // @[ifu_mem_ctl.scala 528:70]
  wire [2:0] _T_2629 = bus_data_beat_count + 3'h1; // @[ifu_mem_ctl.scala 532:115]
  wire [2:0] _T_2631 = bus_inc_data_beat_cnt ? _T_2629 : 3'h0; // @[Mux.scala 27:72]
  wire  _T_2626 = ~bus_inc_data_beat_cnt; // @[ifu_mem_ctl.scala 530:32]
  wire  _T_2627 = ~bus_reset_data_beat_cnt; // @[ifu_mem_ctl.scala 530:57]
  wire  bus_hold_data_beat_cnt = _T_2626 & _T_2627; // @[ifu_mem_ctl.scala 530:55]
  wire [2:0] _T_2632 = bus_hold_data_beat_cnt ? bus_data_beat_count : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] bus_new_data_beat_count = _T_2631 | _T_2632; // @[Mux.scala 27:72]
  wire  _T_15 = &bus_new_data_beat_count; // @[ifu_mem_ctl.scala 99:112]
  wire  _T_16 = _T_14 & _T_15; // @[ifu_mem_ctl.scala 99:85]
  wire  _T_17 = ~uncacheable_miss_ff; // @[ifu_mem_ctl.scala 100:5]
  wire  _T_18 = _T_16 & _T_17; // @[ifu_mem_ctl.scala 99:118]
  wire  _T_19 = miss_state == 3'h5; // @[ifu_mem_ctl.scala 100:41]
  wire  _T_24 = 3'h0 == miss_state; // @[Conditional.scala 37:30]
  wire  _T_26 = ic_act_miss_f & _T_319; // @[ifu_mem_ctl.scala 106:43]
  wire [2:0] _T_28 = _T_26 ? 3'h1 : 3'h2; // @[ifu_mem_ctl.scala 106:27]
  wire  _T_31 = 3'h1 == miss_state; // @[Conditional.scala 37:30]
  wire [4:0] byp_fetch_index = ifu_fetch_addr_int_f[4:0]; // @[ifu_mem_ctl.scala 343:45]
  wire  _T_2155 = byp_fetch_index[4:2] == 3'h0; // @[ifu_mem_ctl.scala 364:127]
  reg [7:0] ic_miss_buff_data_valid; // @[ifu_mem_ctl.scala 320:60]
  wire  _T_2186 = _T_2155 & ic_miss_buff_data_valid[0]; // @[Mux.scala 27:72]
  wire  _T_2159 = byp_fetch_index[4:2] == 3'h1; // @[ifu_mem_ctl.scala 364:127]
  wire  _T_2187 = _T_2159 & ic_miss_buff_data_valid[1]; // @[Mux.scala 27:72]
  wire  _T_2194 = _T_2186 | _T_2187; // @[Mux.scala 27:72]
  wire  _T_2163 = byp_fetch_index[4:2] == 3'h2; // @[ifu_mem_ctl.scala 364:127]
  wire  _T_2188 = _T_2163 & ic_miss_buff_data_valid[2]; // @[Mux.scala 27:72]
  wire  _T_2195 = _T_2194 | _T_2188; // @[Mux.scala 27:72]
  wire  _T_2167 = byp_fetch_index[4:2] == 3'h3; // @[ifu_mem_ctl.scala 364:127]
  wire  _T_2189 = _T_2167 & ic_miss_buff_data_valid[3]; // @[Mux.scala 27:72]
  wire  _T_2196 = _T_2195 | _T_2189; // @[Mux.scala 27:72]
  wire  _T_2171 = byp_fetch_index[4:2] == 3'h4; // @[ifu_mem_ctl.scala 364:127]
  wire  _T_2190 = _T_2171 & ic_miss_buff_data_valid[4]; // @[Mux.scala 27:72]
  wire  _T_2197 = _T_2196 | _T_2190; // @[Mux.scala 27:72]
  wire  _T_2175 = byp_fetch_index[4:2] == 3'h5; // @[ifu_mem_ctl.scala 364:127]
  wire  _T_2191 = _T_2175 & ic_miss_buff_data_valid[5]; // @[Mux.scala 27:72]
  wire  _T_2198 = _T_2197 | _T_2191; // @[Mux.scala 27:72]
  wire  _T_2179 = byp_fetch_index[4:2] == 3'h6; // @[ifu_mem_ctl.scala 364:127]
  wire  _T_2192 = _T_2179 & ic_miss_buff_data_valid[6]; // @[Mux.scala 27:72]
  wire  _T_2199 = _T_2198 | _T_2192; // @[Mux.scala 27:72]
  wire  _T_2183 = byp_fetch_index[4:2] == 3'h7; // @[ifu_mem_ctl.scala 364:127]
  wire  _T_2193 = _T_2183 & ic_miss_buff_data_valid[7]; // @[Mux.scala 27:72]
  wire  ic_miss_buff_data_valid_bypass_index = _T_2199 | _T_2193; // @[Mux.scala 27:72]
  wire  _T_2241 = ~byp_fetch_index[1]; // @[ifu_mem_ctl.scala 366:69]
  wire  _T_2242 = ic_miss_buff_data_valid_bypass_index & _T_2241; // @[ifu_mem_ctl.scala 366:67]
  wire  _T_2244 = ~byp_fetch_index[0]; // @[ifu_mem_ctl.scala 366:91]
  wire  _T_2245 = _T_2242 & _T_2244; // @[ifu_mem_ctl.scala 366:89]
  wire  _T_2250 = _T_2242 & byp_fetch_index[0]; // @[ifu_mem_ctl.scala 367:65]
  wire  _T_2251 = _T_2245 | _T_2250; // @[ifu_mem_ctl.scala 366:112]
  wire  _T_2253 = ic_miss_buff_data_valid_bypass_index & byp_fetch_index[1]; // @[ifu_mem_ctl.scala 368:43]
  wire  _T_2256 = _T_2253 & _T_2244; // @[ifu_mem_ctl.scala 368:65]
  wire  _T_2257 = _T_2251 | _T_2256; // @[ifu_mem_ctl.scala 367:88]
  wire  _T_2261 = _T_2253 & byp_fetch_index[0]; // @[ifu_mem_ctl.scala 369:65]
  wire [2:0] byp_fetch_index_inc = ifu_fetch_addr_int_f[4:2] + 3'h1; // @[ifu_mem_ctl.scala 346:75]
  wire  _T_2201 = byp_fetch_index_inc == 3'h0; // @[ifu_mem_ctl.scala 365:110]
  wire  _T_2225 = _T_2201 & ic_miss_buff_data_valid[0]; // @[Mux.scala 27:72]
  wire  _T_2204 = byp_fetch_index_inc == 3'h1; // @[ifu_mem_ctl.scala 365:110]
  wire  _T_2226 = _T_2204 & ic_miss_buff_data_valid[1]; // @[Mux.scala 27:72]
  wire  _T_2233 = _T_2225 | _T_2226; // @[Mux.scala 27:72]
  wire  _T_2207 = byp_fetch_index_inc == 3'h2; // @[ifu_mem_ctl.scala 365:110]
  wire  _T_2227 = _T_2207 & ic_miss_buff_data_valid[2]; // @[Mux.scala 27:72]
  wire  _T_2234 = _T_2233 | _T_2227; // @[Mux.scala 27:72]
  wire  _T_2210 = byp_fetch_index_inc == 3'h3; // @[ifu_mem_ctl.scala 365:110]
  wire  _T_2228 = _T_2210 & ic_miss_buff_data_valid[3]; // @[Mux.scala 27:72]
  wire  _T_2235 = _T_2234 | _T_2228; // @[Mux.scala 27:72]
  wire  _T_2213 = byp_fetch_index_inc == 3'h4; // @[ifu_mem_ctl.scala 365:110]
  wire  _T_2229 = _T_2213 & ic_miss_buff_data_valid[4]; // @[Mux.scala 27:72]
  wire  _T_2236 = _T_2235 | _T_2229; // @[Mux.scala 27:72]
  wire  _T_2216 = byp_fetch_index_inc == 3'h5; // @[ifu_mem_ctl.scala 365:110]
  wire  _T_2230 = _T_2216 & ic_miss_buff_data_valid[5]; // @[Mux.scala 27:72]
  wire  _T_2237 = _T_2236 | _T_2230; // @[Mux.scala 27:72]
  wire  _T_2219 = byp_fetch_index_inc == 3'h6; // @[ifu_mem_ctl.scala 365:110]
  wire  _T_2231 = _T_2219 & ic_miss_buff_data_valid[6]; // @[Mux.scala 27:72]
  wire  _T_2238 = _T_2237 | _T_2231; // @[Mux.scala 27:72]
  wire  _T_2222 = byp_fetch_index_inc == 3'h7; // @[ifu_mem_ctl.scala 365:110]
  wire  _T_2232 = _T_2222 & ic_miss_buff_data_valid[7]; // @[Mux.scala 27:72]
  wire  ic_miss_buff_data_valid_inc_bypass_index = _T_2238 | _T_2232; // @[Mux.scala 27:72]
  wire  _T_2262 = _T_2261 & ic_miss_buff_data_valid_inc_bypass_index; // @[ifu_mem_ctl.scala 369:87]
  wire  _T_2263 = _T_2257 | _T_2262; // @[ifu_mem_ctl.scala 368:88]
  wire  _T_2267 = ic_miss_buff_data_valid_bypass_index & _T_2183; // @[ifu_mem_ctl.scala 370:43]
  wire  miss_buff_hit_unq_f = _T_2263 | _T_2267; // @[ifu_mem_ctl.scala 369:131]
  wire  _T_2283 = miss_state == 3'h4; // @[ifu_mem_ctl.scala 375:55]
  wire  _T_2284 = miss_state == 3'h1; // @[ifu_mem_ctl.scala 375:87]
  wire  _T_2285 = _T_2283 | _T_2284; // @[ifu_mem_ctl.scala 375:74]
  wire  crit_byp_hit_f = miss_buff_hit_unq_f & _T_2285; // @[ifu_mem_ctl.scala 375:41]
  wire  _T_2268 = miss_state == 3'h6; // @[ifu_mem_ctl.scala 372:30]
  reg [30:0] imb_ff; // @[ifu_mem_ctl.scala 217:49]
  wire  miss_wrap_f = imb_ff[5] != ifu_fetch_addr_int_f[5]; // @[ifu_mem_ctl.scala 363:51]
  wire  _T_2269 = ~miss_wrap_f; // @[ifu_mem_ctl.scala 372:68]
  wire  _T_2270 = miss_buff_hit_unq_f & _T_2269; // @[ifu_mem_ctl.scala 372:66]
  wire  stream_hit_f = _T_2268 & _T_2270; // @[ifu_mem_ctl.scala 372:43]
  wire  _T_215 = crit_byp_hit_f | stream_hit_f; // @[ifu_mem_ctl.scala 184:35]
  wire  _T_216 = _T_215 & fetch_req_icache_f; // @[ifu_mem_ctl.scala 184:52]
  wire  ic_byp_hit_f = _T_216 & miss_pending; // @[ifu_mem_ctl.scala 184:73]
  reg  last_data_recieved_ff; // @[ifu_mem_ctl.scala 535:58]
  wire  last_beat = bus_last_data_beat & bus_ifu_wr_en_ff; // @[ifu_mem_ctl.scala 562:35]
  wire  _T_32 = bus_ifu_wr_en_ff & last_beat; // @[ifu_mem_ctl.scala 110:126]
  wire  _T_33 = last_data_recieved_ff | _T_32; // @[ifu_mem_ctl.scala 110:106]
  wire  _T_34 = ic_byp_hit_f & _T_33; // @[ifu_mem_ctl.scala 110:80]
  wire  _T_35 = _T_34 & uncacheable_miss_ff; // @[ifu_mem_ctl.scala 110:140]
  wire  _T_36 = io_dec_mem_ctrl_dec_tlu_force_halt | _T_35; // @[ifu_mem_ctl.scala 110:64]
  wire  _T_38 = ~last_data_recieved_ff; // @[ifu_mem_ctl.scala 111:30]
  wire  _T_39 = ic_byp_hit_f & _T_38; // @[ifu_mem_ctl.scala 111:27]
  wire  _T_40 = _T_39 & uncacheable_miss_ff; // @[ifu_mem_ctl.scala 111:53]
  wire  _T_42 = ~ic_byp_hit_f; // @[ifu_mem_ctl.scala 112:16]
  wire  _T_44 = _T_42 & _T_319; // @[ifu_mem_ctl.scala 112:30]
  wire  _T_46 = _T_44 & _T_32; // @[ifu_mem_ctl.scala 112:52]
  wire  _T_47 = _T_46 & uncacheable_miss_ff; // @[ifu_mem_ctl.scala 112:85]
  wire  _T_51 = _T_32 & _T_17; // @[ifu_mem_ctl.scala 113:49]
  wire  _T_54 = ic_byp_hit_f & _T_319; // @[ifu_mem_ctl.scala 114:33]
  wire  _T_56 = ~_T_32; // @[ifu_mem_ctl.scala 114:57]
  wire  _T_57 = _T_54 & _T_56; // @[ifu_mem_ctl.scala 114:55]
  wire  ifu_bp_hit_taken_q_f = io_ifu_bp_hit_taken_f & io_ic_hit_f; // @[ifu_mem_ctl.scala 102:52]
  wire  _T_58 = ~ifu_bp_hit_taken_q_f; // @[ifu_mem_ctl.scala 114:91]
  wire  _T_59 = _T_57 & _T_58; // @[ifu_mem_ctl.scala 114:89]
  wire  _T_61 = _T_59 & _T_17; // @[ifu_mem_ctl.scala 114:113]
  wire  _T_64 = bus_ifu_wr_en_ff & _T_319; // @[ifu_mem_ctl.scala 115:39]
  wire  _T_67 = _T_64 & _T_56; // @[ifu_mem_ctl.scala 115:61]
  wire  _T_69 = _T_67 & _T_58; // @[ifu_mem_ctl.scala 115:95]
  wire  _T_71 = _T_69 & _T_17; // @[ifu_mem_ctl.scala 115:119]
  wire  _T_79 = _T_46 & _T_17; // @[ifu_mem_ctl.scala 116:100]
  wire  _T_81 = io_exu_flush_final | ifu_bp_hit_taken_q_f; // @[ifu_mem_ctl.scala 117:44]
  wire  _T_84 = _T_81 & _T_56; // @[ifu_mem_ctl.scala 117:68]
  wire [2:0] _T_86 = _T_84 ? 3'h2 : 3'h0; // @[ifu_mem_ctl.scala 117:22]
  wire [2:0] _T_87 = _T_79 ? 3'h0 : _T_86; // @[ifu_mem_ctl.scala 116:20]
  wire [2:0] _T_88 = _T_71 ? 3'h6 : _T_87; // @[ifu_mem_ctl.scala 115:20]
  wire [2:0] _T_89 = _T_61 ? 3'h6 : _T_88; // @[ifu_mem_ctl.scala 114:18]
  wire [2:0] _T_90 = _T_51 ? 3'h0 : _T_89; // @[ifu_mem_ctl.scala 113:16]
  wire [2:0] _T_91 = _T_47 ? 3'h4 : _T_90; // @[ifu_mem_ctl.scala 112:14]
  wire [2:0] _T_92 = _T_40 ? 3'h3 : _T_91; // @[ifu_mem_ctl.scala 111:12]
  wire [2:0] _T_93 = _T_36 ? 3'h0 : _T_92; // @[ifu_mem_ctl.scala 110:27]
  wire  _T_102 = 3'h4 == miss_state; // @[Conditional.scala 37:30]
  wire  _T_106 = 3'h6 == miss_state; // @[Conditional.scala 37:30]
  wire  _T_2280 = byp_fetch_index[4:1] == 4'hf; // @[ifu_mem_ctl.scala 374:60]
  wire  _T_2281 = _T_2280 & ifc_fetch_req_f; // @[ifu_mem_ctl.scala 374:94]
  wire  stream_eol_f = _T_2281 & stream_hit_f; // @[ifu_mem_ctl.scala 374:112]
  wire  _T_108 = _T_81 | stream_eol_f; // @[ifu_mem_ctl.scala 125:72]
  wire  _T_111 = _T_108 & _T_56; // @[ifu_mem_ctl.scala 125:87]
  wire  _T_113 = _T_111 & _T_2623; // @[ifu_mem_ctl.scala 125:122]
  wire [2:0] _T_115 = _T_113 ? 3'h2 : 3'h0; // @[ifu_mem_ctl.scala 125:27]
  wire  _T_121 = 3'h3 == miss_state; // @[Conditional.scala 37:30]
  wire  _T_124 = io_exu_flush_final & _T_56; // @[ifu_mem_ctl.scala 129:48]
  wire  _T_126 = _T_124 & _T_2623; // @[ifu_mem_ctl.scala 129:82]
  wire [2:0] _T_128 = _T_126 ? 3'h2 : 3'h0; // @[ifu_mem_ctl.scala 129:27]
  wire  _T_132 = 3'h2 == miss_state; // @[Conditional.scala 37:30]
  wire  _T_236 = io_ic_rd_hit == 2'h0; // @[ifu_mem_ctl.scala 190:28]
  wire  _T_237 = _T_236 | reset_all_tags; // @[ifu_mem_ctl.scala 190:42]
  wire  _T_238 = _T_237 & fetch_req_icache_f; // @[ifu_mem_ctl.scala 190:60]
  wire  _T_239 = miss_state == 3'h2; // @[ifu_mem_ctl.scala 190:94]
  wire  _T_240 = _T_238 & _T_239; // @[ifu_mem_ctl.scala 190:81]
  wire  _T_243 = imb_ff[30:5] != ifu_fetch_addr_int_f[30:5]; // @[ifu_mem_ctl.scala 191:39]
  wire  _T_244 = _T_240 & _T_243; // @[ifu_mem_ctl.scala 190:111]
  wire  _T_246 = _T_244 & _T_17; // @[ifu_mem_ctl.scala 191:91]
  reg  sel_mb_addr_ff; // @[ifu_mem_ctl.scala 245:51]
  wire  _T_247 = ~sel_mb_addr_ff; // @[ifu_mem_ctl.scala 191:116]
  wire  _T_248 = _T_246 & _T_247; // @[ifu_mem_ctl.scala 191:114]
  wire  ic_miss_under_miss_f = _T_248 & _T_209; // @[ifu_mem_ctl.scala 191:132]
  wire  _T_135 = ic_miss_under_miss_f & _T_56; // @[ifu_mem_ctl.scala 133:50]
  wire  _T_137 = _T_135 & _T_2623; // @[ifu_mem_ctl.scala 133:84]
  wire  _T_256 = _T_230 & _T_239; // @[ifu_mem_ctl.scala 192:85]
  wire  _T_259 = imb_ff[30:5] == ifu_fetch_addr_int_f[30:5]; // @[ifu_mem_ctl.scala 193:39]
  wire  _T_260 = _T_259 | uncacheable_miss_ff; // @[ifu_mem_ctl.scala 193:91]
  wire  ic_ignore_2nd_miss_f = _T_256 & _T_260; // @[ifu_mem_ctl.scala 192:117]
  wire  _T_141 = ic_ignore_2nd_miss_f & _T_56; // @[ifu_mem_ctl.scala 134:35]
  wire  _T_143 = _T_141 & _T_2623; // @[ifu_mem_ctl.scala 134:69]
  wire [2:0] _T_145 = _T_143 ? 3'h7 : 3'h0; // @[ifu_mem_ctl.scala 134:12]
  wire [2:0] _T_146 = _T_137 ? 3'h5 : _T_145; // @[ifu_mem_ctl.scala 133:27]
  wire  _T_151 = 3'h5 == miss_state; // @[Conditional.scala 37:30]
  wire [2:0] _T_154 = _T_32 ? 3'h0 : 3'h2; // @[ifu_mem_ctl.scala 139:12]
  wire [2:0] _T_155 = io_exu_flush_final ? _T_154 : 3'h1; // @[ifu_mem_ctl.scala 138:75]
  wire [2:0] _T_156 = io_dec_mem_ctrl_dec_tlu_force_halt ? 3'h0 : _T_155; // @[ifu_mem_ctl.scala 138:27]
  wire  _T_160 = 3'h7 == miss_state; // @[Conditional.scala 37:30]
  wire [2:0] _T_164 = io_exu_flush_final ? _T_154 : 3'h0; // @[ifu_mem_ctl.scala 143:75]
  wire [2:0] _T_165 = io_dec_mem_ctrl_dec_tlu_force_halt ? 3'h0 : _T_164; // @[ifu_mem_ctl.scala 143:27]
  wire [2:0] _GEN_0 = _T_160 ? _T_165 : 3'h0; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_2 = _T_151 ? _T_156 : _GEN_0; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_4 = _T_132 ? _T_146 : _GEN_2; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_6 = _T_121 ? _T_128 : _GEN_4; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_8 = _T_106 ? _T_115 : _GEN_6; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_10 = _T_102 ? 3'h0 : _GEN_8; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_12 = _T_31 ? _T_93 : _GEN_10; // @[Conditional.scala 39:67]
  wire [2:0] miss_nxtstate = _T_24 ? _T_28 : _GEN_12; // @[Conditional.scala 40:58]
  wire  _T_20 = miss_nxtstate == 3'h5; // @[ifu_mem_ctl.scala 100:73]
  wire  _T_21 = _T_19 | _T_20; // @[ifu_mem_ctl.scala 100:57]
  wire  _T_22 = _T_18 & _T_21; // @[ifu_mem_ctl.scala 100:26]
  wire  _T_30 = ic_act_miss_f & _T_2623; // @[ifu_mem_ctl.scala 107:38]
  wire  _T_94 = io_dec_mem_ctrl_dec_tlu_force_halt | io_exu_flush_final; // @[ifu_mem_ctl.scala 118:59]
  wire  _T_95 = _T_94 | ic_byp_hit_f; // @[ifu_mem_ctl.scala 118:80]
  wire  _T_96 = _T_95 | ifu_bp_hit_taken_q_f; // @[ifu_mem_ctl.scala 118:95]
  wire  _T_98 = _T_96 | _T_32; // @[ifu_mem_ctl.scala 118:118]
  wire  _T_100 = bus_ifu_wr_en_ff & _T_17; // @[ifu_mem_ctl.scala 118:171]
  wire  _T_101 = _T_98 | _T_100; // @[ifu_mem_ctl.scala 118:151]
  wire  _T_103 = io_exu_flush_final | flush_final_f; // @[ifu_mem_ctl.scala 122:43]
  wire  _T_104 = _T_103 | ic_byp_hit_f; // @[ifu_mem_ctl.scala 122:59]
  wire  _T_105 = _T_104 | io_dec_mem_ctrl_dec_tlu_force_halt; // @[ifu_mem_ctl.scala 122:74]
  wire  _T_119 = _T_108 | _T_32; // @[ifu_mem_ctl.scala 126:84]
  wire  _T_120 = _T_119 | io_dec_mem_ctrl_dec_tlu_force_halt; // @[ifu_mem_ctl.scala 126:118]
  wire  _T_130 = io_exu_flush_final | _T_32; // @[ifu_mem_ctl.scala 130:43]
  wire  _T_131 = _T_130 | io_dec_mem_ctrl_dec_tlu_force_halt; // @[ifu_mem_ctl.scala 130:76]
  wire  _T_148 = _T_32 | ic_miss_under_miss_f; // @[ifu_mem_ctl.scala 135:55]
  wire  _T_149 = _T_148 | ic_ignore_2nd_miss_f; // @[ifu_mem_ctl.scala 135:78]
  wire  _T_150 = _T_149 | io_dec_mem_ctrl_dec_tlu_force_halt; // @[ifu_mem_ctl.scala 135:101]
  wire  _T_158 = _T_32 | io_exu_flush_final; // @[ifu_mem_ctl.scala 140:55]
  wire  _T_159 = _T_158 | io_dec_mem_ctrl_dec_tlu_force_halt; // @[ifu_mem_ctl.scala 140:76]
  wire  _GEN_1 = _T_160 & _T_159; // @[Conditional.scala 39:67]
  wire  _GEN_3 = _T_151 ? _T_159 : _GEN_1; // @[Conditional.scala 39:67]
  wire  _GEN_5 = _T_132 ? _T_150 : _GEN_3; // @[Conditional.scala 39:67]
  wire  _GEN_7 = _T_121 ? _T_131 : _GEN_5; // @[Conditional.scala 39:67]
  wire  _GEN_9 = _T_106 ? _T_120 : _GEN_7; // @[Conditional.scala 39:67]
  wire  _GEN_11 = _T_102 ? _T_105 : _GEN_9; // @[Conditional.scala 39:67]
  wire  _GEN_13 = _T_31 ? _T_101 : _GEN_11; // @[Conditional.scala 39:67]
  wire  miss_state_en = _T_24 ? _T_30 : _GEN_13; // @[Conditional.scala 40:58]
  wire  _T_174 = ~flush_final_f; // @[ifu_mem_ctl.scala 160:95]
  wire  _T_175 = _T_2283 & _T_174; // @[ifu_mem_ctl.scala 160:93]
  wire  crit_wd_byp_ok_ff = _T_2284 | _T_175; // @[ifu_mem_ctl.scala 160:58]
  wire  _T_178 = miss_pending & _T_56; // @[ifu_mem_ctl.scala 161:36]
  wire  _T_180 = _T_2283 & io_exu_flush_final; // @[ifu_mem_ctl.scala 161:106]
  wire  _T_181 = ~_T_180; // @[ifu_mem_ctl.scala 161:72]
  wire  _T_182 = _T_178 & _T_181; // @[ifu_mem_ctl.scala 161:70]
  wire  _T_184 = _T_2283 & crit_byp_hit_f; // @[ifu_mem_ctl.scala 162:57]
  wire  _T_185 = ~_T_184; // @[ifu_mem_ctl.scala 162:23]
  wire  _T_186 = _T_182 & _T_185; // @[ifu_mem_ctl.scala 161:128]
  wire  _T_187 = _T_186 | ic_act_miss_f; // @[ifu_mem_ctl.scala 162:77]
  wire  _T_188 = miss_nxtstate == 3'h4; // @[ifu_mem_ctl.scala 163:36]
  wire  _T_189 = miss_pending & _T_188; // @[ifu_mem_ctl.scala 163:19]
  wire  sel_hold_imb = _T_187 | _T_189; // @[ifu_mem_ctl.scala 162:93]
  wire  _T_191 = _T_19 | ic_miss_under_miss_f; // @[ifu_mem_ctl.scala 165:57]
  wire  sel_hold_imb_scnd = _T_191 & _T_174; // @[ifu_mem_ctl.scala 165:81]
  reg  way_status_mb_scnd_ff; // @[ifu_mem_ctl.scala 173:64]
  reg [6:0] ifu_ic_rw_int_addr_ff; // @[ifu_mem_ctl.scala 669:14]
  wire  _T_4671 = ifu_ic_rw_int_addr_ff == 7'h0; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_0; // @[Reg.scala 27:20]
  wire  _T_4799 = _T_4671 & way_status_out_0; // @[Mux.scala 27:72]
  wire  _T_4672 = ifu_ic_rw_int_addr_ff == 7'h1; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_1; // @[Reg.scala 27:20]
  wire  _T_4800 = _T_4672 & way_status_out_1; // @[Mux.scala 27:72]
  wire  _T_4927 = _T_4799 | _T_4800; // @[Mux.scala 27:72]
  wire  _T_4673 = ifu_ic_rw_int_addr_ff == 7'h2; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_2; // @[Reg.scala 27:20]
  wire  _T_4801 = _T_4673 & way_status_out_2; // @[Mux.scala 27:72]
  wire  _T_4928 = _T_4927 | _T_4801; // @[Mux.scala 27:72]
  wire  _T_4674 = ifu_ic_rw_int_addr_ff == 7'h3; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_3; // @[Reg.scala 27:20]
  wire  _T_4802 = _T_4674 & way_status_out_3; // @[Mux.scala 27:72]
  wire  _T_4929 = _T_4928 | _T_4802; // @[Mux.scala 27:72]
  wire  _T_4675 = ifu_ic_rw_int_addr_ff == 7'h4; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_4; // @[Reg.scala 27:20]
  wire  _T_4803 = _T_4675 & way_status_out_4; // @[Mux.scala 27:72]
  wire  _T_4930 = _T_4929 | _T_4803; // @[Mux.scala 27:72]
  wire  _T_4676 = ifu_ic_rw_int_addr_ff == 7'h5; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_5; // @[Reg.scala 27:20]
  wire  _T_4804 = _T_4676 & way_status_out_5; // @[Mux.scala 27:72]
  wire  _T_4931 = _T_4930 | _T_4804; // @[Mux.scala 27:72]
  wire  _T_4677 = ifu_ic_rw_int_addr_ff == 7'h6; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_6; // @[Reg.scala 27:20]
  wire  _T_4805 = _T_4677 & way_status_out_6; // @[Mux.scala 27:72]
  wire  _T_4932 = _T_4931 | _T_4805; // @[Mux.scala 27:72]
  wire  _T_4678 = ifu_ic_rw_int_addr_ff == 7'h7; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_7; // @[Reg.scala 27:20]
  wire  _T_4806 = _T_4678 & way_status_out_7; // @[Mux.scala 27:72]
  wire  _T_4933 = _T_4932 | _T_4806; // @[Mux.scala 27:72]
  wire  _T_4679 = ifu_ic_rw_int_addr_ff == 7'h8; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_8; // @[Reg.scala 27:20]
  wire  _T_4807 = _T_4679 & way_status_out_8; // @[Mux.scala 27:72]
  wire  _T_4934 = _T_4933 | _T_4807; // @[Mux.scala 27:72]
  wire  _T_4680 = ifu_ic_rw_int_addr_ff == 7'h9; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_9; // @[Reg.scala 27:20]
  wire  _T_4808 = _T_4680 & way_status_out_9; // @[Mux.scala 27:72]
  wire  _T_4935 = _T_4934 | _T_4808; // @[Mux.scala 27:72]
  wire  _T_4681 = ifu_ic_rw_int_addr_ff == 7'ha; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_10; // @[Reg.scala 27:20]
  wire  _T_4809 = _T_4681 & way_status_out_10; // @[Mux.scala 27:72]
  wire  _T_4936 = _T_4935 | _T_4809; // @[Mux.scala 27:72]
  wire  _T_4682 = ifu_ic_rw_int_addr_ff == 7'hb; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_11; // @[Reg.scala 27:20]
  wire  _T_4810 = _T_4682 & way_status_out_11; // @[Mux.scala 27:72]
  wire  _T_4937 = _T_4936 | _T_4810; // @[Mux.scala 27:72]
  wire  _T_4683 = ifu_ic_rw_int_addr_ff == 7'hc; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_12; // @[Reg.scala 27:20]
  wire  _T_4811 = _T_4683 & way_status_out_12; // @[Mux.scala 27:72]
  wire  _T_4938 = _T_4937 | _T_4811; // @[Mux.scala 27:72]
  wire  _T_4684 = ifu_ic_rw_int_addr_ff == 7'hd; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_13; // @[Reg.scala 27:20]
  wire  _T_4812 = _T_4684 & way_status_out_13; // @[Mux.scala 27:72]
  wire  _T_4939 = _T_4938 | _T_4812; // @[Mux.scala 27:72]
  wire  _T_4685 = ifu_ic_rw_int_addr_ff == 7'he; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_14; // @[Reg.scala 27:20]
  wire  _T_4813 = _T_4685 & way_status_out_14; // @[Mux.scala 27:72]
  wire  _T_4940 = _T_4939 | _T_4813; // @[Mux.scala 27:72]
  wire  _T_4686 = ifu_ic_rw_int_addr_ff == 7'hf; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_15; // @[Reg.scala 27:20]
  wire  _T_4814 = _T_4686 & way_status_out_15; // @[Mux.scala 27:72]
  wire  _T_4941 = _T_4940 | _T_4814; // @[Mux.scala 27:72]
  wire  _T_4687 = ifu_ic_rw_int_addr_ff == 7'h10; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_16; // @[Reg.scala 27:20]
  wire  _T_4815 = _T_4687 & way_status_out_16; // @[Mux.scala 27:72]
  wire  _T_4942 = _T_4941 | _T_4815; // @[Mux.scala 27:72]
  wire  _T_4688 = ifu_ic_rw_int_addr_ff == 7'h11; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_17; // @[Reg.scala 27:20]
  wire  _T_4816 = _T_4688 & way_status_out_17; // @[Mux.scala 27:72]
  wire  _T_4943 = _T_4942 | _T_4816; // @[Mux.scala 27:72]
  wire  _T_4689 = ifu_ic_rw_int_addr_ff == 7'h12; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_18; // @[Reg.scala 27:20]
  wire  _T_4817 = _T_4689 & way_status_out_18; // @[Mux.scala 27:72]
  wire  _T_4944 = _T_4943 | _T_4817; // @[Mux.scala 27:72]
  wire  _T_4690 = ifu_ic_rw_int_addr_ff == 7'h13; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_19; // @[Reg.scala 27:20]
  wire  _T_4818 = _T_4690 & way_status_out_19; // @[Mux.scala 27:72]
  wire  _T_4945 = _T_4944 | _T_4818; // @[Mux.scala 27:72]
  wire  _T_4691 = ifu_ic_rw_int_addr_ff == 7'h14; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_20; // @[Reg.scala 27:20]
  wire  _T_4819 = _T_4691 & way_status_out_20; // @[Mux.scala 27:72]
  wire  _T_4946 = _T_4945 | _T_4819; // @[Mux.scala 27:72]
  wire  _T_4692 = ifu_ic_rw_int_addr_ff == 7'h15; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_21; // @[Reg.scala 27:20]
  wire  _T_4820 = _T_4692 & way_status_out_21; // @[Mux.scala 27:72]
  wire  _T_4947 = _T_4946 | _T_4820; // @[Mux.scala 27:72]
  wire  _T_4693 = ifu_ic_rw_int_addr_ff == 7'h16; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_22; // @[Reg.scala 27:20]
  wire  _T_4821 = _T_4693 & way_status_out_22; // @[Mux.scala 27:72]
  wire  _T_4948 = _T_4947 | _T_4821; // @[Mux.scala 27:72]
  wire  _T_4694 = ifu_ic_rw_int_addr_ff == 7'h17; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_23; // @[Reg.scala 27:20]
  wire  _T_4822 = _T_4694 & way_status_out_23; // @[Mux.scala 27:72]
  wire  _T_4949 = _T_4948 | _T_4822; // @[Mux.scala 27:72]
  wire  _T_4695 = ifu_ic_rw_int_addr_ff == 7'h18; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_24; // @[Reg.scala 27:20]
  wire  _T_4823 = _T_4695 & way_status_out_24; // @[Mux.scala 27:72]
  wire  _T_4950 = _T_4949 | _T_4823; // @[Mux.scala 27:72]
  wire  _T_4696 = ifu_ic_rw_int_addr_ff == 7'h19; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_25; // @[Reg.scala 27:20]
  wire  _T_4824 = _T_4696 & way_status_out_25; // @[Mux.scala 27:72]
  wire  _T_4951 = _T_4950 | _T_4824; // @[Mux.scala 27:72]
  wire  _T_4697 = ifu_ic_rw_int_addr_ff == 7'h1a; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_26; // @[Reg.scala 27:20]
  wire  _T_4825 = _T_4697 & way_status_out_26; // @[Mux.scala 27:72]
  wire  _T_4952 = _T_4951 | _T_4825; // @[Mux.scala 27:72]
  wire  _T_4698 = ifu_ic_rw_int_addr_ff == 7'h1b; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_27; // @[Reg.scala 27:20]
  wire  _T_4826 = _T_4698 & way_status_out_27; // @[Mux.scala 27:72]
  wire  _T_4953 = _T_4952 | _T_4826; // @[Mux.scala 27:72]
  wire  _T_4699 = ifu_ic_rw_int_addr_ff == 7'h1c; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_28; // @[Reg.scala 27:20]
  wire  _T_4827 = _T_4699 & way_status_out_28; // @[Mux.scala 27:72]
  wire  _T_4954 = _T_4953 | _T_4827; // @[Mux.scala 27:72]
  wire  _T_4700 = ifu_ic_rw_int_addr_ff == 7'h1d; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_29; // @[Reg.scala 27:20]
  wire  _T_4828 = _T_4700 & way_status_out_29; // @[Mux.scala 27:72]
  wire  _T_4955 = _T_4954 | _T_4828; // @[Mux.scala 27:72]
  wire  _T_4701 = ifu_ic_rw_int_addr_ff == 7'h1e; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_30; // @[Reg.scala 27:20]
  wire  _T_4829 = _T_4701 & way_status_out_30; // @[Mux.scala 27:72]
  wire  _T_4956 = _T_4955 | _T_4829; // @[Mux.scala 27:72]
  wire  _T_4702 = ifu_ic_rw_int_addr_ff == 7'h1f; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_31; // @[Reg.scala 27:20]
  wire  _T_4830 = _T_4702 & way_status_out_31; // @[Mux.scala 27:72]
  wire  _T_4957 = _T_4956 | _T_4830; // @[Mux.scala 27:72]
  wire  _T_4703 = ifu_ic_rw_int_addr_ff == 7'h20; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_32; // @[Reg.scala 27:20]
  wire  _T_4831 = _T_4703 & way_status_out_32; // @[Mux.scala 27:72]
  wire  _T_4958 = _T_4957 | _T_4831; // @[Mux.scala 27:72]
  wire  _T_4704 = ifu_ic_rw_int_addr_ff == 7'h21; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_33; // @[Reg.scala 27:20]
  wire  _T_4832 = _T_4704 & way_status_out_33; // @[Mux.scala 27:72]
  wire  _T_4959 = _T_4958 | _T_4832; // @[Mux.scala 27:72]
  wire  _T_4705 = ifu_ic_rw_int_addr_ff == 7'h22; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_34; // @[Reg.scala 27:20]
  wire  _T_4833 = _T_4705 & way_status_out_34; // @[Mux.scala 27:72]
  wire  _T_4960 = _T_4959 | _T_4833; // @[Mux.scala 27:72]
  wire  _T_4706 = ifu_ic_rw_int_addr_ff == 7'h23; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_35; // @[Reg.scala 27:20]
  wire  _T_4834 = _T_4706 & way_status_out_35; // @[Mux.scala 27:72]
  wire  _T_4961 = _T_4960 | _T_4834; // @[Mux.scala 27:72]
  wire  _T_4707 = ifu_ic_rw_int_addr_ff == 7'h24; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_36; // @[Reg.scala 27:20]
  wire  _T_4835 = _T_4707 & way_status_out_36; // @[Mux.scala 27:72]
  wire  _T_4962 = _T_4961 | _T_4835; // @[Mux.scala 27:72]
  wire  _T_4708 = ifu_ic_rw_int_addr_ff == 7'h25; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_37; // @[Reg.scala 27:20]
  wire  _T_4836 = _T_4708 & way_status_out_37; // @[Mux.scala 27:72]
  wire  _T_4963 = _T_4962 | _T_4836; // @[Mux.scala 27:72]
  wire  _T_4709 = ifu_ic_rw_int_addr_ff == 7'h26; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_38; // @[Reg.scala 27:20]
  wire  _T_4837 = _T_4709 & way_status_out_38; // @[Mux.scala 27:72]
  wire  _T_4964 = _T_4963 | _T_4837; // @[Mux.scala 27:72]
  wire  _T_4710 = ifu_ic_rw_int_addr_ff == 7'h27; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_39; // @[Reg.scala 27:20]
  wire  _T_4838 = _T_4710 & way_status_out_39; // @[Mux.scala 27:72]
  wire  _T_4965 = _T_4964 | _T_4838; // @[Mux.scala 27:72]
  wire  _T_4711 = ifu_ic_rw_int_addr_ff == 7'h28; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_40; // @[Reg.scala 27:20]
  wire  _T_4839 = _T_4711 & way_status_out_40; // @[Mux.scala 27:72]
  wire  _T_4966 = _T_4965 | _T_4839; // @[Mux.scala 27:72]
  wire  _T_4712 = ifu_ic_rw_int_addr_ff == 7'h29; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_41; // @[Reg.scala 27:20]
  wire  _T_4840 = _T_4712 & way_status_out_41; // @[Mux.scala 27:72]
  wire  _T_4967 = _T_4966 | _T_4840; // @[Mux.scala 27:72]
  wire  _T_4713 = ifu_ic_rw_int_addr_ff == 7'h2a; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_42; // @[Reg.scala 27:20]
  wire  _T_4841 = _T_4713 & way_status_out_42; // @[Mux.scala 27:72]
  wire  _T_4968 = _T_4967 | _T_4841; // @[Mux.scala 27:72]
  wire  _T_4714 = ifu_ic_rw_int_addr_ff == 7'h2b; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_43; // @[Reg.scala 27:20]
  wire  _T_4842 = _T_4714 & way_status_out_43; // @[Mux.scala 27:72]
  wire  _T_4969 = _T_4968 | _T_4842; // @[Mux.scala 27:72]
  wire  _T_4715 = ifu_ic_rw_int_addr_ff == 7'h2c; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_44; // @[Reg.scala 27:20]
  wire  _T_4843 = _T_4715 & way_status_out_44; // @[Mux.scala 27:72]
  wire  _T_4970 = _T_4969 | _T_4843; // @[Mux.scala 27:72]
  wire  _T_4716 = ifu_ic_rw_int_addr_ff == 7'h2d; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_45; // @[Reg.scala 27:20]
  wire  _T_4844 = _T_4716 & way_status_out_45; // @[Mux.scala 27:72]
  wire  _T_4971 = _T_4970 | _T_4844; // @[Mux.scala 27:72]
  wire  _T_4717 = ifu_ic_rw_int_addr_ff == 7'h2e; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_46; // @[Reg.scala 27:20]
  wire  _T_4845 = _T_4717 & way_status_out_46; // @[Mux.scala 27:72]
  wire  _T_4972 = _T_4971 | _T_4845; // @[Mux.scala 27:72]
  wire  _T_4718 = ifu_ic_rw_int_addr_ff == 7'h2f; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_47; // @[Reg.scala 27:20]
  wire  _T_4846 = _T_4718 & way_status_out_47; // @[Mux.scala 27:72]
  wire  _T_4973 = _T_4972 | _T_4846; // @[Mux.scala 27:72]
  wire  _T_4719 = ifu_ic_rw_int_addr_ff == 7'h30; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_48; // @[Reg.scala 27:20]
  wire  _T_4847 = _T_4719 & way_status_out_48; // @[Mux.scala 27:72]
  wire  _T_4974 = _T_4973 | _T_4847; // @[Mux.scala 27:72]
  wire  _T_4720 = ifu_ic_rw_int_addr_ff == 7'h31; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_49; // @[Reg.scala 27:20]
  wire  _T_4848 = _T_4720 & way_status_out_49; // @[Mux.scala 27:72]
  wire  _T_4975 = _T_4974 | _T_4848; // @[Mux.scala 27:72]
  wire  _T_4721 = ifu_ic_rw_int_addr_ff == 7'h32; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_50; // @[Reg.scala 27:20]
  wire  _T_4849 = _T_4721 & way_status_out_50; // @[Mux.scala 27:72]
  wire  _T_4976 = _T_4975 | _T_4849; // @[Mux.scala 27:72]
  wire  _T_4722 = ifu_ic_rw_int_addr_ff == 7'h33; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_51; // @[Reg.scala 27:20]
  wire  _T_4850 = _T_4722 & way_status_out_51; // @[Mux.scala 27:72]
  wire  _T_4977 = _T_4976 | _T_4850; // @[Mux.scala 27:72]
  wire  _T_4723 = ifu_ic_rw_int_addr_ff == 7'h34; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_52; // @[Reg.scala 27:20]
  wire  _T_4851 = _T_4723 & way_status_out_52; // @[Mux.scala 27:72]
  wire  _T_4978 = _T_4977 | _T_4851; // @[Mux.scala 27:72]
  wire  _T_4724 = ifu_ic_rw_int_addr_ff == 7'h35; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_53; // @[Reg.scala 27:20]
  wire  _T_4852 = _T_4724 & way_status_out_53; // @[Mux.scala 27:72]
  wire  _T_4979 = _T_4978 | _T_4852; // @[Mux.scala 27:72]
  wire  _T_4725 = ifu_ic_rw_int_addr_ff == 7'h36; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_54; // @[Reg.scala 27:20]
  wire  _T_4853 = _T_4725 & way_status_out_54; // @[Mux.scala 27:72]
  wire  _T_4980 = _T_4979 | _T_4853; // @[Mux.scala 27:72]
  wire  _T_4726 = ifu_ic_rw_int_addr_ff == 7'h37; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_55; // @[Reg.scala 27:20]
  wire  _T_4854 = _T_4726 & way_status_out_55; // @[Mux.scala 27:72]
  wire  _T_4981 = _T_4980 | _T_4854; // @[Mux.scala 27:72]
  wire  _T_4727 = ifu_ic_rw_int_addr_ff == 7'h38; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_56; // @[Reg.scala 27:20]
  wire  _T_4855 = _T_4727 & way_status_out_56; // @[Mux.scala 27:72]
  wire  _T_4982 = _T_4981 | _T_4855; // @[Mux.scala 27:72]
  wire  _T_4728 = ifu_ic_rw_int_addr_ff == 7'h39; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_57; // @[Reg.scala 27:20]
  wire  _T_4856 = _T_4728 & way_status_out_57; // @[Mux.scala 27:72]
  wire  _T_4983 = _T_4982 | _T_4856; // @[Mux.scala 27:72]
  wire  _T_4729 = ifu_ic_rw_int_addr_ff == 7'h3a; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_58; // @[Reg.scala 27:20]
  wire  _T_4857 = _T_4729 & way_status_out_58; // @[Mux.scala 27:72]
  wire  _T_4984 = _T_4983 | _T_4857; // @[Mux.scala 27:72]
  wire  _T_4730 = ifu_ic_rw_int_addr_ff == 7'h3b; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_59; // @[Reg.scala 27:20]
  wire  _T_4858 = _T_4730 & way_status_out_59; // @[Mux.scala 27:72]
  wire  _T_4985 = _T_4984 | _T_4858; // @[Mux.scala 27:72]
  wire  _T_4731 = ifu_ic_rw_int_addr_ff == 7'h3c; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_60; // @[Reg.scala 27:20]
  wire  _T_4859 = _T_4731 & way_status_out_60; // @[Mux.scala 27:72]
  wire  _T_4986 = _T_4985 | _T_4859; // @[Mux.scala 27:72]
  wire  _T_4732 = ifu_ic_rw_int_addr_ff == 7'h3d; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_61; // @[Reg.scala 27:20]
  wire  _T_4860 = _T_4732 & way_status_out_61; // @[Mux.scala 27:72]
  wire  _T_4987 = _T_4986 | _T_4860; // @[Mux.scala 27:72]
  wire  _T_4733 = ifu_ic_rw_int_addr_ff == 7'h3e; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_62; // @[Reg.scala 27:20]
  wire  _T_4861 = _T_4733 & way_status_out_62; // @[Mux.scala 27:72]
  wire  _T_4988 = _T_4987 | _T_4861; // @[Mux.scala 27:72]
  wire  _T_4734 = ifu_ic_rw_int_addr_ff == 7'h3f; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_63; // @[Reg.scala 27:20]
  wire  _T_4862 = _T_4734 & way_status_out_63; // @[Mux.scala 27:72]
  wire  _T_4989 = _T_4988 | _T_4862; // @[Mux.scala 27:72]
  wire  _T_4735 = ifu_ic_rw_int_addr_ff == 7'h40; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_64; // @[Reg.scala 27:20]
  wire  _T_4863 = _T_4735 & way_status_out_64; // @[Mux.scala 27:72]
  wire  _T_4990 = _T_4989 | _T_4863; // @[Mux.scala 27:72]
  wire  _T_4736 = ifu_ic_rw_int_addr_ff == 7'h41; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_65; // @[Reg.scala 27:20]
  wire  _T_4864 = _T_4736 & way_status_out_65; // @[Mux.scala 27:72]
  wire  _T_4991 = _T_4990 | _T_4864; // @[Mux.scala 27:72]
  wire  _T_4737 = ifu_ic_rw_int_addr_ff == 7'h42; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_66; // @[Reg.scala 27:20]
  wire  _T_4865 = _T_4737 & way_status_out_66; // @[Mux.scala 27:72]
  wire  _T_4992 = _T_4991 | _T_4865; // @[Mux.scala 27:72]
  wire  _T_4738 = ifu_ic_rw_int_addr_ff == 7'h43; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_67; // @[Reg.scala 27:20]
  wire  _T_4866 = _T_4738 & way_status_out_67; // @[Mux.scala 27:72]
  wire  _T_4993 = _T_4992 | _T_4866; // @[Mux.scala 27:72]
  wire  _T_4739 = ifu_ic_rw_int_addr_ff == 7'h44; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_68; // @[Reg.scala 27:20]
  wire  _T_4867 = _T_4739 & way_status_out_68; // @[Mux.scala 27:72]
  wire  _T_4994 = _T_4993 | _T_4867; // @[Mux.scala 27:72]
  wire  _T_4740 = ifu_ic_rw_int_addr_ff == 7'h45; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_69; // @[Reg.scala 27:20]
  wire  _T_4868 = _T_4740 & way_status_out_69; // @[Mux.scala 27:72]
  wire  _T_4995 = _T_4994 | _T_4868; // @[Mux.scala 27:72]
  wire  _T_4741 = ifu_ic_rw_int_addr_ff == 7'h46; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_70; // @[Reg.scala 27:20]
  wire  _T_4869 = _T_4741 & way_status_out_70; // @[Mux.scala 27:72]
  wire  _T_4996 = _T_4995 | _T_4869; // @[Mux.scala 27:72]
  wire  _T_4742 = ifu_ic_rw_int_addr_ff == 7'h47; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_71; // @[Reg.scala 27:20]
  wire  _T_4870 = _T_4742 & way_status_out_71; // @[Mux.scala 27:72]
  wire  _T_4997 = _T_4996 | _T_4870; // @[Mux.scala 27:72]
  wire  _T_4743 = ifu_ic_rw_int_addr_ff == 7'h48; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_72; // @[Reg.scala 27:20]
  wire  _T_4871 = _T_4743 & way_status_out_72; // @[Mux.scala 27:72]
  wire  _T_4998 = _T_4997 | _T_4871; // @[Mux.scala 27:72]
  wire  _T_4744 = ifu_ic_rw_int_addr_ff == 7'h49; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_73; // @[Reg.scala 27:20]
  wire  _T_4872 = _T_4744 & way_status_out_73; // @[Mux.scala 27:72]
  wire  _T_4999 = _T_4998 | _T_4872; // @[Mux.scala 27:72]
  wire  _T_4745 = ifu_ic_rw_int_addr_ff == 7'h4a; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_74; // @[Reg.scala 27:20]
  wire  _T_4873 = _T_4745 & way_status_out_74; // @[Mux.scala 27:72]
  wire  _T_5000 = _T_4999 | _T_4873; // @[Mux.scala 27:72]
  wire  _T_4746 = ifu_ic_rw_int_addr_ff == 7'h4b; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_75; // @[Reg.scala 27:20]
  wire  _T_4874 = _T_4746 & way_status_out_75; // @[Mux.scala 27:72]
  wire  _T_5001 = _T_5000 | _T_4874; // @[Mux.scala 27:72]
  wire  _T_4747 = ifu_ic_rw_int_addr_ff == 7'h4c; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_76; // @[Reg.scala 27:20]
  wire  _T_4875 = _T_4747 & way_status_out_76; // @[Mux.scala 27:72]
  wire  _T_5002 = _T_5001 | _T_4875; // @[Mux.scala 27:72]
  wire  _T_4748 = ifu_ic_rw_int_addr_ff == 7'h4d; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_77; // @[Reg.scala 27:20]
  wire  _T_4876 = _T_4748 & way_status_out_77; // @[Mux.scala 27:72]
  wire  _T_5003 = _T_5002 | _T_4876; // @[Mux.scala 27:72]
  wire  _T_4749 = ifu_ic_rw_int_addr_ff == 7'h4e; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_78; // @[Reg.scala 27:20]
  wire  _T_4877 = _T_4749 & way_status_out_78; // @[Mux.scala 27:72]
  wire  _T_5004 = _T_5003 | _T_4877; // @[Mux.scala 27:72]
  wire  _T_4750 = ifu_ic_rw_int_addr_ff == 7'h4f; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_79; // @[Reg.scala 27:20]
  wire  _T_4878 = _T_4750 & way_status_out_79; // @[Mux.scala 27:72]
  wire  _T_5005 = _T_5004 | _T_4878; // @[Mux.scala 27:72]
  wire  _T_4751 = ifu_ic_rw_int_addr_ff == 7'h50; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_80; // @[Reg.scala 27:20]
  wire  _T_4879 = _T_4751 & way_status_out_80; // @[Mux.scala 27:72]
  wire  _T_5006 = _T_5005 | _T_4879; // @[Mux.scala 27:72]
  wire  _T_4752 = ifu_ic_rw_int_addr_ff == 7'h51; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_81; // @[Reg.scala 27:20]
  wire  _T_4880 = _T_4752 & way_status_out_81; // @[Mux.scala 27:72]
  wire  _T_5007 = _T_5006 | _T_4880; // @[Mux.scala 27:72]
  wire  _T_4753 = ifu_ic_rw_int_addr_ff == 7'h52; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_82; // @[Reg.scala 27:20]
  wire  _T_4881 = _T_4753 & way_status_out_82; // @[Mux.scala 27:72]
  wire  _T_5008 = _T_5007 | _T_4881; // @[Mux.scala 27:72]
  wire  _T_4754 = ifu_ic_rw_int_addr_ff == 7'h53; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_83; // @[Reg.scala 27:20]
  wire  _T_4882 = _T_4754 & way_status_out_83; // @[Mux.scala 27:72]
  wire  _T_5009 = _T_5008 | _T_4882; // @[Mux.scala 27:72]
  wire  _T_4755 = ifu_ic_rw_int_addr_ff == 7'h54; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_84; // @[Reg.scala 27:20]
  wire  _T_4883 = _T_4755 & way_status_out_84; // @[Mux.scala 27:72]
  wire  _T_5010 = _T_5009 | _T_4883; // @[Mux.scala 27:72]
  wire  _T_4756 = ifu_ic_rw_int_addr_ff == 7'h55; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_85; // @[Reg.scala 27:20]
  wire  _T_4884 = _T_4756 & way_status_out_85; // @[Mux.scala 27:72]
  wire  _T_5011 = _T_5010 | _T_4884; // @[Mux.scala 27:72]
  wire  _T_4757 = ifu_ic_rw_int_addr_ff == 7'h56; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_86; // @[Reg.scala 27:20]
  wire  _T_4885 = _T_4757 & way_status_out_86; // @[Mux.scala 27:72]
  wire  _T_5012 = _T_5011 | _T_4885; // @[Mux.scala 27:72]
  wire  _T_4758 = ifu_ic_rw_int_addr_ff == 7'h57; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_87; // @[Reg.scala 27:20]
  wire  _T_4886 = _T_4758 & way_status_out_87; // @[Mux.scala 27:72]
  wire  _T_5013 = _T_5012 | _T_4886; // @[Mux.scala 27:72]
  wire  _T_4759 = ifu_ic_rw_int_addr_ff == 7'h58; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_88; // @[Reg.scala 27:20]
  wire  _T_4887 = _T_4759 & way_status_out_88; // @[Mux.scala 27:72]
  wire  _T_5014 = _T_5013 | _T_4887; // @[Mux.scala 27:72]
  wire  _T_4760 = ifu_ic_rw_int_addr_ff == 7'h59; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_89; // @[Reg.scala 27:20]
  wire  _T_4888 = _T_4760 & way_status_out_89; // @[Mux.scala 27:72]
  wire  _T_5015 = _T_5014 | _T_4888; // @[Mux.scala 27:72]
  wire  _T_4761 = ifu_ic_rw_int_addr_ff == 7'h5a; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_90; // @[Reg.scala 27:20]
  wire  _T_4889 = _T_4761 & way_status_out_90; // @[Mux.scala 27:72]
  wire  _T_5016 = _T_5015 | _T_4889; // @[Mux.scala 27:72]
  wire  _T_4762 = ifu_ic_rw_int_addr_ff == 7'h5b; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_91; // @[Reg.scala 27:20]
  wire  _T_4890 = _T_4762 & way_status_out_91; // @[Mux.scala 27:72]
  wire  _T_5017 = _T_5016 | _T_4890; // @[Mux.scala 27:72]
  wire  _T_4763 = ifu_ic_rw_int_addr_ff == 7'h5c; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_92; // @[Reg.scala 27:20]
  wire  _T_4891 = _T_4763 & way_status_out_92; // @[Mux.scala 27:72]
  wire  _T_5018 = _T_5017 | _T_4891; // @[Mux.scala 27:72]
  wire  _T_4764 = ifu_ic_rw_int_addr_ff == 7'h5d; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_93; // @[Reg.scala 27:20]
  wire  _T_4892 = _T_4764 & way_status_out_93; // @[Mux.scala 27:72]
  wire  _T_5019 = _T_5018 | _T_4892; // @[Mux.scala 27:72]
  wire  _T_4765 = ifu_ic_rw_int_addr_ff == 7'h5e; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_94; // @[Reg.scala 27:20]
  wire  _T_4893 = _T_4765 & way_status_out_94; // @[Mux.scala 27:72]
  wire  _T_5020 = _T_5019 | _T_4893; // @[Mux.scala 27:72]
  wire  _T_4766 = ifu_ic_rw_int_addr_ff == 7'h5f; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_95; // @[Reg.scala 27:20]
  wire  _T_4894 = _T_4766 & way_status_out_95; // @[Mux.scala 27:72]
  wire  _T_5021 = _T_5020 | _T_4894; // @[Mux.scala 27:72]
  wire  _T_4767 = ifu_ic_rw_int_addr_ff == 7'h60; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_96; // @[Reg.scala 27:20]
  wire  _T_4895 = _T_4767 & way_status_out_96; // @[Mux.scala 27:72]
  wire  _T_5022 = _T_5021 | _T_4895; // @[Mux.scala 27:72]
  wire  _T_4768 = ifu_ic_rw_int_addr_ff == 7'h61; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_97; // @[Reg.scala 27:20]
  wire  _T_4896 = _T_4768 & way_status_out_97; // @[Mux.scala 27:72]
  wire  _T_5023 = _T_5022 | _T_4896; // @[Mux.scala 27:72]
  wire  _T_4769 = ifu_ic_rw_int_addr_ff == 7'h62; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_98; // @[Reg.scala 27:20]
  wire  _T_4897 = _T_4769 & way_status_out_98; // @[Mux.scala 27:72]
  wire  _T_5024 = _T_5023 | _T_4897; // @[Mux.scala 27:72]
  wire  _T_4770 = ifu_ic_rw_int_addr_ff == 7'h63; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_99; // @[Reg.scala 27:20]
  wire  _T_4898 = _T_4770 & way_status_out_99; // @[Mux.scala 27:72]
  wire  _T_5025 = _T_5024 | _T_4898; // @[Mux.scala 27:72]
  wire  _T_4771 = ifu_ic_rw_int_addr_ff == 7'h64; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_100; // @[Reg.scala 27:20]
  wire  _T_4899 = _T_4771 & way_status_out_100; // @[Mux.scala 27:72]
  wire  _T_5026 = _T_5025 | _T_4899; // @[Mux.scala 27:72]
  wire  _T_4772 = ifu_ic_rw_int_addr_ff == 7'h65; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_101; // @[Reg.scala 27:20]
  wire  _T_4900 = _T_4772 & way_status_out_101; // @[Mux.scala 27:72]
  wire  _T_5027 = _T_5026 | _T_4900; // @[Mux.scala 27:72]
  wire  _T_4773 = ifu_ic_rw_int_addr_ff == 7'h66; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_102; // @[Reg.scala 27:20]
  wire  _T_4901 = _T_4773 & way_status_out_102; // @[Mux.scala 27:72]
  wire  _T_5028 = _T_5027 | _T_4901; // @[Mux.scala 27:72]
  wire  _T_4774 = ifu_ic_rw_int_addr_ff == 7'h67; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_103; // @[Reg.scala 27:20]
  wire  _T_4902 = _T_4774 & way_status_out_103; // @[Mux.scala 27:72]
  wire  _T_5029 = _T_5028 | _T_4902; // @[Mux.scala 27:72]
  wire  _T_4775 = ifu_ic_rw_int_addr_ff == 7'h68; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_104; // @[Reg.scala 27:20]
  wire  _T_4903 = _T_4775 & way_status_out_104; // @[Mux.scala 27:72]
  wire  _T_5030 = _T_5029 | _T_4903; // @[Mux.scala 27:72]
  wire  _T_4776 = ifu_ic_rw_int_addr_ff == 7'h69; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_105; // @[Reg.scala 27:20]
  wire  _T_4904 = _T_4776 & way_status_out_105; // @[Mux.scala 27:72]
  wire  _T_5031 = _T_5030 | _T_4904; // @[Mux.scala 27:72]
  wire  _T_4777 = ifu_ic_rw_int_addr_ff == 7'h6a; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_106; // @[Reg.scala 27:20]
  wire  _T_4905 = _T_4777 & way_status_out_106; // @[Mux.scala 27:72]
  wire  _T_5032 = _T_5031 | _T_4905; // @[Mux.scala 27:72]
  wire  _T_4778 = ifu_ic_rw_int_addr_ff == 7'h6b; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_107; // @[Reg.scala 27:20]
  wire  _T_4906 = _T_4778 & way_status_out_107; // @[Mux.scala 27:72]
  wire  _T_5033 = _T_5032 | _T_4906; // @[Mux.scala 27:72]
  wire  _T_4779 = ifu_ic_rw_int_addr_ff == 7'h6c; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_108; // @[Reg.scala 27:20]
  wire  _T_4907 = _T_4779 & way_status_out_108; // @[Mux.scala 27:72]
  wire  _T_5034 = _T_5033 | _T_4907; // @[Mux.scala 27:72]
  wire  _T_4780 = ifu_ic_rw_int_addr_ff == 7'h6d; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_109; // @[Reg.scala 27:20]
  wire  _T_4908 = _T_4780 & way_status_out_109; // @[Mux.scala 27:72]
  wire  _T_5035 = _T_5034 | _T_4908; // @[Mux.scala 27:72]
  wire  _T_4781 = ifu_ic_rw_int_addr_ff == 7'h6e; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_110; // @[Reg.scala 27:20]
  wire  _T_4909 = _T_4781 & way_status_out_110; // @[Mux.scala 27:72]
  wire  _T_5036 = _T_5035 | _T_4909; // @[Mux.scala 27:72]
  wire  _T_4782 = ifu_ic_rw_int_addr_ff == 7'h6f; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_111; // @[Reg.scala 27:20]
  wire  _T_4910 = _T_4782 & way_status_out_111; // @[Mux.scala 27:72]
  wire  _T_5037 = _T_5036 | _T_4910; // @[Mux.scala 27:72]
  wire  _T_4783 = ifu_ic_rw_int_addr_ff == 7'h70; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_112; // @[Reg.scala 27:20]
  wire  _T_4911 = _T_4783 & way_status_out_112; // @[Mux.scala 27:72]
  wire  _T_5038 = _T_5037 | _T_4911; // @[Mux.scala 27:72]
  wire  _T_4784 = ifu_ic_rw_int_addr_ff == 7'h71; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_113; // @[Reg.scala 27:20]
  wire  _T_4912 = _T_4784 & way_status_out_113; // @[Mux.scala 27:72]
  wire  _T_5039 = _T_5038 | _T_4912; // @[Mux.scala 27:72]
  wire  _T_4785 = ifu_ic_rw_int_addr_ff == 7'h72; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_114; // @[Reg.scala 27:20]
  wire  _T_4913 = _T_4785 & way_status_out_114; // @[Mux.scala 27:72]
  wire  _T_5040 = _T_5039 | _T_4913; // @[Mux.scala 27:72]
  wire  _T_4786 = ifu_ic_rw_int_addr_ff == 7'h73; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_115; // @[Reg.scala 27:20]
  wire  _T_4914 = _T_4786 & way_status_out_115; // @[Mux.scala 27:72]
  wire  _T_5041 = _T_5040 | _T_4914; // @[Mux.scala 27:72]
  wire  _T_4787 = ifu_ic_rw_int_addr_ff == 7'h74; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_116; // @[Reg.scala 27:20]
  wire  _T_4915 = _T_4787 & way_status_out_116; // @[Mux.scala 27:72]
  wire  _T_5042 = _T_5041 | _T_4915; // @[Mux.scala 27:72]
  wire  _T_4788 = ifu_ic_rw_int_addr_ff == 7'h75; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_117; // @[Reg.scala 27:20]
  wire  _T_4916 = _T_4788 & way_status_out_117; // @[Mux.scala 27:72]
  wire  _T_5043 = _T_5042 | _T_4916; // @[Mux.scala 27:72]
  wire  _T_4789 = ifu_ic_rw_int_addr_ff == 7'h76; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_118; // @[Reg.scala 27:20]
  wire  _T_4917 = _T_4789 & way_status_out_118; // @[Mux.scala 27:72]
  wire  _T_5044 = _T_5043 | _T_4917; // @[Mux.scala 27:72]
  wire  _T_4790 = ifu_ic_rw_int_addr_ff == 7'h77; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_119; // @[Reg.scala 27:20]
  wire  _T_4918 = _T_4790 & way_status_out_119; // @[Mux.scala 27:72]
  wire  _T_5045 = _T_5044 | _T_4918; // @[Mux.scala 27:72]
  wire  _T_4791 = ifu_ic_rw_int_addr_ff == 7'h78; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_120; // @[Reg.scala 27:20]
  wire  _T_4919 = _T_4791 & way_status_out_120; // @[Mux.scala 27:72]
  wire  _T_5046 = _T_5045 | _T_4919; // @[Mux.scala 27:72]
  wire  _T_4792 = ifu_ic_rw_int_addr_ff == 7'h79; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_121; // @[Reg.scala 27:20]
  wire  _T_4920 = _T_4792 & way_status_out_121; // @[Mux.scala 27:72]
  wire  _T_5047 = _T_5046 | _T_4920; // @[Mux.scala 27:72]
  wire  _T_4793 = ifu_ic_rw_int_addr_ff == 7'h7a; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_122; // @[Reg.scala 27:20]
  wire  _T_4921 = _T_4793 & way_status_out_122; // @[Mux.scala 27:72]
  wire  _T_5048 = _T_5047 | _T_4921; // @[Mux.scala 27:72]
  wire  _T_4794 = ifu_ic_rw_int_addr_ff == 7'h7b; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_123; // @[Reg.scala 27:20]
  wire  _T_4922 = _T_4794 & way_status_out_123; // @[Mux.scala 27:72]
  wire  _T_5049 = _T_5048 | _T_4922; // @[Mux.scala 27:72]
  wire  _T_4795 = ifu_ic_rw_int_addr_ff == 7'h7c; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_124; // @[Reg.scala 27:20]
  wire  _T_4923 = _T_4795 & way_status_out_124; // @[Mux.scala 27:72]
  wire  _T_5050 = _T_5049 | _T_4923; // @[Mux.scala 27:72]
  wire  _T_4796 = ifu_ic_rw_int_addr_ff == 7'h7d; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_125; // @[Reg.scala 27:20]
  wire  _T_4924 = _T_4796 & way_status_out_125; // @[Mux.scala 27:72]
  wire  _T_5051 = _T_5050 | _T_4924; // @[Mux.scala 27:72]
  wire  _T_4797 = ifu_ic_rw_int_addr_ff == 7'h7e; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_126; // @[Reg.scala 27:20]
  wire  _T_4925 = _T_4797 & way_status_out_126; // @[Mux.scala 27:72]
  wire  _T_5052 = _T_5051 | _T_4925; // @[Mux.scala 27:72]
  wire  _T_4798 = ifu_ic_rw_int_addr_ff == 7'h7f; // @[ifu_mem_ctl.scala 665:80]
  reg  way_status_out_127; // @[Reg.scala 27:20]
  wire  _T_4926 = _T_4798 & way_status_out_127; // @[Mux.scala 27:72]
  wire  way_status = _T_5052 | _T_4926; // @[Mux.scala 27:72]
  wire  _T_195 = ~reset_all_tags; // @[ifu_mem_ctl.scala 168:96]
  wire [1:0] _T_197 = _T_195 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [1:0] _T_198 = _T_197 & io_ic_tag_valid; // @[ifu_mem_ctl.scala 168:113]
  reg [1:0] tagv_mb_scnd_ff; // @[ifu_mem_ctl.scala 174:58]
  reg  uncacheable_miss_scnd_ff; // @[ifu_mem_ctl.scala 170:67]
  reg [30:0] imb_scnd_ff; // @[ifu_mem_ctl.scala 172:54]
  wire [2:0] _T_206 = bus_ifu_wr_en_ff ? 3'h7 : 3'h0; // @[Bitwise.scala 72:12]
  reg [2:0] ifu_bus_rid_ff; // @[ifu_mem_ctl.scala 514:46]
  wire [2:0] ic_wr_addr_bits_hi_3 = ifu_bus_rid_ff & _T_206; // @[ifu_mem_ctl.scala 177:45]
  wire  _T_212 = _T_231 | _T_239; // @[ifu_mem_ctl.scala 182:59]
  wire  _T_214 = _T_212 | _T_2268; // @[ifu_mem_ctl.scala 182:91]
  wire  ic_iccm_hit_f = fetch_req_iccm_f & _T_214; // @[ifu_mem_ctl.scala 182:41]
  wire  _T_219 = _T_227 & fetch_req_icache_f; // @[ifu_mem_ctl.scala 188:39]
  wire  _T_221 = _T_219 & _T_195; // @[ifu_mem_ctl.scala 188:60]
  wire  _T_225 = _T_221 & _T_212; // @[ifu_mem_ctl.scala 188:78]
  wire  ic_act_hit_f = _T_225 & _T_247; // @[ifu_mem_ctl.scala 188:126]
  wire  _T_262 = ic_act_hit_f | ic_byp_hit_f; // @[ifu_mem_ctl.scala 195:31]
  wire  _T_263 = _T_262 | ic_iccm_hit_f; // @[ifu_mem_ctl.scala 195:46]
  wire  _T_264 = ifc_region_acc_fault_final_f & ifc_fetch_req_f; // @[ifu_mem_ctl.scala 195:94]
  wire  _T_268 = sel_hold_imb ? uncacheable_miss_ff : io_ifc_fetch_uncacheable_bf; // @[ifu_mem_ctl.scala 196:84]
  wire  uncacheable_miss_in = scnd_miss_req ? uncacheable_miss_scnd_ff : _T_268; // @[ifu_mem_ctl.scala 196:32]
  wire  _T_274 = imb_ff[11:5] == imb_scnd_ff[11:5]; // @[ifu_mem_ctl.scala 199:79]
  wire  _T_275 = _T_274 & scnd_miss_req; // @[ifu_mem_ctl.scala 199:135]
  reg [1:0] ifu_bus_rresp_ff; // @[ifu_mem_ctl.scala 512:51]
  wire  _T_2693 = |ifu_bus_rresp_ff; // @[ifu_mem_ctl.scala 558:48]
  wire  _T_2694 = _T_2693 & ifu_bus_rvalid_ff; // @[ifu_mem_ctl.scala 558:52]
  wire  bus_ifu_wr_data_error_ff = _T_2694 & miss_pending; // @[ifu_mem_ctl.scala 558:73]
  reg  ifu_wr_data_comb_err_ff; // @[ifu_mem_ctl.scala 276:61]
  wire  ifu_wr_cumulative_err_data = bus_ifu_wr_data_error_ff | ifu_wr_data_comb_err_ff; // @[ifu_mem_ctl.scala 275:55]
  wire  _T_276 = ~ifu_wr_cumulative_err_data; // @[ifu_mem_ctl.scala 199:153]
  wire  scnd_miss_index_match = _T_275 & _T_276; // @[ifu_mem_ctl.scala 199:151]
  wire  _T_277 = ~scnd_miss_index_match; // @[ifu_mem_ctl.scala 202:47]
  wire  _T_278 = scnd_miss_req & _T_277; // @[ifu_mem_ctl.scala 202:45]
  wire  _T_280 = scnd_miss_req & scnd_miss_index_match; // @[ifu_mem_ctl.scala 203:26]
  reg  way_status_mb_ff; // @[ifu_mem_ctl.scala 223:59]
  wire  _T_9756 = ~way_status_mb_ff; // @[ifu_mem_ctl.scala 720:33]
  reg [1:0] tagv_mb_ff; // @[ifu_mem_ctl.scala 224:53]
  wire  _T_9758 = _T_9756 & tagv_mb_ff[0]; // @[ifu_mem_ctl.scala 720:51]
  wire  _T_9760 = _T_9758 & tagv_mb_ff[1]; // @[ifu_mem_ctl.scala 720:67]
  wire  _T_9762 = ~tagv_mb_ff[0]; // @[ifu_mem_ctl.scala 720:86]
  wire  replace_way_mb_any_0 = _T_9760 | _T_9762; // @[ifu_mem_ctl.scala 720:84]
  wire [1:0] _T_287 = scnd_miss_index_match ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire  _T_9765 = way_status_mb_ff & tagv_mb_ff[0]; // @[ifu_mem_ctl.scala 721:50]
  wire  _T_9767 = _T_9765 & tagv_mb_ff[1]; // @[ifu_mem_ctl.scala 721:66]
  wire  _T_9769 = ~tagv_mb_ff[1]; // @[ifu_mem_ctl.scala 721:85]
  wire  _T_9771 = _T_9769 & tagv_mb_ff[0]; // @[ifu_mem_ctl.scala 721:100]
  wire  replace_way_mb_any_1 = _T_9767 | _T_9771; // @[ifu_mem_ctl.scala 721:83]
  wire [1:0] _T_288 = {replace_way_mb_any_1,replace_way_mb_any_0}; // @[Cat.scala 29:58]
  wire [1:0] _T_289 = _T_287 & _T_288; // @[ifu_mem_ctl.scala 207:110]
  wire [1:0] _T_290 = tagv_mb_scnd_ff | _T_289; // @[ifu_mem_ctl.scala 207:62]
  wire [1:0] _T_295 = io_ic_tag_valid & _T_197; // @[ifu_mem_ctl.scala 208:56]
  wire  _T_297 = ~scnd_miss_req_q; // @[ifu_mem_ctl.scala 211:36]
  wire  _T_298 = miss_pending & _T_297; // @[ifu_mem_ctl.scala 211:34]
  reg  reset_ic_ff; // @[ifu_mem_ctl.scala 212:48]
  wire  _T_299 = reset_all_tags | reset_ic_ff; // @[ifu_mem_ctl.scala 211:72]
  wire  reset_ic_in = _T_298 & _T_299; // @[ifu_mem_ctl.scala 211:53]
  reg  fetch_uncacheable_ff; // @[ifu_mem_ctl.scala 213:62]
  reg [25:0] miss_addr; // @[ifu_mem_ctl.scala 222:48]
  wire  _T_309 = io_ifu_bus_clk_en | ic_act_miss_f; // @[ifu_mem_ctl.scala 221:57]
  wire  _T_315 = _T_2283 & flush_final_f; // @[ifu_mem_ctl.scala 226:87]
  wire  _T_316 = ~_T_315; // @[ifu_mem_ctl.scala 226:55]
  wire  _T_317 = io_ifc_fetch_req_bf & _T_316; // @[ifu_mem_ctl.scala 226:53]
  wire  _T_2275 = ~_T_2270; // @[ifu_mem_ctl.scala 373:46]
  wire  _T_2276 = _T_2268 & _T_2275; // @[ifu_mem_ctl.scala 373:44]
  wire  stream_miss_f = _T_2276 & ifc_fetch_req_f; // @[ifu_mem_ctl.scala 373:84]
  wire  _T_318 = ~stream_miss_f; // @[ifu_mem_ctl.scala 226:106]
  reg  ifc_region_acc_fault_f; // @[ifu_mem_ctl.scala 232:68]
  reg [2:0] bus_rd_addr_count; // @[ifu_mem_ctl.scala 540:55]
  wire [28:0] ifu_ic_req_addr_f = {miss_addr,bus_rd_addr_count}; // @[Cat.scala 29:58]
  wire  _T_325 = _T_239 | _T_2268; // @[ifu_mem_ctl.scala 234:55]
  wire  _T_328 = _T_325 & _T_56; // @[ifu_mem_ctl.scala 234:82]
  wire  _T_2289 = ~ifu_bus_rid_ff[0]; // @[ifu_mem_ctl.scala 378:55]
  wire [2:0] other_tag = {ifu_bus_rid_ff[2:1],_T_2289}; // @[Cat.scala 29:58]
  wire  _T_2290 = other_tag == 3'h0; // @[ifu_mem_ctl.scala 379:81]
  wire  _T_2314 = _T_2290 & ic_miss_buff_data_valid[0]; // @[Mux.scala 27:72]
  wire  _T_2293 = other_tag == 3'h1; // @[ifu_mem_ctl.scala 379:81]
  wire  _T_2315 = _T_2293 & ic_miss_buff_data_valid[1]; // @[Mux.scala 27:72]
  wire  _T_2322 = _T_2314 | _T_2315; // @[Mux.scala 27:72]
  wire  _T_2296 = other_tag == 3'h2; // @[ifu_mem_ctl.scala 379:81]
  wire  _T_2316 = _T_2296 & ic_miss_buff_data_valid[2]; // @[Mux.scala 27:72]
  wire  _T_2323 = _T_2322 | _T_2316; // @[Mux.scala 27:72]
  wire  _T_2299 = other_tag == 3'h3; // @[ifu_mem_ctl.scala 379:81]
  wire  _T_2317 = _T_2299 & ic_miss_buff_data_valid[3]; // @[Mux.scala 27:72]
  wire  _T_2324 = _T_2323 | _T_2317; // @[Mux.scala 27:72]
  wire  _T_2302 = other_tag == 3'h4; // @[ifu_mem_ctl.scala 379:81]
  wire  _T_2318 = _T_2302 & ic_miss_buff_data_valid[4]; // @[Mux.scala 27:72]
  wire  _T_2325 = _T_2324 | _T_2318; // @[Mux.scala 27:72]
  wire  _T_2305 = other_tag == 3'h5; // @[ifu_mem_ctl.scala 379:81]
  wire  _T_2319 = _T_2305 & ic_miss_buff_data_valid[5]; // @[Mux.scala 27:72]
  wire  _T_2326 = _T_2325 | _T_2319; // @[Mux.scala 27:72]
  wire  _T_2308 = other_tag == 3'h6; // @[ifu_mem_ctl.scala 379:81]
  wire  _T_2320 = _T_2308 & ic_miss_buff_data_valid[6]; // @[Mux.scala 27:72]
  wire  _T_2327 = _T_2326 | _T_2320; // @[Mux.scala 27:72]
  wire  _T_2311 = other_tag == 3'h7; // @[ifu_mem_ctl.scala 379:81]
  wire  _T_2321 = _T_2311 & ic_miss_buff_data_valid[7]; // @[Mux.scala 27:72]
  wire  second_half_available = _T_2327 | _T_2321; // @[Mux.scala 27:72]
  wire  write_ic_16_bytes = second_half_available & bus_ifu_wr_en_ff; // @[ifu_mem_ctl.scala 380:46]
  wire  _T_332 = miss_pending & write_ic_16_bytes; // @[ifu_mem_ctl.scala 238:35]
  wire  _T_334 = _T_332 & _T_17; // @[ifu_mem_ctl.scala 238:55]
  reg  ic_act_miss_f_delayed; // @[ifu_mem_ctl.scala 555:61]
  wire  _T_2687 = ic_act_miss_f_delayed & _T_2284; // @[ifu_mem_ctl.scala 556:53]
  wire  reset_tag_valid_for_miss = _T_2687 & _T_17; // @[ifu_mem_ctl.scala 556:84]
  wire  sel_mb_addr = _T_334 | reset_tag_valid_for_miss; // @[ifu_mem_ctl.scala 238:79]
  wire [30:0] _T_338 = {imb_ff[30:5],ic_wr_addr_bits_hi_3,imb_ff[1:0]}; // @[Cat.scala 29:58]
  wire  _T_339 = ~sel_mb_addr; // @[ifu_mem_ctl.scala 240:37]
  wire [30:0] _T_340 = sel_mb_addr ? _T_338 : 31'h0; // @[Mux.scala 27:72]
  wire [30:0] _T_341 = _T_339 ? io_ifc_fetch_addr_bf : 31'h0; // @[Mux.scala 27:72]
  wire [30:0] ifu_ic_rw_int_addr = _T_340 | _T_341; // @[Mux.scala 27:72]
  wire  _T_346 = _T_334 & last_beat; // @[ifu_mem_ctl.scala 242:85]
  wire  _T_2681 = ~_T_2693; // @[ifu_mem_ctl.scala 553:84]
  wire  _T_2682 = _T_100 & _T_2681; // @[ifu_mem_ctl.scala 553:82]
  wire  bus_ifu_wr_en_ff_q = _T_2682 & write_ic_16_bytes; // @[ifu_mem_ctl.scala 553:108]
  wire  _T_347 = _T_346 & bus_ifu_wr_en_ff_q; // @[ifu_mem_ctl.scala 242:97]
  wire  sel_mb_status_addr = _T_347 | reset_tag_valid_for_miss; // @[ifu_mem_ctl.scala 242:119]
  wire [30:0] ifu_status_wr_addr = sel_mb_status_addr ? _T_338 : ifu_fetch_addr_int_f; // @[ifu_mem_ctl.scala 243:31]
  reg [63:0] ifu_bus_rdata_ff; // @[ifu_mem_ctl.scala 513:48]
  wire [6:0] _T_570 = {ifu_bus_rdata_ff[63],ifu_bus_rdata_ff[62],ifu_bus_rdata_ff[61],ifu_bus_rdata_ff[60],ifu_bus_rdata_ff[59],ifu_bus_rdata_ff[58],ifu_bus_rdata_ff[57]}; // @[lib.scala 276:13]
  wire  _T_571 = ^_T_570; // @[lib.scala 276:20]
  wire [6:0] _T_577 = {ifu_bus_rdata_ff[32],ifu_bus_rdata_ff[31],ifu_bus_rdata_ff[30],ifu_bus_rdata_ff[29],ifu_bus_rdata_ff[28],ifu_bus_rdata_ff[27],ifu_bus_rdata_ff[26]}; // @[lib.scala 276:30]
  wire [7:0] _T_584 = {ifu_bus_rdata_ff[40],ifu_bus_rdata_ff[39],ifu_bus_rdata_ff[38],ifu_bus_rdata_ff[37],ifu_bus_rdata_ff[36],ifu_bus_rdata_ff[35],ifu_bus_rdata_ff[34],ifu_bus_rdata_ff[33]}; // @[lib.scala 276:30]
  wire [14:0] _T_585 = {ifu_bus_rdata_ff[40],ifu_bus_rdata_ff[39],ifu_bus_rdata_ff[38],ifu_bus_rdata_ff[37],ifu_bus_rdata_ff[36],ifu_bus_rdata_ff[35],ifu_bus_rdata_ff[34],ifu_bus_rdata_ff[33],_T_577}; // @[lib.scala 276:30]
  wire [7:0] _T_592 = {ifu_bus_rdata_ff[48],ifu_bus_rdata_ff[47],ifu_bus_rdata_ff[46],ifu_bus_rdata_ff[45],ifu_bus_rdata_ff[44],ifu_bus_rdata_ff[43],ifu_bus_rdata_ff[42],ifu_bus_rdata_ff[41]}; // @[lib.scala 276:30]
  wire [30:0] _T_601 = {ifu_bus_rdata_ff[56],ifu_bus_rdata_ff[55],ifu_bus_rdata_ff[54],ifu_bus_rdata_ff[53],ifu_bus_rdata_ff[52],ifu_bus_rdata_ff[51],ifu_bus_rdata_ff[50],ifu_bus_rdata_ff[49],_T_592,_T_585}; // @[lib.scala 276:30]
  wire  _T_602 = ^_T_601; // @[lib.scala 276:37]
  wire [6:0] _T_608 = {ifu_bus_rdata_ff[17],ifu_bus_rdata_ff[16],ifu_bus_rdata_ff[15],ifu_bus_rdata_ff[14],ifu_bus_rdata_ff[13],ifu_bus_rdata_ff[12],ifu_bus_rdata_ff[11]}; // @[lib.scala 276:47]
  wire [14:0] _T_616 = {ifu_bus_rdata_ff[25],ifu_bus_rdata_ff[24],ifu_bus_rdata_ff[23],ifu_bus_rdata_ff[22],ifu_bus_rdata_ff[21],ifu_bus_rdata_ff[20],ifu_bus_rdata_ff[19],ifu_bus_rdata_ff[18],_T_608}; // @[lib.scala 276:47]
  wire [30:0] _T_632 = {ifu_bus_rdata_ff[56],ifu_bus_rdata_ff[55],ifu_bus_rdata_ff[54],ifu_bus_rdata_ff[53],ifu_bus_rdata_ff[52],ifu_bus_rdata_ff[51],ifu_bus_rdata_ff[50],ifu_bus_rdata_ff[49],_T_592,_T_616}; // @[lib.scala 276:47]
  wire  _T_633 = ^_T_632; // @[lib.scala 276:54]
  wire [6:0] _T_639 = {ifu_bus_rdata_ff[10],ifu_bus_rdata_ff[9],ifu_bus_rdata_ff[8],ifu_bus_rdata_ff[7],ifu_bus_rdata_ff[6],ifu_bus_rdata_ff[5],ifu_bus_rdata_ff[4]}; // @[lib.scala 276:64]
  wire [14:0] _T_647 = {ifu_bus_rdata_ff[25],ifu_bus_rdata_ff[24],ifu_bus_rdata_ff[23],ifu_bus_rdata_ff[22],ifu_bus_rdata_ff[21],ifu_bus_rdata_ff[20],ifu_bus_rdata_ff[19],ifu_bus_rdata_ff[18],_T_639}; // @[lib.scala 276:64]
  wire [30:0] _T_663 = {ifu_bus_rdata_ff[56],ifu_bus_rdata_ff[55],ifu_bus_rdata_ff[54],ifu_bus_rdata_ff[53],ifu_bus_rdata_ff[52],ifu_bus_rdata_ff[51],ifu_bus_rdata_ff[50],ifu_bus_rdata_ff[49],_T_584,_T_647}; // @[lib.scala 276:64]
  wire  _T_664 = ^_T_663; // @[lib.scala 276:71]
  wire [7:0] _T_671 = {ifu_bus_rdata_ff[14],ifu_bus_rdata_ff[10],ifu_bus_rdata_ff[9],ifu_bus_rdata_ff[8],ifu_bus_rdata_ff[7],ifu_bus_rdata_ff[3],ifu_bus_rdata_ff[2],ifu_bus_rdata_ff[1]}; // @[lib.scala 276:81]
  wire [16:0] _T_680 = {ifu_bus_rdata_ff[30],ifu_bus_rdata_ff[29],ifu_bus_rdata_ff[25],ifu_bus_rdata_ff[24],ifu_bus_rdata_ff[23],ifu_bus_rdata_ff[22],ifu_bus_rdata_ff[17],ifu_bus_rdata_ff[16],ifu_bus_rdata_ff[15],_T_671}; // @[lib.scala 276:81]
  wire [8:0] _T_688 = {ifu_bus_rdata_ff[47],ifu_bus_rdata_ff[46],ifu_bus_rdata_ff[45],ifu_bus_rdata_ff[40],ifu_bus_rdata_ff[39],ifu_bus_rdata_ff[38],ifu_bus_rdata_ff[37],ifu_bus_rdata_ff[32],ifu_bus_rdata_ff[31]}; // @[lib.scala 276:81]
  wire [17:0] _T_697 = {ifu_bus_rdata_ff[63],ifu_bus_rdata_ff[62],ifu_bus_rdata_ff[61],ifu_bus_rdata_ff[60],ifu_bus_rdata_ff[56],ifu_bus_rdata_ff[55],ifu_bus_rdata_ff[54],ifu_bus_rdata_ff[53],ifu_bus_rdata_ff[48],_T_688}; // @[lib.scala 276:81]
  wire [34:0] _T_698 = {_T_697,_T_680}; // @[lib.scala 276:81]
  wire  _T_699 = ^_T_698; // @[lib.scala 276:88]
  wire [7:0] _T_706 = {ifu_bus_rdata_ff[12],ifu_bus_rdata_ff[10],ifu_bus_rdata_ff[9],ifu_bus_rdata_ff[6],ifu_bus_rdata_ff[5],ifu_bus_rdata_ff[3],ifu_bus_rdata_ff[2],ifu_bus_rdata_ff[0]}; // @[lib.scala 276:98]
  wire [16:0] _T_715 = {ifu_bus_rdata_ff[28],ifu_bus_rdata_ff[27],ifu_bus_rdata_ff[25],ifu_bus_rdata_ff[24],ifu_bus_rdata_ff[21],ifu_bus_rdata_ff[20],ifu_bus_rdata_ff[17],ifu_bus_rdata_ff[16],ifu_bus_rdata_ff[13],_T_706}; // @[lib.scala 276:98]
  wire [8:0] _T_723 = {ifu_bus_rdata_ff[47],ifu_bus_rdata_ff[44],ifu_bus_rdata_ff[43],ifu_bus_rdata_ff[40],ifu_bus_rdata_ff[39],ifu_bus_rdata_ff[36],ifu_bus_rdata_ff[35],ifu_bus_rdata_ff[32],ifu_bus_rdata_ff[31]}; // @[lib.scala 276:98]
  wire [17:0] _T_732 = {ifu_bus_rdata_ff[63],ifu_bus_rdata_ff[62],ifu_bus_rdata_ff[59],ifu_bus_rdata_ff[58],ifu_bus_rdata_ff[56],ifu_bus_rdata_ff[55],ifu_bus_rdata_ff[52],ifu_bus_rdata_ff[51],ifu_bus_rdata_ff[48],_T_723}; // @[lib.scala 276:98]
  wire [34:0] _T_733 = {_T_732,_T_715}; // @[lib.scala 276:98]
  wire  _T_734 = ^_T_733; // @[lib.scala 276:105]
  wire [7:0] _T_741 = {ifu_bus_rdata_ff[11],ifu_bus_rdata_ff[10],ifu_bus_rdata_ff[8],ifu_bus_rdata_ff[6],ifu_bus_rdata_ff[4],ifu_bus_rdata_ff[3],ifu_bus_rdata_ff[1],ifu_bus_rdata_ff[0]}; // @[lib.scala 276:115]
  wire [16:0] _T_750 = {ifu_bus_rdata_ff[28],ifu_bus_rdata_ff[26],ifu_bus_rdata_ff[25],ifu_bus_rdata_ff[23],ifu_bus_rdata_ff[21],ifu_bus_rdata_ff[19],ifu_bus_rdata_ff[17],ifu_bus_rdata_ff[15],ifu_bus_rdata_ff[13],_T_741}; // @[lib.scala 276:115]
  wire [8:0] _T_758 = {ifu_bus_rdata_ff[46],ifu_bus_rdata_ff[44],ifu_bus_rdata_ff[42],ifu_bus_rdata_ff[40],ifu_bus_rdata_ff[38],ifu_bus_rdata_ff[36],ifu_bus_rdata_ff[34],ifu_bus_rdata_ff[32],ifu_bus_rdata_ff[30]}; // @[lib.scala 276:115]
  wire [17:0] _T_767 = {ifu_bus_rdata_ff[63],ifu_bus_rdata_ff[61],ifu_bus_rdata_ff[59],ifu_bus_rdata_ff[57],ifu_bus_rdata_ff[56],ifu_bus_rdata_ff[54],ifu_bus_rdata_ff[52],ifu_bus_rdata_ff[50],ifu_bus_rdata_ff[48],_T_758}; // @[lib.scala 276:115]
  wire [34:0] _T_768 = {_T_767,_T_750}; // @[lib.scala 276:115]
  wire  _T_769 = ^_T_768; // @[lib.scala 276:122]
  wire [3:0] _T_2330 = {ifu_bus_rid_ff[2:1],_T_2289,1'h1}; // @[Cat.scala 29:58]
  wire  _T_2331 = _T_2330 == 4'h0; // @[ifu_mem_ctl.scala 381:89]
  reg [31:0] ic_miss_buff_data_0; // @[ifu_mem_ctl.scala 316:65]
  wire [31:0] _T_2378 = _T_2331 ? ic_miss_buff_data_0 : 32'h0; // @[Mux.scala 27:72]
  wire  _T_2334 = _T_2330 == 4'h1; // @[ifu_mem_ctl.scala 381:89]
  reg [31:0] ic_miss_buff_data_1; // @[ifu_mem_ctl.scala 317:67]
  wire [31:0] _T_2379 = _T_2334 ? ic_miss_buff_data_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2394 = _T_2378 | _T_2379; // @[Mux.scala 27:72]
  wire  _T_2337 = _T_2330 == 4'h2; // @[ifu_mem_ctl.scala 381:89]
  reg [31:0] ic_miss_buff_data_2; // @[ifu_mem_ctl.scala 316:65]
  wire [31:0] _T_2380 = _T_2337 ? ic_miss_buff_data_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2395 = _T_2394 | _T_2380; // @[Mux.scala 27:72]
  wire  _T_2340 = _T_2330 == 4'h3; // @[ifu_mem_ctl.scala 381:89]
  reg [31:0] ic_miss_buff_data_3; // @[ifu_mem_ctl.scala 317:67]
  wire [31:0] _T_2381 = _T_2340 ? ic_miss_buff_data_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2396 = _T_2395 | _T_2381; // @[Mux.scala 27:72]
  wire  _T_2343 = _T_2330 == 4'h4; // @[ifu_mem_ctl.scala 381:89]
  reg [31:0] ic_miss_buff_data_4; // @[ifu_mem_ctl.scala 316:65]
  wire [31:0] _T_2382 = _T_2343 ? ic_miss_buff_data_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2397 = _T_2396 | _T_2382; // @[Mux.scala 27:72]
  wire  _T_2346 = _T_2330 == 4'h5; // @[ifu_mem_ctl.scala 381:89]
  reg [31:0] ic_miss_buff_data_5; // @[ifu_mem_ctl.scala 317:67]
  wire [31:0] _T_2383 = _T_2346 ? ic_miss_buff_data_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2398 = _T_2397 | _T_2383; // @[Mux.scala 27:72]
  wire  _T_2349 = _T_2330 == 4'h6; // @[ifu_mem_ctl.scala 381:89]
  reg [31:0] ic_miss_buff_data_6; // @[ifu_mem_ctl.scala 316:65]
  wire [31:0] _T_2384 = _T_2349 ? ic_miss_buff_data_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2399 = _T_2398 | _T_2384; // @[Mux.scala 27:72]
  wire  _T_2352 = _T_2330 == 4'h7; // @[ifu_mem_ctl.scala 381:89]
  reg [31:0] ic_miss_buff_data_7; // @[ifu_mem_ctl.scala 317:67]
  wire [31:0] _T_2385 = _T_2352 ? ic_miss_buff_data_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2400 = _T_2399 | _T_2385; // @[Mux.scala 27:72]
  wire  _T_2355 = _T_2330 == 4'h8; // @[ifu_mem_ctl.scala 381:89]
  reg [31:0] ic_miss_buff_data_8; // @[ifu_mem_ctl.scala 316:65]
  wire [31:0] _T_2386 = _T_2355 ? ic_miss_buff_data_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2401 = _T_2400 | _T_2386; // @[Mux.scala 27:72]
  wire  _T_2358 = _T_2330 == 4'h9; // @[ifu_mem_ctl.scala 381:89]
  reg [31:0] ic_miss_buff_data_9; // @[ifu_mem_ctl.scala 317:67]
  wire [31:0] _T_2387 = _T_2358 ? ic_miss_buff_data_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2402 = _T_2401 | _T_2387; // @[Mux.scala 27:72]
  wire  _T_2361 = _T_2330 == 4'ha; // @[ifu_mem_ctl.scala 381:89]
  reg [31:0] ic_miss_buff_data_10; // @[ifu_mem_ctl.scala 316:65]
  wire [31:0] _T_2388 = _T_2361 ? ic_miss_buff_data_10 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2403 = _T_2402 | _T_2388; // @[Mux.scala 27:72]
  wire  _T_2364 = _T_2330 == 4'hb; // @[ifu_mem_ctl.scala 381:89]
  reg [31:0] ic_miss_buff_data_11; // @[ifu_mem_ctl.scala 317:67]
  wire [31:0] _T_2389 = _T_2364 ? ic_miss_buff_data_11 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2404 = _T_2403 | _T_2389; // @[Mux.scala 27:72]
  wire  _T_2367 = _T_2330 == 4'hc; // @[ifu_mem_ctl.scala 381:89]
  reg [31:0] ic_miss_buff_data_12; // @[ifu_mem_ctl.scala 316:65]
  wire [31:0] _T_2390 = _T_2367 ? ic_miss_buff_data_12 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2405 = _T_2404 | _T_2390; // @[Mux.scala 27:72]
  wire  _T_2370 = _T_2330 == 4'hd; // @[ifu_mem_ctl.scala 381:89]
  reg [31:0] ic_miss_buff_data_13; // @[ifu_mem_ctl.scala 317:67]
  wire [31:0] _T_2391 = _T_2370 ? ic_miss_buff_data_13 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2406 = _T_2405 | _T_2391; // @[Mux.scala 27:72]
  wire  _T_2373 = _T_2330 == 4'he; // @[ifu_mem_ctl.scala 381:89]
  reg [31:0] ic_miss_buff_data_14; // @[ifu_mem_ctl.scala 316:65]
  wire [31:0] _T_2392 = _T_2373 ? ic_miss_buff_data_14 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2407 = _T_2406 | _T_2392; // @[Mux.scala 27:72]
  wire  _T_2376 = _T_2330 == 4'hf; // @[ifu_mem_ctl.scala 381:89]
  reg [31:0] ic_miss_buff_data_15; // @[ifu_mem_ctl.scala 317:67]
  wire [31:0] _T_2393 = _T_2376 ? ic_miss_buff_data_15 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2408 = _T_2407 | _T_2393; // @[Mux.scala 27:72]
  wire [3:0] _T_2410 = {ifu_bus_rid_ff[2:1],_T_2289,1'h0}; // @[Cat.scala 29:58]
  wire  _T_2411 = _T_2410 == 4'h0; // @[ifu_mem_ctl.scala 382:66]
  wire [31:0] _T_2458 = _T_2411 ? ic_miss_buff_data_0 : 32'h0; // @[Mux.scala 27:72]
  wire  _T_2414 = _T_2410 == 4'h1; // @[ifu_mem_ctl.scala 382:66]
  wire [31:0] _T_2459 = _T_2414 ? ic_miss_buff_data_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2474 = _T_2458 | _T_2459; // @[Mux.scala 27:72]
  wire  _T_2417 = _T_2410 == 4'h2; // @[ifu_mem_ctl.scala 382:66]
  wire [31:0] _T_2460 = _T_2417 ? ic_miss_buff_data_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2475 = _T_2474 | _T_2460; // @[Mux.scala 27:72]
  wire  _T_2420 = _T_2410 == 4'h3; // @[ifu_mem_ctl.scala 382:66]
  wire [31:0] _T_2461 = _T_2420 ? ic_miss_buff_data_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2476 = _T_2475 | _T_2461; // @[Mux.scala 27:72]
  wire  _T_2423 = _T_2410 == 4'h4; // @[ifu_mem_ctl.scala 382:66]
  wire [31:0] _T_2462 = _T_2423 ? ic_miss_buff_data_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2477 = _T_2476 | _T_2462; // @[Mux.scala 27:72]
  wire  _T_2426 = _T_2410 == 4'h5; // @[ifu_mem_ctl.scala 382:66]
  wire [31:0] _T_2463 = _T_2426 ? ic_miss_buff_data_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2478 = _T_2477 | _T_2463; // @[Mux.scala 27:72]
  wire  _T_2429 = _T_2410 == 4'h6; // @[ifu_mem_ctl.scala 382:66]
  wire [31:0] _T_2464 = _T_2429 ? ic_miss_buff_data_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2479 = _T_2478 | _T_2464; // @[Mux.scala 27:72]
  wire  _T_2432 = _T_2410 == 4'h7; // @[ifu_mem_ctl.scala 382:66]
  wire [31:0] _T_2465 = _T_2432 ? ic_miss_buff_data_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2480 = _T_2479 | _T_2465; // @[Mux.scala 27:72]
  wire  _T_2435 = _T_2410 == 4'h8; // @[ifu_mem_ctl.scala 382:66]
  wire [31:0] _T_2466 = _T_2435 ? ic_miss_buff_data_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2481 = _T_2480 | _T_2466; // @[Mux.scala 27:72]
  wire  _T_2438 = _T_2410 == 4'h9; // @[ifu_mem_ctl.scala 382:66]
  wire [31:0] _T_2467 = _T_2438 ? ic_miss_buff_data_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2482 = _T_2481 | _T_2467; // @[Mux.scala 27:72]
  wire  _T_2441 = _T_2410 == 4'ha; // @[ifu_mem_ctl.scala 382:66]
  wire [31:0] _T_2468 = _T_2441 ? ic_miss_buff_data_10 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2483 = _T_2482 | _T_2468; // @[Mux.scala 27:72]
  wire  _T_2444 = _T_2410 == 4'hb; // @[ifu_mem_ctl.scala 382:66]
  wire [31:0] _T_2469 = _T_2444 ? ic_miss_buff_data_11 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2484 = _T_2483 | _T_2469; // @[Mux.scala 27:72]
  wire  _T_2447 = _T_2410 == 4'hc; // @[ifu_mem_ctl.scala 382:66]
  wire [31:0] _T_2470 = _T_2447 ? ic_miss_buff_data_12 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2485 = _T_2484 | _T_2470; // @[Mux.scala 27:72]
  wire  _T_2450 = _T_2410 == 4'hd; // @[ifu_mem_ctl.scala 382:66]
  wire [31:0] _T_2471 = _T_2450 ? ic_miss_buff_data_13 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2486 = _T_2485 | _T_2471; // @[Mux.scala 27:72]
  wire  _T_2453 = _T_2410 == 4'he; // @[ifu_mem_ctl.scala 382:66]
  wire [31:0] _T_2472 = _T_2453 ? ic_miss_buff_data_14 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2487 = _T_2486 | _T_2472; // @[Mux.scala 27:72]
  wire  _T_2456 = _T_2410 == 4'hf; // @[ifu_mem_ctl.scala 382:66]
  wire [31:0] _T_2473 = _T_2456 ? ic_miss_buff_data_15 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2488 = _T_2487 | _T_2473; // @[Mux.scala 27:72]
  wire [63:0] ic_miss_buff_half = {_T_2408,_T_2488}; // @[Cat.scala 29:58]
  wire [6:0] _T_992 = {ic_miss_buff_half[63],ic_miss_buff_half[62],ic_miss_buff_half[61],ic_miss_buff_half[60],ic_miss_buff_half[59],ic_miss_buff_half[58],ic_miss_buff_half[57]}; // @[lib.scala 276:13]
  wire  _T_993 = ^_T_992; // @[lib.scala 276:20]
  wire [6:0] _T_999 = {ic_miss_buff_half[32],ic_miss_buff_half[31],ic_miss_buff_half[30],ic_miss_buff_half[29],ic_miss_buff_half[28],ic_miss_buff_half[27],ic_miss_buff_half[26]}; // @[lib.scala 276:30]
  wire [7:0] _T_1006 = {ic_miss_buff_half[40],ic_miss_buff_half[39],ic_miss_buff_half[38],ic_miss_buff_half[37],ic_miss_buff_half[36],ic_miss_buff_half[35],ic_miss_buff_half[34],ic_miss_buff_half[33]}; // @[lib.scala 276:30]
  wire [14:0] _T_1007 = {ic_miss_buff_half[40],ic_miss_buff_half[39],ic_miss_buff_half[38],ic_miss_buff_half[37],ic_miss_buff_half[36],ic_miss_buff_half[35],ic_miss_buff_half[34],ic_miss_buff_half[33],_T_999}; // @[lib.scala 276:30]
  wire [7:0] _T_1014 = {ic_miss_buff_half[48],ic_miss_buff_half[47],ic_miss_buff_half[46],ic_miss_buff_half[45],ic_miss_buff_half[44],ic_miss_buff_half[43],ic_miss_buff_half[42],ic_miss_buff_half[41]}; // @[lib.scala 276:30]
  wire [30:0] _T_1023 = {ic_miss_buff_half[56],ic_miss_buff_half[55],ic_miss_buff_half[54],ic_miss_buff_half[53],ic_miss_buff_half[52],ic_miss_buff_half[51],ic_miss_buff_half[50],ic_miss_buff_half[49],_T_1014,_T_1007}; // @[lib.scala 276:30]
  wire  _T_1024 = ^_T_1023; // @[lib.scala 276:37]
  wire [6:0] _T_1030 = {ic_miss_buff_half[17],ic_miss_buff_half[16],ic_miss_buff_half[15],ic_miss_buff_half[14],ic_miss_buff_half[13],ic_miss_buff_half[12],ic_miss_buff_half[11]}; // @[lib.scala 276:47]
  wire [14:0] _T_1038 = {ic_miss_buff_half[25],ic_miss_buff_half[24],ic_miss_buff_half[23],ic_miss_buff_half[22],ic_miss_buff_half[21],ic_miss_buff_half[20],ic_miss_buff_half[19],ic_miss_buff_half[18],_T_1030}; // @[lib.scala 276:47]
  wire [30:0] _T_1054 = {ic_miss_buff_half[56],ic_miss_buff_half[55],ic_miss_buff_half[54],ic_miss_buff_half[53],ic_miss_buff_half[52],ic_miss_buff_half[51],ic_miss_buff_half[50],ic_miss_buff_half[49],_T_1014,_T_1038}; // @[lib.scala 276:47]
  wire  _T_1055 = ^_T_1054; // @[lib.scala 276:54]
  wire [6:0] _T_1061 = {ic_miss_buff_half[10],ic_miss_buff_half[9],ic_miss_buff_half[8],ic_miss_buff_half[7],ic_miss_buff_half[6],ic_miss_buff_half[5],ic_miss_buff_half[4]}; // @[lib.scala 276:64]
  wire [14:0] _T_1069 = {ic_miss_buff_half[25],ic_miss_buff_half[24],ic_miss_buff_half[23],ic_miss_buff_half[22],ic_miss_buff_half[21],ic_miss_buff_half[20],ic_miss_buff_half[19],ic_miss_buff_half[18],_T_1061}; // @[lib.scala 276:64]
  wire [30:0] _T_1085 = {ic_miss_buff_half[56],ic_miss_buff_half[55],ic_miss_buff_half[54],ic_miss_buff_half[53],ic_miss_buff_half[52],ic_miss_buff_half[51],ic_miss_buff_half[50],ic_miss_buff_half[49],_T_1006,_T_1069}; // @[lib.scala 276:64]
  wire  _T_1086 = ^_T_1085; // @[lib.scala 276:71]
  wire [7:0] _T_1093 = {ic_miss_buff_half[14],ic_miss_buff_half[10],ic_miss_buff_half[9],ic_miss_buff_half[8],ic_miss_buff_half[7],ic_miss_buff_half[3],ic_miss_buff_half[2],ic_miss_buff_half[1]}; // @[lib.scala 276:81]
  wire [16:0] _T_1102 = {ic_miss_buff_half[30],ic_miss_buff_half[29],ic_miss_buff_half[25],ic_miss_buff_half[24],ic_miss_buff_half[23],ic_miss_buff_half[22],ic_miss_buff_half[17],ic_miss_buff_half[16],ic_miss_buff_half[15],_T_1093}; // @[lib.scala 276:81]
  wire [8:0] _T_1110 = {ic_miss_buff_half[47],ic_miss_buff_half[46],ic_miss_buff_half[45],ic_miss_buff_half[40],ic_miss_buff_half[39],ic_miss_buff_half[38],ic_miss_buff_half[37],ic_miss_buff_half[32],ic_miss_buff_half[31]}; // @[lib.scala 276:81]
  wire [17:0] _T_1119 = {ic_miss_buff_half[63],ic_miss_buff_half[62],ic_miss_buff_half[61],ic_miss_buff_half[60],ic_miss_buff_half[56],ic_miss_buff_half[55],ic_miss_buff_half[54],ic_miss_buff_half[53],ic_miss_buff_half[48],_T_1110}; // @[lib.scala 276:81]
  wire [34:0] _T_1120 = {_T_1119,_T_1102}; // @[lib.scala 276:81]
  wire  _T_1121 = ^_T_1120; // @[lib.scala 276:88]
  wire [7:0] _T_1128 = {ic_miss_buff_half[12],ic_miss_buff_half[10],ic_miss_buff_half[9],ic_miss_buff_half[6],ic_miss_buff_half[5],ic_miss_buff_half[3],ic_miss_buff_half[2],ic_miss_buff_half[0]}; // @[lib.scala 276:98]
  wire [16:0] _T_1137 = {ic_miss_buff_half[28],ic_miss_buff_half[27],ic_miss_buff_half[25],ic_miss_buff_half[24],ic_miss_buff_half[21],ic_miss_buff_half[20],ic_miss_buff_half[17],ic_miss_buff_half[16],ic_miss_buff_half[13],_T_1128}; // @[lib.scala 276:98]
  wire [8:0] _T_1145 = {ic_miss_buff_half[47],ic_miss_buff_half[44],ic_miss_buff_half[43],ic_miss_buff_half[40],ic_miss_buff_half[39],ic_miss_buff_half[36],ic_miss_buff_half[35],ic_miss_buff_half[32],ic_miss_buff_half[31]}; // @[lib.scala 276:98]
  wire [17:0] _T_1154 = {ic_miss_buff_half[63],ic_miss_buff_half[62],ic_miss_buff_half[59],ic_miss_buff_half[58],ic_miss_buff_half[56],ic_miss_buff_half[55],ic_miss_buff_half[52],ic_miss_buff_half[51],ic_miss_buff_half[48],_T_1145}; // @[lib.scala 276:98]
  wire [34:0] _T_1155 = {_T_1154,_T_1137}; // @[lib.scala 276:98]
  wire  _T_1156 = ^_T_1155; // @[lib.scala 276:105]
  wire [7:0] _T_1163 = {ic_miss_buff_half[11],ic_miss_buff_half[10],ic_miss_buff_half[8],ic_miss_buff_half[6],ic_miss_buff_half[4],ic_miss_buff_half[3],ic_miss_buff_half[1],ic_miss_buff_half[0]}; // @[lib.scala 276:115]
  wire [16:0] _T_1172 = {ic_miss_buff_half[28],ic_miss_buff_half[26],ic_miss_buff_half[25],ic_miss_buff_half[23],ic_miss_buff_half[21],ic_miss_buff_half[19],ic_miss_buff_half[17],ic_miss_buff_half[15],ic_miss_buff_half[13],_T_1163}; // @[lib.scala 276:115]
  wire [8:0] _T_1180 = {ic_miss_buff_half[46],ic_miss_buff_half[44],ic_miss_buff_half[42],ic_miss_buff_half[40],ic_miss_buff_half[38],ic_miss_buff_half[36],ic_miss_buff_half[34],ic_miss_buff_half[32],ic_miss_buff_half[30]}; // @[lib.scala 276:115]
  wire [17:0] _T_1189 = {ic_miss_buff_half[63],ic_miss_buff_half[61],ic_miss_buff_half[59],ic_miss_buff_half[57],ic_miss_buff_half[56],ic_miss_buff_half[54],ic_miss_buff_half[52],ic_miss_buff_half[50],ic_miss_buff_half[48],_T_1180}; // @[lib.scala 276:115]
  wire [34:0] _T_1190 = {_T_1189,_T_1172}; // @[lib.scala 276:115]
  wire  _T_1191 = ^_T_1190; // @[lib.scala 276:122]
  wire [70:0] _T_1236 = {_T_571,_T_602,_T_633,_T_664,_T_699,_T_734,_T_769,ifu_bus_rdata_ff}; // @[Cat.scala 29:58]
  wire [70:0] _T_1235 = {_T_993,_T_1024,_T_1055,_T_1086,_T_1121,_T_1156,_T_1191,_T_2408,_T_2488}; // @[Cat.scala 29:58]
  wire [141:0] _T_1237 = {_T_571,_T_602,_T_633,_T_664,_T_699,_T_734,_T_769,ifu_bus_rdata_ff,_T_1235}; // @[Cat.scala 29:58]
  wire [141:0] _T_1240 = {_T_993,_T_1024,_T_1055,_T_1086,_T_1121,_T_1156,_T_1191,_T_2408,_T_2488,_T_1236}; // @[Cat.scala 29:58]
  wire [141:0] ic_wr_16bytes_data = ifu_bus_rid_ff[0] ? _T_1237 : _T_1240; // @[ifu_mem_ctl.scala 267:28]
  wire  _T_1199 = |io_ic_eccerr; // @[ifu_mem_ctl.scala 256:73]
  wire  _T_1200 = _T_1199 & ic_act_hit_f; // @[ifu_mem_ctl.scala 256:100]
  wire [4:0] bypass_index = imb_ff[4:0]; // @[ifu_mem_ctl.scala 328:28]
  wire  _T_1404 = bypass_index[4:2] == 3'h0; // @[ifu_mem_ctl.scala 330:114]
  wire  bus_ifu_wr_en = _T_13 & miss_pending; // @[ifu_mem_ctl.scala 551:35]
  wire  _T_1289 = io_ifu_axi_r_bits_id == 3'h0; // @[ifu_mem_ctl.scala 312:91]
  wire  write_fill_data_0 = bus_ifu_wr_en & _T_1289; // @[ifu_mem_ctl.scala 312:73]
  wire  _T_1330 = ~ic_act_miss_f; // @[ifu_mem_ctl.scala 319:118]
  wire  _T_1331 = ic_miss_buff_data_valid[0] & _T_1330; // @[ifu_mem_ctl.scala 319:116]
  wire  ic_miss_buff_data_valid_in_0 = write_fill_data_0 | _T_1331; // @[ifu_mem_ctl.scala 319:88]
  wire  _T_1427 = _T_1404 & ic_miss_buff_data_valid_in_0; // @[Mux.scala 27:72]
  wire  _T_1407 = bypass_index[4:2] == 3'h1; // @[ifu_mem_ctl.scala 330:114]
  wire  _T_1290 = io_ifu_axi_r_bits_id == 3'h1; // @[ifu_mem_ctl.scala 312:91]
  wire  write_fill_data_1 = bus_ifu_wr_en & _T_1290; // @[ifu_mem_ctl.scala 312:73]
  wire  _T_1334 = ic_miss_buff_data_valid[1] & _T_1330; // @[ifu_mem_ctl.scala 319:116]
  wire  ic_miss_buff_data_valid_in_1 = write_fill_data_1 | _T_1334; // @[ifu_mem_ctl.scala 319:88]
  wire  _T_1428 = _T_1407 & ic_miss_buff_data_valid_in_1; // @[Mux.scala 27:72]
  wire  _T_1435 = _T_1427 | _T_1428; // @[Mux.scala 27:72]
  wire  _T_1410 = bypass_index[4:2] == 3'h2; // @[ifu_mem_ctl.scala 330:114]
  wire  _T_1291 = io_ifu_axi_r_bits_id == 3'h2; // @[ifu_mem_ctl.scala 312:91]
  wire  write_fill_data_2 = bus_ifu_wr_en & _T_1291; // @[ifu_mem_ctl.scala 312:73]
  wire  _T_1337 = ic_miss_buff_data_valid[2] & _T_1330; // @[ifu_mem_ctl.scala 319:116]
  wire  ic_miss_buff_data_valid_in_2 = write_fill_data_2 | _T_1337; // @[ifu_mem_ctl.scala 319:88]
  wire  _T_1429 = _T_1410 & ic_miss_buff_data_valid_in_2; // @[Mux.scala 27:72]
  wire  _T_1436 = _T_1435 | _T_1429; // @[Mux.scala 27:72]
  wire  _T_1413 = bypass_index[4:2] == 3'h3; // @[ifu_mem_ctl.scala 330:114]
  wire  _T_1292 = io_ifu_axi_r_bits_id == 3'h3; // @[ifu_mem_ctl.scala 312:91]
  wire  write_fill_data_3 = bus_ifu_wr_en & _T_1292; // @[ifu_mem_ctl.scala 312:73]
  wire  _T_1340 = ic_miss_buff_data_valid[3] & _T_1330; // @[ifu_mem_ctl.scala 319:116]
  wire  ic_miss_buff_data_valid_in_3 = write_fill_data_3 | _T_1340; // @[ifu_mem_ctl.scala 319:88]
  wire  _T_1430 = _T_1413 & ic_miss_buff_data_valid_in_3; // @[Mux.scala 27:72]
  wire  _T_1437 = _T_1436 | _T_1430; // @[Mux.scala 27:72]
  wire  _T_1416 = bypass_index[4:2] == 3'h4; // @[ifu_mem_ctl.scala 330:114]
  wire  _T_1293 = io_ifu_axi_r_bits_id == 3'h4; // @[ifu_mem_ctl.scala 312:91]
  wire  write_fill_data_4 = bus_ifu_wr_en & _T_1293; // @[ifu_mem_ctl.scala 312:73]
  wire  _T_1343 = ic_miss_buff_data_valid[4] & _T_1330; // @[ifu_mem_ctl.scala 319:116]
  wire  ic_miss_buff_data_valid_in_4 = write_fill_data_4 | _T_1343; // @[ifu_mem_ctl.scala 319:88]
  wire  _T_1431 = _T_1416 & ic_miss_buff_data_valid_in_4; // @[Mux.scala 27:72]
  wire  _T_1438 = _T_1437 | _T_1431; // @[Mux.scala 27:72]
  wire  _T_1419 = bypass_index[4:2] == 3'h5; // @[ifu_mem_ctl.scala 330:114]
  wire  _T_1294 = io_ifu_axi_r_bits_id == 3'h5; // @[ifu_mem_ctl.scala 312:91]
  wire  write_fill_data_5 = bus_ifu_wr_en & _T_1294; // @[ifu_mem_ctl.scala 312:73]
  wire  _T_1346 = ic_miss_buff_data_valid[5] & _T_1330; // @[ifu_mem_ctl.scala 319:116]
  wire  ic_miss_buff_data_valid_in_5 = write_fill_data_5 | _T_1346; // @[ifu_mem_ctl.scala 319:88]
  wire  _T_1432 = _T_1419 & ic_miss_buff_data_valid_in_5; // @[Mux.scala 27:72]
  wire  _T_1439 = _T_1438 | _T_1432; // @[Mux.scala 27:72]
  wire  _T_1422 = bypass_index[4:2] == 3'h6; // @[ifu_mem_ctl.scala 330:114]
  wire  _T_1295 = io_ifu_axi_r_bits_id == 3'h6; // @[ifu_mem_ctl.scala 312:91]
  wire  write_fill_data_6 = bus_ifu_wr_en & _T_1295; // @[ifu_mem_ctl.scala 312:73]
  wire  _T_1349 = ic_miss_buff_data_valid[6] & _T_1330; // @[ifu_mem_ctl.scala 319:116]
  wire  ic_miss_buff_data_valid_in_6 = write_fill_data_6 | _T_1349; // @[ifu_mem_ctl.scala 319:88]
  wire  _T_1433 = _T_1422 & ic_miss_buff_data_valid_in_6; // @[Mux.scala 27:72]
  wire  _T_1440 = _T_1439 | _T_1433; // @[Mux.scala 27:72]
  wire  _T_1425 = bypass_index[4:2] == 3'h7; // @[ifu_mem_ctl.scala 330:114]
  wire  _T_1296 = io_ifu_axi_r_bits_id == 3'h7; // @[ifu_mem_ctl.scala 312:91]
  wire  write_fill_data_7 = bus_ifu_wr_en & _T_1296; // @[ifu_mem_ctl.scala 312:73]
  wire  _T_1352 = ic_miss_buff_data_valid[7] & _T_1330; // @[ifu_mem_ctl.scala 319:116]
  wire  ic_miss_buff_data_valid_in_7 = write_fill_data_7 | _T_1352; // @[ifu_mem_ctl.scala 319:88]
  wire  _T_1434 = _T_1425 & ic_miss_buff_data_valid_in_7; // @[Mux.scala 27:72]
  wire  bypass_valid_value_check = _T_1440 | _T_1434; // @[Mux.scala 27:72]
  wire  _T_1443 = ~bypass_index[1]; // @[ifu_mem_ctl.scala 331:58]
  wire  _T_1444 = bypass_valid_value_check & _T_1443; // @[ifu_mem_ctl.scala 331:56]
  wire  _T_1446 = ~bypass_index[0]; // @[ifu_mem_ctl.scala 331:77]
  wire  _T_1447 = _T_1444 & _T_1446; // @[ifu_mem_ctl.scala 331:75]
  wire  _T_1452 = _T_1444 & bypass_index[0]; // @[ifu_mem_ctl.scala 332:75]
  wire  _T_1453 = _T_1447 | _T_1452; // @[ifu_mem_ctl.scala 331:95]
  wire  _T_1455 = bypass_valid_value_check & bypass_index[1]; // @[ifu_mem_ctl.scala 333:56]
  wire  _T_1458 = _T_1455 & _T_1446; // @[ifu_mem_ctl.scala 333:74]
  wire  _T_1459 = _T_1453 | _T_1458; // @[ifu_mem_ctl.scala 332:94]
  wire  _T_1463 = _T_1455 & bypass_index[0]; // @[ifu_mem_ctl.scala 334:51]
  wire [2:0] bypass_index_5_3_inc = bypass_index[4:2] + 3'h1; // @[ifu_mem_ctl.scala 329:70]
  wire  _T_1464 = bypass_index_5_3_inc == 3'h0; // @[ifu_mem_ctl.scala 334:132]
  wire  _T_1480 = _T_1464 & ic_miss_buff_data_valid_in_0; // @[Mux.scala 27:72]
  wire  _T_1466 = bypass_index_5_3_inc == 3'h1; // @[ifu_mem_ctl.scala 334:132]
  wire  _T_1481 = _T_1466 & ic_miss_buff_data_valid_in_1; // @[Mux.scala 27:72]
  wire  _T_1488 = _T_1480 | _T_1481; // @[Mux.scala 27:72]
  wire  _T_1468 = bypass_index_5_3_inc == 3'h2; // @[ifu_mem_ctl.scala 334:132]
  wire  _T_1482 = _T_1468 & ic_miss_buff_data_valid_in_2; // @[Mux.scala 27:72]
  wire  _T_1489 = _T_1488 | _T_1482; // @[Mux.scala 27:72]
  wire  _T_1470 = bypass_index_5_3_inc == 3'h3; // @[ifu_mem_ctl.scala 334:132]
  wire  _T_1483 = _T_1470 & ic_miss_buff_data_valid_in_3; // @[Mux.scala 27:72]
  wire  _T_1490 = _T_1489 | _T_1483; // @[Mux.scala 27:72]
  wire  _T_1472 = bypass_index_5_3_inc == 3'h4; // @[ifu_mem_ctl.scala 334:132]
  wire  _T_1484 = _T_1472 & ic_miss_buff_data_valid_in_4; // @[Mux.scala 27:72]
  wire  _T_1491 = _T_1490 | _T_1484; // @[Mux.scala 27:72]
  wire  _T_1474 = bypass_index_5_3_inc == 3'h5; // @[ifu_mem_ctl.scala 334:132]
  wire  _T_1485 = _T_1474 & ic_miss_buff_data_valid_in_5; // @[Mux.scala 27:72]
  wire  _T_1492 = _T_1491 | _T_1485; // @[Mux.scala 27:72]
  wire  _T_1476 = bypass_index_5_3_inc == 3'h6; // @[ifu_mem_ctl.scala 334:132]
  wire  _T_1486 = _T_1476 & ic_miss_buff_data_valid_in_6; // @[Mux.scala 27:72]
  wire  _T_1493 = _T_1492 | _T_1486; // @[Mux.scala 27:72]
  wire  _T_1478 = bypass_index_5_3_inc == 3'h7; // @[ifu_mem_ctl.scala 334:132]
  wire  _T_1487 = _T_1478 & ic_miss_buff_data_valid_in_7; // @[Mux.scala 27:72]
  wire  _T_1494 = _T_1493 | _T_1487; // @[Mux.scala 27:72]
  wire  _T_1496 = _T_1463 & _T_1494; // @[ifu_mem_ctl.scala 334:69]
  wire  _T_1497 = _T_1459 | _T_1496; // @[ifu_mem_ctl.scala 333:94]
  wire [4:0] _GEN_436 = {{2'd0}, bypass_index[4:2]}; // @[ifu_mem_ctl.scala 335:95]
  wire  _T_1500 = _GEN_436 == 5'h1f; // @[ifu_mem_ctl.scala 335:95]
  wire  _T_1501 = bypass_valid_value_check & _T_1500; // @[ifu_mem_ctl.scala 335:56]
  wire  bypass_data_ready_in = _T_1497 | _T_1501; // @[ifu_mem_ctl.scala 334:181]
  wire  _T_1502 = bypass_data_ready_in & crit_wd_byp_ok_ff; // @[ifu_mem_ctl.scala 339:53]
  wire  _T_1503 = _T_1502 & uncacheable_miss_ff; // @[ifu_mem_ctl.scala 339:73]
  wire  _T_1505 = _T_1503 & _T_319; // @[ifu_mem_ctl.scala 339:96]
  wire  _T_1507 = _T_1505 & _T_58; // @[ifu_mem_ctl.scala 339:118]
  wire  _T_1509 = crit_wd_byp_ok_ff & _T_17; // @[ifu_mem_ctl.scala 340:73]
  wire  _T_1511 = _T_1509 & _T_319; // @[ifu_mem_ctl.scala 340:96]
  wire  _T_1513 = _T_1511 & _T_58; // @[ifu_mem_ctl.scala 340:118]
  wire  _T_1514 = _T_1507 | _T_1513; // @[ifu_mem_ctl.scala 339:143]
  reg  ic_crit_wd_rdy_new_ff; // @[ifu_mem_ctl.scala 342:58]
  wire  _T_1515 = ic_crit_wd_rdy_new_ff & crit_wd_byp_ok_ff; // @[ifu_mem_ctl.scala 341:54]
  wire  _T_1516 = ~fetch_req_icache_f; // @[ifu_mem_ctl.scala 341:76]
  wire  _T_1517 = _T_1515 & _T_1516; // @[ifu_mem_ctl.scala 341:74]
  wire  _T_1519 = _T_1517 & _T_319; // @[ifu_mem_ctl.scala 341:96]
  wire  ic_crit_wd_rdy_new_in = _T_1514 | _T_1519; // @[ifu_mem_ctl.scala 340:143]
  wire  ic_crit_wd_rdy = ic_crit_wd_rdy_new_in | ic_crit_wd_rdy_new_ff; // @[ifu_mem_ctl.scala 561:43]
  wire  _T_1252 = ic_crit_wd_rdy | _T_2268; // @[ifu_mem_ctl.scala 280:38]
  wire  _T_1254 = _T_1252 | _T_2284; // @[ifu_mem_ctl.scala 280:64]
  wire  _T_1255 = ~_T_1254; // @[ifu_mem_ctl.scala 280:21]
  wire  _T_1256 = ~fetch_req_iccm_f; // @[ifu_mem_ctl.scala 280:98]
  wire  sel_ic_data = _T_1255 & _T_1256; // @[ifu_mem_ctl.scala 280:96]
  wire  _T_2491 = io_ic_tag_perr & sel_ic_data; // @[ifu_mem_ctl.scala 385:44]
  wire  _T_1612 = ~ifu_fetch_addr_int_f[1]; // @[ifu_mem_ctl.scala 351:30]
  wire  _T_1614 = ~ifu_fetch_addr_int_f[0]; // @[ifu_mem_ctl.scala 351:57]
  wire  _T_1615 = _T_1612 & _T_1614; // @[ifu_mem_ctl.scala 351:55]
  reg [7:0] ic_miss_buff_data_error; // @[ifu_mem_ctl.scala 325:60]
  wire [7:0] _T_1617 = ic_miss_buff_data_error >> byp_fetch_index[4:2]; // @[ifu_mem_ctl.scala 351:107]
  wire  _T_1619 = _T_1615 & _T_1617[0]; // @[ifu_mem_ctl.scala 351:82]
  wire  _T_1623 = _T_1612 & ifu_fetch_addr_int_f[0]; // @[ifu_mem_ctl.scala 352:33]
  wire  _T_1627 = _T_1623 & _T_1617[0]; // @[ifu_mem_ctl.scala 352:60]
  wire  _T_1628 = _T_1619 | _T_1627; // @[ifu_mem_ctl.scala 351:151]
  wire  _T_1637 = _T_1628 | _T_1627; // @[ifu_mem_ctl.scala 352:129]
  wire  _T_1641 = ifu_fetch_addr_int_f[1] & _T_1614; // @[ifu_mem_ctl.scala 354:33]
  wire  _T_1645 = _T_1641 & _T_1617[0]; // @[ifu_mem_ctl.scala 354:60]
  wire  _T_1646 = _T_1637 | _T_1645; // @[ifu_mem_ctl.scala 353:129]
  wire  _T_1649 = ifu_fetch_addr_int_f[1] & ifu_fetch_addr_int_f[0]; // @[ifu_mem_ctl.scala 355:32]
  wire [7:0] _T_1654 = ic_miss_buff_data_error >> byp_fetch_index_inc; // @[ifu_mem_ctl.scala 356:32]
  wire  _T_1656 = _T_1617[0] | _T_1654[0]; // @[ifu_mem_ctl.scala 355:127]
  wire  _T_1657 = _T_1649 & _T_1656; // @[ifu_mem_ctl.scala 355:58]
  wire  ifu_byp_data_err_new = _T_1646 | _T_1657; // @[ifu_mem_ctl.scala 354:129]
  wire  ifc_bus_acc_fault_f = ic_byp_hit_f & ifu_byp_data_err_new; // @[ifu_mem_ctl.scala 297:42]
  wire  _T_2492 = ifc_region_acc_fault_final_f | ifc_bus_acc_fault_f; // @[ifu_mem_ctl.scala 385:91]
  wire  _T_2493 = ~_T_2492; // @[ifu_mem_ctl.scala 385:60]
  wire  ic_rd_parity_final_err = _T_2491 & _T_2493; // @[ifu_mem_ctl.scala 385:58]
  reg  ic_debug_ict_array_sel_ff; // @[ifu_mem_ctl.scala 768:63]
  reg  ic_tag_valid_out_1_0; // @[Reg.scala 27:20]
  wire  _T_9374 = _T_4671 & ic_tag_valid_out_1_0; // @[ifu_mem_ctl.scala 696:10]
  reg  ic_tag_valid_out_1_1; // @[Reg.scala 27:20]
  wire  _T_9376 = _T_4672 & ic_tag_valid_out_1_1; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9629 = _T_9374 | _T_9376; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_2; // @[Reg.scala 27:20]
  wire  _T_9378 = _T_4673 & ic_tag_valid_out_1_2; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9630 = _T_9629 | _T_9378; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_3; // @[Reg.scala 27:20]
  wire  _T_9380 = _T_4674 & ic_tag_valid_out_1_3; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9631 = _T_9630 | _T_9380; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_4; // @[Reg.scala 27:20]
  wire  _T_9382 = _T_4675 & ic_tag_valid_out_1_4; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9632 = _T_9631 | _T_9382; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_5; // @[Reg.scala 27:20]
  wire  _T_9384 = _T_4676 & ic_tag_valid_out_1_5; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9633 = _T_9632 | _T_9384; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_6; // @[Reg.scala 27:20]
  wire  _T_9386 = _T_4677 & ic_tag_valid_out_1_6; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9634 = _T_9633 | _T_9386; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_7; // @[Reg.scala 27:20]
  wire  _T_9388 = _T_4678 & ic_tag_valid_out_1_7; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9635 = _T_9634 | _T_9388; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_8; // @[Reg.scala 27:20]
  wire  _T_9390 = _T_4679 & ic_tag_valid_out_1_8; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9636 = _T_9635 | _T_9390; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_9; // @[Reg.scala 27:20]
  wire  _T_9392 = _T_4680 & ic_tag_valid_out_1_9; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9637 = _T_9636 | _T_9392; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_10; // @[Reg.scala 27:20]
  wire  _T_9394 = _T_4681 & ic_tag_valid_out_1_10; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9638 = _T_9637 | _T_9394; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_11; // @[Reg.scala 27:20]
  wire  _T_9396 = _T_4682 & ic_tag_valid_out_1_11; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9639 = _T_9638 | _T_9396; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_12; // @[Reg.scala 27:20]
  wire  _T_9398 = _T_4683 & ic_tag_valid_out_1_12; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9640 = _T_9639 | _T_9398; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_13; // @[Reg.scala 27:20]
  wire  _T_9400 = _T_4684 & ic_tag_valid_out_1_13; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9641 = _T_9640 | _T_9400; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_14; // @[Reg.scala 27:20]
  wire  _T_9402 = _T_4685 & ic_tag_valid_out_1_14; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9642 = _T_9641 | _T_9402; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_15; // @[Reg.scala 27:20]
  wire  _T_9404 = _T_4686 & ic_tag_valid_out_1_15; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9643 = _T_9642 | _T_9404; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_16; // @[Reg.scala 27:20]
  wire  _T_9406 = _T_4687 & ic_tag_valid_out_1_16; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9644 = _T_9643 | _T_9406; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_17; // @[Reg.scala 27:20]
  wire  _T_9408 = _T_4688 & ic_tag_valid_out_1_17; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9645 = _T_9644 | _T_9408; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_18; // @[Reg.scala 27:20]
  wire  _T_9410 = _T_4689 & ic_tag_valid_out_1_18; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9646 = _T_9645 | _T_9410; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_19; // @[Reg.scala 27:20]
  wire  _T_9412 = _T_4690 & ic_tag_valid_out_1_19; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9647 = _T_9646 | _T_9412; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_20; // @[Reg.scala 27:20]
  wire  _T_9414 = _T_4691 & ic_tag_valid_out_1_20; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9648 = _T_9647 | _T_9414; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_21; // @[Reg.scala 27:20]
  wire  _T_9416 = _T_4692 & ic_tag_valid_out_1_21; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9649 = _T_9648 | _T_9416; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_22; // @[Reg.scala 27:20]
  wire  _T_9418 = _T_4693 & ic_tag_valid_out_1_22; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9650 = _T_9649 | _T_9418; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_23; // @[Reg.scala 27:20]
  wire  _T_9420 = _T_4694 & ic_tag_valid_out_1_23; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9651 = _T_9650 | _T_9420; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_24; // @[Reg.scala 27:20]
  wire  _T_9422 = _T_4695 & ic_tag_valid_out_1_24; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9652 = _T_9651 | _T_9422; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_25; // @[Reg.scala 27:20]
  wire  _T_9424 = _T_4696 & ic_tag_valid_out_1_25; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9653 = _T_9652 | _T_9424; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_26; // @[Reg.scala 27:20]
  wire  _T_9426 = _T_4697 & ic_tag_valid_out_1_26; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9654 = _T_9653 | _T_9426; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_27; // @[Reg.scala 27:20]
  wire  _T_9428 = _T_4698 & ic_tag_valid_out_1_27; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9655 = _T_9654 | _T_9428; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_28; // @[Reg.scala 27:20]
  wire  _T_9430 = _T_4699 & ic_tag_valid_out_1_28; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9656 = _T_9655 | _T_9430; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_29; // @[Reg.scala 27:20]
  wire  _T_9432 = _T_4700 & ic_tag_valid_out_1_29; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9657 = _T_9656 | _T_9432; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_30; // @[Reg.scala 27:20]
  wire  _T_9434 = _T_4701 & ic_tag_valid_out_1_30; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9658 = _T_9657 | _T_9434; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_31; // @[Reg.scala 27:20]
  wire  _T_9436 = _T_4702 & ic_tag_valid_out_1_31; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9659 = _T_9658 | _T_9436; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_32; // @[Reg.scala 27:20]
  wire  _T_9438 = _T_4703 & ic_tag_valid_out_1_32; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9660 = _T_9659 | _T_9438; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_33; // @[Reg.scala 27:20]
  wire  _T_9440 = _T_4704 & ic_tag_valid_out_1_33; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9661 = _T_9660 | _T_9440; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_34; // @[Reg.scala 27:20]
  wire  _T_9442 = _T_4705 & ic_tag_valid_out_1_34; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9662 = _T_9661 | _T_9442; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_35; // @[Reg.scala 27:20]
  wire  _T_9444 = _T_4706 & ic_tag_valid_out_1_35; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9663 = _T_9662 | _T_9444; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_36; // @[Reg.scala 27:20]
  wire  _T_9446 = _T_4707 & ic_tag_valid_out_1_36; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9664 = _T_9663 | _T_9446; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_37; // @[Reg.scala 27:20]
  wire  _T_9448 = _T_4708 & ic_tag_valid_out_1_37; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9665 = _T_9664 | _T_9448; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_38; // @[Reg.scala 27:20]
  wire  _T_9450 = _T_4709 & ic_tag_valid_out_1_38; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9666 = _T_9665 | _T_9450; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_39; // @[Reg.scala 27:20]
  wire  _T_9452 = _T_4710 & ic_tag_valid_out_1_39; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9667 = _T_9666 | _T_9452; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_40; // @[Reg.scala 27:20]
  wire  _T_9454 = _T_4711 & ic_tag_valid_out_1_40; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9668 = _T_9667 | _T_9454; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_41; // @[Reg.scala 27:20]
  wire  _T_9456 = _T_4712 & ic_tag_valid_out_1_41; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9669 = _T_9668 | _T_9456; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_42; // @[Reg.scala 27:20]
  wire  _T_9458 = _T_4713 & ic_tag_valid_out_1_42; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9670 = _T_9669 | _T_9458; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_43; // @[Reg.scala 27:20]
  wire  _T_9460 = _T_4714 & ic_tag_valid_out_1_43; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9671 = _T_9670 | _T_9460; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_44; // @[Reg.scala 27:20]
  wire  _T_9462 = _T_4715 & ic_tag_valid_out_1_44; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9672 = _T_9671 | _T_9462; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_45; // @[Reg.scala 27:20]
  wire  _T_9464 = _T_4716 & ic_tag_valid_out_1_45; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9673 = _T_9672 | _T_9464; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_46; // @[Reg.scala 27:20]
  wire  _T_9466 = _T_4717 & ic_tag_valid_out_1_46; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9674 = _T_9673 | _T_9466; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_47; // @[Reg.scala 27:20]
  wire  _T_9468 = _T_4718 & ic_tag_valid_out_1_47; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9675 = _T_9674 | _T_9468; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_48; // @[Reg.scala 27:20]
  wire  _T_9470 = _T_4719 & ic_tag_valid_out_1_48; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9676 = _T_9675 | _T_9470; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_49; // @[Reg.scala 27:20]
  wire  _T_9472 = _T_4720 & ic_tag_valid_out_1_49; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9677 = _T_9676 | _T_9472; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_50; // @[Reg.scala 27:20]
  wire  _T_9474 = _T_4721 & ic_tag_valid_out_1_50; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9678 = _T_9677 | _T_9474; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_51; // @[Reg.scala 27:20]
  wire  _T_9476 = _T_4722 & ic_tag_valid_out_1_51; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9679 = _T_9678 | _T_9476; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_52; // @[Reg.scala 27:20]
  wire  _T_9478 = _T_4723 & ic_tag_valid_out_1_52; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9680 = _T_9679 | _T_9478; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_53; // @[Reg.scala 27:20]
  wire  _T_9480 = _T_4724 & ic_tag_valid_out_1_53; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9681 = _T_9680 | _T_9480; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_54; // @[Reg.scala 27:20]
  wire  _T_9482 = _T_4725 & ic_tag_valid_out_1_54; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9682 = _T_9681 | _T_9482; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_55; // @[Reg.scala 27:20]
  wire  _T_9484 = _T_4726 & ic_tag_valid_out_1_55; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9683 = _T_9682 | _T_9484; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_56; // @[Reg.scala 27:20]
  wire  _T_9486 = _T_4727 & ic_tag_valid_out_1_56; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9684 = _T_9683 | _T_9486; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_57; // @[Reg.scala 27:20]
  wire  _T_9488 = _T_4728 & ic_tag_valid_out_1_57; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9685 = _T_9684 | _T_9488; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_58; // @[Reg.scala 27:20]
  wire  _T_9490 = _T_4729 & ic_tag_valid_out_1_58; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9686 = _T_9685 | _T_9490; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_59; // @[Reg.scala 27:20]
  wire  _T_9492 = _T_4730 & ic_tag_valid_out_1_59; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9687 = _T_9686 | _T_9492; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_60; // @[Reg.scala 27:20]
  wire  _T_9494 = _T_4731 & ic_tag_valid_out_1_60; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9688 = _T_9687 | _T_9494; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_61; // @[Reg.scala 27:20]
  wire  _T_9496 = _T_4732 & ic_tag_valid_out_1_61; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9689 = _T_9688 | _T_9496; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_62; // @[Reg.scala 27:20]
  wire  _T_9498 = _T_4733 & ic_tag_valid_out_1_62; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9690 = _T_9689 | _T_9498; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_63; // @[Reg.scala 27:20]
  wire  _T_9500 = _T_4734 & ic_tag_valid_out_1_63; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9691 = _T_9690 | _T_9500; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_64; // @[Reg.scala 27:20]
  wire  _T_9502 = _T_4735 & ic_tag_valid_out_1_64; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9692 = _T_9691 | _T_9502; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_65; // @[Reg.scala 27:20]
  wire  _T_9504 = _T_4736 & ic_tag_valid_out_1_65; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9693 = _T_9692 | _T_9504; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_66; // @[Reg.scala 27:20]
  wire  _T_9506 = _T_4737 & ic_tag_valid_out_1_66; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9694 = _T_9693 | _T_9506; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_67; // @[Reg.scala 27:20]
  wire  _T_9508 = _T_4738 & ic_tag_valid_out_1_67; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9695 = _T_9694 | _T_9508; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_68; // @[Reg.scala 27:20]
  wire  _T_9510 = _T_4739 & ic_tag_valid_out_1_68; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9696 = _T_9695 | _T_9510; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_69; // @[Reg.scala 27:20]
  wire  _T_9512 = _T_4740 & ic_tag_valid_out_1_69; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9697 = _T_9696 | _T_9512; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_70; // @[Reg.scala 27:20]
  wire  _T_9514 = _T_4741 & ic_tag_valid_out_1_70; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9698 = _T_9697 | _T_9514; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_71; // @[Reg.scala 27:20]
  wire  _T_9516 = _T_4742 & ic_tag_valid_out_1_71; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9699 = _T_9698 | _T_9516; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_72; // @[Reg.scala 27:20]
  wire  _T_9518 = _T_4743 & ic_tag_valid_out_1_72; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9700 = _T_9699 | _T_9518; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_73; // @[Reg.scala 27:20]
  wire  _T_9520 = _T_4744 & ic_tag_valid_out_1_73; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9701 = _T_9700 | _T_9520; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_74; // @[Reg.scala 27:20]
  wire  _T_9522 = _T_4745 & ic_tag_valid_out_1_74; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9702 = _T_9701 | _T_9522; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_75; // @[Reg.scala 27:20]
  wire  _T_9524 = _T_4746 & ic_tag_valid_out_1_75; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9703 = _T_9702 | _T_9524; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_76; // @[Reg.scala 27:20]
  wire  _T_9526 = _T_4747 & ic_tag_valid_out_1_76; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9704 = _T_9703 | _T_9526; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_77; // @[Reg.scala 27:20]
  wire  _T_9528 = _T_4748 & ic_tag_valid_out_1_77; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9705 = _T_9704 | _T_9528; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_78; // @[Reg.scala 27:20]
  wire  _T_9530 = _T_4749 & ic_tag_valid_out_1_78; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9706 = _T_9705 | _T_9530; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_79; // @[Reg.scala 27:20]
  wire  _T_9532 = _T_4750 & ic_tag_valid_out_1_79; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9707 = _T_9706 | _T_9532; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_80; // @[Reg.scala 27:20]
  wire  _T_9534 = _T_4751 & ic_tag_valid_out_1_80; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9708 = _T_9707 | _T_9534; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_81; // @[Reg.scala 27:20]
  wire  _T_9536 = _T_4752 & ic_tag_valid_out_1_81; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9709 = _T_9708 | _T_9536; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_82; // @[Reg.scala 27:20]
  wire  _T_9538 = _T_4753 & ic_tag_valid_out_1_82; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9710 = _T_9709 | _T_9538; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_83; // @[Reg.scala 27:20]
  wire  _T_9540 = _T_4754 & ic_tag_valid_out_1_83; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9711 = _T_9710 | _T_9540; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_84; // @[Reg.scala 27:20]
  wire  _T_9542 = _T_4755 & ic_tag_valid_out_1_84; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9712 = _T_9711 | _T_9542; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_85; // @[Reg.scala 27:20]
  wire  _T_9544 = _T_4756 & ic_tag_valid_out_1_85; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9713 = _T_9712 | _T_9544; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_86; // @[Reg.scala 27:20]
  wire  _T_9546 = _T_4757 & ic_tag_valid_out_1_86; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9714 = _T_9713 | _T_9546; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_87; // @[Reg.scala 27:20]
  wire  _T_9548 = _T_4758 & ic_tag_valid_out_1_87; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9715 = _T_9714 | _T_9548; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_88; // @[Reg.scala 27:20]
  wire  _T_9550 = _T_4759 & ic_tag_valid_out_1_88; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9716 = _T_9715 | _T_9550; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_89; // @[Reg.scala 27:20]
  wire  _T_9552 = _T_4760 & ic_tag_valid_out_1_89; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9717 = _T_9716 | _T_9552; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_90; // @[Reg.scala 27:20]
  wire  _T_9554 = _T_4761 & ic_tag_valid_out_1_90; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9718 = _T_9717 | _T_9554; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_91; // @[Reg.scala 27:20]
  wire  _T_9556 = _T_4762 & ic_tag_valid_out_1_91; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9719 = _T_9718 | _T_9556; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_92; // @[Reg.scala 27:20]
  wire  _T_9558 = _T_4763 & ic_tag_valid_out_1_92; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9720 = _T_9719 | _T_9558; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_93; // @[Reg.scala 27:20]
  wire  _T_9560 = _T_4764 & ic_tag_valid_out_1_93; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9721 = _T_9720 | _T_9560; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_94; // @[Reg.scala 27:20]
  wire  _T_9562 = _T_4765 & ic_tag_valid_out_1_94; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9722 = _T_9721 | _T_9562; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_95; // @[Reg.scala 27:20]
  wire  _T_9564 = _T_4766 & ic_tag_valid_out_1_95; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9723 = _T_9722 | _T_9564; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_96; // @[Reg.scala 27:20]
  wire  _T_9566 = _T_4767 & ic_tag_valid_out_1_96; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9724 = _T_9723 | _T_9566; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_97; // @[Reg.scala 27:20]
  wire  _T_9568 = _T_4768 & ic_tag_valid_out_1_97; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9725 = _T_9724 | _T_9568; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_98; // @[Reg.scala 27:20]
  wire  _T_9570 = _T_4769 & ic_tag_valid_out_1_98; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9726 = _T_9725 | _T_9570; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_99; // @[Reg.scala 27:20]
  wire  _T_9572 = _T_4770 & ic_tag_valid_out_1_99; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9727 = _T_9726 | _T_9572; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_100; // @[Reg.scala 27:20]
  wire  _T_9574 = _T_4771 & ic_tag_valid_out_1_100; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9728 = _T_9727 | _T_9574; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_101; // @[Reg.scala 27:20]
  wire  _T_9576 = _T_4772 & ic_tag_valid_out_1_101; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9729 = _T_9728 | _T_9576; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_102; // @[Reg.scala 27:20]
  wire  _T_9578 = _T_4773 & ic_tag_valid_out_1_102; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9730 = _T_9729 | _T_9578; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_103; // @[Reg.scala 27:20]
  wire  _T_9580 = _T_4774 & ic_tag_valid_out_1_103; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9731 = _T_9730 | _T_9580; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_104; // @[Reg.scala 27:20]
  wire  _T_9582 = _T_4775 & ic_tag_valid_out_1_104; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9732 = _T_9731 | _T_9582; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_105; // @[Reg.scala 27:20]
  wire  _T_9584 = _T_4776 & ic_tag_valid_out_1_105; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9733 = _T_9732 | _T_9584; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_106; // @[Reg.scala 27:20]
  wire  _T_9586 = _T_4777 & ic_tag_valid_out_1_106; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9734 = _T_9733 | _T_9586; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_107; // @[Reg.scala 27:20]
  wire  _T_9588 = _T_4778 & ic_tag_valid_out_1_107; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9735 = _T_9734 | _T_9588; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_108; // @[Reg.scala 27:20]
  wire  _T_9590 = _T_4779 & ic_tag_valid_out_1_108; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9736 = _T_9735 | _T_9590; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_109; // @[Reg.scala 27:20]
  wire  _T_9592 = _T_4780 & ic_tag_valid_out_1_109; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9737 = _T_9736 | _T_9592; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_110; // @[Reg.scala 27:20]
  wire  _T_9594 = _T_4781 & ic_tag_valid_out_1_110; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9738 = _T_9737 | _T_9594; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_111; // @[Reg.scala 27:20]
  wire  _T_9596 = _T_4782 & ic_tag_valid_out_1_111; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9739 = _T_9738 | _T_9596; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_112; // @[Reg.scala 27:20]
  wire  _T_9598 = _T_4783 & ic_tag_valid_out_1_112; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9740 = _T_9739 | _T_9598; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_113; // @[Reg.scala 27:20]
  wire  _T_9600 = _T_4784 & ic_tag_valid_out_1_113; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9741 = _T_9740 | _T_9600; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_114; // @[Reg.scala 27:20]
  wire  _T_9602 = _T_4785 & ic_tag_valid_out_1_114; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9742 = _T_9741 | _T_9602; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_115; // @[Reg.scala 27:20]
  wire  _T_9604 = _T_4786 & ic_tag_valid_out_1_115; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9743 = _T_9742 | _T_9604; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_116; // @[Reg.scala 27:20]
  wire  _T_9606 = _T_4787 & ic_tag_valid_out_1_116; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9744 = _T_9743 | _T_9606; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_117; // @[Reg.scala 27:20]
  wire  _T_9608 = _T_4788 & ic_tag_valid_out_1_117; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9745 = _T_9744 | _T_9608; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_118; // @[Reg.scala 27:20]
  wire  _T_9610 = _T_4789 & ic_tag_valid_out_1_118; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9746 = _T_9745 | _T_9610; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_119; // @[Reg.scala 27:20]
  wire  _T_9612 = _T_4790 & ic_tag_valid_out_1_119; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9747 = _T_9746 | _T_9612; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_120; // @[Reg.scala 27:20]
  wire  _T_9614 = _T_4791 & ic_tag_valid_out_1_120; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9748 = _T_9747 | _T_9614; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_121; // @[Reg.scala 27:20]
  wire  _T_9616 = _T_4792 & ic_tag_valid_out_1_121; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9749 = _T_9748 | _T_9616; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_122; // @[Reg.scala 27:20]
  wire  _T_9618 = _T_4793 & ic_tag_valid_out_1_122; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9750 = _T_9749 | _T_9618; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_123; // @[Reg.scala 27:20]
  wire  _T_9620 = _T_4794 & ic_tag_valid_out_1_123; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9751 = _T_9750 | _T_9620; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_124; // @[Reg.scala 27:20]
  wire  _T_9622 = _T_4795 & ic_tag_valid_out_1_124; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9752 = _T_9751 | _T_9622; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_125; // @[Reg.scala 27:20]
  wire  _T_9624 = _T_4796 & ic_tag_valid_out_1_125; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9753 = _T_9752 | _T_9624; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_126; // @[Reg.scala 27:20]
  wire  _T_9626 = _T_4797 & ic_tag_valid_out_1_126; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9754 = _T_9753 | _T_9626; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_1_127; // @[Reg.scala 27:20]
  wire  _T_9628 = _T_4798 & ic_tag_valid_out_1_127; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9755 = _T_9754 | _T_9628; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_0; // @[Reg.scala 27:20]
  wire  _T_8991 = _T_4671 & ic_tag_valid_out_0_0; // @[ifu_mem_ctl.scala 696:10]
  reg  ic_tag_valid_out_0_1; // @[Reg.scala 27:20]
  wire  _T_8993 = _T_4672 & ic_tag_valid_out_0_1; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9246 = _T_8991 | _T_8993; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_2; // @[Reg.scala 27:20]
  wire  _T_8995 = _T_4673 & ic_tag_valid_out_0_2; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9247 = _T_9246 | _T_8995; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_3; // @[Reg.scala 27:20]
  wire  _T_8997 = _T_4674 & ic_tag_valid_out_0_3; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9248 = _T_9247 | _T_8997; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_4; // @[Reg.scala 27:20]
  wire  _T_8999 = _T_4675 & ic_tag_valid_out_0_4; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9249 = _T_9248 | _T_8999; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_5; // @[Reg.scala 27:20]
  wire  _T_9001 = _T_4676 & ic_tag_valid_out_0_5; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9250 = _T_9249 | _T_9001; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_6; // @[Reg.scala 27:20]
  wire  _T_9003 = _T_4677 & ic_tag_valid_out_0_6; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9251 = _T_9250 | _T_9003; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_7; // @[Reg.scala 27:20]
  wire  _T_9005 = _T_4678 & ic_tag_valid_out_0_7; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9252 = _T_9251 | _T_9005; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_8; // @[Reg.scala 27:20]
  wire  _T_9007 = _T_4679 & ic_tag_valid_out_0_8; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9253 = _T_9252 | _T_9007; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_9; // @[Reg.scala 27:20]
  wire  _T_9009 = _T_4680 & ic_tag_valid_out_0_9; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9254 = _T_9253 | _T_9009; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_10; // @[Reg.scala 27:20]
  wire  _T_9011 = _T_4681 & ic_tag_valid_out_0_10; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9255 = _T_9254 | _T_9011; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_11; // @[Reg.scala 27:20]
  wire  _T_9013 = _T_4682 & ic_tag_valid_out_0_11; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9256 = _T_9255 | _T_9013; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_12; // @[Reg.scala 27:20]
  wire  _T_9015 = _T_4683 & ic_tag_valid_out_0_12; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9257 = _T_9256 | _T_9015; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_13; // @[Reg.scala 27:20]
  wire  _T_9017 = _T_4684 & ic_tag_valid_out_0_13; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9258 = _T_9257 | _T_9017; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_14; // @[Reg.scala 27:20]
  wire  _T_9019 = _T_4685 & ic_tag_valid_out_0_14; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9259 = _T_9258 | _T_9019; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_15; // @[Reg.scala 27:20]
  wire  _T_9021 = _T_4686 & ic_tag_valid_out_0_15; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9260 = _T_9259 | _T_9021; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_16; // @[Reg.scala 27:20]
  wire  _T_9023 = _T_4687 & ic_tag_valid_out_0_16; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9261 = _T_9260 | _T_9023; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_17; // @[Reg.scala 27:20]
  wire  _T_9025 = _T_4688 & ic_tag_valid_out_0_17; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9262 = _T_9261 | _T_9025; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_18; // @[Reg.scala 27:20]
  wire  _T_9027 = _T_4689 & ic_tag_valid_out_0_18; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9263 = _T_9262 | _T_9027; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_19; // @[Reg.scala 27:20]
  wire  _T_9029 = _T_4690 & ic_tag_valid_out_0_19; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9264 = _T_9263 | _T_9029; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_20; // @[Reg.scala 27:20]
  wire  _T_9031 = _T_4691 & ic_tag_valid_out_0_20; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9265 = _T_9264 | _T_9031; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_21; // @[Reg.scala 27:20]
  wire  _T_9033 = _T_4692 & ic_tag_valid_out_0_21; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9266 = _T_9265 | _T_9033; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_22; // @[Reg.scala 27:20]
  wire  _T_9035 = _T_4693 & ic_tag_valid_out_0_22; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9267 = _T_9266 | _T_9035; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_23; // @[Reg.scala 27:20]
  wire  _T_9037 = _T_4694 & ic_tag_valid_out_0_23; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9268 = _T_9267 | _T_9037; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_24; // @[Reg.scala 27:20]
  wire  _T_9039 = _T_4695 & ic_tag_valid_out_0_24; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9269 = _T_9268 | _T_9039; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_25; // @[Reg.scala 27:20]
  wire  _T_9041 = _T_4696 & ic_tag_valid_out_0_25; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9270 = _T_9269 | _T_9041; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_26; // @[Reg.scala 27:20]
  wire  _T_9043 = _T_4697 & ic_tag_valid_out_0_26; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9271 = _T_9270 | _T_9043; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_27; // @[Reg.scala 27:20]
  wire  _T_9045 = _T_4698 & ic_tag_valid_out_0_27; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9272 = _T_9271 | _T_9045; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_28; // @[Reg.scala 27:20]
  wire  _T_9047 = _T_4699 & ic_tag_valid_out_0_28; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9273 = _T_9272 | _T_9047; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_29; // @[Reg.scala 27:20]
  wire  _T_9049 = _T_4700 & ic_tag_valid_out_0_29; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9274 = _T_9273 | _T_9049; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_30; // @[Reg.scala 27:20]
  wire  _T_9051 = _T_4701 & ic_tag_valid_out_0_30; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9275 = _T_9274 | _T_9051; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_31; // @[Reg.scala 27:20]
  wire  _T_9053 = _T_4702 & ic_tag_valid_out_0_31; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9276 = _T_9275 | _T_9053; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_32; // @[Reg.scala 27:20]
  wire  _T_9055 = _T_4703 & ic_tag_valid_out_0_32; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9277 = _T_9276 | _T_9055; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_33; // @[Reg.scala 27:20]
  wire  _T_9057 = _T_4704 & ic_tag_valid_out_0_33; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9278 = _T_9277 | _T_9057; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_34; // @[Reg.scala 27:20]
  wire  _T_9059 = _T_4705 & ic_tag_valid_out_0_34; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9279 = _T_9278 | _T_9059; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_35; // @[Reg.scala 27:20]
  wire  _T_9061 = _T_4706 & ic_tag_valid_out_0_35; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9280 = _T_9279 | _T_9061; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_36; // @[Reg.scala 27:20]
  wire  _T_9063 = _T_4707 & ic_tag_valid_out_0_36; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9281 = _T_9280 | _T_9063; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_37; // @[Reg.scala 27:20]
  wire  _T_9065 = _T_4708 & ic_tag_valid_out_0_37; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9282 = _T_9281 | _T_9065; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_38; // @[Reg.scala 27:20]
  wire  _T_9067 = _T_4709 & ic_tag_valid_out_0_38; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9283 = _T_9282 | _T_9067; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_39; // @[Reg.scala 27:20]
  wire  _T_9069 = _T_4710 & ic_tag_valid_out_0_39; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9284 = _T_9283 | _T_9069; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_40; // @[Reg.scala 27:20]
  wire  _T_9071 = _T_4711 & ic_tag_valid_out_0_40; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9285 = _T_9284 | _T_9071; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_41; // @[Reg.scala 27:20]
  wire  _T_9073 = _T_4712 & ic_tag_valid_out_0_41; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9286 = _T_9285 | _T_9073; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_42; // @[Reg.scala 27:20]
  wire  _T_9075 = _T_4713 & ic_tag_valid_out_0_42; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9287 = _T_9286 | _T_9075; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_43; // @[Reg.scala 27:20]
  wire  _T_9077 = _T_4714 & ic_tag_valid_out_0_43; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9288 = _T_9287 | _T_9077; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_44; // @[Reg.scala 27:20]
  wire  _T_9079 = _T_4715 & ic_tag_valid_out_0_44; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9289 = _T_9288 | _T_9079; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_45; // @[Reg.scala 27:20]
  wire  _T_9081 = _T_4716 & ic_tag_valid_out_0_45; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9290 = _T_9289 | _T_9081; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_46; // @[Reg.scala 27:20]
  wire  _T_9083 = _T_4717 & ic_tag_valid_out_0_46; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9291 = _T_9290 | _T_9083; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_47; // @[Reg.scala 27:20]
  wire  _T_9085 = _T_4718 & ic_tag_valid_out_0_47; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9292 = _T_9291 | _T_9085; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_48; // @[Reg.scala 27:20]
  wire  _T_9087 = _T_4719 & ic_tag_valid_out_0_48; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9293 = _T_9292 | _T_9087; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_49; // @[Reg.scala 27:20]
  wire  _T_9089 = _T_4720 & ic_tag_valid_out_0_49; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9294 = _T_9293 | _T_9089; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_50; // @[Reg.scala 27:20]
  wire  _T_9091 = _T_4721 & ic_tag_valid_out_0_50; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9295 = _T_9294 | _T_9091; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_51; // @[Reg.scala 27:20]
  wire  _T_9093 = _T_4722 & ic_tag_valid_out_0_51; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9296 = _T_9295 | _T_9093; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_52; // @[Reg.scala 27:20]
  wire  _T_9095 = _T_4723 & ic_tag_valid_out_0_52; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9297 = _T_9296 | _T_9095; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_53; // @[Reg.scala 27:20]
  wire  _T_9097 = _T_4724 & ic_tag_valid_out_0_53; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9298 = _T_9297 | _T_9097; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_54; // @[Reg.scala 27:20]
  wire  _T_9099 = _T_4725 & ic_tag_valid_out_0_54; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9299 = _T_9298 | _T_9099; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_55; // @[Reg.scala 27:20]
  wire  _T_9101 = _T_4726 & ic_tag_valid_out_0_55; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9300 = _T_9299 | _T_9101; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_56; // @[Reg.scala 27:20]
  wire  _T_9103 = _T_4727 & ic_tag_valid_out_0_56; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9301 = _T_9300 | _T_9103; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_57; // @[Reg.scala 27:20]
  wire  _T_9105 = _T_4728 & ic_tag_valid_out_0_57; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9302 = _T_9301 | _T_9105; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_58; // @[Reg.scala 27:20]
  wire  _T_9107 = _T_4729 & ic_tag_valid_out_0_58; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9303 = _T_9302 | _T_9107; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_59; // @[Reg.scala 27:20]
  wire  _T_9109 = _T_4730 & ic_tag_valid_out_0_59; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9304 = _T_9303 | _T_9109; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_60; // @[Reg.scala 27:20]
  wire  _T_9111 = _T_4731 & ic_tag_valid_out_0_60; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9305 = _T_9304 | _T_9111; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_61; // @[Reg.scala 27:20]
  wire  _T_9113 = _T_4732 & ic_tag_valid_out_0_61; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9306 = _T_9305 | _T_9113; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_62; // @[Reg.scala 27:20]
  wire  _T_9115 = _T_4733 & ic_tag_valid_out_0_62; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9307 = _T_9306 | _T_9115; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_63; // @[Reg.scala 27:20]
  wire  _T_9117 = _T_4734 & ic_tag_valid_out_0_63; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9308 = _T_9307 | _T_9117; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_64; // @[Reg.scala 27:20]
  wire  _T_9119 = _T_4735 & ic_tag_valid_out_0_64; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9309 = _T_9308 | _T_9119; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_65; // @[Reg.scala 27:20]
  wire  _T_9121 = _T_4736 & ic_tag_valid_out_0_65; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9310 = _T_9309 | _T_9121; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_66; // @[Reg.scala 27:20]
  wire  _T_9123 = _T_4737 & ic_tag_valid_out_0_66; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9311 = _T_9310 | _T_9123; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_67; // @[Reg.scala 27:20]
  wire  _T_9125 = _T_4738 & ic_tag_valid_out_0_67; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9312 = _T_9311 | _T_9125; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_68; // @[Reg.scala 27:20]
  wire  _T_9127 = _T_4739 & ic_tag_valid_out_0_68; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9313 = _T_9312 | _T_9127; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_69; // @[Reg.scala 27:20]
  wire  _T_9129 = _T_4740 & ic_tag_valid_out_0_69; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9314 = _T_9313 | _T_9129; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_70; // @[Reg.scala 27:20]
  wire  _T_9131 = _T_4741 & ic_tag_valid_out_0_70; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9315 = _T_9314 | _T_9131; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_71; // @[Reg.scala 27:20]
  wire  _T_9133 = _T_4742 & ic_tag_valid_out_0_71; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9316 = _T_9315 | _T_9133; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_72; // @[Reg.scala 27:20]
  wire  _T_9135 = _T_4743 & ic_tag_valid_out_0_72; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9317 = _T_9316 | _T_9135; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_73; // @[Reg.scala 27:20]
  wire  _T_9137 = _T_4744 & ic_tag_valid_out_0_73; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9318 = _T_9317 | _T_9137; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_74; // @[Reg.scala 27:20]
  wire  _T_9139 = _T_4745 & ic_tag_valid_out_0_74; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9319 = _T_9318 | _T_9139; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_75; // @[Reg.scala 27:20]
  wire  _T_9141 = _T_4746 & ic_tag_valid_out_0_75; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9320 = _T_9319 | _T_9141; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_76; // @[Reg.scala 27:20]
  wire  _T_9143 = _T_4747 & ic_tag_valid_out_0_76; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9321 = _T_9320 | _T_9143; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_77; // @[Reg.scala 27:20]
  wire  _T_9145 = _T_4748 & ic_tag_valid_out_0_77; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9322 = _T_9321 | _T_9145; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_78; // @[Reg.scala 27:20]
  wire  _T_9147 = _T_4749 & ic_tag_valid_out_0_78; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9323 = _T_9322 | _T_9147; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_79; // @[Reg.scala 27:20]
  wire  _T_9149 = _T_4750 & ic_tag_valid_out_0_79; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9324 = _T_9323 | _T_9149; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_80; // @[Reg.scala 27:20]
  wire  _T_9151 = _T_4751 & ic_tag_valid_out_0_80; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9325 = _T_9324 | _T_9151; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_81; // @[Reg.scala 27:20]
  wire  _T_9153 = _T_4752 & ic_tag_valid_out_0_81; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9326 = _T_9325 | _T_9153; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_82; // @[Reg.scala 27:20]
  wire  _T_9155 = _T_4753 & ic_tag_valid_out_0_82; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9327 = _T_9326 | _T_9155; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_83; // @[Reg.scala 27:20]
  wire  _T_9157 = _T_4754 & ic_tag_valid_out_0_83; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9328 = _T_9327 | _T_9157; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_84; // @[Reg.scala 27:20]
  wire  _T_9159 = _T_4755 & ic_tag_valid_out_0_84; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9329 = _T_9328 | _T_9159; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_85; // @[Reg.scala 27:20]
  wire  _T_9161 = _T_4756 & ic_tag_valid_out_0_85; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9330 = _T_9329 | _T_9161; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_86; // @[Reg.scala 27:20]
  wire  _T_9163 = _T_4757 & ic_tag_valid_out_0_86; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9331 = _T_9330 | _T_9163; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_87; // @[Reg.scala 27:20]
  wire  _T_9165 = _T_4758 & ic_tag_valid_out_0_87; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9332 = _T_9331 | _T_9165; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_88; // @[Reg.scala 27:20]
  wire  _T_9167 = _T_4759 & ic_tag_valid_out_0_88; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9333 = _T_9332 | _T_9167; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_89; // @[Reg.scala 27:20]
  wire  _T_9169 = _T_4760 & ic_tag_valid_out_0_89; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9334 = _T_9333 | _T_9169; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_90; // @[Reg.scala 27:20]
  wire  _T_9171 = _T_4761 & ic_tag_valid_out_0_90; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9335 = _T_9334 | _T_9171; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_91; // @[Reg.scala 27:20]
  wire  _T_9173 = _T_4762 & ic_tag_valid_out_0_91; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9336 = _T_9335 | _T_9173; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_92; // @[Reg.scala 27:20]
  wire  _T_9175 = _T_4763 & ic_tag_valid_out_0_92; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9337 = _T_9336 | _T_9175; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_93; // @[Reg.scala 27:20]
  wire  _T_9177 = _T_4764 & ic_tag_valid_out_0_93; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9338 = _T_9337 | _T_9177; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_94; // @[Reg.scala 27:20]
  wire  _T_9179 = _T_4765 & ic_tag_valid_out_0_94; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9339 = _T_9338 | _T_9179; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_95; // @[Reg.scala 27:20]
  wire  _T_9181 = _T_4766 & ic_tag_valid_out_0_95; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9340 = _T_9339 | _T_9181; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_96; // @[Reg.scala 27:20]
  wire  _T_9183 = _T_4767 & ic_tag_valid_out_0_96; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9341 = _T_9340 | _T_9183; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_97; // @[Reg.scala 27:20]
  wire  _T_9185 = _T_4768 & ic_tag_valid_out_0_97; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9342 = _T_9341 | _T_9185; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_98; // @[Reg.scala 27:20]
  wire  _T_9187 = _T_4769 & ic_tag_valid_out_0_98; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9343 = _T_9342 | _T_9187; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_99; // @[Reg.scala 27:20]
  wire  _T_9189 = _T_4770 & ic_tag_valid_out_0_99; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9344 = _T_9343 | _T_9189; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_100; // @[Reg.scala 27:20]
  wire  _T_9191 = _T_4771 & ic_tag_valid_out_0_100; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9345 = _T_9344 | _T_9191; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_101; // @[Reg.scala 27:20]
  wire  _T_9193 = _T_4772 & ic_tag_valid_out_0_101; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9346 = _T_9345 | _T_9193; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_102; // @[Reg.scala 27:20]
  wire  _T_9195 = _T_4773 & ic_tag_valid_out_0_102; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9347 = _T_9346 | _T_9195; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_103; // @[Reg.scala 27:20]
  wire  _T_9197 = _T_4774 & ic_tag_valid_out_0_103; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9348 = _T_9347 | _T_9197; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_104; // @[Reg.scala 27:20]
  wire  _T_9199 = _T_4775 & ic_tag_valid_out_0_104; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9349 = _T_9348 | _T_9199; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_105; // @[Reg.scala 27:20]
  wire  _T_9201 = _T_4776 & ic_tag_valid_out_0_105; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9350 = _T_9349 | _T_9201; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_106; // @[Reg.scala 27:20]
  wire  _T_9203 = _T_4777 & ic_tag_valid_out_0_106; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9351 = _T_9350 | _T_9203; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_107; // @[Reg.scala 27:20]
  wire  _T_9205 = _T_4778 & ic_tag_valid_out_0_107; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9352 = _T_9351 | _T_9205; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_108; // @[Reg.scala 27:20]
  wire  _T_9207 = _T_4779 & ic_tag_valid_out_0_108; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9353 = _T_9352 | _T_9207; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_109; // @[Reg.scala 27:20]
  wire  _T_9209 = _T_4780 & ic_tag_valid_out_0_109; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9354 = _T_9353 | _T_9209; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_110; // @[Reg.scala 27:20]
  wire  _T_9211 = _T_4781 & ic_tag_valid_out_0_110; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9355 = _T_9354 | _T_9211; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_111; // @[Reg.scala 27:20]
  wire  _T_9213 = _T_4782 & ic_tag_valid_out_0_111; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9356 = _T_9355 | _T_9213; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_112; // @[Reg.scala 27:20]
  wire  _T_9215 = _T_4783 & ic_tag_valid_out_0_112; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9357 = _T_9356 | _T_9215; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_113; // @[Reg.scala 27:20]
  wire  _T_9217 = _T_4784 & ic_tag_valid_out_0_113; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9358 = _T_9357 | _T_9217; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_114; // @[Reg.scala 27:20]
  wire  _T_9219 = _T_4785 & ic_tag_valid_out_0_114; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9359 = _T_9358 | _T_9219; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_115; // @[Reg.scala 27:20]
  wire  _T_9221 = _T_4786 & ic_tag_valid_out_0_115; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9360 = _T_9359 | _T_9221; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_116; // @[Reg.scala 27:20]
  wire  _T_9223 = _T_4787 & ic_tag_valid_out_0_116; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9361 = _T_9360 | _T_9223; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_117; // @[Reg.scala 27:20]
  wire  _T_9225 = _T_4788 & ic_tag_valid_out_0_117; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9362 = _T_9361 | _T_9225; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_118; // @[Reg.scala 27:20]
  wire  _T_9227 = _T_4789 & ic_tag_valid_out_0_118; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9363 = _T_9362 | _T_9227; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_119; // @[Reg.scala 27:20]
  wire  _T_9229 = _T_4790 & ic_tag_valid_out_0_119; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9364 = _T_9363 | _T_9229; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_120; // @[Reg.scala 27:20]
  wire  _T_9231 = _T_4791 & ic_tag_valid_out_0_120; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9365 = _T_9364 | _T_9231; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_121; // @[Reg.scala 27:20]
  wire  _T_9233 = _T_4792 & ic_tag_valid_out_0_121; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9366 = _T_9365 | _T_9233; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_122; // @[Reg.scala 27:20]
  wire  _T_9235 = _T_4793 & ic_tag_valid_out_0_122; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9367 = _T_9366 | _T_9235; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_123; // @[Reg.scala 27:20]
  wire  _T_9237 = _T_4794 & ic_tag_valid_out_0_123; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9368 = _T_9367 | _T_9237; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_124; // @[Reg.scala 27:20]
  wire  _T_9239 = _T_4795 & ic_tag_valid_out_0_124; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9369 = _T_9368 | _T_9239; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_125; // @[Reg.scala 27:20]
  wire  _T_9241 = _T_4796 & ic_tag_valid_out_0_125; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9370 = _T_9369 | _T_9241; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_126; // @[Reg.scala 27:20]
  wire  _T_9243 = _T_4797 & ic_tag_valid_out_0_126; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9371 = _T_9370 | _T_9243; // @[ifu_mem_ctl.scala 696:91]
  reg  ic_tag_valid_out_0_127; // @[Reg.scala 27:20]
  wire  _T_9245 = _T_4798 & ic_tag_valid_out_0_127; // @[ifu_mem_ctl.scala 696:10]
  wire  _T_9372 = _T_9371 | _T_9245; // @[ifu_mem_ctl.scala 696:91]
  wire [1:0] ic_tag_valid_unq = {_T_9755,_T_9372}; // @[Cat.scala 29:58]
  reg [1:0] ic_debug_way_ff; // @[ifu_mem_ctl.scala 767:53]
  reg  ic_debug_rd_en_ff; // @[ifu_mem_ctl.scala 769:54]
  wire [1:0] _T_9795 = ic_debug_rd_en_ff ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [1:0] _T_9796 = ic_debug_way_ff & _T_9795; // @[ifu_mem_ctl.scala 750:67]
  wire [1:0] _T_9797 = ic_tag_valid_unq & _T_9796; // @[ifu_mem_ctl.scala 750:48]
  wire  ic_debug_tag_val_rd_out = |_T_9797; // @[ifu_mem_ctl.scala 750:115]
  wire [70:0] _T_1211 = {2'h0,io_ic_tag_debug_rd_data[25:21],32'h0,io_ic_tag_debug_rd_data[20:0],6'h0,way_status,3'h0,ic_debug_tag_val_rd_out}; // @[Cat.scala 29:58]
  reg [70:0] _T_1212; // @[ifu_mem_ctl.scala 263:76]
  wire  _T_1250 = ~ifu_byp_data_err_new; // @[ifu_mem_ctl.scala 279:98]
  wire  sel_byp_data = _T_1254 & _T_1250; // @[ifu_mem_ctl.scala 279:96]
  wire  _T_1257 = sel_byp_data | fetch_req_iccm_f; // @[ifu_mem_ctl.scala 284:46]
  wire  final_data_sel1_0 = _T_1257 | sel_ic_data; // @[ifu_mem_ctl.scala 284:62]
  wire [63:0] _T_1263 = final_data_sel1_0 ? 64'hffffffffffffffff : 64'h0; // @[Bitwise.scala 72:12]
  wire [63:0] ic_final_data = _T_1263 & io_ic_rd_data; // @[ifu_mem_ctl.scala 288:92]
  wire [63:0] _T_1265 = fetch_req_iccm_f ? 64'hffffffffffffffff : 64'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_1266 = _T_1265 & io_iccm_rd_data; // @[ifu_mem_ctl.scala 292:69]
  wire [63:0] _T_1268 = sel_byp_data ? 64'hffffffffffffffff : 64'h0; // @[Bitwise.scala 72:12]
  wire [3:0] byp_fetch_index_inc_0 = {byp_fetch_index_inc,1'h0}; // @[Cat.scala 29:58]
  wire  _T_1662 = byp_fetch_index_inc_0 == 4'h0; // @[ifu_mem_ctl.scala 358:73]
  wire [15:0] _T_1710 = _T_1662 ? ic_miss_buff_data_0[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire  _T_1665 = byp_fetch_index_inc_0 == 4'h1; // @[ifu_mem_ctl.scala 358:73]
  wire [15:0] _T_1711 = _T_1665 ? ic_miss_buff_data_1[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1726 = _T_1710 | _T_1711; // @[Mux.scala 27:72]
  wire  _T_1668 = byp_fetch_index_inc_0 == 4'h2; // @[ifu_mem_ctl.scala 358:73]
  wire [15:0] _T_1712 = _T_1668 ? ic_miss_buff_data_2[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1727 = _T_1726 | _T_1712; // @[Mux.scala 27:72]
  wire  _T_1671 = byp_fetch_index_inc_0 == 4'h3; // @[ifu_mem_ctl.scala 358:73]
  wire [15:0] _T_1713 = _T_1671 ? ic_miss_buff_data_3[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1728 = _T_1727 | _T_1713; // @[Mux.scala 27:72]
  wire  _T_1674 = byp_fetch_index_inc_0 == 4'h4; // @[ifu_mem_ctl.scala 358:73]
  wire [15:0] _T_1714 = _T_1674 ? ic_miss_buff_data_4[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1729 = _T_1728 | _T_1714; // @[Mux.scala 27:72]
  wire  _T_1677 = byp_fetch_index_inc_0 == 4'h5; // @[ifu_mem_ctl.scala 358:73]
  wire [15:0] _T_1715 = _T_1677 ? ic_miss_buff_data_5[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1730 = _T_1729 | _T_1715; // @[Mux.scala 27:72]
  wire  _T_1680 = byp_fetch_index_inc_0 == 4'h6; // @[ifu_mem_ctl.scala 358:73]
  wire [15:0] _T_1716 = _T_1680 ? ic_miss_buff_data_6[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1731 = _T_1730 | _T_1716; // @[Mux.scala 27:72]
  wire  _T_1683 = byp_fetch_index_inc_0 == 4'h7; // @[ifu_mem_ctl.scala 358:73]
  wire [15:0] _T_1717 = _T_1683 ? ic_miss_buff_data_7[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1732 = _T_1731 | _T_1717; // @[Mux.scala 27:72]
  wire  _T_1686 = byp_fetch_index_inc_0 == 4'h8; // @[ifu_mem_ctl.scala 358:73]
  wire [15:0] _T_1718 = _T_1686 ? ic_miss_buff_data_8[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1733 = _T_1732 | _T_1718; // @[Mux.scala 27:72]
  wire  _T_1689 = byp_fetch_index_inc_0 == 4'h9; // @[ifu_mem_ctl.scala 358:73]
  wire [15:0] _T_1719 = _T_1689 ? ic_miss_buff_data_9[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1734 = _T_1733 | _T_1719; // @[Mux.scala 27:72]
  wire  _T_1692 = byp_fetch_index_inc_0 == 4'ha; // @[ifu_mem_ctl.scala 358:73]
  wire [15:0] _T_1720 = _T_1692 ? ic_miss_buff_data_10[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1735 = _T_1734 | _T_1720; // @[Mux.scala 27:72]
  wire  _T_1695 = byp_fetch_index_inc_0 == 4'hb; // @[ifu_mem_ctl.scala 358:73]
  wire [15:0] _T_1721 = _T_1695 ? ic_miss_buff_data_11[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1736 = _T_1735 | _T_1721; // @[Mux.scala 27:72]
  wire  _T_1698 = byp_fetch_index_inc_0 == 4'hc; // @[ifu_mem_ctl.scala 358:73]
  wire [15:0] _T_1722 = _T_1698 ? ic_miss_buff_data_12[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1737 = _T_1736 | _T_1722; // @[Mux.scala 27:72]
  wire  _T_1701 = byp_fetch_index_inc_0 == 4'hd; // @[ifu_mem_ctl.scala 358:73]
  wire [15:0] _T_1723 = _T_1701 ? ic_miss_buff_data_13[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1738 = _T_1737 | _T_1723; // @[Mux.scala 27:72]
  wire  _T_1704 = byp_fetch_index_inc_0 == 4'he; // @[ifu_mem_ctl.scala 358:73]
  wire [15:0] _T_1724 = _T_1704 ? ic_miss_buff_data_14[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1739 = _T_1738 | _T_1724; // @[Mux.scala 27:72]
  wire  _T_1707 = byp_fetch_index_inc_0 == 4'hf; // @[ifu_mem_ctl.scala 358:73]
  wire [15:0] _T_1725 = _T_1707 ? ic_miss_buff_data_15[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1740 = _T_1739 | _T_1725; // @[Mux.scala 27:72]
  wire [3:0] byp_fetch_index_1 = {ifu_fetch_addr_int_f[4:2],1'h1}; // @[Cat.scala 29:58]
  wire  _T_1742 = byp_fetch_index_1 == 4'h0; // @[ifu_mem_ctl.scala 358:179]
  wire [31:0] _T_1790 = _T_1742 ? ic_miss_buff_data_0 : 32'h0; // @[Mux.scala 27:72]
  wire  _T_1745 = byp_fetch_index_1 == 4'h1; // @[ifu_mem_ctl.scala 358:179]
  wire [31:0] _T_1791 = _T_1745 ? ic_miss_buff_data_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1806 = _T_1790 | _T_1791; // @[Mux.scala 27:72]
  wire  _T_1748 = byp_fetch_index_1 == 4'h2; // @[ifu_mem_ctl.scala 358:179]
  wire [31:0] _T_1792 = _T_1748 ? ic_miss_buff_data_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1807 = _T_1806 | _T_1792; // @[Mux.scala 27:72]
  wire  _T_1751 = byp_fetch_index_1 == 4'h3; // @[ifu_mem_ctl.scala 358:179]
  wire [31:0] _T_1793 = _T_1751 ? ic_miss_buff_data_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1808 = _T_1807 | _T_1793; // @[Mux.scala 27:72]
  wire  _T_1754 = byp_fetch_index_1 == 4'h4; // @[ifu_mem_ctl.scala 358:179]
  wire [31:0] _T_1794 = _T_1754 ? ic_miss_buff_data_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1809 = _T_1808 | _T_1794; // @[Mux.scala 27:72]
  wire  _T_1757 = byp_fetch_index_1 == 4'h5; // @[ifu_mem_ctl.scala 358:179]
  wire [31:0] _T_1795 = _T_1757 ? ic_miss_buff_data_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1810 = _T_1809 | _T_1795; // @[Mux.scala 27:72]
  wire  _T_1760 = byp_fetch_index_1 == 4'h6; // @[ifu_mem_ctl.scala 358:179]
  wire [31:0] _T_1796 = _T_1760 ? ic_miss_buff_data_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1811 = _T_1810 | _T_1796; // @[Mux.scala 27:72]
  wire  _T_1763 = byp_fetch_index_1 == 4'h7; // @[ifu_mem_ctl.scala 358:179]
  wire [31:0] _T_1797 = _T_1763 ? ic_miss_buff_data_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1812 = _T_1811 | _T_1797; // @[Mux.scala 27:72]
  wire  _T_1766 = byp_fetch_index_1 == 4'h8; // @[ifu_mem_ctl.scala 358:179]
  wire [31:0] _T_1798 = _T_1766 ? ic_miss_buff_data_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1813 = _T_1812 | _T_1798; // @[Mux.scala 27:72]
  wire  _T_1769 = byp_fetch_index_1 == 4'h9; // @[ifu_mem_ctl.scala 358:179]
  wire [31:0] _T_1799 = _T_1769 ? ic_miss_buff_data_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1814 = _T_1813 | _T_1799; // @[Mux.scala 27:72]
  wire  _T_1772 = byp_fetch_index_1 == 4'ha; // @[ifu_mem_ctl.scala 358:179]
  wire [31:0] _T_1800 = _T_1772 ? ic_miss_buff_data_10 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1815 = _T_1814 | _T_1800; // @[Mux.scala 27:72]
  wire  _T_1775 = byp_fetch_index_1 == 4'hb; // @[ifu_mem_ctl.scala 358:179]
  wire [31:0] _T_1801 = _T_1775 ? ic_miss_buff_data_11 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1816 = _T_1815 | _T_1801; // @[Mux.scala 27:72]
  wire  _T_1778 = byp_fetch_index_1 == 4'hc; // @[ifu_mem_ctl.scala 358:179]
  wire [31:0] _T_1802 = _T_1778 ? ic_miss_buff_data_12 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1817 = _T_1816 | _T_1802; // @[Mux.scala 27:72]
  wire  _T_1781 = byp_fetch_index_1 == 4'hd; // @[ifu_mem_ctl.scala 358:179]
  wire [31:0] _T_1803 = _T_1781 ? ic_miss_buff_data_13 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1818 = _T_1817 | _T_1803; // @[Mux.scala 27:72]
  wire  _T_1784 = byp_fetch_index_1 == 4'he; // @[ifu_mem_ctl.scala 358:179]
  wire [31:0] _T_1804 = _T_1784 ? ic_miss_buff_data_14 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1819 = _T_1818 | _T_1804; // @[Mux.scala 27:72]
  wire  _T_1787 = byp_fetch_index_1 == 4'hf; // @[ifu_mem_ctl.scala 358:179]
  wire [31:0] _T_1805 = _T_1787 ? ic_miss_buff_data_15 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1820 = _T_1819 | _T_1805; // @[Mux.scala 27:72]
  wire [3:0] byp_fetch_index_0 = {ifu_fetch_addr_int_f[4:2],1'h0}; // @[Cat.scala 29:58]
  wire  _T_1822 = byp_fetch_index_0 == 4'h0; // @[ifu_mem_ctl.scala 358:285]
  wire [31:0] _T_1870 = _T_1822 ? ic_miss_buff_data_0 : 32'h0; // @[Mux.scala 27:72]
  wire  _T_1825 = byp_fetch_index_0 == 4'h1; // @[ifu_mem_ctl.scala 358:285]
  wire [31:0] _T_1871 = _T_1825 ? ic_miss_buff_data_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1886 = _T_1870 | _T_1871; // @[Mux.scala 27:72]
  wire  _T_1828 = byp_fetch_index_0 == 4'h2; // @[ifu_mem_ctl.scala 358:285]
  wire [31:0] _T_1872 = _T_1828 ? ic_miss_buff_data_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1887 = _T_1886 | _T_1872; // @[Mux.scala 27:72]
  wire  _T_1831 = byp_fetch_index_0 == 4'h3; // @[ifu_mem_ctl.scala 358:285]
  wire [31:0] _T_1873 = _T_1831 ? ic_miss_buff_data_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1888 = _T_1887 | _T_1873; // @[Mux.scala 27:72]
  wire  _T_1834 = byp_fetch_index_0 == 4'h4; // @[ifu_mem_ctl.scala 358:285]
  wire [31:0] _T_1874 = _T_1834 ? ic_miss_buff_data_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1889 = _T_1888 | _T_1874; // @[Mux.scala 27:72]
  wire  _T_1837 = byp_fetch_index_0 == 4'h5; // @[ifu_mem_ctl.scala 358:285]
  wire [31:0] _T_1875 = _T_1837 ? ic_miss_buff_data_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1890 = _T_1889 | _T_1875; // @[Mux.scala 27:72]
  wire  _T_1840 = byp_fetch_index_0 == 4'h6; // @[ifu_mem_ctl.scala 358:285]
  wire [31:0] _T_1876 = _T_1840 ? ic_miss_buff_data_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1891 = _T_1890 | _T_1876; // @[Mux.scala 27:72]
  wire  _T_1843 = byp_fetch_index_0 == 4'h7; // @[ifu_mem_ctl.scala 358:285]
  wire [31:0] _T_1877 = _T_1843 ? ic_miss_buff_data_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1892 = _T_1891 | _T_1877; // @[Mux.scala 27:72]
  wire  _T_1846 = byp_fetch_index_0 == 4'h8; // @[ifu_mem_ctl.scala 358:285]
  wire [31:0] _T_1878 = _T_1846 ? ic_miss_buff_data_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1893 = _T_1892 | _T_1878; // @[Mux.scala 27:72]
  wire  _T_1849 = byp_fetch_index_0 == 4'h9; // @[ifu_mem_ctl.scala 358:285]
  wire [31:0] _T_1879 = _T_1849 ? ic_miss_buff_data_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1894 = _T_1893 | _T_1879; // @[Mux.scala 27:72]
  wire  _T_1852 = byp_fetch_index_0 == 4'ha; // @[ifu_mem_ctl.scala 358:285]
  wire [31:0] _T_1880 = _T_1852 ? ic_miss_buff_data_10 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1895 = _T_1894 | _T_1880; // @[Mux.scala 27:72]
  wire  _T_1855 = byp_fetch_index_0 == 4'hb; // @[ifu_mem_ctl.scala 358:285]
  wire [31:0] _T_1881 = _T_1855 ? ic_miss_buff_data_11 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1896 = _T_1895 | _T_1881; // @[Mux.scala 27:72]
  wire  _T_1858 = byp_fetch_index_0 == 4'hc; // @[ifu_mem_ctl.scala 358:285]
  wire [31:0] _T_1882 = _T_1858 ? ic_miss_buff_data_12 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1897 = _T_1896 | _T_1882; // @[Mux.scala 27:72]
  wire  _T_1861 = byp_fetch_index_0 == 4'hd; // @[ifu_mem_ctl.scala 358:285]
  wire [31:0] _T_1883 = _T_1861 ? ic_miss_buff_data_13 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1898 = _T_1897 | _T_1883; // @[Mux.scala 27:72]
  wire  _T_1864 = byp_fetch_index_0 == 4'he; // @[ifu_mem_ctl.scala 358:285]
  wire [31:0] _T_1884 = _T_1864 ? ic_miss_buff_data_14 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1899 = _T_1898 | _T_1884; // @[Mux.scala 27:72]
  wire  _T_1867 = byp_fetch_index_0 == 4'hf; // @[ifu_mem_ctl.scala 358:285]
  wire [31:0] _T_1885 = _T_1867 ? ic_miss_buff_data_15 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1900 = _T_1899 | _T_1885; // @[Mux.scala 27:72]
  wire [79:0] _T_1903 = {_T_1740,_T_1820,_T_1900}; // @[Cat.scala 29:58]
  wire [3:0] byp_fetch_index_inc_1 = {byp_fetch_index_inc,1'h1}; // @[Cat.scala 29:58]
  wire  _T_1904 = byp_fetch_index_inc_1 == 4'h0; // @[ifu_mem_ctl.scala 359:73]
  wire [15:0] _T_1952 = _T_1904 ? ic_miss_buff_data_0[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire  _T_1907 = byp_fetch_index_inc_1 == 4'h1; // @[ifu_mem_ctl.scala 359:73]
  wire [15:0] _T_1953 = _T_1907 ? ic_miss_buff_data_1[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1968 = _T_1952 | _T_1953; // @[Mux.scala 27:72]
  wire  _T_1910 = byp_fetch_index_inc_1 == 4'h2; // @[ifu_mem_ctl.scala 359:73]
  wire [15:0] _T_1954 = _T_1910 ? ic_miss_buff_data_2[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1969 = _T_1968 | _T_1954; // @[Mux.scala 27:72]
  wire  _T_1913 = byp_fetch_index_inc_1 == 4'h3; // @[ifu_mem_ctl.scala 359:73]
  wire [15:0] _T_1955 = _T_1913 ? ic_miss_buff_data_3[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1970 = _T_1969 | _T_1955; // @[Mux.scala 27:72]
  wire  _T_1916 = byp_fetch_index_inc_1 == 4'h4; // @[ifu_mem_ctl.scala 359:73]
  wire [15:0] _T_1956 = _T_1916 ? ic_miss_buff_data_4[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1971 = _T_1970 | _T_1956; // @[Mux.scala 27:72]
  wire  _T_1919 = byp_fetch_index_inc_1 == 4'h5; // @[ifu_mem_ctl.scala 359:73]
  wire [15:0] _T_1957 = _T_1919 ? ic_miss_buff_data_5[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1972 = _T_1971 | _T_1957; // @[Mux.scala 27:72]
  wire  _T_1922 = byp_fetch_index_inc_1 == 4'h6; // @[ifu_mem_ctl.scala 359:73]
  wire [15:0] _T_1958 = _T_1922 ? ic_miss_buff_data_6[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1973 = _T_1972 | _T_1958; // @[Mux.scala 27:72]
  wire  _T_1925 = byp_fetch_index_inc_1 == 4'h7; // @[ifu_mem_ctl.scala 359:73]
  wire [15:0] _T_1959 = _T_1925 ? ic_miss_buff_data_7[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1974 = _T_1973 | _T_1959; // @[Mux.scala 27:72]
  wire  _T_1928 = byp_fetch_index_inc_1 == 4'h8; // @[ifu_mem_ctl.scala 359:73]
  wire [15:0] _T_1960 = _T_1928 ? ic_miss_buff_data_8[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1975 = _T_1974 | _T_1960; // @[Mux.scala 27:72]
  wire  _T_1931 = byp_fetch_index_inc_1 == 4'h9; // @[ifu_mem_ctl.scala 359:73]
  wire [15:0] _T_1961 = _T_1931 ? ic_miss_buff_data_9[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1976 = _T_1975 | _T_1961; // @[Mux.scala 27:72]
  wire  _T_1934 = byp_fetch_index_inc_1 == 4'ha; // @[ifu_mem_ctl.scala 359:73]
  wire [15:0] _T_1962 = _T_1934 ? ic_miss_buff_data_10[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1977 = _T_1976 | _T_1962; // @[Mux.scala 27:72]
  wire  _T_1937 = byp_fetch_index_inc_1 == 4'hb; // @[ifu_mem_ctl.scala 359:73]
  wire [15:0] _T_1963 = _T_1937 ? ic_miss_buff_data_11[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1978 = _T_1977 | _T_1963; // @[Mux.scala 27:72]
  wire  _T_1940 = byp_fetch_index_inc_1 == 4'hc; // @[ifu_mem_ctl.scala 359:73]
  wire [15:0] _T_1964 = _T_1940 ? ic_miss_buff_data_12[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1979 = _T_1978 | _T_1964; // @[Mux.scala 27:72]
  wire  _T_1943 = byp_fetch_index_inc_1 == 4'hd; // @[ifu_mem_ctl.scala 359:73]
  wire [15:0] _T_1965 = _T_1943 ? ic_miss_buff_data_13[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1980 = _T_1979 | _T_1965; // @[Mux.scala 27:72]
  wire  _T_1946 = byp_fetch_index_inc_1 == 4'he; // @[ifu_mem_ctl.scala 359:73]
  wire [15:0] _T_1966 = _T_1946 ? ic_miss_buff_data_14[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1981 = _T_1980 | _T_1966; // @[Mux.scala 27:72]
  wire  _T_1949 = byp_fetch_index_inc_1 == 4'hf; // @[ifu_mem_ctl.scala 359:73]
  wire [15:0] _T_1967 = _T_1949 ? ic_miss_buff_data_15[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1982 = _T_1981 | _T_1967; // @[Mux.scala 27:72]
  wire [31:0] _T_2032 = _T_1662 ? ic_miss_buff_data_0 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2033 = _T_1665 ? ic_miss_buff_data_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2048 = _T_2032 | _T_2033; // @[Mux.scala 27:72]
  wire [31:0] _T_2034 = _T_1668 ? ic_miss_buff_data_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2049 = _T_2048 | _T_2034; // @[Mux.scala 27:72]
  wire [31:0] _T_2035 = _T_1671 ? ic_miss_buff_data_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2050 = _T_2049 | _T_2035; // @[Mux.scala 27:72]
  wire [31:0] _T_2036 = _T_1674 ? ic_miss_buff_data_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2051 = _T_2050 | _T_2036; // @[Mux.scala 27:72]
  wire [31:0] _T_2037 = _T_1677 ? ic_miss_buff_data_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2052 = _T_2051 | _T_2037; // @[Mux.scala 27:72]
  wire [31:0] _T_2038 = _T_1680 ? ic_miss_buff_data_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2053 = _T_2052 | _T_2038; // @[Mux.scala 27:72]
  wire [31:0] _T_2039 = _T_1683 ? ic_miss_buff_data_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2054 = _T_2053 | _T_2039; // @[Mux.scala 27:72]
  wire [31:0] _T_2040 = _T_1686 ? ic_miss_buff_data_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2055 = _T_2054 | _T_2040; // @[Mux.scala 27:72]
  wire [31:0] _T_2041 = _T_1689 ? ic_miss_buff_data_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2056 = _T_2055 | _T_2041; // @[Mux.scala 27:72]
  wire [31:0] _T_2042 = _T_1692 ? ic_miss_buff_data_10 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2057 = _T_2056 | _T_2042; // @[Mux.scala 27:72]
  wire [31:0] _T_2043 = _T_1695 ? ic_miss_buff_data_11 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2058 = _T_2057 | _T_2043; // @[Mux.scala 27:72]
  wire [31:0] _T_2044 = _T_1698 ? ic_miss_buff_data_12 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2059 = _T_2058 | _T_2044; // @[Mux.scala 27:72]
  wire [31:0] _T_2045 = _T_1701 ? ic_miss_buff_data_13 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2060 = _T_2059 | _T_2045; // @[Mux.scala 27:72]
  wire [31:0] _T_2046 = _T_1704 ? ic_miss_buff_data_14 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2061 = _T_2060 | _T_2046; // @[Mux.scala 27:72]
  wire [31:0] _T_2047 = _T_1707 ? ic_miss_buff_data_15 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2062 = _T_2061 | _T_2047; // @[Mux.scala 27:72]
  wire [79:0] _T_2145 = {_T_1982,_T_2062,_T_1820}; // @[Cat.scala 29:58]
  wire [79:0] ic_byp_data_only_pre_new = _T_1612 ? _T_1903 : _T_2145; // @[ifu_mem_ctl.scala 357:37]
  wire [79:0] _T_2150 = {16'h0,ic_byp_data_only_pre_new[79:16]}; // @[Cat.scala 29:58]
  wire [79:0] ic_byp_data_only_new = _T_1614 ? ic_byp_data_only_pre_new : _T_2150; // @[ifu_mem_ctl.scala 361:30]
  wire [79:0] _GEN_437 = {{16'd0}, _T_1268}; // @[ifu_mem_ctl.scala 292:114]
  wire [79:0] _T_1269 = _GEN_437 & ic_byp_data_only_new; // @[ifu_mem_ctl.scala 292:114]
  wire [79:0] _GEN_438 = {{16'd0}, _T_1266}; // @[ifu_mem_ctl.scala 292:88]
  wire [79:0] ic_premux_data_temp = _GEN_438 | _T_1269; // @[ifu_mem_ctl.scala 292:88]
  wire  fetch_req_f_qual = io_ic_hit_f & _T_319; // @[ifu_mem_ctl.scala 299:38]
  reg  ifc_region_acc_fault_memory_f; // @[ifu_mem_ctl.scala 783:66]
  wire [1:0] _T_1277 = ifc_region_acc_fault_memory_f ? 2'h3 : 2'h0; // @[ifu_mem_ctl.scala 304:10]
  wire [1:0] _T_1278 = ifc_region_acc_fault_f ? 2'h2 : _T_1277; // @[ifu_mem_ctl.scala 303:8]
  wire  _T_1280 = fetch_req_f_qual & io_ifu_bp_inst_mask_f; // @[ifu_mem_ctl.scala 305:45]
  wire  _T_1282 = byp_fetch_index == 5'h1f; // @[ifu_mem_ctl.scala 305:80]
  wire  _T_1283 = ~_T_1282; // @[ifu_mem_ctl.scala 305:71]
  wire  _T_1284 = _T_1280 & _T_1283; // @[ifu_mem_ctl.scala 305:69]
  wire  _T_1285 = err_stop_state != 2'h2; // @[ifu_mem_ctl.scala 305:131]
  wire  _T_1286 = _T_1284 & _T_1285; // @[ifu_mem_ctl.scala 305:114]
  wire [6:0] _T_1358 = {ic_miss_buff_data_valid_in_7,ic_miss_buff_data_valid_in_6,ic_miss_buff_data_valid_in_5,ic_miss_buff_data_valid_in_4,ic_miss_buff_data_valid_in_3,ic_miss_buff_data_valid_in_2,ic_miss_buff_data_valid_in_1}; // @[Cat.scala 29:58]
  wire  _T_1364 = ic_miss_buff_data_error[0] & _T_1330; // @[ifu_mem_ctl.scala 324:32]
  wire  _T_2690 = |io_ifu_axi_r_bits_resp; // @[ifu_mem_ctl.scala 557:47]
  wire  _T_2691 = _T_2690 & _T_13; // @[ifu_mem_ctl.scala 557:50]
  wire  bus_ifu_wr_data_error = _T_2691 & miss_pending; // @[ifu_mem_ctl.scala 557:68]
  wire  ic_miss_buff_data_error_in_0 = write_fill_data_0 ? bus_ifu_wr_data_error : _T_1364; // @[ifu_mem_ctl.scala 323:72]
  wire  _T_1368 = ic_miss_buff_data_error[1] & _T_1330; // @[ifu_mem_ctl.scala 324:32]
  wire  ic_miss_buff_data_error_in_1 = write_fill_data_1 ? bus_ifu_wr_data_error : _T_1368; // @[ifu_mem_ctl.scala 323:72]
  wire  _T_1372 = ic_miss_buff_data_error[2] & _T_1330; // @[ifu_mem_ctl.scala 324:32]
  wire  ic_miss_buff_data_error_in_2 = write_fill_data_2 ? bus_ifu_wr_data_error : _T_1372; // @[ifu_mem_ctl.scala 323:72]
  wire  _T_1376 = ic_miss_buff_data_error[3] & _T_1330; // @[ifu_mem_ctl.scala 324:32]
  wire  ic_miss_buff_data_error_in_3 = write_fill_data_3 ? bus_ifu_wr_data_error : _T_1376; // @[ifu_mem_ctl.scala 323:72]
  wire  _T_1380 = ic_miss_buff_data_error[4] & _T_1330; // @[ifu_mem_ctl.scala 324:32]
  wire  ic_miss_buff_data_error_in_4 = write_fill_data_4 ? bus_ifu_wr_data_error : _T_1380; // @[ifu_mem_ctl.scala 323:72]
  wire  _T_1384 = ic_miss_buff_data_error[5] & _T_1330; // @[ifu_mem_ctl.scala 324:32]
  wire  ic_miss_buff_data_error_in_5 = write_fill_data_5 ? bus_ifu_wr_data_error : _T_1384; // @[ifu_mem_ctl.scala 323:72]
  wire  _T_1388 = ic_miss_buff_data_error[6] & _T_1330; // @[ifu_mem_ctl.scala 324:32]
  wire  ic_miss_buff_data_error_in_6 = write_fill_data_6 ? bus_ifu_wr_data_error : _T_1388; // @[ifu_mem_ctl.scala 323:72]
  wire  _T_1392 = ic_miss_buff_data_error[7] & _T_1330; // @[ifu_mem_ctl.scala 324:32]
  wire  ic_miss_buff_data_error_in_7 = write_fill_data_7 ? bus_ifu_wr_data_error : _T_1392; // @[ifu_mem_ctl.scala 323:72]
  wire [6:0] _T_1398 = {ic_miss_buff_data_error_in_7,ic_miss_buff_data_error_in_6,ic_miss_buff_data_error_in_5,ic_miss_buff_data_error_in_4,ic_miss_buff_data_error_in_3,ic_miss_buff_data_error_in_2,ic_miss_buff_data_error_in_1}; // @[Cat.scala 29:58]
  reg [6:0] perr_ic_index_ff; // @[Reg.scala 27:20]
  wire  _T_2500 = 3'h0 == perr_state; // @[Conditional.scala 37:30]
  wire  _T_2508 = _T_6 & _T_319; // @[ifu_mem_ctl.scala 405:82]
  wire  _T_2509 = _T_2508 | io_iccm_dma_sb_error; // @[ifu_mem_ctl.scala 405:105]
  wire  _T_2511 = _T_2509 & _T_2623; // @[ifu_mem_ctl.scala 405:129]
  wire  _T_2512 = 3'h1 == perr_state; // @[Conditional.scala 37:30]
  wire  _T_2513 = io_dec_tlu_flush_lower_wb | io_dec_mem_ctrl_dec_tlu_force_halt; // @[ifu_mem_ctl.scala 410:50]
  wire  _T_2515 = 3'h2 == perr_state; // @[Conditional.scala 37:30]
  wire  _T_2522 = 3'h4 == perr_state; // @[Conditional.scala 37:30]
  wire  _T_2524 = 3'h3 == perr_state; // @[Conditional.scala 37:30]
  wire  _GEN_21 = _T_2522 | _T_2524; // @[Conditional.scala 39:67]
  wire  _GEN_23 = _T_2515 ? _T_2513 : _GEN_21; // @[Conditional.scala 39:67]
  wire  _GEN_25 = _T_2512 ? _T_2513 : _GEN_23; // @[Conditional.scala 39:67]
  wire  perr_state_en = _T_2500 ? _T_2511 : _GEN_25; // @[Conditional.scala 40:58]
  wire  perr_sb_write_status = _T_2500 & perr_state_en; // @[Conditional.scala 40:58]
  wire  _T_2514 = io_dec_tlu_flush_lower_wb & io_dec_mem_ctrl_dec_tlu_flush_err_wb; // @[ifu_mem_ctl.scala 411:56]
  wire  _GEN_26 = _T_2512 & _T_2514; // @[Conditional.scala 39:67]
  wire  perr_sel_invalidate = _T_2500 ? 1'h0 : _GEN_26; // @[Conditional.scala 40:58]
  wire [1:0] perr_err_inv_way = perr_sel_invalidate ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  reg  dma_sb_err_state_ff; // @[ifu_mem_ctl.scala 396:58]
  wire  _T_2497 = ~dma_sb_err_state_ff; // @[ifu_mem_ctl.scala 395:49]
  wire  _T_2502 = io_dec_mem_ctrl_ifu_ic_error_start & _T_319; // @[ifu_mem_ctl.scala 404:104]
  wire  _T_2516 = ~io_dec_mem_ctrl_dec_tlu_flush_err_wb; // @[ifu_mem_ctl.scala 414:30]
  wire  _T_2517 = _T_2516 & io_dec_tlu_flush_lower_wb; // @[ifu_mem_ctl.scala 414:68]
  wire  _T_2518 = _T_2517 | io_dec_mem_ctrl_dec_tlu_force_halt; // @[ifu_mem_ctl.scala 414:98]
  wire  _T_2527 = perr_state == 3'h2; // @[ifu_mem_ctl.scala 434:79]
  wire  _T_2528 = io_dec_mem_ctrl_dec_tlu_flush_err_wb & _T_2527; // @[ifu_mem_ctl.scala 434:65]
  wire  _T_2530 = _T_2528 & _T_2623; // @[ifu_mem_ctl.scala 434:94]
  wire  _T_2532 = io_dec_tlu_flush_lower_wb | io_dec_mem_ctrl_dec_tlu_i0_commit_cmt; // @[ifu_mem_ctl.scala 437:59]
  wire  _T_2533 = _T_2532 | io_dec_mem_ctrl_dec_tlu_force_halt; // @[ifu_mem_ctl.scala 437:99]
  wire  _T_2547 = _T_2532 | io_ifu_fetch_val[0]; // @[ifu_mem_ctl.scala 440:94]
  wire  _T_2548 = _T_2547 | ifu_bp_hit_taken_q_f; // @[ifu_mem_ctl.scala 440:116]
  wire  _T_2549 = _T_2548 | io_dec_mem_ctrl_dec_tlu_force_halt; // @[ifu_mem_ctl.scala 440:139]
  wire  _T_2569 = _T_2547 | io_dec_mem_ctrl_dec_tlu_force_halt; // @[ifu_mem_ctl.scala 447:116]
  wire  _T_2577 = io_dec_tlu_flush_lower_wb & _T_2516; // @[ifu_mem_ctl.scala 452:60]
  wire  _T_2578 = _T_2577 | io_dec_mem_ctrl_dec_tlu_i0_commit_cmt; // @[ifu_mem_ctl.scala 452:101]
  wire  _T_2579 = _T_2578 | io_dec_mem_ctrl_dec_tlu_force_halt; // @[ifu_mem_ctl.scala 452:141]
  wire  _GEN_33 = _T_2575 & _T_2533; // @[Conditional.scala 39:67]
  wire  _GEN_36 = _T_2558 ? _T_2569 : _GEN_33; // @[Conditional.scala 39:67]
  wire  _GEN_38 = _T_2558 | _T_2575; // @[Conditional.scala 39:67]
  wire  _GEN_40 = _T_2531 ? _T_2549 : _GEN_36; // @[Conditional.scala 39:67]
  wire  _GEN_42 = _T_2531 | _GEN_38; // @[Conditional.scala 39:67]
  wire  err_stop_state_en = _T_2526 ? _T_2530 : _GEN_40; // @[Conditional.scala 40:58]
  reg  bus_cmd_req_hold; // @[ifu_mem_ctl.scala 475:53]
  wire  _T_2591 = ic_act_miss_f | bus_cmd_req_hold; // @[ifu_mem_ctl.scala 471:45]
  reg  ifu_bus_cmd_valid; // @[ifu_mem_ctl.scala 472:55]
  wire  _T_2592 = _T_2591 | ifu_bus_cmd_valid; // @[ifu_mem_ctl.scala 471:64]
  wire  _T_2594 = _T_2592 & _T_2623; // @[ifu_mem_ctl.scala 471:85]
  reg [2:0] bus_cmd_beat_count; // @[Reg.scala 27:20]
  wire  _T_2596 = bus_cmd_beat_count == 3'h7; // @[ifu_mem_ctl.scala 471:146]
  wire  _T_2597 = _T_2596 & ifu_bus_cmd_valid; // @[ifu_mem_ctl.scala 471:177]
  wire  _T_2598 = _T_2597 & io_ifu_axi_ar_ready; // @[ifu_mem_ctl.scala 471:197]
  wire  _T_2599 = _T_2598 & miss_pending; // @[ifu_mem_ctl.scala 471:217]
  wire  _T_2600 = ~_T_2599; // @[ifu_mem_ctl.scala 471:125]
  wire  ifu_bus_arready = io_ifu_axi_ar_ready & io_ifu_bus_clk_en; // @[ifu_mem_ctl.scala 522:45]
  wire  _T_2617 = io_ifu_axi_ar_valid & ifu_bus_arready; // @[ifu_mem_ctl.scala 526:35]
  wire  _T_2618 = _T_2617 & miss_pending; // @[ifu_mem_ctl.scala 526:53]
  wire  bus_cmd_sent = _T_2618 & _T_2623; // @[ifu_mem_ctl.scala 526:68]
  wire  _T_2603 = ~bus_cmd_sent; // @[ifu_mem_ctl.scala 474:61]
  wire  _T_2604 = _T_2591 & _T_2603; // @[ifu_mem_ctl.scala 474:59]
  wire [2:0] _T_2608 = ifu_bus_cmd_valid ? 3'h7 : 3'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_2610 = {miss_addr,bus_rd_addr_count,3'h0}; // @[Cat.scala 29:58]
  wire [31:0] _T_2612 = ifu_bus_cmd_valid ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  reg  ifu_bus_arready_unq_ff; // @[ifu_mem_ctl.scala 509:57]
  reg  ifu_bus_arvalid_ff; // @[ifu_mem_ctl.scala 511:53]
  wire  ifu_bus_arready_ff = ifu_bus_arready_unq_ff & bus_ifu_bus_clk_en_ff; // @[ifu_mem_ctl.scala 523:51]
  wire  _T_2638 = ~scnd_miss_req; // @[ifu_mem_ctl.scala 534:73]
  wire  _T_2639 = _T_2624 & _T_2638; // @[ifu_mem_ctl.scala 534:71]
  wire  _T_2641 = last_data_recieved_ff & _T_1330; // @[ifu_mem_ctl.scala 534:114]
  wire [2:0] _T_2647 = bus_rd_addr_count + 3'h1; // @[ifu_mem_ctl.scala 539:45]
  wire  _T_2651 = ifu_bus_cmd_valid & io_ifu_axi_ar_ready; // @[ifu_mem_ctl.scala 542:48]
  wire  _T_2652 = _T_2651 & miss_pending; // @[ifu_mem_ctl.scala 542:68]
  wire  bus_inc_cmd_beat_cnt = _T_2652 & _T_2623; // @[ifu_mem_ctl.scala 542:83]
  wire  bus_reset_cmd_beat_cnt_secondlast = ic_act_miss_f & uncacheable_miss_in; // @[ifu_mem_ctl.scala 544:57]
  wire  _T_2656 = ~bus_inc_cmd_beat_cnt; // @[ifu_mem_ctl.scala 545:31]
  wire  _T_2657 = ic_act_miss_f | scnd_miss_req; // @[ifu_mem_ctl.scala 545:71]
  wire  _T_2658 = _T_2657 | io_dec_mem_ctrl_dec_tlu_force_halt; // @[ifu_mem_ctl.scala 545:87]
  wire  _T_2659 = ~_T_2658; // @[ifu_mem_ctl.scala 545:55]
  wire  bus_hold_cmd_beat_cnt = _T_2656 & _T_2659; // @[ifu_mem_ctl.scala 545:53]
  wire  _T_2660 = bus_inc_cmd_beat_cnt | ic_act_miss_f; // @[ifu_mem_ctl.scala 546:46]
  wire  bus_cmd_beat_en = _T_2660 | io_dec_mem_ctrl_dec_tlu_force_halt; // @[ifu_mem_ctl.scala 546:62]
  wire [2:0] _T_2663 = bus_cmd_beat_count + 3'h1; // @[ifu_mem_ctl.scala 548:46]
  wire [2:0] _T_2665 = bus_reset_cmd_beat_cnt_secondlast ? 3'h6 : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_2666 = bus_inc_cmd_beat_cnt ? _T_2663 : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_2667 = bus_hold_cmd_beat_cnt ? bus_cmd_beat_count : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_2669 = _T_2665 | _T_2666; // @[Mux.scala 27:72]
  wire [2:0] bus_new_cmd_beat_count = _T_2669 | _T_2667; // @[Mux.scala 27:72]
  reg  ifc_dma_access_ok_prev; // @[ifu_mem_ctl.scala 560:62]
  wire  _T_2698 = ~iccm_correct_ecc; // @[ifu_mem_ctl.scala 565:50]
  wire  _T_2699 = io_ifc_dma_access_ok & _T_2698; // @[ifu_mem_ctl.scala 565:47]
  wire  _T_2700 = ~io_iccm_dma_sb_error; // @[ifu_mem_ctl.scala 565:70]
  wire  _T_2704 = _T_2699 & ifc_dma_access_ok_prev; // @[ifu_mem_ctl.scala 566:72]
  wire  _T_2705 = perr_state == 3'h0; // @[ifu_mem_ctl.scala 566:111]
  wire  _T_2706 = _T_2704 & _T_2705; // @[ifu_mem_ctl.scala 566:97]
  wire  ifc_dma_access_q_ok = _T_2706 & _T_2700; // @[ifu_mem_ctl.scala 566:127]
  wire  _T_2709 = ifc_dma_access_q_ok & io_dma_mem_ctl_dma_iccm_req; // @[ifu_mem_ctl.scala 569:40]
  wire  _T_2710 = _T_2709 & io_dma_mem_ctl_dma_mem_write; // @[ifu_mem_ctl.scala 569:70]
  wire  _T_2713 = ~io_dma_mem_ctl_dma_mem_write; // @[ifu_mem_ctl.scala 570:72]
  wire  _T_2714 = _T_2709 & _T_2713; // @[ifu_mem_ctl.scala 570:70]
  wire  _T_2715 = io_ifc_iccm_access_bf & io_ifc_fetch_req_bf; // @[ifu_mem_ctl.scala 570:128]
  wire [2:0] _T_2720 = io_dma_mem_ctl_dma_iccm_req ? 3'h7 : 3'h0; // @[Bitwise.scala 72:12]
  wire  _T_2741 = io_dma_mem_ctl_dma_mem_wdata[32] ^ io_dma_mem_ctl_dma_mem_wdata[33]; // @[lib.scala 119:74]
  wire  _T_2742 = _T_2741 ^ io_dma_mem_ctl_dma_mem_wdata[35]; // @[lib.scala 119:74]
  wire  _T_2743 = _T_2742 ^ io_dma_mem_ctl_dma_mem_wdata[36]; // @[lib.scala 119:74]
  wire  _T_2744 = _T_2743 ^ io_dma_mem_ctl_dma_mem_wdata[38]; // @[lib.scala 119:74]
  wire  _T_2745 = _T_2744 ^ io_dma_mem_ctl_dma_mem_wdata[40]; // @[lib.scala 119:74]
  wire  _T_2746 = _T_2745 ^ io_dma_mem_ctl_dma_mem_wdata[42]; // @[lib.scala 119:74]
  wire  _T_2747 = _T_2746 ^ io_dma_mem_ctl_dma_mem_wdata[43]; // @[lib.scala 119:74]
  wire  _T_2748 = _T_2747 ^ io_dma_mem_ctl_dma_mem_wdata[45]; // @[lib.scala 119:74]
  wire  _T_2749 = _T_2748 ^ io_dma_mem_ctl_dma_mem_wdata[47]; // @[lib.scala 119:74]
  wire  _T_2750 = _T_2749 ^ io_dma_mem_ctl_dma_mem_wdata[49]; // @[lib.scala 119:74]
  wire  _T_2751 = _T_2750 ^ io_dma_mem_ctl_dma_mem_wdata[51]; // @[lib.scala 119:74]
  wire  _T_2752 = _T_2751 ^ io_dma_mem_ctl_dma_mem_wdata[53]; // @[lib.scala 119:74]
  wire  _T_2753 = _T_2752 ^ io_dma_mem_ctl_dma_mem_wdata[55]; // @[lib.scala 119:74]
  wire  _T_2754 = _T_2753 ^ io_dma_mem_ctl_dma_mem_wdata[57]; // @[lib.scala 119:74]
  wire  _T_2755 = _T_2754 ^ io_dma_mem_ctl_dma_mem_wdata[58]; // @[lib.scala 119:74]
  wire  _T_2756 = _T_2755 ^ io_dma_mem_ctl_dma_mem_wdata[60]; // @[lib.scala 119:74]
  wire  _T_2757 = _T_2756 ^ io_dma_mem_ctl_dma_mem_wdata[62]; // @[lib.scala 119:74]
  wire  _T_2776 = io_dma_mem_ctl_dma_mem_wdata[32] ^ io_dma_mem_ctl_dma_mem_wdata[34]; // @[lib.scala 119:74]
  wire  _T_2777 = _T_2776 ^ io_dma_mem_ctl_dma_mem_wdata[35]; // @[lib.scala 119:74]
  wire  _T_2778 = _T_2777 ^ io_dma_mem_ctl_dma_mem_wdata[37]; // @[lib.scala 119:74]
  wire  _T_2779 = _T_2778 ^ io_dma_mem_ctl_dma_mem_wdata[38]; // @[lib.scala 119:74]
  wire  _T_2780 = _T_2779 ^ io_dma_mem_ctl_dma_mem_wdata[41]; // @[lib.scala 119:74]
  wire  _T_2781 = _T_2780 ^ io_dma_mem_ctl_dma_mem_wdata[42]; // @[lib.scala 119:74]
  wire  _T_2782 = _T_2781 ^ io_dma_mem_ctl_dma_mem_wdata[44]; // @[lib.scala 119:74]
  wire  _T_2783 = _T_2782 ^ io_dma_mem_ctl_dma_mem_wdata[45]; // @[lib.scala 119:74]
  wire  _T_2784 = _T_2783 ^ io_dma_mem_ctl_dma_mem_wdata[48]; // @[lib.scala 119:74]
  wire  _T_2785 = _T_2784 ^ io_dma_mem_ctl_dma_mem_wdata[49]; // @[lib.scala 119:74]
  wire  _T_2786 = _T_2785 ^ io_dma_mem_ctl_dma_mem_wdata[52]; // @[lib.scala 119:74]
  wire  _T_2787 = _T_2786 ^ io_dma_mem_ctl_dma_mem_wdata[53]; // @[lib.scala 119:74]
  wire  _T_2788 = _T_2787 ^ io_dma_mem_ctl_dma_mem_wdata[56]; // @[lib.scala 119:74]
  wire  _T_2789 = _T_2788 ^ io_dma_mem_ctl_dma_mem_wdata[57]; // @[lib.scala 119:74]
  wire  _T_2790 = _T_2789 ^ io_dma_mem_ctl_dma_mem_wdata[59]; // @[lib.scala 119:74]
  wire  _T_2791 = _T_2790 ^ io_dma_mem_ctl_dma_mem_wdata[60]; // @[lib.scala 119:74]
  wire  _T_2792 = _T_2791 ^ io_dma_mem_ctl_dma_mem_wdata[63]; // @[lib.scala 119:74]
  wire  _T_2811 = io_dma_mem_ctl_dma_mem_wdata[33] ^ io_dma_mem_ctl_dma_mem_wdata[34]; // @[lib.scala 119:74]
  wire  _T_2812 = _T_2811 ^ io_dma_mem_ctl_dma_mem_wdata[35]; // @[lib.scala 119:74]
  wire  _T_2813 = _T_2812 ^ io_dma_mem_ctl_dma_mem_wdata[39]; // @[lib.scala 119:74]
  wire  _T_2814 = _T_2813 ^ io_dma_mem_ctl_dma_mem_wdata[40]; // @[lib.scala 119:74]
  wire  _T_2815 = _T_2814 ^ io_dma_mem_ctl_dma_mem_wdata[41]; // @[lib.scala 119:74]
  wire  _T_2816 = _T_2815 ^ io_dma_mem_ctl_dma_mem_wdata[42]; // @[lib.scala 119:74]
  wire  _T_2817 = _T_2816 ^ io_dma_mem_ctl_dma_mem_wdata[46]; // @[lib.scala 119:74]
  wire  _T_2818 = _T_2817 ^ io_dma_mem_ctl_dma_mem_wdata[47]; // @[lib.scala 119:74]
  wire  _T_2819 = _T_2818 ^ io_dma_mem_ctl_dma_mem_wdata[48]; // @[lib.scala 119:74]
  wire  _T_2820 = _T_2819 ^ io_dma_mem_ctl_dma_mem_wdata[49]; // @[lib.scala 119:74]
  wire  _T_2821 = _T_2820 ^ io_dma_mem_ctl_dma_mem_wdata[54]; // @[lib.scala 119:74]
  wire  _T_2822 = _T_2821 ^ io_dma_mem_ctl_dma_mem_wdata[55]; // @[lib.scala 119:74]
  wire  _T_2823 = _T_2822 ^ io_dma_mem_ctl_dma_mem_wdata[56]; // @[lib.scala 119:74]
  wire  _T_2824 = _T_2823 ^ io_dma_mem_ctl_dma_mem_wdata[57]; // @[lib.scala 119:74]
  wire  _T_2825 = _T_2824 ^ io_dma_mem_ctl_dma_mem_wdata[61]; // @[lib.scala 119:74]
  wire  _T_2826 = _T_2825 ^ io_dma_mem_ctl_dma_mem_wdata[62]; // @[lib.scala 119:74]
  wire  _T_2827 = _T_2826 ^ io_dma_mem_ctl_dma_mem_wdata[63]; // @[lib.scala 119:74]
  wire  _T_2843 = io_dma_mem_ctl_dma_mem_wdata[36] ^ io_dma_mem_ctl_dma_mem_wdata[37]; // @[lib.scala 119:74]
  wire  _T_2844 = _T_2843 ^ io_dma_mem_ctl_dma_mem_wdata[38]; // @[lib.scala 119:74]
  wire  _T_2845 = _T_2844 ^ io_dma_mem_ctl_dma_mem_wdata[39]; // @[lib.scala 119:74]
  wire  _T_2846 = _T_2845 ^ io_dma_mem_ctl_dma_mem_wdata[40]; // @[lib.scala 119:74]
  wire  _T_2847 = _T_2846 ^ io_dma_mem_ctl_dma_mem_wdata[41]; // @[lib.scala 119:74]
  wire  _T_2848 = _T_2847 ^ io_dma_mem_ctl_dma_mem_wdata[42]; // @[lib.scala 119:74]
  wire  _T_2849 = _T_2848 ^ io_dma_mem_ctl_dma_mem_wdata[50]; // @[lib.scala 119:74]
  wire  _T_2850 = _T_2849 ^ io_dma_mem_ctl_dma_mem_wdata[51]; // @[lib.scala 119:74]
  wire  _T_2851 = _T_2850 ^ io_dma_mem_ctl_dma_mem_wdata[52]; // @[lib.scala 119:74]
  wire  _T_2852 = _T_2851 ^ io_dma_mem_ctl_dma_mem_wdata[53]; // @[lib.scala 119:74]
  wire  _T_2853 = _T_2852 ^ io_dma_mem_ctl_dma_mem_wdata[54]; // @[lib.scala 119:74]
  wire  _T_2854 = _T_2853 ^ io_dma_mem_ctl_dma_mem_wdata[55]; // @[lib.scala 119:74]
  wire  _T_2855 = _T_2854 ^ io_dma_mem_ctl_dma_mem_wdata[56]; // @[lib.scala 119:74]
  wire  _T_2856 = _T_2855 ^ io_dma_mem_ctl_dma_mem_wdata[57]; // @[lib.scala 119:74]
  wire  _T_2872 = io_dma_mem_ctl_dma_mem_wdata[43] ^ io_dma_mem_ctl_dma_mem_wdata[44]; // @[lib.scala 119:74]
  wire  _T_2873 = _T_2872 ^ io_dma_mem_ctl_dma_mem_wdata[45]; // @[lib.scala 119:74]
  wire  _T_2874 = _T_2873 ^ io_dma_mem_ctl_dma_mem_wdata[46]; // @[lib.scala 119:74]
  wire  _T_2875 = _T_2874 ^ io_dma_mem_ctl_dma_mem_wdata[47]; // @[lib.scala 119:74]
  wire  _T_2876 = _T_2875 ^ io_dma_mem_ctl_dma_mem_wdata[48]; // @[lib.scala 119:74]
  wire  _T_2877 = _T_2876 ^ io_dma_mem_ctl_dma_mem_wdata[49]; // @[lib.scala 119:74]
  wire  _T_2878 = _T_2877 ^ io_dma_mem_ctl_dma_mem_wdata[50]; // @[lib.scala 119:74]
  wire  _T_2879 = _T_2878 ^ io_dma_mem_ctl_dma_mem_wdata[51]; // @[lib.scala 119:74]
  wire  _T_2880 = _T_2879 ^ io_dma_mem_ctl_dma_mem_wdata[52]; // @[lib.scala 119:74]
  wire  _T_2881 = _T_2880 ^ io_dma_mem_ctl_dma_mem_wdata[53]; // @[lib.scala 119:74]
  wire  _T_2882 = _T_2881 ^ io_dma_mem_ctl_dma_mem_wdata[54]; // @[lib.scala 119:74]
  wire  _T_2883 = _T_2882 ^ io_dma_mem_ctl_dma_mem_wdata[55]; // @[lib.scala 119:74]
  wire  _T_2884 = _T_2883 ^ io_dma_mem_ctl_dma_mem_wdata[56]; // @[lib.scala 119:74]
  wire  _T_2885 = _T_2884 ^ io_dma_mem_ctl_dma_mem_wdata[57]; // @[lib.scala 119:74]
  wire  _T_2892 = io_dma_mem_ctl_dma_mem_wdata[58] ^ io_dma_mem_ctl_dma_mem_wdata[59]; // @[lib.scala 119:74]
  wire  _T_2893 = _T_2892 ^ io_dma_mem_ctl_dma_mem_wdata[60]; // @[lib.scala 119:74]
  wire  _T_2894 = _T_2893 ^ io_dma_mem_ctl_dma_mem_wdata[61]; // @[lib.scala 119:74]
  wire  _T_2895 = _T_2894 ^ io_dma_mem_ctl_dma_mem_wdata[62]; // @[lib.scala 119:74]
  wire  _T_2896 = _T_2895 ^ io_dma_mem_ctl_dma_mem_wdata[63]; // @[lib.scala 119:74]
  wire [5:0] _T_2901 = {_T_2896,_T_2885,_T_2856,_T_2827,_T_2792,_T_2757}; // @[Cat.scala 29:58]
  wire  _T_2902 = ^io_dma_mem_ctl_dma_mem_wdata[63:32]; // @[lib.scala 127:13]
  wire  _T_2903 = ^_T_2901; // @[lib.scala 127:23]
  wire  _T_2904 = _T_2902 ^ _T_2903; // @[lib.scala 127:18]
  wire  _T_2925 = io_dma_mem_ctl_dma_mem_wdata[0] ^ io_dma_mem_ctl_dma_mem_wdata[1]; // @[lib.scala 119:74]
  wire  _T_2926 = _T_2925 ^ io_dma_mem_ctl_dma_mem_wdata[3]; // @[lib.scala 119:74]
  wire  _T_2927 = _T_2926 ^ io_dma_mem_ctl_dma_mem_wdata[4]; // @[lib.scala 119:74]
  wire  _T_2928 = _T_2927 ^ io_dma_mem_ctl_dma_mem_wdata[6]; // @[lib.scala 119:74]
  wire  _T_2929 = _T_2928 ^ io_dma_mem_ctl_dma_mem_wdata[8]; // @[lib.scala 119:74]
  wire  _T_2930 = _T_2929 ^ io_dma_mem_ctl_dma_mem_wdata[10]; // @[lib.scala 119:74]
  wire  _T_2931 = _T_2930 ^ io_dma_mem_ctl_dma_mem_wdata[11]; // @[lib.scala 119:74]
  wire  _T_2932 = _T_2931 ^ io_dma_mem_ctl_dma_mem_wdata[13]; // @[lib.scala 119:74]
  wire  _T_2933 = _T_2932 ^ io_dma_mem_ctl_dma_mem_wdata[15]; // @[lib.scala 119:74]
  wire  _T_2934 = _T_2933 ^ io_dma_mem_ctl_dma_mem_wdata[17]; // @[lib.scala 119:74]
  wire  _T_2935 = _T_2934 ^ io_dma_mem_ctl_dma_mem_wdata[19]; // @[lib.scala 119:74]
  wire  _T_2936 = _T_2935 ^ io_dma_mem_ctl_dma_mem_wdata[21]; // @[lib.scala 119:74]
  wire  _T_2937 = _T_2936 ^ io_dma_mem_ctl_dma_mem_wdata[23]; // @[lib.scala 119:74]
  wire  _T_2938 = _T_2937 ^ io_dma_mem_ctl_dma_mem_wdata[25]; // @[lib.scala 119:74]
  wire  _T_2939 = _T_2938 ^ io_dma_mem_ctl_dma_mem_wdata[26]; // @[lib.scala 119:74]
  wire  _T_2940 = _T_2939 ^ io_dma_mem_ctl_dma_mem_wdata[28]; // @[lib.scala 119:74]
  wire  _T_2941 = _T_2940 ^ io_dma_mem_ctl_dma_mem_wdata[30]; // @[lib.scala 119:74]
  wire  _T_2960 = io_dma_mem_ctl_dma_mem_wdata[0] ^ io_dma_mem_ctl_dma_mem_wdata[2]; // @[lib.scala 119:74]
  wire  _T_2961 = _T_2960 ^ io_dma_mem_ctl_dma_mem_wdata[3]; // @[lib.scala 119:74]
  wire  _T_2962 = _T_2961 ^ io_dma_mem_ctl_dma_mem_wdata[5]; // @[lib.scala 119:74]
  wire  _T_2963 = _T_2962 ^ io_dma_mem_ctl_dma_mem_wdata[6]; // @[lib.scala 119:74]
  wire  _T_2964 = _T_2963 ^ io_dma_mem_ctl_dma_mem_wdata[9]; // @[lib.scala 119:74]
  wire  _T_2965 = _T_2964 ^ io_dma_mem_ctl_dma_mem_wdata[10]; // @[lib.scala 119:74]
  wire  _T_2966 = _T_2965 ^ io_dma_mem_ctl_dma_mem_wdata[12]; // @[lib.scala 119:74]
  wire  _T_2967 = _T_2966 ^ io_dma_mem_ctl_dma_mem_wdata[13]; // @[lib.scala 119:74]
  wire  _T_2968 = _T_2967 ^ io_dma_mem_ctl_dma_mem_wdata[16]; // @[lib.scala 119:74]
  wire  _T_2969 = _T_2968 ^ io_dma_mem_ctl_dma_mem_wdata[17]; // @[lib.scala 119:74]
  wire  _T_2970 = _T_2969 ^ io_dma_mem_ctl_dma_mem_wdata[20]; // @[lib.scala 119:74]
  wire  _T_2971 = _T_2970 ^ io_dma_mem_ctl_dma_mem_wdata[21]; // @[lib.scala 119:74]
  wire  _T_2972 = _T_2971 ^ io_dma_mem_ctl_dma_mem_wdata[24]; // @[lib.scala 119:74]
  wire  _T_2973 = _T_2972 ^ io_dma_mem_ctl_dma_mem_wdata[25]; // @[lib.scala 119:74]
  wire  _T_2974 = _T_2973 ^ io_dma_mem_ctl_dma_mem_wdata[27]; // @[lib.scala 119:74]
  wire  _T_2975 = _T_2974 ^ io_dma_mem_ctl_dma_mem_wdata[28]; // @[lib.scala 119:74]
  wire  _T_2976 = _T_2975 ^ io_dma_mem_ctl_dma_mem_wdata[31]; // @[lib.scala 119:74]
  wire  _T_2995 = io_dma_mem_ctl_dma_mem_wdata[1] ^ io_dma_mem_ctl_dma_mem_wdata[2]; // @[lib.scala 119:74]
  wire  _T_2996 = _T_2995 ^ io_dma_mem_ctl_dma_mem_wdata[3]; // @[lib.scala 119:74]
  wire  _T_2997 = _T_2996 ^ io_dma_mem_ctl_dma_mem_wdata[7]; // @[lib.scala 119:74]
  wire  _T_2998 = _T_2997 ^ io_dma_mem_ctl_dma_mem_wdata[8]; // @[lib.scala 119:74]
  wire  _T_2999 = _T_2998 ^ io_dma_mem_ctl_dma_mem_wdata[9]; // @[lib.scala 119:74]
  wire  _T_3000 = _T_2999 ^ io_dma_mem_ctl_dma_mem_wdata[10]; // @[lib.scala 119:74]
  wire  _T_3001 = _T_3000 ^ io_dma_mem_ctl_dma_mem_wdata[14]; // @[lib.scala 119:74]
  wire  _T_3002 = _T_3001 ^ io_dma_mem_ctl_dma_mem_wdata[15]; // @[lib.scala 119:74]
  wire  _T_3003 = _T_3002 ^ io_dma_mem_ctl_dma_mem_wdata[16]; // @[lib.scala 119:74]
  wire  _T_3004 = _T_3003 ^ io_dma_mem_ctl_dma_mem_wdata[17]; // @[lib.scala 119:74]
  wire  _T_3005 = _T_3004 ^ io_dma_mem_ctl_dma_mem_wdata[22]; // @[lib.scala 119:74]
  wire  _T_3006 = _T_3005 ^ io_dma_mem_ctl_dma_mem_wdata[23]; // @[lib.scala 119:74]
  wire  _T_3007 = _T_3006 ^ io_dma_mem_ctl_dma_mem_wdata[24]; // @[lib.scala 119:74]
  wire  _T_3008 = _T_3007 ^ io_dma_mem_ctl_dma_mem_wdata[25]; // @[lib.scala 119:74]
  wire  _T_3009 = _T_3008 ^ io_dma_mem_ctl_dma_mem_wdata[29]; // @[lib.scala 119:74]
  wire  _T_3010 = _T_3009 ^ io_dma_mem_ctl_dma_mem_wdata[30]; // @[lib.scala 119:74]
  wire  _T_3011 = _T_3010 ^ io_dma_mem_ctl_dma_mem_wdata[31]; // @[lib.scala 119:74]
  wire  _T_3027 = io_dma_mem_ctl_dma_mem_wdata[4] ^ io_dma_mem_ctl_dma_mem_wdata[5]; // @[lib.scala 119:74]
  wire  _T_3028 = _T_3027 ^ io_dma_mem_ctl_dma_mem_wdata[6]; // @[lib.scala 119:74]
  wire  _T_3029 = _T_3028 ^ io_dma_mem_ctl_dma_mem_wdata[7]; // @[lib.scala 119:74]
  wire  _T_3030 = _T_3029 ^ io_dma_mem_ctl_dma_mem_wdata[8]; // @[lib.scala 119:74]
  wire  _T_3031 = _T_3030 ^ io_dma_mem_ctl_dma_mem_wdata[9]; // @[lib.scala 119:74]
  wire  _T_3032 = _T_3031 ^ io_dma_mem_ctl_dma_mem_wdata[10]; // @[lib.scala 119:74]
  wire  _T_3033 = _T_3032 ^ io_dma_mem_ctl_dma_mem_wdata[18]; // @[lib.scala 119:74]
  wire  _T_3034 = _T_3033 ^ io_dma_mem_ctl_dma_mem_wdata[19]; // @[lib.scala 119:74]
  wire  _T_3035 = _T_3034 ^ io_dma_mem_ctl_dma_mem_wdata[20]; // @[lib.scala 119:74]
  wire  _T_3036 = _T_3035 ^ io_dma_mem_ctl_dma_mem_wdata[21]; // @[lib.scala 119:74]
  wire  _T_3037 = _T_3036 ^ io_dma_mem_ctl_dma_mem_wdata[22]; // @[lib.scala 119:74]
  wire  _T_3038 = _T_3037 ^ io_dma_mem_ctl_dma_mem_wdata[23]; // @[lib.scala 119:74]
  wire  _T_3039 = _T_3038 ^ io_dma_mem_ctl_dma_mem_wdata[24]; // @[lib.scala 119:74]
  wire  _T_3040 = _T_3039 ^ io_dma_mem_ctl_dma_mem_wdata[25]; // @[lib.scala 119:74]
  wire  _T_3056 = io_dma_mem_ctl_dma_mem_wdata[11] ^ io_dma_mem_ctl_dma_mem_wdata[12]; // @[lib.scala 119:74]
  wire  _T_3057 = _T_3056 ^ io_dma_mem_ctl_dma_mem_wdata[13]; // @[lib.scala 119:74]
  wire  _T_3058 = _T_3057 ^ io_dma_mem_ctl_dma_mem_wdata[14]; // @[lib.scala 119:74]
  wire  _T_3059 = _T_3058 ^ io_dma_mem_ctl_dma_mem_wdata[15]; // @[lib.scala 119:74]
  wire  _T_3060 = _T_3059 ^ io_dma_mem_ctl_dma_mem_wdata[16]; // @[lib.scala 119:74]
  wire  _T_3061 = _T_3060 ^ io_dma_mem_ctl_dma_mem_wdata[17]; // @[lib.scala 119:74]
  wire  _T_3062 = _T_3061 ^ io_dma_mem_ctl_dma_mem_wdata[18]; // @[lib.scala 119:74]
  wire  _T_3063 = _T_3062 ^ io_dma_mem_ctl_dma_mem_wdata[19]; // @[lib.scala 119:74]
  wire  _T_3064 = _T_3063 ^ io_dma_mem_ctl_dma_mem_wdata[20]; // @[lib.scala 119:74]
  wire  _T_3065 = _T_3064 ^ io_dma_mem_ctl_dma_mem_wdata[21]; // @[lib.scala 119:74]
  wire  _T_3066 = _T_3065 ^ io_dma_mem_ctl_dma_mem_wdata[22]; // @[lib.scala 119:74]
  wire  _T_3067 = _T_3066 ^ io_dma_mem_ctl_dma_mem_wdata[23]; // @[lib.scala 119:74]
  wire  _T_3068 = _T_3067 ^ io_dma_mem_ctl_dma_mem_wdata[24]; // @[lib.scala 119:74]
  wire  _T_3069 = _T_3068 ^ io_dma_mem_ctl_dma_mem_wdata[25]; // @[lib.scala 119:74]
  wire  _T_3076 = io_dma_mem_ctl_dma_mem_wdata[26] ^ io_dma_mem_ctl_dma_mem_wdata[27]; // @[lib.scala 119:74]
  wire  _T_3077 = _T_3076 ^ io_dma_mem_ctl_dma_mem_wdata[28]; // @[lib.scala 119:74]
  wire  _T_3078 = _T_3077 ^ io_dma_mem_ctl_dma_mem_wdata[29]; // @[lib.scala 119:74]
  wire  _T_3079 = _T_3078 ^ io_dma_mem_ctl_dma_mem_wdata[30]; // @[lib.scala 119:74]
  wire  _T_3080 = _T_3079 ^ io_dma_mem_ctl_dma_mem_wdata[31]; // @[lib.scala 119:74]
  wire [5:0] _T_3085 = {_T_3080,_T_3069,_T_3040,_T_3011,_T_2976,_T_2941}; // @[Cat.scala 29:58]
  wire  _T_3086 = ^io_dma_mem_ctl_dma_mem_wdata[31:0]; // @[lib.scala 127:13]
  wire  _T_3087 = ^_T_3085; // @[lib.scala 127:23]
  wire  _T_3088 = _T_3086 ^ _T_3087; // @[lib.scala 127:18]
  wire [6:0] _T_3089 = {_T_3088,_T_3080,_T_3069,_T_3040,_T_3011,_T_2976,_T_2941}; // @[Cat.scala 29:58]
  wire [13:0] dma_mem_ecc = {_T_2904,_T_2896,_T_2885,_T_2856,_T_2827,_T_2792,_T_2757,_T_3089}; // @[Cat.scala 29:58]
  wire  _T_3091 = ~_T_2709; // @[ifu_mem_ctl.scala 576:45]
  wire  _T_3092 = iccm_correct_ecc & _T_3091; // @[ifu_mem_ctl.scala 576:43]
  reg [38:0] iccm_ecc_corr_data_ff; // @[Reg.scala 27:20]
  wire [77:0] _T_3093 = {iccm_ecc_corr_data_ff,iccm_ecc_corr_data_ff}; // @[Cat.scala 29:58]
  wire [77:0] _T_3100 = {dma_mem_ecc[13:7],io_dma_mem_ctl_dma_mem_wdata[63:32],dma_mem_ecc[6:0],io_dma_mem_ctl_dma_mem_wdata[31:0]}; // @[Cat.scala 29:58]
  reg [1:0] dma_mem_addr_ff; // @[ifu_mem_ctl.scala 590:53]
  wire  _T_3435 = _T_3347[5:0] == 6'h27; // @[lib.scala 199:41]
  wire  _T_3433 = _T_3347[5:0] == 6'h26; // @[lib.scala 199:41]
  wire  _T_3431 = _T_3347[5:0] == 6'h25; // @[lib.scala 199:41]
  wire  _T_3429 = _T_3347[5:0] == 6'h24; // @[lib.scala 199:41]
  wire  _T_3427 = _T_3347[5:0] == 6'h23; // @[lib.scala 199:41]
  wire  _T_3425 = _T_3347[5:0] == 6'h22; // @[lib.scala 199:41]
  wire  _T_3423 = _T_3347[5:0] == 6'h21; // @[lib.scala 199:41]
  wire  _T_3421 = _T_3347[5:0] == 6'h20; // @[lib.scala 199:41]
  wire  _T_3419 = _T_3347[5:0] == 6'h1f; // @[lib.scala 199:41]
  wire  _T_3417 = _T_3347[5:0] == 6'h1e; // @[lib.scala 199:41]
  wire [9:0] _T_3493 = {_T_3435,_T_3433,_T_3431,_T_3429,_T_3427,_T_3425,_T_3423,_T_3421,_T_3419,_T_3417}; // @[lib.scala 202:69]
  wire  _T_3415 = _T_3347[5:0] == 6'h1d; // @[lib.scala 199:41]
  wire  _T_3413 = _T_3347[5:0] == 6'h1c; // @[lib.scala 199:41]
  wire  _T_3411 = _T_3347[5:0] == 6'h1b; // @[lib.scala 199:41]
  wire  _T_3409 = _T_3347[5:0] == 6'h1a; // @[lib.scala 199:41]
  wire  _T_3407 = _T_3347[5:0] == 6'h19; // @[lib.scala 199:41]
  wire  _T_3405 = _T_3347[5:0] == 6'h18; // @[lib.scala 199:41]
  wire  _T_3403 = _T_3347[5:0] == 6'h17; // @[lib.scala 199:41]
  wire  _T_3401 = _T_3347[5:0] == 6'h16; // @[lib.scala 199:41]
  wire  _T_3399 = _T_3347[5:0] == 6'h15; // @[lib.scala 199:41]
  wire  _T_3397 = _T_3347[5:0] == 6'h14; // @[lib.scala 199:41]
  wire [9:0] _T_3484 = {_T_3415,_T_3413,_T_3411,_T_3409,_T_3407,_T_3405,_T_3403,_T_3401,_T_3399,_T_3397}; // @[lib.scala 202:69]
  wire  _T_3395 = _T_3347[5:0] == 6'h13; // @[lib.scala 199:41]
  wire  _T_3393 = _T_3347[5:0] == 6'h12; // @[lib.scala 199:41]
  wire  _T_3391 = _T_3347[5:0] == 6'h11; // @[lib.scala 199:41]
  wire  _T_3389 = _T_3347[5:0] == 6'h10; // @[lib.scala 199:41]
  wire  _T_3387 = _T_3347[5:0] == 6'hf; // @[lib.scala 199:41]
  wire  _T_3385 = _T_3347[5:0] == 6'he; // @[lib.scala 199:41]
  wire  _T_3383 = _T_3347[5:0] == 6'hd; // @[lib.scala 199:41]
  wire  _T_3381 = _T_3347[5:0] == 6'hc; // @[lib.scala 199:41]
  wire  _T_3379 = _T_3347[5:0] == 6'hb; // @[lib.scala 199:41]
  wire  _T_3377 = _T_3347[5:0] == 6'ha; // @[lib.scala 199:41]
  wire [9:0] _T_3474 = {_T_3395,_T_3393,_T_3391,_T_3389,_T_3387,_T_3385,_T_3383,_T_3381,_T_3379,_T_3377}; // @[lib.scala 202:69]
  wire  _T_3375 = _T_3347[5:0] == 6'h9; // @[lib.scala 199:41]
  wire  _T_3373 = _T_3347[5:0] == 6'h8; // @[lib.scala 199:41]
  wire  _T_3371 = _T_3347[5:0] == 6'h7; // @[lib.scala 199:41]
  wire  _T_3369 = _T_3347[5:0] == 6'h6; // @[lib.scala 199:41]
  wire  _T_3367 = _T_3347[5:0] == 6'h5; // @[lib.scala 199:41]
  wire  _T_3365 = _T_3347[5:0] == 6'h4; // @[lib.scala 199:41]
  wire  _T_3363 = _T_3347[5:0] == 6'h3; // @[lib.scala 199:41]
  wire  _T_3361 = _T_3347[5:0] == 6'h2; // @[lib.scala 199:41]
  wire  _T_3359 = _T_3347[5:0] == 6'h1; // @[lib.scala 199:41]
  wire [18:0] _T_3475 = {_T_3474,_T_3375,_T_3373,_T_3371,_T_3369,_T_3367,_T_3365,_T_3363,_T_3361,_T_3359}; // @[lib.scala 202:69]
  wire [38:0] _T_3495 = {_T_3493,_T_3484,_T_3475}; // @[lib.scala 202:69]
  wire [7:0] _T_3450 = {io_iccm_rd_data_ecc[35],io_iccm_rd_data_ecc[3:1],io_iccm_rd_data_ecc[34],io_iccm_rd_data_ecc[0],io_iccm_rd_data_ecc[33:32]}; // @[Cat.scala 29:58]
  wire [38:0] _T_3456 = {io_iccm_rd_data_ecc[38],io_iccm_rd_data_ecc[31:26],io_iccm_rd_data_ecc[37],io_iccm_rd_data_ecc[25:11],io_iccm_rd_data_ecc[36],io_iccm_rd_data_ecc[10:4],_T_3450}; // @[Cat.scala 29:58]
  wire [38:0] _T_3496 = _T_3495 ^ _T_3456; // @[lib.scala 202:76]
  wire [38:0] _T_3497 = _T_3351 ? _T_3496 : _T_3456; // @[lib.scala 202:31]
  wire [31:0] iccm_corrected_data_0 = {_T_3497[37:32],_T_3497[30:16],_T_3497[14:8],_T_3497[6:4],_T_3497[2]}; // @[Cat.scala 29:58]
  wire  _T_3820 = _T_3732[5:0] == 6'h27; // @[lib.scala 199:41]
  wire  _T_3818 = _T_3732[5:0] == 6'h26; // @[lib.scala 199:41]
  wire  _T_3816 = _T_3732[5:0] == 6'h25; // @[lib.scala 199:41]
  wire  _T_3814 = _T_3732[5:0] == 6'h24; // @[lib.scala 199:41]
  wire  _T_3812 = _T_3732[5:0] == 6'h23; // @[lib.scala 199:41]
  wire  _T_3810 = _T_3732[5:0] == 6'h22; // @[lib.scala 199:41]
  wire  _T_3808 = _T_3732[5:0] == 6'h21; // @[lib.scala 199:41]
  wire  _T_3806 = _T_3732[5:0] == 6'h20; // @[lib.scala 199:41]
  wire  _T_3804 = _T_3732[5:0] == 6'h1f; // @[lib.scala 199:41]
  wire  _T_3802 = _T_3732[5:0] == 6'h1e; // @[lib.scala 199:41]
  wire [9:0] _T_3878 = {_T_3820,_T_3818,_T_3816,_T_3814,_T_3812,_T_3810,_T_3808,_T_3806,_T_3804,_T_3802}; // @[lib.scala 202:69]
  wire  _T_3800 = _T_3732[5:0] == 6'h1d; // @[lib.scala 199:41]
  wire  _T_3798 = _T_3732[5:0] == 6'h1c; // @[lib.scala 199:41]
  wire  _T_3796 = _T_3732[5:0] == 6'h1b; // @[lib.scala 199:41]
  wire  _T_3794 = _T_3732[5:0] == 6'h1a; // @[lib.scala 199:41]
  wire  _T_3792 = _T_3732[5:0] == 6'h19; // @[lib.scala 199:41]
  wire  _T_3790 = _T_3732[5:0] == 6'h18; // @[lib.scala 199:41]
  wire  _T_3788 = _T_3732[5:0] == 6'h17; // @[lib.scala 199:41]
  wire  _T_3786 = _T_3732[5:0] == 6'h16; // @[lib.scala 199:41]
  wire  _T_3784 = _T_3732[5:0] == 6'h15; // @[lib.scala 199:41]
  wire  _T_3782 = _T_3732[5:0] == 6'h14; // @[lib.scala 199:41]
  wire [9:0] _T_3869 = {_T_3800,_T_3798,_T_3796,_T_3794,_T_3792,_T_3790,_T_3788,_T_3786,_T_3784,_T_3782}; // @[lib.scala 202:69]
  wire  _T_3780 = _T_3732[5:0] == 6'h13; // @[lib.scala 199:41]
  wire  _T_3778 = _T_3732[5:0] == 6'h12; // @[lib.scala 199:41]
  wire  _T_3776 = _T_3732[5:0] == 6'h11; // @[lib.scala 199:41]
  wire  _T_3774 = _T_3732[5:0] == 6'h10; // @[lib.scala 199:41]
  wire  _T_3772 = _T_3732[5:0] == 6'hf; // @[lib.scala 199:41]
  wire  _T_3770 = _T_3732[5:0] == 6'he; // @[lib.scala 199:41]
  wire  _T_3768 = _T_3732[5:0] == 6'hd; // @[lib.scala 199:41]
  wire  _T_3766 = _T_3732[5:0] == 6'hc; // @[lib.scala 199:41]
  wire  _T_3764 = _T_3732[5:0] == 6'hb; // @[lib.scala 199:41]
  wire  _T_3762 = _T_3732[5:0] == 6'ha; // @[lib.scala 199:41]
  wire [9:0] _T_3859 = {_T_3780,_T_3778,_T_3776,_T_3774,_T_3772,_T_3770,_T_3768,_T_3766,_T_3764,_T_3762}; // @[lib.scala 202:69]
  wire  _T_3760 = _T_3732[5:0] == 6'h9; // @[lib.scala 199:41]
  wire  _T_3758 = _T_3732[5:0] == 6'h8; // @[lib.scala 199:41]
  wire  _T_3756 = _T_3732[5:0] == 6'h7; // @[lib.scala 199:41]
  wire  _T_3754 = _T_3732[5:0] == 6'h6; // @[lib.scala 199:41]
  wire  _T_3752 = _T_3732[5:0] == 6'h5; // @[lib.scala 199:41]
  wire  _T_3750 = _T_3732[5:0] == 6'h4; // @[lib.scala 199:41]
  wire  _T_3748 = _T_3732[5:0] == 6'h3; // @[lib.scala 199:41]
  wire  _T_3746 = _T_3732[5:0] == 6'h2; // @[lib.scala 199:41]
  wire  _T_3744 = _T_3732[5:0] == 6'h1; // @[lib.scala 199:41]
  wire [18:0] _T_3860 = {_T_3859,_T_3760,_T_3758,_T_3756,_T_3754,_T_3752,_T_3750,_T_3748,_T_3746,_T_3744}; // @[lib.scala 202:69]
  wire [38:0] _T_3880 = {_T_3878,_T_3869,_T_3860}; // @[lib.scala 202:69]
  wire [7:0] _T_3835 = {io_iccm_rd_data_ecc[74],io_iccm_rd_data_ecc[42:40],io_iccm_rd_data_ecc[73],io_iccm_rd_data_ecc[39],io_iccm_rd_data_ecc[72:71]}; // @[Cat.scala 29:58]
  wire [38:0] _T_3841 = {io_iccm_rd_data_ecc[77],io_iccm_rd_data_ecc[70:65],io_iccm_rd_data_ecc[76],io_iccm_rd_data_ecc[64:50],io_iccm_rd_data_ecc[75],io_iccm_rd_data_ecc[49:43],_T_3835}; // @[Cat.scala 29:58]
  wire [38:0] _T_3881 = _T_3880 ^ _T_3841; // @[lib.scala 202:76]
  wire [38:0] _T_3882 = _T_3736 ? _T_3881 : _T_3841; // @[lib.scala 202:31]
  wire [31:0] iccm_corrected_data_1 = {_T_3882[37:32],_T_3882[30:16],_T_3882[14:8],_T_3882[6:4],_T_3882[2]}; // @[Cat.scala 29:58]
  wire [31:0] iccm_dma_rdata_1_muxed = dma_mem_addr_ff[0] ? iccm_corrected_data_0 : iccm_corrected_data_1; // @[ifu_mem_ctl.scala 582:35]
  wire  _T_3740 = ~_T_3732[6]; // @[lib.scala 195:55]
  wire  _T_3741 = _T_3734 & _T_3740; // @[lib.scala 195:53]
  wire  _T_3355 = ~_T_3347[6]; // @[lib.scala 195:55]
  wire  _T_3356 = _T_3349 & _T_3355; // @[lib.scala 195:53]
  wire [1:0] iccm_double_ecc_error = {_T_3741,_T_3356}; // @[Cat.scala 29:58]
  wire  iccm_dma_ecc_error_in = |iccm_double_ecc_error; // @[ifu_mem_ctl.scala 584:53]
  wire [63:0] _T_3104 = {io_dma_mem_ctl_dma_mem_addr,io_dma_mem_ctl_dma_mem_addr}; // @[Cat.scala 29:58]
  wire [63:0] _T_3105 = {iccm_dma_rdata_1_muxed,_T_3497[37:32],_T_3497[30:16],_T_3497[14:8],_T_3497[6:4],_T_3497[2]}; // @[Cat.scala 29:58]
  reg [2:0] dma_mem_tag_ff; // @[ifu_mem_ctl.scala 586:54]
  reg [2:0] iccm_dma_rtag_temp; // @[ifu_mem_ctl.scala 587:74]
  reg  iccm_dma_rvalid_temp; // @[ifu_mem_ctl.scala 592:76]
  reg  iccm_dma_ecc_error; // @[ifu_mem_ctl.scala 594:74]
  reg [63:0] iccm_dma_rdata_temp; // @[ifu_mem_ctl.scala 596:75]
  wire  _T_3110 = _T_2709 & _T_2698; // @[ifu_mem_ctl.scala 599:77]
  wire  _T_3114 = _T_3091 & iccm_correct_ecc; // @[ifu_mem_ctl.scala 600:62]
  reg [13:0] iccm_ecc_corr_index_ff; // @[Reg.scala 27:20]
  wire [14:0] _T_3115 = {iccm_ecc_corr_index_ff,1'h0}; // @[Cat.scala 29:58]
  wire [14:0] _T_3117 = _T_3114 ? _T_3115 : io_ifc_fetch_addr_bf[14:0]; // @[ifu_mem_ctl.scala 600:8]
  wire  _T_3509 = _T_3347 == 7'h40; // @[lib.scala 205:62]
  wire  _T_3510 = _T_3497[38] ^ _T_3509; // @[lib.scala 205:44]
  wire [6:0] iccm_corrected_ecc_0 = {_T_3510,_T_3497[31],_T_3497[15],_T_3497[7],_T_3497[3],_T_3497[1:0]}; // @[Cat.scala 29:58]
  wire  _T_3894 = _T_3732 == 7'h40; // @[lib.scala 205:62]
  wire  _T_3895 = _T_3882[38] ^ _T_3894; // @[lib.scala 205:44]
  wire [6:0] iccm_corrected_ecc_1 = {_T_3895,_T_3882[31],_T_3882[15],_T_3882[7],_T_3882[3],_T_3882[1:0]}; // @[Cat.scala 29:58]
  wire  _T_3911 = _T_3 & ifc_iccm_access_f; // @[ifu_mem_ctl.scala 612:75]
  wire [31:0] iccm_corrected_data_f_mux = iccm_single_ecc_error[0] ? iccm_corrected_data_0 : iccm_corrected_data_1; // @[ifu_mem_ctl.scala 614:38]
  wire [6:0] iccm_corrected_ecc_f_mux = iccm_single_ecc_error[0] ? iccm_corrected_ecc_0 : iccm_corrected_ecc_1; // @[ifu_mem_ctl.scala 615:37]
  reg  iccm_rd_ecc_single_err_ff; // @[ifu_mem_ctl.scala 623:62]
  wire  _T_3919 = ~iccm_rd_ecc_single_err_ff; // @[ifu_mem_ctl.scala 617:93]
  wire  _T_3920 = io_dec_mem_ctrl_ifu_iccm_rd_ecc_single_err & _T_3919; // @[ifu_mem_ctl.scala 617:91]
  wire  _T_3922 = _T_3920 & _T_319; // @[ifu_mem_ctl.scala 617:121]
  wire  iccm_ecc_write_status = _T_3922 | io_iccm_dma_sb_error; // @[ifu_mem_ctl.scala 617:144]
  wire  _T_3923 = io_dec_mem_ctrl_ifu_iccm_rd_ecc_single_err | iccm_rd_ecc_single_err_ff; // @[ifu_mem_ctl.scala 618:84]
  reg [13:0] iccm_rw_addr_f; // @[ifu_mem_ctl.scala 622:51]
  wire [13:0] _T_3928 = iccm_rw_addr_f + 14'h1; // @[ifu_mem_ctl.scala 621:102]
  wire [38:0] _T_3932 = {iccm_corrected_ecc_f_mux,iccm_corrected_data_f_mux}; // @[Cat.scala 29:58]
  wire  _T_3937 = ~io_ifc_fetch_uncacheable_bf; // @[ifu_mem_ctl.scala 626:41]
  wire  _T_3938 = io_ifc_fetch_req_bf & _T_3937; // @[ifu_mem_ctl.scala 626:39]
  wire  _T_3939 = ~io_ifc_iccm_access_bf; // @[ifu_mem_ctl.scala 626:72]
  wire  _T_3940 = _T_3938 & _T_3939; // @[ifu_mem_ctl.scala 626:70]
  wire  _T_3942 = ~miss_state_en; // @[ifu_mem_ctl.scala 627:34]
  wire  _T_3943 = _T_2268 & _T_3942; // @[ifu_mem_ctl.scala 627:32]
  wire  _T_3946 = _T_2284 & _T_3942; // @[ifu_mem_ctl.scala 628:37]
  wire  _T_3947 = _T_3943 | _T_3946; // @[ifu_mem_ctl.scala 627:88]
  wire  _T_3948 = miss_state == 3'h7; // @[ifu_mem_ctl.scala 629:19]
  wire  _T_3950 = _T_3948 & _T_3942; // @[ifu_mem_ctl.scala 629:41]
  wire  _T_3951 = _T_3947 | _T_3950; // @[ifu_mem_ctl.scala 628:88]
  wire  _T_3952 = miss_state == 3'h3; // @[ifu_mem_ctl.scala 630:19]
  wire  _T_3954 = _T_3952 & _T_3942; // @[ifu_mem_ctl.scala 630:35]
  wire  _T_3955 = _T_3951 | _T_3954; // @[ifu_mem_ctl.scala 629:88]
  wire  _T_3958 = _T_2283 & _T_3942; // @[ifu_mem_ctl.scala 631:38]
  wire  _T_3959 = _T_3955 | _T_3958; // @[ifu_mem_ctl.scala 630:88]
  wire  _T_3961 = _T_2284 & miss_state_en; // @[ifu_mem_ctl.scala 632:37]
  wire  _T_3962 = miss_nxtstate == 3'h3; // @[ifu_mem_ctl.scala 632:71]
  wire  _T_3963 = _T_3961 & _T_3962; // @[ifu_mem_ctl.scala 632:54]
  wire  _T_3964 = _T_3959 | _T_3963; // @[ifu_mem_ctl.scala 631:57]
  wire  _T_3965 = ~_T_3964; // @[ifu_mem_ctl.scala 627:5]
  wire  _T_3966 = _T_3940 & _T_3965; // @[ifu_mem_ctl.scala 626:96]
  wire  _T_3967 = io_ifc_fetch_req_bf & io_exu_flush_final; // @[ifu_mem_ctl.scala 633:28]
  wire  _T_3969 = _T_3967 & _T_3937; // @[ifu_mem_ctl.scala 633:50]
  wire  _T_3971 = _T_3969 & _T_3939; // @[ifu_mem_ctl.scala 633:81]
  wire [1:0] _T_3974 = write_ic_16_bytes ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire  _T_9780 = bus_ifu_wr_en_ff_q & replace_way_mb_any_1; // @[ifu_mem_ctl.scala 727:74]
  wire  bus_wren_1 = _T_9780 & miss_pending; // @[ifu_mem_ctl.scala 727:98]
  wire  _T_9779 = bus_ifu_wr_en_ff_q & replace_way_mb_any_0; // @[ifu_mem_ctl.scala 727:74]
  wire  bus_wren_0 = _T_9779 & miss_pending; // @[ifu_mem_ctl.scala 727:98]
  wire [1:0] bus_ic_wr_en = {bus_wren_1,bus_wren_0}; // @[Cat.scala 29:58]
  wire  _T_3980 = ~_T_108; // @[ifu_mem_ctl.scala 636:106]
  wire  _T_3981 = _T_2268 & _T_3980; // @[ifu_mem_ctl.scala 636:104]
  wire  _T_3982 = _T_2284 | _T_3981; // @[ifu_mem_ctl.scala 636:77]
  wire  _T_3986 = ~_T_51; // @[ifu_mem_ctl.scala 636:172]
  wire  _T_3987 = _T_3982 & _T_3986; // @[ifu_mem_ctl.scala 636:170]
  wire  _T_3988 = ~_T_3987; // @[ifu_mem_ctl.scala 636:44]
  wire  _T_3992 = reset_ic_in | reset_ic_ff; // @[ifu_mem_ctl.scala 639:64]
  wire  _T_3993 = ~_T_3992; // @[ifu_mem_ctl.scala 639:50]
  wire  _T_3994 = _T_276 & _T_3993; // @[ifu_mem_ctl.scala 639:48]
  wire  _T_3995 = ~reset_tag_valid_for_miss; // @[ifu_mem_ctl.scala 639:81]
  wire  ic_valid = _T_3994 & _T_3995; // @[ifu_mem_ctl.scala 639:79]
  wire  _T_3997 = debug_c1_clken & io_ic_debug_tag_array; // @[ifu_mem_ctl.scala 640:82]
  reg [6:0] ifu_status_wr_addr_ff; // @[ifu_mem_ctl.scala 643:14]
  wire  _T_4000 = io_ic_debug_wr_en & io_ic_debug_tag_array; // @[ifu_mem_ctl.scala 646:74]
  wire  _T_9777 = bus_ifu_wr_en_ff_q & last_beat; // @[ifu_mem_ctl.scala 726:45]
  wire  way_status_wr_en = _T_9777 | ic_act_hit_f; // @[ifu_mem_ctl.scala 726:58]
  reg  way_status_wr_en_ff; // @[ifu_mem_ctl.scala 648:14]
  wire  way_status_hit_new = io_ic_rd_hit[0]; // @[ifu_mem_ctl.scala 722:41]
  reg  way_status_new_ff; // @[ifu_mem_ctl.scala 654:14]
  wire  _T_4020 = ifu_status_wr_addr_ff[2:0] == 3'h0; // @[ifu_mem_ctl.scala 660:128]
  wire  _T_4021 = _T_4020 & way_status_wr_en_ff; // @[ifu_mem_ctl.scala 660:136]
  wire  _T_4024 = ifu_status_wr_addr_ff[2:0] == 3'h1; // @[ifu_mem_ctl.scala 660:128]
  wire  _T_4025 = _T_4024 & way_status_wr_en_ff; // @[ifu_mem_ctl.scala 660:136]
  wire  _T_4028 = ifu_status_wr_addr_ff[2:0] == 3'h2; // @[ifu_mem_ctl.scala 660:128]
  wire  _T_4029 = _T_4028 & way_status_wr_en_ff; // @[ifu_mem_ctl.scala 660:136]
  wire  _T_4032 = ifu_status_wr_addr_ff[2:0] == 3'h3; // @[ifu_mem_ctl.scala 660:128]
  wire  _T_4033 = _T_4032 & way_status_wr_en_ff; // @[ifu_mem_ctl.scala 660:136]
  wire  _T_4036 = ifu_status_wr_addr_ff[2:0] == 3'h4; // @[ifu_mem_ctl.scala 660:128]
  wire  _T_4037 = _T_4036 & way_status_wr_en_ff; // @[ifu_mem_ctl.scala 660:136]
  wire  _T_4040 = ifu_status_wr_addr_ff[2:0] == 3'h5; // @[ifu_mem_ctl.scala 660:128]
  wire  _T_4041 = _T_4040 & way_status_wr_en_ff; // @[ifu_mem_ctl.scala 660:136]
  wire  _T_4044 = ifu_status_wr_addr_ff[2:0] == 3'h6; // @[ifu_mem_ctl.scala 660:128]
  wire  _T_4045 = _T_4044 & way_status_wr_en_ff; // @[ifu_mem_ctl.scala 660:136]
  wire  _T_4048 = ifu_status_wr_addr_ff[2:0] == 3'h7; // @[ifu_mem_ctl.scala 660:128]
  wire  _T_4049 = _T_4048 & way_status_wr_en_ff; // @[ifu_mem_ctl.scala 660:136]
  wire  _T_9783 = _T_100 & replace_way_mb_any_1; // @[ifu_mem_ctl.scala 729:84]
  wire  _T_9784 = _T_9783 & miss_pending; // @[ifu_mem_ctl.scala 729:108]
  wire  bus_wren_last_1 = _T_9784 & bus_last_data_beat; // @[ifu_mem_ctl.scala 729:123]
  wire  wren_reset_miss_1 = replace_way_mb_any_1 & reset_tag_valid_for_miss; // @[ifu_mem_ctl.scala 730:84]
  wire  _T_9786 = bus_wren_last_1 | wren_reset_miss_1; // @[ifu_mem_ctl.scala 731:73]
  wire  _T_9781 = _T_100 & replace_way_mb_any_0; // @[ifu_mem_ctl.scala 729:84]
  wire  _T_9782 = _T_9781 & miss_pending; // @[ifu_mem_ctl.scala 729:108]
  wire  bus_wren_last_0 = _T_9782 & bus_last_data_beat; // @[ifu_mem_ctl.scala 729:123]
  wire  wren_reset_miss_0 = replace_way_mb_any_0 & reset_tag_valid_for_miss; // @[ifu_mem_ctl.scala 730:84]
  wire  _T_9785 = bus_wren_last_0 | wren_reset_miss_0; // @[ifu_mem_ctl.scala 731:73]
  wire [1:0] ifu_tag_wren = {_T_9786,_T_9785}; // @[Cat.scala 29:58]
  wire [1:0] _T_9821 = _T_4000 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [1:0] ic_debug_tag_wr_en = _T_9821 & io_ic_debug_way; // @[ifu_mem_ctl.scala 765:90]
  reg [1:0] ifu_tag_wren_ff; // @[ifu_mem_ctl.scala 675:14]
  reg  ic_valid_ff; // @[ifu_mem_ctl.scala 679:14]
  wire  _T_5063 = ifu_ic_rw_int_addr_ff[6:5] == 2'h0; // @[ifu_mem_ctl.scala 683:78]
  wire  _T_5065 = _T_5063 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 683:87]
  wire  _T_5067 = perr_ic_index_ff[6:5] == 2'h0; // @[ifu_mem_ctl.scala 684:70]
  wire  _T_5069 = _T_5067 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 684:79]
  wire  _T_5070 = _T_5065 | _T_5069; // @[ifu_mem_ctl.scala 683:109]
  wire  _T_5071 = _T_5070 | reset_all_tags; // @[ifu_mem_ctl.scala 684:102]
  wire  _T_5075 = _T_5063 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 683:87]
  wire  _T_5079 = _T_5067 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 684:79]
  wire  _T_5080 = _T_5075 | _T_5079; // @[ifu_mem_ctl.scala 683:109]
  wire  _T_5081 = _T_5080 | reset_all_tags; // @[ifu_mem_ctl.scala 684:102]
  wire [1:0] tag_valid_clken_0 = {_T_5081,_T_5071}; // @[Cat.scala 29:58]
  wire  _T_5083 = ifu_ic_rw_int_addr_ff[6:5] == 2'h1; // @[ifu_mem_ctl.scala 683:78]
  wire  _T_5085 = _T_5083 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 683:87]
  wire  _T_5087 = perr_ic_index_ff[6:5] == 2'h1; // @[ifu_mem_ctl.scala 684:70]
  wire  _T_5089 = _T_5087 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 684:79]
  wire  _T_5090 = _T_5085 | _T_5089; // @[ifu_mem_ctl.scala 683:109]
  wire  _T_5091 = _T_5090 | reset_all_tags; // @[ifu_mem_ctl.scala 684:102]
  wire  _T_5095 = _T_5083 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 683:87]
  wire  _T_5099 = _T_5087 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 684:79]
  wire  _T_5100 = _T_5095 | _T_5099; // @[ifu_mem_ctl.scala 683:109]
  wire  _T_5101 = _T_5100 | reset_all_tags; // @[ifu_mem_ctl.scala 684:102]
  wire [1:0] tag_valid_clken_1 = {_T_5101,_T_5091}; // @[Cat.scala 29:58]
  wire  _T_5103 = ifu_ic_rw_int_addr_ff[6:5] == 2'h2; // @[ifu_mem_ctl.scala 683:78]
  wire  _T_5105 = _T_5103 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 683:87]
  wire  _T_5107 = perr_ic_index_ff[6:5] == 2'h2; // @[ifu_mem_ctl.scala 684:70]
  wire  _T_5109 = _T_5107 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 684:79]
  wire  _T_5110 = _T_5105 | _T_5109; // @[ifu_mem_ctl.scala 683:109]
  wire  _T_5111 = _T_5110 | reset_all_tags; // @[ifu_mem_ctl.scala 684:102]
  wire  _T_5115 = _T_5103 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 683:87]
  wire  _T_5119 = _T_5107 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 684:79]
  wire  _T_5120 = _T_5115 | _T_5119; // @[ifu_mem_ctl.scala 683:109]
  wire  _T_5121 = _T_5120 | reset_all_tags; // @[ifu_mem_ctl.scala 684:102]
  wire [1:0] tag_valid_clken_2 = {_T_5121,_T_5111}; // @[Cat.scala 29:58]
  wire  _T_5123 = ifu_ic_rw_int_addr_ff[6:5] == 2'h3; // @[ifu_mem_ctl.scala 683:78]
  wire  _T_5125 = _T_5123 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 683:87]
  wire  _T_5127 = perr_ic_index_ff[6:5] == 2'h3; // @[ifu_mem_ctl.scala 684:70]
  wire  _T_5129 = _T_5127 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 684:79]
  wire  _T_5130 = _T_5125 | _T_5129; // @[ifu_mem_ctl.scala 683:109]
  wire  _T_5131 = _T_5130 | reset_all_tags; // @[ifu_mem_ctl.scala 684:102]
  wire  _T_5135 = _T_5123 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 683:87]
  wire  _T_5139 = _T_5127 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 684:79]
  wire  _T_5140 = _T_5135 | _T_5139; // @[ifu_mem_ctl.scala 683:109]
  wire  _T_5141 = _T_5140 | reset_all_tags; // @[ifu_mem_ctl.scala 684:102]
  wire [1:0] tag_valid_clken_3 = {_T_5141,_T_5131}; // @[Cat.scala 29:58]
  wire  _T_5152 = ic_valid_ff & _T_195; // @[ifu_mem_ctl.scala 692:97]
  wire  _T_5153 = ~perr_sel_invalidate; // @[ifu_mem_ctl.scala 692:124]
  wire  _T_5154 = _T_5152 & _T_5153; // @[ifu_mem_ctl.scala 692:122]
  wire  _T_5157 = _T_4671 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_5158 = perr_ic_index_ff == 7'h0; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_5160 = _T_5158 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_5161 = _T_5157 | _T_5160; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_5162 = _T_5161 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_5172 = _T_4672 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_5173 = perr_ic_index_ff == 7'h1; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_5175 = _T_5173 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_5176 = _T_5172 | _T_5175; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_5177 = _T_5176 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_5187 = _T_4673 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_5188 = perr_ic_index_ff == 7'h2; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_5190 = _T_5188 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_5191 = _T_5187 | _T_5190; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_5192 = _T_5191 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_5202 = _T_4674 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_5203 = perr_ic_index_ff == 7'h3; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_5205 = _T_5203 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_5206 = _T_5202 | _T_5205; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_5207 = _T_5206 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_5217 = _T_4675 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_5218 = perr_ic_index_ff == 7'h4; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_5220 = _T_5218 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_5221 = _T_5217 | _T_5220; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_5222 = _T_5221 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_5232 = _T_4676 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_5233 = perr_ic_index_ff == 7'h5; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_5235 = _T_5233 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_5236 = _T_5232 | _T_5235; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_5237 = _T_5236 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_5247 = _T_4677 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_5248 = perr_ic_index_ff == 7'h6; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_5250 = _T_5248 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_5251 = _T_5247 | _T_5250; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_5252 = _T_5251 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_5262 = _T_4678 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_5263 = perr_ic_index_ff == 7'h7; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_5265 = _T_5263 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_5266 = _T_5262 | _T_5265; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_5267 = _T_5266 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_5277 = _T_4679 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_5278 = perr_ic_index_ff == 7'h8; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_5280 = _T_5278 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_5281 = _T_5277 | _T_5280; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_5282 = _T_5281 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_5292 = _T_4680 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_5293 = perr_ic_index_ff == 7'h9; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_5295 = _T_5293 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_5296 = _T_5292 | _T_5295; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_5297 = _T_5296 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_5307 = _T_4681 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_5308 = perr_ic_index_ff == 7'ha; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_5310 = _T_5308 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_5311 = _T_5307 | _T_5310; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_5312 = _T_5311 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_5322 = _T_4682 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_5323 = perr_ic_index_ff == 7'hb; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_5325 = _T_5323 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_5326 = _T_5322 | _T_5325; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_5327 = _T_5326 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_5337 = _T_4683 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_5338 = perr_ic_index_ff == 7'hc; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_5340 = _T_5338 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_5341 = _T_5337 | _T_5340; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_5342 = _T_5341 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_5352 = _T_4684 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_5353 = perr_ic_index_ff == 7'hd; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_5355 = _T_5353 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_5356 = _T_5352 | _T_5355; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_5357 = _T_5356 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_5367 = _T_4685 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_5368 = perr_ic_index_ff == 7'he; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_5370 = _T_5368 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_5371 = _T_5367 | _T_5370; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_5372 = _T_5371 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_5382 = _T_4686 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_5383 = perr_ic_index_ff == 7'hf; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_5385 = _T_5383 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_5386 = _T_5382 | _T_5385; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_5387 = _T_5386 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_5397 = _T_4687 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_5398 = perr_ic_index_ff == 7'h10; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_5400 = _T_5398 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_5401 = _T_5397 | _T_5400; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_5402 = _T_5401 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_5412 = _T_4688 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_5413 = perr_ic_index_ff == 7'h11; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_5415 = _T_5413 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_5416 = _T_5412 | _T_5415; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_5417 = _T_5416 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_5427 = _T_4689 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_5428 = perr_ic_index_ff == 7'h12; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_5430 = _T_5428 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_5431 = _T_5427 | _T_5430; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_5432 = _T_5431 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_5442 = _T_4690 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_5443 = perr_ic_index_ff == 7'h13; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_5445 = _T_5443 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_5446 = _T_5442 | _T_5445; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_5447 = _T_5446 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_5457 = _T_4691 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_5458 = perr_ic_index_ff == 7'h14; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_5460 = _T_5458 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_5461 = _T_5457 | _T_5460; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_5462 = _T_5461 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_5472 = _T_4692 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_5473 = perr_ic_index_ff == 7'h15; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_5475 = _T_5473 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_5476 = _T_5472 | _T_5475; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_5477 = _T_5476 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_5487 = _T_4693 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_5488 = perr_ic_index_ff == 7'h16; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_5490 = _T_5488 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_5491 = _T_5487 | _T_5490; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_5492 = _T_5491 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_5502 = _T_4694 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_5503 = perr_ic_index_ff == 7'h17; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_5505 = _T_5503 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_5506 = _T_5502 | _T_5505; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_5507 = _T_5506 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_5517 = _T_4695 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_5518 = perr_ic_index_ff == 7'h18; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_5520 = _T_5518 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_5521 = _T_5517 | _T_5520; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_5522 = _T_5521 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_5532 = _T_4696 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_5533 = perr_ic_index_ff == 7'h19; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_5535 = _T_5533 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_5536 = _T_5532 | _T_5535; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_5537 = _T_5536 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_5547 = _T_4697 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_5548 = perr_ic_index_ff == 7'h1a; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_5550 = _T_5548 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_5551 = _T_5547 | _T_5550; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_5552 = _T_5551 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_5562 = _T_4698 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_5563 = perr_ic_index_ff == 7'h1b; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_5565 = _T_5563 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_5566 = _T_5562 | _T_5565; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_5567 = _T_5566 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_5577 = _T_4699 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_5578 = perr_ic_index_ff == 7'h1c; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_5580 = _T_5578 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_5581 = _T_5577 | _T_5580; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_5582 = _T_5581 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_5592 = _T_4700 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_5593 = perr_ic_index_ff == 7'h1d; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_5595 = _T_5593 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_5596 = _T_5592 | _T_5595; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_5597 = _T_5596 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_5607 = _T_4701 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_5608 = perr_ic_index_ff == 7'h1e; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_5610 = _T_5608 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_5611 = _T_5607 | _T_5610; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_5612 = _T_5611 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_5622 = _T_4702 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_5623 = perr_ic_index_ff == 7'h1f; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_5625 = _T_5623 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_5626 = _T_5622 | _T_5625; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_5627 = _T_5626 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_5637 = _T_4671 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_5640 = _T_5158 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_5641 = _T_5637 | _T_5640; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_5642 = _T_5641 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_5652 = _T_4672 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_5655 = _T_5173 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_5656 = _T_5652 | _T_5655; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_5657 = _T_5656 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_5667 = _T_4673 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_5670 = _T_5188 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_5671 = _T_5667 | _T_5670; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_5672 = _T_5671 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_5682 = _T_4674 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_5685 = _T_5203 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_5686 = _T_5682 | _T_5685; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_5687 = _T_5686 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_5697 = _T_4675 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_5700 = _T_5218 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_5701 = _T_5697 | _T_5700; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_5702 = _T_5701 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_5712 = _T_4676 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_5715 = _T_5233 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_5716 = _T_5712 | _T_5715; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_5717 = _T_5716 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_5727 = _T_4677 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_5730 = _T_5248 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_5731 = _T_5727 | _T_5730; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_5732 = _T_5731 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_5742 = _T_4678 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_5745 = _T_5263 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_5746 = _T_5742 | _T_5745; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_5747 = _T_5746 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_5757 = _T_4679 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_5760 = _T_5278 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_5761 = _T_5757 | _T_5760; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_5762 = _T_5761 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_5772 = _T_4680 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_5775 = _T_5293 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_5776 = _T_5772 | _T_5775; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_5777 = _T_5776 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_5787 = _T_4681 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_5790 = _T_5308 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_5791 = _T_5787 | _T_5790; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_5792 = _T_5791 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_5802 = _T_4682 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_5805 = _T_5323 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_5806 = _T_5802 | _T_5805; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_5807 = _T_5806 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_5817 = _T_4683 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_5820 = _T_5338 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_5821 = _T_5817 | _T_5820; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_5822 = _T_5821 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_5832 = _T_4684 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_5835 = _T_5353 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_5836 = _T_5832 | _T_5835; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_5837 = _T_5836 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_5847 = _T_4685 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_5850 = _T_5368 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_5851 = _T_5847 | _T_5850; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_5852 = _T_5851 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_5862 = _T_4686 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_5865 = _T_5383 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_5866 = _T_5862 | _T_5865; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_5867 = _T_5866 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_5877 = _T_4687 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_5880 = _T_5398 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_5881 = _T_5877 | _T_5880; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_5882 = _T_5881 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_5892 = _T_4688 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_5895 = _T_5413 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_5896 = _T_5892 | _T_5895; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_5897 = _T_5896 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_5907 = _T_4689 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_5910 = _T_5428 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_5911 = _T_5907 | _T_5910; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_5912 = _T_5911 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_5922 = _T_4690 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_5925 = _T_5443 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_5926 = _T_5922 | _T_5925; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_5927 = _T_5926 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_5937 = _T_4691 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_5940 = _T_5458 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_5941 = _T_5937 | _T_5940; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_5942 = _T_5941 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_5952 = _T_4692 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_5955 = _T_5473 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_5956 = _T_5952 | _T_5955; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_5957 = _T_5956 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_5967 = _T_4693 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_5970 = _T_5488 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_5971 = _T_5967 | _T_5970; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_5972 = _T_5971 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_5982 = _T_4694 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_5985 = _T_5503 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_5986 = _T_5982 | _T_5985; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_5987 = _T_5986 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_5997 = _T_4695 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6000 = _T_5518 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6001 = _T_5997 | _T_6000; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6002 = _T_6001 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6012 = _T_4696 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6015 = _T_5533 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6016 = _T_6012 | _T_6015; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6017 = _T_6016 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6027 = _T_4697 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6030 = _T_5548 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6031 = _T_6027 | _T_6030; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6032 = _T_6031 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6042 = _T_4698 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6045 = _T_5563 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6046 = _T_6042 | _T_6045; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6047 = _T_6046 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6057 = _T_4699 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6060 = _T_5578 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6061 = _T_6057 | _T_6060; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6062 = _T_6061 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6072 = _T_4700 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6075 = _T_5593 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6076 = _T_6072 | _T_6075; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6077 = _T_6076 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6087 = _T_4701 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6090 = _T_5608 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6091 = _T_6087 | _T_6090; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6092 = _T_6091 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6102 = _T_4702 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6105 = _T_5623 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6106 = _T_6102 | _T_6105; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6107 = _T_6106 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6117 = _T_4703 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6118 = perr_ic_index_ff == 7'h20; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_6120 = _T_6118 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6121 = _T_6117 | _T_6120; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6122 = _T_6121 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6132 = _T_4704 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6133 = perr_ic_index_ff == 7'h21; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_6135 = _T_6133 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6136 = _T_6132 | _T_6135; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6137 = _T_6136 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6147 = _T_4705 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6148 = perr_ic_index_ff == 7'h22; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_6150 = _T_6148 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6151 = _T_6147 | _T_6150; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6152 = _T_6151 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6162 = _T_4706 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6163 = perr_ic_index_ff == 7'h23; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_6165 = _T_6163 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6166 = _T_6162 | _T_6165; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6167 = _T_6166 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6177 = _T_4707 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6178 = perr_ic_index_ff == 7'h24; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_6180 = _T_6178 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6181 = _T_6177 | _T_6180; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6182 = _T_6181 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6192 = _T_4708 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6193 = perr_ic_index_ff == 7'h25; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_6195 = _T_6193 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6196 = _T_6192 | _T_6195; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6197 = _T_6196 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6207 = _T_4709 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6208 = perr_ic_index_ff == 7'h26; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_6210 = _T_6208 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6211 = _T_6207 | _T_6210; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6212 = _T_6211 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6222 = _T_4710 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6223 = perr_ic_index_ff == 7'h27; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_6225 = _T_6223 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6226 = _T_6222 | _T_6225; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6227 = _T_6226 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6237 = _T_4711 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6238 = perr_ic_index_ff == 7'h28; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_6240 = _T_6238 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6241 = _T_6237 | _T_6240; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6242 = _T_6241 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6252 = _T_4712 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6253 = perr_ic_index_ff == 7'h29; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_6255 = _T_6253 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6256 = _T_6252 | _T_6255; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6257 = _T_6256 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6267 = _T_4713 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6268 = perr_ic_index_ff == 7'h2a; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_6270 = _T_6268 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6271 = _T_6267 | _T_6270; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6272 = _T_6271 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6282 = _T_4714 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6283 = perr_ic_index_ff == 7'h2b; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_6285 = _T_6283 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6286 = _T_6282 | _T_6285; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6287 = _T_6286 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6297 = _T_4715 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6298 = perr_ic_index_ff == 7'h2c; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_6300 = _T_6298 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6301 = _T_6297 | _T_6300; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6302 = _T_6301 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6312 = _T_4716 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6313 = perr_ic_index_ff == 7'h2d; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_6315 = _T_6313 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6316 = _T_6312 | _T_6315; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6317 = _T_6316 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6327 = _T_4717 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6328 = perr_ic_index_ff == 7'h2e; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_6330 = _T_6328 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6331 = _T_6327 | _T_6330; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6332 = _T_6331 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6342 = _T_4718 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6343 = perr_ic_index_ff == 7'h2f; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_6345 = _T_6343 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6346 = _T_6342 | _T_6345; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6347 = _T_6346 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6357 = _T_4719 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6358 = perr_ic_index_ff == 7'h30; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_6360 = _T_6358 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6361 = _T_6357 | _T_6360; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6362 = _T_6361 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6372 = _T_4720 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6373 = perr_ic_index_ff == 7'h31; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_6375 = _T_6373 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6376 = _T_6372 | _T_6375; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6377 = _T_6376 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6387 = _T_4721 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6388 = perr_ic_index_ff == 7'h32; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_6390 = _T_6388 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6391 = _T_6387 | _T_6390; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6392 = _T_6391 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6402 = _T_4722 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6403 = perr_ic_index_ff == 7'h33; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_6405 = _T_6403 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6406 = _T_6402 | _T_6405; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6407 = _T_6406 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6417 = _T_4723 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6418 = perr_ic_index_ff == 7'h34; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_6420 = _T_6418 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6421 = _T_6417 | _T_6420; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6422 = _T_6421 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6432 = _T_4724 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6433 = perr_ic_index_ff == 7'h35; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_6435 = _T_6433 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6436 = _T_6432 | _T_6435; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6437 = _T_6436 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6447 = _T_4725 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6448 = perr_ic_index_ff == 7'h36; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_6450 = _T_6448 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6451 = _T_6447 | _T_6450; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6452 = _T_6451 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6462 = _T_4726 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6463 = perr_ic_index_ff == 7'h37; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_6465 = _T_6463 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6466 = _T_6462 | _T_6465; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6467 = _T_6466 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6477 = _T_4727 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6478 = perr_ic_index_ff == 7'h38; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_6480 = _T_6478 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6481 = _T_6477 | _T_6480; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6482 = _T_6481 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6492 = _T_4728 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6493 = perr_ic_index_ff == 7'h39; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_6495 = _T_6493 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6496 = _T_6492 | _T_6495; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6497 = _T_6496 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6507 = _T_4729 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6508 = perr_ic_index_ff == 7'h3a; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_6510 = _T_6508 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6511 = _T_6507 | _T_6510; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6512 = _T_6511 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6522 = _T_4730 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6523 = perr_ic_index_ff == 7'h3b; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_6525 = _T_6523 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6526 = _T_6522 | _T_6525; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6527 = _T_6526 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6537 = _T_4731 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6538 = perr_ic_index_ff == 7'h3c; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_6540 = _T_6538 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6541 = _T_6537 | _T_6540; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6542 = _T_6541 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6552 = _T_4732 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6553 = perr_ic_index_ff == 7'h3d; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_6555 = _T_6553 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6556 = _T_6552 | _T_6555; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6557 = _T_6556 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6567 = _T_4733 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6568 = perr_ic_index_ff == 7'h3e; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_6570 = _T_6568 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6571 = _T_6567 | _T_6570; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6572 = _T_6571 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6582 = _T_4734 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6583 = perr_ic_index_ff == 7'h3f; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_6585 = _T_6583 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6586 = _T_6582 | _T_6585; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6587 = _T_6586 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6597 = _T_4703 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6600 = _T_6118 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6601 = _T_6597 | _T_6600; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6602 = _T_6601 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6612 = _T_4704 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6615 = _T_6133 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6616 = _T_6612 | _T_6615; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6617 = _T_6616 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6627 = _T_4705 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6630 = _T_6148 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6631 = _T_6627 | _T_6630; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6632 = _T_6631 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6642 = _T_4706 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6645 = _T_6163 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6646 = _T_6642 | _T_6645; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6647 = _T_6646 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6657 = _T_4707 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6660 = _T_6178 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6661 = _T_6657 | _T_6660; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6662 = _T_6661 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6672 = _T_4708 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6675 = _T_6193 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6676 = _T_6672 | _T_6675; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6677 = _T_6676 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6687 = _T_4709 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6690 = _T_6208 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6691 = _T_6687 | _T_6690; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6692 = _T_6691 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6702 = _T_4710 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6705 = _T_6223 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6706 = _T_6702 | _T_6705; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6707 = _T_6706 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6717 = _T_4711 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6720 = _T_6238 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6721 = _T_6717 | _T_6720; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6722 = _T_6721 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6732 = _T_4712 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6735 = _T_6253 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6736 = _T_6732 | _T_6735; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6737 = _T_6736 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6747 = _T_4713 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6750 = _T_6268 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6751 = _T_6747 | _T_6750; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6752 = _T_6751 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6762 = _T_4714 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6765 = _T_6283 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6766 = _T_6762 | _T_6765; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6767 = _T_6766 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6777 = _T_4715 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6780 = _T_6298 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6781 = _T_6777 | _T_6780; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6782 = _T_6781 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6792 = _T_4716 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6795 = _T_6313 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6796 = _T_6792 | _T_6795; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6797 = _T_6796 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6807 = _T_4717 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6810 = _T_6328 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6811 = _T_6807 | _T_6810; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6812 = _T_6811 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6822 = _T_4718 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6825 = _T_6343 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6826 = _T_6822 | _T_6825; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6827 = _T_6826 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6837 = _T_4719 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6840 = _T_6358 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6841 = _T_6837 | _T_6840; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6842 = _T_6841 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6852 = _T_4720 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6855 = _T_6373 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6856 = _T_6852 | _T_6855; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6857 = _T_6856 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6867 = _T_4721 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6870 = _T_6388 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6871 = _T_6867 | _T_6870; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6872 = _T_6871 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6882 = _T_4722 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6885 = _T_6403 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6886 = _T_6882 | _T_6885; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6887 = _T_6886 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6897 = _T_4723 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6900 = _T_6418 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6901 = _T_6897 | _T_6900; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6902 = _T_6901 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6912 = _T_4724 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6915 = _T_6433 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6916 = _T_6912 | _T_6915; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6917 = _T_6916 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6927 = _T_4725 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6930 = _T_6448 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6931 = _T_6927 | _T_6930; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6932 = _T_6931 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6942 = _T_4726 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6945 = _T_6463 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6946 = _T_6942 | _T_6945; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6947 = _T_6946 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6957 = _T_4727 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6960 = _T_6478 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6961 = _T_6957 | _T_6960; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6962 = _T_6961 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6972 = _T_4728 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6975 = _T_6493 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6976 = _T_6972 | _T_6975; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6977 = _T_6976 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_6987 = _T_4729 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_6990 = _T_6508 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_6991 = _T_6987 | _T_6990; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_6992 = _T_6991 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7002 = _T_4730 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7005 = _T_6523 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7006 = _T_7002 | _T_7005; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7007 = _T_7006 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7017 = _T_4731 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7020 = _T_6538 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7021 = _T_7017 | _T_7020; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7022 = _T_7021 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7032 = _T_4732 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7035 = _T_6553 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7036 = _T_7032 | _T_7035; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7037 = _T_7036 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7047 = _T_4733 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7050 = _T_6568 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7051 = _T_7047 | _T_7050; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7052 = _T_7051 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7062 = _T_4734 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7065 = _T_6583 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7066 = _T_7062 | _T_7065; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7067 = _T_7066 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7077 = _T_4735 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7078 = perr_ic_index_ff == 7'h40; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_7080 = _T_7078 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7081 = _T_7077 | _T_7080; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7082 = _T_7081 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7092 = _T_4736 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7093 = perr_ic_index_ff == 7'h41; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_7095 = _T_7093 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7096 = _T_7092 | _T_7095; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7097 = _T_7096 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7107 = _T_4737 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7108 = perr_ic_index_ff == 7'h42; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_7110 = _T_7108 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7111 = _T_7107 | _T_7110; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7112 = _T_7111 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7122 = _T_4738 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7123 = perr_ic_index_ff == 7'h43; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_7125 = _T_7123 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7126 = _T_7122 | _T_7125; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7127 = _T_7126 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7137 = _T_4739 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7138 = perr_ic_index_ff == 7'h44; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_7140 = _T_7138 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7141 = _T_7137 | _T_7140; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7142 = _T_7141 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7152 = _T_4740 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7153 = perr_ic_index_ff == 7'h45; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_7155 = _T_7153 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7156 = _T_7152 | _T_7155; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7157 = _T_7156 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7167 = _T_4741 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7168 = perr_ic_index_ff == 7'h46; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_7170 = _T_7168 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7171 = _T_7167 | _T_7170; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7172 = _T_7171 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7182 = _T_4742 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7183 = perr_ic_index_ff == 7'h47; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_7185 = _T_7183 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7186 = _T_7182 | _T_7185; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7187 = _T_7186 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7197 = _T_4743 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7198 = perr_ic_index_ff == 7'h48; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_7200 = _T_7198 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7201 = _T_7197 | _T_7200; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7202 = _T_7201 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7212 = _T_4744 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7213 = perr_ic_index_ff == 7'h49; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_7215 = _T_7213 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7216 = _T_7212 | _T_7215; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7217 = _T_7216 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7227 = _T_4745 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7228 = perr_ic_index_ff == 7'h4a; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_7230 = _T_7228 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7231 = _T_7227 | _T_7230; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7232 = _T_7231 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7242 = _T_4746 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7243 = perr_ic_index_ff == 7'h4b; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_7245 = _T_7243 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7246 = _T_7242 | _T_7245; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7247 = _T_7246 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7257 = _T_4747 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7258 = perr_ic_index_ff == 7'h4c; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_7260 = _T_7258 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7261 = _T_7257 | _T_7260; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7262 = _T_7261 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7272 = _T_4748 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7273 = perr_ic_index_ff == 7'h4d; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_7275 = _T_7273 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7276 = _T_7272 | _T_7275; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7277 = _T_7276 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7287 = _T_4749 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7288 = perr_ic_index_ff == 7'h4e; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_7290 = _T_7288 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7291 = _T_7287 | _T_7290; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7292 = _T_7291 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7302 = _T_4750 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7303 = perr_ic_index_ff == 7'h4f; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_7305 = _T_7303 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7306 = _T_7302 | _T_7305; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7307 = _T_7306 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7317 = _T_4751 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7318 = perr_ic_index_ff == 7'h50; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_7320 = _T_7318 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7321 = _T_7317 | _T_7320; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7322 = _T_7321 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7332 = _T_4752 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7333 = perr_ic_index_ff == 7'h51; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_7335 = _T_7333 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7336 = _T_7332 | _T_7335; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7337 = _T_7336 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7347 = _T_4753 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7348 = perr_ic_index_ff == 7'h52; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_7350 = _T_7348 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7351 = _T_7347 | _T_7350; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7352 = _T_7351 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7362 = _T_4754 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7363 = perr_ic_index_ff == 7'h53; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_7365 = _T_7363 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7366 = _T_7362 | _T_7365; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7367 = _T_7366 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7377 = _T_4755 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7378 = perr_ic_index_ff == 7'h54; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_7380 = _T_7378 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7381 = _T_7377 | _T_7380; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7382 = _T_7381 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7392 = _T_4756 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7393 = perr_ic_index_ff == 7'h55; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_7395 = _T_7393 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7396 = _T_7392 | _T_7395; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7397 = _T_7396 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7407 = _T_4757 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7408 = perr_ic_index_ff == 7'h56; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_7410 = _T_7408 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7411 = _T_7407 | _T_7410; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7412 = _T_7411 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7422 = _T_4758 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7423 = perr_ic_index_ff == 7'h57; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_7425 = _T_7423 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7426 = _T_7422 | _T_7425; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7427 = _T_7426 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7437 = _T_4759 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7438 = perr_ic_index_ff == 7'h58; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_7440 = _T_7438 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7441 = _T_7437 | _T_7440; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7442 = _T_7441 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7452 = _T_4760 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7453 = perr_ic_index_ff == 7'h59; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_7455 = _T_7453 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7456 = _T_7452 | _T_7455; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7457 = _T_7456 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7467 = _T_4761 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7468 = perr_ic_index_ff == 7'h5a; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_7470 = _T_7468 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7471 = _T_7467 | _T_7470; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7472 = _T_7471 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7482 = _T_4762 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7483 = perr_ic_index_ff == 7'h5b; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_7485 = _T_7483 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7486 = _T_7482 | _T_7485; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7487 = _T_7486 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7497 = _T_4763 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7498 = perr_ic_index_ff == 7'h5c; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_7500 = _T_7498 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7501 = _T_7497 | _T_7500; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7502 = _T_7501 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7512 = _T_4764 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7513 = perr_ic_index_ff == 7'h5d; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_7515 = _T_7513 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7516 = _T_7512 | _T_7515; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7517 = _T_7516 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7527 = _T_4765 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7528 = perr_ic_index_ff == 7'h5e; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_7530 = _T_7528 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7531 = _T_7527 | _T_7530; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7532 = _T_7531 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7542 = _T_4766 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7543 = perr_ic_index_ff == 7'h5f; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_7545 = _T_7543 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7546 = _T_7542 | _T_7545; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7547 = _T_7546 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7557 = _T_4735 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7560 = _T_7078 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7561 = _T_7557 | _T_7560; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7562 = _T_7561 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7572 = _T_4736 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7575 = _T_7093 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7576 = _T_7572 | _T_7575; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7577 = _T_7576 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7587 = _T_4737 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7590 = _T_7108 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7591 = _T_7587 | _T_7590; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7592 = _T_7591 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7602 = _T_4738 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7605 = _T_7123 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7606 = _T_7602 | _T_7605; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7607 = _T_7606 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7617 = _T_4739 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7620 = _T_7138 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7621 = _T_7617 | _T_7620; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7622 = _T_7621 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7632 = _T_4740 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7635 = _T_7153 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7636 = _T_7632 | _T_7635; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7637 = _T_7636 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7647 = _T_4741 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7650 = _T_7168 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7651 = _T_7647 | _T_7650; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7652 = _T_7651 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7662 = _T_4742 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7665 = _T_7183 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7666 = _T_7662 | _T_7665; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7667 = _T_7666 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7677 = _T_4743 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7680 = _T_7198 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7681 = _T_7677 | _T_7680; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7682 = _T_7681 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7692 = _T_4744 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7695 = _T_7213 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7696 = _T_7692 | _T_7695; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7697 = _T_7696 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7707 = _T_4745 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7710 = _T_7228 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7711 = _T_7707 | _T_7710; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7712 = _T_7711 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7722 = _T_4746 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7725 = _T_7243 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7726 = _T_7722 | _T_7725; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7727 = _T_7726 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7737 = _T_4747 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7740 = _T_7258 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7741 = _T_7737 | _T_7740; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7742 = _T_7741 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7752 = _T_4748 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7755 = _T_7273 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7756 = _T_7752 | _T_7755; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7757 = _T_7756 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7767 = _T_4749 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7770 = _T_7288 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7771 = _T_7767 | _T_7770; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7772 = _T_7771 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7782 = _T_4750 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7785 = _T_7303 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7786 = _T_7782 | _T_7785; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7787 = _T_7786 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7797 = _T_4751 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7800 = _T_7318 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7801 = _T_7797 | _T_7800; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7802 = _T_7801 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7812 = _T_4752 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7815 = _T_7333 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7816 = _T_7812 | _T_7815; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7817 = _T_7816 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7827 = _T_4753 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7830 = _T_7348 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7831 = _T_7827 | _T_7830; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7832 = _T_7831 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7842 = _T_4754 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7845 = _T_7363 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7846 = _T_7842 | _T_7845; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7847 = _T_7846 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7857 = _T_4755 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7860 = _T_7378 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7861 = _T_7857 | _T_7860; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7862 = _T_7861 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7872 = _T_4756 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7875 = _T_7393 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7876 = _T_7872 | _T_7875; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7877 = _T_7876 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7887 = _T_4757 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7890 = _T_7408 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7891 = _T_7887 | _T_7890; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7892 = _T_7891 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7902 = _T_4758 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7905 = _T_7423 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7906 = _T_7902 | _T_7905; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7907 = _T_7906 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7917 = _T_4759 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7920 = _T_7438 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7921 = _T_7917 | _T_7920; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7922 = _T_7921 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7932 = _T_4760 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7935 = _T_7453 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7936 = _T_7932 | _T_7935; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7937 = _T_7936 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7947 = _T_4761 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7950 = _T_7468 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7951 = _T_7947 | _T_7950; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7952 = _T_7951 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7962 = _T_4762 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7965 = _T_7483 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7966 = _T_7962 | _T_7965; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7967 = _T_7966 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7977 = _T_4763 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7980 = _T_7498 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7981 = _T_7977 | _T_7980; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7982 = _T_7981 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_7992 = _T_4764 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_7995 = _T_7513 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_7996 = _T_7992 | _T_7995; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_7997 = _T_7996 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8007 = _T_4765 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8010 = _T_7528 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8011 = _T_8007 | _T_8010; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8012 = _T_8011 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8022 = _T_4766 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8025 = _T_7543 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8026 = _T_8022 | _T_8025; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8027 = _T_8026 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8037 = _T_4767 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8038 = perr_ic_index_ff == 7'h60; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_8040 = _T_8038 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8041 = _T_8037 | _T_8040; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8042 = _T_8041 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8052 = _T_4768 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8053 = perr_ic_index_ff == 7'h61; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_8055 = _T_8053 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8056 = _T_8052 | _T_8055; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8057 = _T_8056 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8067 = _T_4769 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8068 = perr_ic_index_ff == 7'h62; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_8070 = _T_8068 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8071 = _T_8067 | _T_8070; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8072 = _T_8071 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8082 = _T_4770 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8083 = perr_ic_index_ff == 7'h63; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_8085 = _T_8083 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8086 = _T_8082 | _T_8085; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8087 = _T_8086 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8097 = _T_4771 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8098 = perr_ic_index_ff == 7'h64; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_8100 = _T_8098 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8101 = _T_8097 | _T_8100; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8102 = _T_8101 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8112 = _T_4772 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8113 = perr_ic_index_ff == 7'h65; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_8115 = _T_8113 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8116 = _T_8112 | _T_8115; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8117 = _T_8116 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8127 = _T_4773 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8128 = perr_ic_index_ff == 7'h66; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_8130 = _T_8128 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8131 = _T_8127 | _T_8130; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8132 = _T_8131 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8142 = _T_4774 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8143 = perr_ic_index_ff == 7'h67; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_8145 = _T_8143 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8146 = _T_8142 | _T_8145; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8147 = _T_8146 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8157 = _T_4775 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8158 = perr_ic_index_ff == 7'h68; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_8160 = _T_8158 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8161 = _T_8157 | _T_8160; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8162 = _T_8161 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8172 = _T_4776 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8173 = perr_ic_index_ff == 7'h69; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_8175 = _T_8173 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8176 = _T_8172 | _T_8175; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8177 = _T_8176 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8187 = _T_4777 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8188 = perr_ic_index_ff == 7'h6a; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_8190 = _T_8188 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8191 = _T_8187 | _T_8190; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8192 = _T_8191 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8202 = _T_4778 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8203 = perr_ic_index_ff == 7'h6b; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_8205 = _T_8203 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8206 = _T_8202 | _T_8205; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8207 = _T_8206 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8217 = _T_4779 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8218 = perr_ic_index_ff == 7'h6c; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_8220 = _T_8218 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8221 = _T_8217 | _T_8220; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8222 = _T_8221 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8232 = _T_4780 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8233 = perr_ic_index_ff == 7'h6d; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_8235 = _T_8233 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8236 = _T_8232 | _T_8235; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8237 = _T_8236 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8247 = _T_4781 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8248 = perr_ic_index_ff == 7'h6e; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_8250 = _T_8248 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8251 = _T_8247 | _T_8250; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8252 = _T_8251 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8262 = _T_4782 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8263 = perr_ic_index_ff == 7'h6f; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_8265 = _T_8263 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8266 = _T_8262 | _T_8265; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8267 = _T_8266 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8277 = _T_4783 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8278 = perr_ic_index_ff == 7'h70; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_8280 = _T_8278 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8281 = _T_8277 | _T_8280; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8282 = _T_8281 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8292 = _T_4784 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8293 = perr_ic_index_ff == 7'h71; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_8295 = _T_8293 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8296 = _T_8292 | _T_8295; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8297 = _T_8296 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8307 = _T_4785 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8308 = perr_ic_index_ff == 7'h72; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_8310 = _T_8308 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8311 = _T_8307 | _T_8310; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8312 = _T_8311 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8322 = _T_4786 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8323 = perr_ic_index_ff == 7'h73; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_8325 = _T_8323 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8326 = _T_8322 | _T_8325; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8327 = _T_8326 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8337 = _T_4787 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8338 = perr_ic_index_ff == 7'h74; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_8340 = _T_8338 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8341 = _T_8337 | _T_8340; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8342 = _T_8341 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8352 = _T_4788 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8353 = perr_ic_index_ff == 7'h75; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_8355 = _T_8353 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8356 = _T_8352 | _T_8355; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8357 = _T_8356 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8367 = _T_4789 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8368 = perr_ic_index_ff == 7'h76; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_8370 = _T_8368 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8371 = _T_8367 | _T_8370; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8372 = _T_8371 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8382 = _T_4790 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8383 = perr_ic_index_ff == 7'h77; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_8385 = _T_8383 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8386 = _T_8382 | _T_8385; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8387 = _T_8386 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8397 = _T_4791 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8398 = perr_ic_index_ff == 7'h78; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_8400 = _T_8398 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8401 = _T_8397 | _T_8400; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8402 = _T_8401 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8412 = _T_4792 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8413 = perr_ic_index_ff == 7'h79; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_8415 = _T_8413 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8416 = _T_8412 | _T_8415; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8417 = _T_8416 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8427 = _T_4793 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8428 = perr_ic_index_ff == 7'h7a; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_8430 = _T_8428 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8431 = _T_8427 | _T_8430; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8432 = _T_8431 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8442 = _T_4794 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8443 = perr_ic_index_ff == 7'h7b; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_8445 = _T_8443 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8446 = _T_8442 | _T_8445; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8447 = _T_8446 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8457 = _T_4795 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8458 = perr_ic_index_ff == 7'h7c; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_8460 = _T_8458 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8461 = _T_8457 | _T_8460; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8462 = _T_8461 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8472 = _T_4796 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8473 = perr_ic_index_ff == 7'h7d; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_8475 = _T_8473 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8476 = _T_8472 | _T_8475; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8477 = _T_8476 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8487 = _T_4797 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8488 = perr_ic_index_ff == 7'h7e; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_8490 = _T_8488 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8491 = _T_8487 | _T_8490; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8492 = _T_8491 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8502 = _T_4798 & ifu_tag_wren_ff[0]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8503 = perr_ic_index_ff == 7'h7f; // @[ifu_mem_ctl.scala 693:102]
  wire  _T_8505 = _T_8503 & perr_err_inv_way[0]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8506 = _T_8502 | _T_8505; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8507 = _T_8506 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8517 = _T_4767 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8520 = _T_8038 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8521 = _T_8517 | _T_8520; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8522 = _T_8521 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8532 = _T_4768 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8535 = _T_8053 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8536 = _T_8532 | _T_8535; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8537 = _T_8536 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8547 = _T_4769 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8550 = _T_8068 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8551 = _T_8547 | _T_8550; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8552 = _T_8551 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8562 = _T_4770 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8565 = _T_8083 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8566 = _T_8562 | _T_8565; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8567 = _T_8566 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8577 = _T_4771 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8580 = _T_8098 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8581 = _T_8577 | _T_8580; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8582 = _T_8581 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8592 = _T_4772 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8595 = _T_8113 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8596 = _T_8592 | _T_8595; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8597 = _T_8596 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8607 = _T_4773 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8610 = _T_8128 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8611 = _T_8607 | _T_8610; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8612 = _T_8611 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8622 = _T_4774 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8625 = _T_8143 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8626 = _T_8622 | _T_8625; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8627 = _T_8626 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8637 = _T_4775 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8640 = _T_8158 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8641 = _T_8637 | _T_8640; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8642 = _T_8641 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8652 = _T_4776 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8655 = _T_8173 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8656 = _T_8652 | _T_8655; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8657 = _T_8656 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8667 = _T_4777 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8670 = _T_8188 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8671 = _T_8667 | _T_8670; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8672 = _T_8671 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8682 = _T_4778 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8685 = _T_8203 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8686 = _T_8682 | _T_8685; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8687 = _T_8686 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8697 = _T_4779 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8700 = _T_8218 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8701 = _T_8697 | _T_8700; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8702 = _T_8701 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8712 = _T_4780 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8715 = _T_8233 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8716 = _T_8712 | _T_8715; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8717 = _T_8716 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8727 = _T_4781 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8730 = _T_8248 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8731 = _T_8727 | _T_8730; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8732 = _T_8731 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8742 = _T_4782 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8745 = _T_8263 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8746 = _T_8742 | _T_8745; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8747 = _T_8746 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8757 = _T_4783 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8760 = _T_8278 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8761 = _T_8757 | _T_8760; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8762 = _T_8761 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8772 = _T_4784 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8775 = _T_8293 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8776 = _T_8772 | _T_8775; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8777 = _T_8776 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8787 = _T_4785 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8790 = _T_8308 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8791 = _T_8787 | _T_8790; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8792 = _T_8791 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8802 = _T_4786 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8805 = _T_8323 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8806 = _T_8802 | _T_8805; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8807 = _T_8806 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8817 = _T_4787 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8820 = _T_8338 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8821 = _T_8817 | _T_8820; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8822 = _T_8821 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8832 = _T_4788 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8835 = _T_8353 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8836 = _T_8832 | _T_8835; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8837 = _T_8836 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8847 = _T_4789 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8850 = _T_8368 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8851 = _T_8847 | _T_8850; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8852 = _T_8851 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8862 = _T_4790 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8865 = _T_8383 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8866 = _T_8862 | _T_8865; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8867 = _T_8866 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8877 = _T_4791 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8880 = _T_8398 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8881 = _T_8877 | _T_8880; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8882 = _T_8881 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8892 = _T_4792 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8895 = _T_8413 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8896 = _T_8892 | _T_8895; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8897 = _T_8896 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8907 = _T_4793 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8910 = _T_8428 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8911 = _T_8907 | _T_8910; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8912 = _T_8911 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8922 = _T_4794 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8925 = _T_8443 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8926 = _T_8922 | _T_8925; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8927 = _T_8926 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8937 = _T_4795 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8940 = _T_8458 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8941 = _T_8937 | _T_8940; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8942 = _T_8941 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8952 = _T_4796 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8955 = _T_8473 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8956 = _T_8952 | _T_8955; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8957 = _T_8956 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8967 = _T_4797 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8970 = _T_8488 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8971 = _T_8967 | _T_8970; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8972 = _T_8971 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_8982 = _T_4798 & ifu_tag_wren_ff[1]; // @[ifu_mem_ctl.scala 693:59]
  wire  _T_8985 = _T_8503 & perr_err_inv_way[1]; // @[ifu_mem_ctl.scala 693:124]
  wire  _T_8986 = _T_8982 | _T_8985; // @[ifu_mem_ctl.scala 693:81]
  wire  _T_8987 = _T_8986 | reset_all_tags; // @[ifu_mem_ctl.scala 693:147]
  wire  _T_9789 = ~fetch_uncacheable_ff; // @[ifu_mem_ctl.scala 747:63]
  wire  _T_9790 = _T_9789 & ifc_fetch_req_f; // @[ifu_mem_ctl.scala 747:85]
  wire [1:0] _T_9792 = _T_9790 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  reg  _T_9799; // @[ifu_mem_ctl.scala 752:70]
  reg  _T_9800; // @[ifu_mem_ctl.scala 753:69]
  reg  _T_9801; // @[ifu_mem_ctl.scala 754:72]
  wire  _T_9802 = ~ifu_bus_arready_ff; // @[ifu_mem_ctl.scala 755:93]
  wire  _T_9803 = ifu_bus_arvalid_ff & _T_9802; // @[ifu_mem_ctl.scala 755:91]
  reg  _T_9805; // @[ifu_mem_ctl.scala 755:71]
  reg  _T_9806; // @[ifu_mem_ctl.scala 756:71]
  wire  _T_9809 = io_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_dicawics[15:14] == 2'h3; // @[ifu_mem_ctl.scala 763:84]
  wire  _T_9811 = io_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_dicawics[15:14] == 2'h2; // @[ifu_mem_ctl.scala 763:150]
  wire  _T_9813 = io_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_dicawics[15:14] == 2'h1; // @[ifu_mem_ctl.scala 764:63]
  wire  _T_9815 = io_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_dicawics[15:14] == 2'h0; // @[ifu_mem_ctl.scala 764:129]
  wire [3:0] _T_9818 = {_T_9809,_T_9811,_T_9813,_T_9815}; // @[Cat.scala 29:58]
  reg  _T_9826; // @[ifu_mem_ctl.scala 770:79]
  wire [31:0] _T_9836 = {io_ifc_fetch_addr_bf,1'h0}; // @[Cat.scala 29:58]
  wire [31:0] _T_9837 = _T_9836 | 32'h7fffffff; // @[ifu_mem_ctl.scala 773:65]
  wire  _T_9839 = _T_9837 == 32'h7fffffff; // @[ifu_mem_ctl.scala 773:96]
  wire [31:0] _T_9843 = _T_9836 | 32'h3fffffff; // @[ifu_mem_ctl.scala 774:65]
  wire  _T_9845 = _T_9843 == 32'hffffffff; // @[ifu_mem_ctl.scala 774:96]
  wire  _T_9847 = _T_9839 | _T_9845; // @[ifu_mem_ctl.scala 773:162]
  wire [31:0] _T_9849 = _T_9836 | 32'h1fffffff; // @[ifu_mem_ctl.scala 775:65]
  wire  _T_9851 = _T_9849 == 32'hbfffffff; // @[ifu_mem_ctl.scala 775:96]
  wire  _T_9853 = _T_9847 | _T_9851; // @[ifu_mem_ctl.scala 774:162]
  wire [31:0] _T_9855 = _T_9836 | 32'hfffffff; // @[ifu_mem_ctl.scala 776:65]
  wire  _T_9857 = _T_9855 == 32'h8fffffff; // @[ifu_mem_ctl.scala 776:96]
  wire  ifc_region_acc_okay = _T_9853 | _T_9857; // @[ifu_mem_ctl.scala 775:162]
  wire  _T_9884 = ~ifc_region_acc_okay; // @[ifu_mem_ctl.scala 781:65]
  wire  _T_9885 = _T_3939 & _T_9884; // @[ifu_mem_ctl.scala 781:63]
  wire  ifc_region_acc_fault_memory_bf = _T_9885 & io_ifc_fetch_req_bf; // @[ifu_mem_ctl.scala 781:86]
  rvclkhdr rvclkhdr ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_io_l1clk),
    .io_clk(rvclkhdr_io_clk),
    .io_en(rvclkhdr_io_en),
    .io_scan_mode(rvclkhdr_io_scan_mode)
  );
  rvclkhdr rvclkhdr_1 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_1_io_l1clk),
    .io_clk(rvclkhdr_1_io_clk),
    .io_en(rvclkhdr_1_io_en),
    .io_scan_mode(rvclkhdr_1_io_scan_mode)
  );
  rvclkhdr rvclkhdr_2 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_2_io_l1clk),
    .io_clk(rvclkhdr_2_io_clk),
    .io_en(rvclkhdr_2_io_en),
    .io_scan_mode(rvclkhdr_2_io_scan_mode)
  );
  rvclkhdr rvclkhdr_3 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_3_io_l1clk),
    .io_clk(rvclkhdr_3_io_clk),
    .io_en(rvclkhdr_3_io_en),
    .io_scan_mode(rvclkhdr_3_io_scan_mode)
  );
  rvclkhdr rvclkhdr_4 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_4_io_l1clk),
    .io_clk(rvclkhdr_4_io_clk),
    .io_en(rvclkhdr_4_io_en),
    .io_scan_mode(rvclkhdr_4_io_scan_mode)
  );
  rvclkhdr rvclkhdr_5 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_5_io_l1clk),
    .io_clk(rvclkhdr_5_io_clk),
    .io_en(rvclkhdr_5_io_en),
    .io_scan_mode(rvclkhdr_5_io_scan_mode)
  );
  rvclkhdr rvclkhdr_6 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_6_io_l1clk),
    .io_clk(rvclkhdr_6_io_clk),
    .io_en(rvclkhdr_6_io_en),
    .io_scan_mode(rvclkhdr_6_io_scan_mode)
  );
  rvclkhdr rvclkhdr_7 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_7_io_l1clk),
    .io_clk(rvclkhdr_7_io_clk),
    .io_en(rvclkhdr_7_io_en),
    .io_scan_mode(rvclkhdr_7_io_scan_mode)
  );
  rvclkhdr rvclkhdr_8 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_8_io_l1clk),
    .io_clk(rvclkhdr_8_io_clk),
    .io_en(rvclkhdr_8_io_en),
    .io_scan_mode(rvclkhdr_8_io_scan_mode)
  );
  rvclkhdr rvclkhdr_9 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_9_io_l1clk),
    .io_clk(rvclkhdr_9_io_clk),
    .io_en(rvclkhdr_9_io_en),
    .io_scan_mode(rvclkhdr_9_io_scan_mode)
  );
  rvclkhdr rvclkhdr_10 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_10_io_l1clk),
    .io_clk(rvclkhdr_10_io_clk),
    .io_en(rvclkhdr_10_io_en),
    .io_scan_mode(rvclkhdr_10_io_scan_mode)
  );
  rvclkhdr rvclkhdr_11 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_11_io_l1clk),
    .io_clk(rvclkhdr_11_io_clk),
    .io_en(rvclkhdr_11_io_en),
    .io_scan_mode(rvclkhdr_11_io_scan_mode)
  );
  rvclkhdr rvclkhdr_12 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_12_io_l1clk),
    .io_clk(rvclkhdr_12_io_clk),
    .io_en(rvclkhdr_12_io_en),
    .io_scan_mode(rvclkhdr_12_io_scan_mode)
  );
  rvclkhdr rvclkhdr_13 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_13_io_l1clk),
    .io_clk(rvclkhdr_13_io_clk),
    .io_en(rvclkhdr_13_io_en),
    .io_scan_mode(rvclkhdr_13_io_scan_mode)
  );
  rvclkhdr rvclkhdr_14 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_14_io_l1clk),
    .io_clk(rvclkhdr_14_io_clk),
    .io_en(rvclkhdr_14_io_en),
    .io_scan_mode(rvclkhdr_14_io_scan_mode)
  );
  rvclkhdr rvclkhdr_15 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_15_io_l1clk),
    .io_clk(rvclkhdr_15_io_clk),
    .io_en(rvclkhdr_15_io_en),
    .io_scan_mode(rvclkhdr_15_io_scan_mode)
  );
  rvclkhdr rvclkhdr_16 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_16_io_l1clk),
    .io_clk(rvclkhdr_16_io_clk),
    .io_en(rvclkhdr_16_io_en),
    .io_scan_mode(rvclkhdr_16_io_scan_mode)
  );
  rvclkhdr rvclkhdr_17 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_17_io_l1clk),
    .io_clk(rvclkhdr_17_io_clk),
    .io_en(rvclkhdr_17_io_en),
    .io_scan_mode(rvclkhdr_17_io_scan_mode)
  );
  rvclkhdr rvclkhdr_18 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_18_io_l1clk),
    .io_clk(rvclkhdr_18_io_clk),
    .io_en(rvclkhdr_18_io_en),
    .io_scan_mode(rvclkhdr_18_io_scan_mode)
  );
  rvclkhdr rvclkhdr_19 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_19_io_l1clk),
    .io_clk(rvclkhdr_19_io_clk),
    .io_en(rvclkhdr_19_io_en),
    .io_scan_mode(rvclkhdr_19_io_scan_mode)
  );
  rvclkhdr rvclkhdr_20 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_20_io_l1clk),
    .io_clk(rvclkhdr_20_io_clk),
    .io_en(rvclkhdr_20_io_en),
    .io_scan_mode(rvclkhdr_20_io_scan_mode)
  );
  rvclkhdr rvclkhdr_21 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_21_io_l1clk),
    .io_clk(rvclkhdr_21_io_clk),
    .io_en(rvclkhdr_21_io_en),
    .io_scan_mode(rvclkhdr_21_io_scan_mode)
  );
  rvclkhdr rvclkhdr_22 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_22_io_l1clk),
    .io_clk(rvclkhdr_22_io_clk),
    .io_en(rvclkhdr_22_io_en),
    .io_scan_mode(rvclkhdr_22_io_scan_mode)
  );
  rvclkhdr rvclkhdr_23 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_23_io_l1clk),
    .io_clk(rvclkhdr_23_io_clk),
    .io_en(rvclkhdr_23_io_en),
    .io_scan_mode(rvclkhdr_23_io_scan_mode)
  );
  rvclkhdr rvclkhdr_24 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_24_io_l1clk),
    .io_clk(rvclkhdr_24_io_clk),
    .io_en(rvclkhdr_24_io_en),
    .io_scan_mode(rvclkhdr_24_io_scan_mode)
  );
  rvclkhdr rvclkhdr_25 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_25_io_l1clk),
    .io_clk(rvclkhdr_25_io_clk),
    .io_en(rvclkhdr_25_io_en),
    .io_scan_mode(rvclkhdr_25_io_scan_mode)
  );
  rvclkhdr rvclkhdr_26 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_26_io_l1clk),
    .io_clk(rvclkhdr_26_io_clk),
    .io_en(rvclkhdr_26_io_en),
    .io_scan_mode(rvclkhdr_26_io_scan_mode)
  );
  rvclkhdr rvclkhdr_27 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_27_io_l1clk),
    .io_clk(rvclkhdr_27_io_clk),
    .io_en(rvclkhdr_27_io_en),
    .io_scan_mode(rvclkhdr_27_io_scan_mode)
  );
  rvclkhdr rvclkhdr_28 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_28_io_l1clk),
    .io_clk(rvclkhdr_28_io_clk),
    .io_en(rvclkhdr_28_io_en),
    .io_scan_mode(rvclkhdr_28_io_scan_mode)
  );
  rvclkhdr rvclkhdr_29 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_29_io_l1clk),
    .io_clk(rvclkhdr_29_io_clk),
    .io_en(rvclkhdr_29_io_en),
    .io_scan_mode(rvclkhdr_29_io_scan_mode)
  );
  rvclkhdr rvclkhdr_30 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_30_io_l1clk),
    .io_clk(rvclkhdr_30_io_clk),
    .io_en(rvclkhdr_30_io_en),
    .io_scan_mode(rvclkhdr_30_io_scan_mode)
  );
  rvclkhdr rvclkhdr_31 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_31_io_l1clk),
    .io_clk(rvclkhdr_31_io_clk),
    .io_en(rvclkhdr_31_io_en),
    .io_scan_mode(rvclkhdr_31_io_scan_mode)
  );
  rvclkhdr rvclkhdr_32 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_32_io_l1clk),
    .io_clk(rvclkhdr_32_io_clk),
    .io_en(rvclkhdr_32_io_en),
    .io_scan_mode(rvclkhdr_32_io_scan_mode)
  );
  rvclkhdr rvclkhdr_33 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_33_io_l1clk),
    .io_clk(rvclkhdr_33_io_clk),
    .io_en(rvclkhdr_33_io_en),
    .io_scan_mode(rvclkhdr_33_io_scan_mode)
  );
  rvclkhdr rvclkhdr_34 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_34_io_l1clk),
    .io_clk(rvclkhdr_34_io_clk),
    .io_en(rvclkhdr_34_io_en),
    .io_scan_mode(rvclkhdr_34_io_scan_mode)
  );
  rvclkhdr rvclkhdr_35 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_35_io_l1clk),
    .io_clk(rvclkhdr_35_io_clk),
    .io_en(rvclkhdr_35_io_en),
    .io_scan_mode(rvclkhdr_35_io_scan_mode)
  );
  rvclkhdr rvclkhdr_36 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_36_io_l1clk),
    .io_clk(rvclkhdr_36_io_clk),
    .io_en(rvclkhdr_36_io_en),
    .io_scan_mode(rvclkhdr_36_io_scan_mode)
  );
  rvclkhdr rvclkhdr_37 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_37_io_l1clk),
    .io_clk(rvclkhdr_37_io_clk),
    .io_en(rvclkhdr_37_io_en),
    .io_scan_mode(rvclkhdr_37_io_scan_mode)
  );
  rvclkhdr rvclkhdr_38 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_38_io_l1clk),
    .io_clk(rvclkhdr_38_io_clk),
    .io_en(rvclkhdr_38_io_en),
    .io_scan_mode(rvclkhdr_38_io_scan_mode)
  );
  rvclkhdr rvclkhdr_39 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_39_io_l1clk),
    .io_clk(rvclkhdr_39_io_clk),
    .io_en(rvclkhdr_39_io_en),
    .io_scan_mode(rvclkhdr_39_io_scan_mode)
  );
  rvclkhdr rvclkhdr_40 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_40_io_l1clk),
    .io_clk(rvclkhdr_40_io_clk),
    .io_en(rvclkhdr_40_io_en),
    .io_scan_mode(rvclkhdr_40_io_scan_mode)
  );
  rvclkhdr rvclkhdr_41 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_41_io_l1clk),
    .io_clk(rvclkhdr_41_io_clk),
    .io_en(rvclkhdr_41_io_en),
    .io_scan_mode(rvclkhdr_41_io_scan_mode)
  );
  rvclkhdr rvclkhdr_42 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_42_io_l1clk),
    .io_clk(rvclkhdr_42_io_clk),
    .io_en(rvclkhdr_42_io_en),
    .io_scan_mode(rvclkhdr_42_io_scan_mode)
  );
  rvclkhdr rvclkhdr_43 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_43_io_l1clk),
    .io_clk(rvclkhdr_43_io_clk),
    .io_en(rvclkhdr_43_io_en),
    .io_scan_mode(rvclkhdr_43_io_scan_mode)
  );
  rvclkhdr rvclkhdr_44 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_44_io_l1clk),
    .io_clk(rvclkhdr_44_io_clk),
    .io_en(rvclkhdr_44_io_en),
    .io_scan_mode(rvclkhdr_44_io_scan_mode)
  );
  rvclkhdr rvclkhdr_45 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_45_io_l1clk),
    .io_clk(rvclkhdr_45_io_clk),
    .io_en(rvclkhdr_45_io_en),
    .io_scan_mode(rvclkhdr_45_io_scan_mode)
  );
  rvclkhdr rvclkhdr_46 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_46_io_l1clk),
    .io_clk(rvclkhdr_46_io_clk),
    .io_en(rvclkhdr_46_io_en),
    .io_scan_mode(rvclkhdr_46_io_scan_mode)
  );
  rvclkhdr rvclkhdr_47 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_47_io_l1clk),
    .io_clk(rvclkhdr_47_io_clk),
    .io_en(rvclkhdr_47_io_en),
    .io_scan_mode(rvclkhdr_47_io_scan_mode)
  );
  rvclkhdr rvclkhdr_48 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_48_io_l1clk),
    .io_clk(rvclkhdr_48_io_clk),
    .io_en(rvclkhdr_48_io_en),
    .io_scan_mode(rvclkhdr_48_io_scan_mode)
  );
  rvclkhdr rvclkhdr_49 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_49_io_l1clk),
    .io_clk(rvclkhdr_49_io_clk),
    .io_en(rvclkhdr_49_io_en),
    .io_scan_mode(rvclkhdr_49_io_scan_mode)
  );
  rvclkhdr rvclkhdr_50 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_50_io_l1clk),
    .io_clk(rvclkhdr_50_io_clk),
    .io_en(rvclkhdr_50_io_en),
    .io_scan_mode(rvclkhdr_50_io_scan_mode)
  );
  rvclkhdr rvclkhdr_51 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_51_io_l1clk),
    .io_clk(rvclkhdr_51_io_clk),
    .io_en(rvclkhdr_51_io_en),
    .io_scan_mode(rvclkhdr_51_io_scan_mode)
  );
  rvclkhdr rvclkhdr_52 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_52_io_l1clk),
    .io_clk(rvclkhdr_52_io_clk),
    .io_en(rvclkhdr_52_io_en),
    .io_scan_mode(rvclkhdr_52_io_scan_mode)
  );
  rvclkhdr rvclkhdr_53 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_53_io_l1clk),
    .io_clk(rvclkhdr_53_io_clk),
    .io_en(rvclkhdr_53_io_en),
    .io_scan_mode(rvclkhdr_53_io_scan_mode)
  );
  rvclkhdr rvclkhdr_54 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_54_io_l1clk),
    .io_clk(rvclkhdr_54_io_clk),
    .io_en(rvclkhdr_54_io_en),
    .io_scan_mode(rvclkhdr_54_io_scan_mode)
  );
  rvclkhdr rvclkhdr_55 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_55_io_l1clk),
    .io_clk(rvclkhdr_55_io_clk),
    .io_en(rvclkhdr_55_io_en),
    .io_scan_mode(rvclkhdr_55_io_scan_mode)
  );
  rvclkhdr rvclkhdr_56 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_56_io_l1clk),
    .io_clk(rvclkhdr_56_io_clk),
    .io_en(rvclkhdr_56_io_en),
    .io_scan_mode(rvclkhdr_56_io_scan_mode)
  );
  rvclkhdr rvclkhdr_57 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_57_io_l1clk),
    .io_clk(rvclkhdr_57_io_clk),
    .io_en(rvclkhdr_57_io_en),
    .io_scan_mode(rvclkhdr_57_io_scan_mode)
  );
  rvclkhdr rvclkhdr_58 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_58_io_l1clk),
    .io_clk(rvclkhdr_58_io_clk),
    .io_en(rvclkhdr_58_io_en),
    .io_scan_mode(rvclkhdr_58_io_scan_mode)
  );
  rvclkhdr rvclkhdr_59 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_59_io_l1clk),
    .io_clk(rvclkhdr_59_io_clk),
    .io_en(rvclkhdr_59_io_en),
    .io_scan_mode(rvclkhdr_59_io_scan_mode)
  );
  rvclkhdr rvclkhdr_60 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_60_io_l1clk),
    .io_clk(rvclkhdr_60_io_clk),
    .io_en(rvclkhdr_60_io_en),
    .io_scan_mode(rvclkhdr_60_io_scan_mode)
  );
  rvclkhdr rvclkhdr_61 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_61_io_l1clk),
    .io_clk(rvclkhdr_61_io_clk),
    .io_en(rvclkhdr_61_io_en),
    .io_scan_mode(rvclkhdr_61_io_scan_mode)
  );
  rvclkhdr rvclkhdr_62 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_62_io_l1clk),
    .io_clk(rvclkhdr_62_io_clk),
    .io_en(rvclkhdr_62_io_en),
    .io_scan_mode(rvclkhdr_62_io_scan_mode)
  );
  rvclkhdr rvclkhdr_63 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_63_io_l1clk),
    .io_clk(rvclkhdr_63_io_clk),
    .io_en(rvclkhdr_63_io_en),
    .io_scan_mode(rvclkhdr_63_io_scan_mode)
  );
  rvclkhdr rvclkhdr_64 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_64_io_l1clk),
    .io_clk(rvclkhdr_64_io_clk),
    .io_en(rvclkhdr_64_io_en),
    .io_scan_mode(rvclkhdr_64_io_scan_mode)
  );
  rvclkhdr rvclkhdr_65 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_65_io_l1clk),
    .io_clk(rvclkhdr_65_io_clk),
    .io_en(rvclkhdr_65_io_en),
    .io_scan_mode(rvclkhdr_65_io_scan_mode)
  );
  rvclkhdr rvclkhdr_66 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_66_io_l1clk),
    .io_clk(rvclkhdr_66_io_clk),
    .io_en(rvclkhdr_66_io_en),
    .io_scan_mode(rvclkhdr_66_io_scan_mode)
  );
  rvclkhdr rvclkhdr_67 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_67_io_l1clk),
    .io_clk(rvclkhdr_67_io_clk),
    .io_en(rvclkhdr_67_io_en),
    .io_scan_mode(rvclkhdr_67_io_scan_mode)
  );
  rvclkhdr rvclkhdr_68 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_68_io_l1clk),
    .io_clk(rvclkhdr_68_io_clk),
    .io_en(rvclkhdr_68_io_en),
    .io_scan_mode(rvclkhdr_68_io_scan_mode)
  );
  rvclkhdr rvclkhdr_69 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_69_io_l1clk),
    .io_clk(rvclkhdr_69_io_clk),
    .io_en(rvclkhdr_69_io_en),
    .io_scan_mode(rvclkhdr_69_io_scan_mode)
  );
  rvclkhdr rvclkhdr_70 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_70_io_l1clk),
    .io_clk(rvclkhdr_70_io_clk),
    .io_en(rvclkhdr_70_io_en),
    .io_scan_mode(rvclkhdr_70_io_scan_mode)
  );
  rvclkhdr rvclkhdr_71 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_71_io_l1clk),
    .io_clk(rvclkhdr_71_io_clk),
    .io_en(rvclkhdr_71_io_en),
    .io_scan_mode(rvclkhdr_71_io_scan_mode)
  );
  rvclkhdr rvclkhdr_72 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_72_io_l1clk),
    .io_clk(rvclkhdr_72_io_clk),
    .io_en(rvclkhdr_72_io_en),
    .io_scan_mode(rvclkhdr_72_io_scan_mode)
  );
  rvclkhdr rvclkhdr_73 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_73_io_l1clk),
    .io_clk(rvclkhdr_73_io_clk),
    .io_en(rvclkhdr_73_io_en),
    .io_scan_mode(rvclkhdr_73_io_scan_mode)
  );
  rvclkhdr rvclkhdr_74 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_74_io_l1clk),
    .io_clk(rvclkhdr_74_io_clk),
    .io_en(rvclkhdr_74_io_en),
    .io_scan_mode(rvclkhdr_74_io_scan_mode)
  );
  rvclkhdr rvclkhdr_75 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_75_io_l1clk),
    .io_clk(rvclkhdr_75_io_clk),
    .io_en(rvclkhdr_75_io_en),
    .io_scan_mode(rvclkhdr_75_io_scan_mode)
  );
  rvclkhdr rvclkhdr_76 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_76_io_l1clk),
    .io_clk(rvclkhdr_76_io_clk),
    .io_en(rvclkhdr_76_io_en),
    .io_scan_mode(rvclkhdr_76_io_scan_mode)
  );
  rvclkhdr rvclkhdr_77 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_77_io_l1clk),
    .io_clk(rvclkhdr_77_io_clk),
    .io_en(rvclkhdr_77_io_en),
    .io_scan_mode(rvclkhdr_77_io_scan_mode)
  );
  rvclkhdr rvclkhdr_78 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_78_io_l1clk),
    .io_clk(rvclkhdr_78_io_clk),
    .io_en(rvclkhdr_78_io_en),
    .io_scan_mode(rvclkhdr_78_io_scan_mode)
  );
  rvclkhdr rvclkhdr_79 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_79_io_l1clk),
    .io_clk(rvclkhdr_79_io_clk),
    .io_en(rvclkhdr_79_io_en),
    .io_scan_mode(rvclkhdr_79_io_scan_mode)
  );
  rvclkhdr rvclkhdr_80 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_80_io_l1clk),
    .io_clk(rvclkhdr_80_io_clk),
    .io_en(rvclkhdr_80_io_en),
    .io_scan_mode(rvclkhdr_80_io_scan_mode)
  );
  rvclkhdr rvclkhdr_81 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_81_io_l1clk),
    .io_clk(rvclkhdr_81_io_clk),
    .io_en(rvclkhdr_81_io_en),
    .io_scan_mode(rvclkhdr_81_io_scan_mode)
  );
  rvclkhdr rvclkhdr_82 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_82_io_l1clk),
    .io_clk(rvclkhdr_82_io_clk),
    .io_en(rvclkhdr_82_io_en),
    .io_scan_mode(rvclkhdr_82_io_scan_mode)
  );
  rvclkhdr rvclkhdr_83 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_83_io_l1clk),
    .io_clk(rvclkhdr_83_io_clk),
    .io_en(rvclkhdr_83_io_en),
    .io_scan_mode(rvclkhdr_83_io_scan_mode)
  );
  rvclkhdr rvclkhdr_84 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_84_io_l1clk),
    .io_clk(rvclkhdr_84_io_clk),
    .io_en(rvclkhdr_84_io_en),
    .io_scan_mode(rvclkhdr_84_io_scan_mode)
  );
  rvclkhdr rvclkhdr_85 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_85_io_l1clk),
    .io_clk(rvclkhdr_85_io_clk),
    .io_en(rvclkhdr_85_io_en),
    .io_scan_mode(rvclkhdr_85_io_scan_mode)
  );
  rvclkhdr rvclkhdr_86 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_86_io_l1clk),
    .io_clk(rvclkhdr_86_io_clk),
    .io_en(rvclkhdr_86_io_en),
    .io_scan_mode(rvclkhdr_86_io_scan_mode)
  );
  rvclkhdr rvclkhdr_87 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_87_io_l1clk),
    .io_clk(rvclkhdr_87_io_clk),
    .io_en(rvclkhdr_87_io_en),
    .io_scan_mode(rvclkhdr_87_io_scan_mode)
  );
  rvclkhdr rvclkhdr_88 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_88_io_l1clk),
    .io_clk(rvclkhdr_88_io_clk),
    .io_en(rvclkhdr_88_io_en),
    .io_scan_mode(rvclkhdr_88_io_scan_mode)
  );
  rvclkhdr rvclkhdr_89 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_89_io_l1clk),
    .io_clk(rvclkhdr_89_io_clk),
    .io_en(rvclkhdr_89_io_en),
    .io_scan_mode(rvclkhdr_89_io_scan_mode)
  );
  rvclkhdr rvclkhdr_90 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_90_io_l1clk),
    .io_clk(rvclkhdr_90_io_clk),
    .io_en(rvclkhdr_90_io_en),
    .io_scan_mode(rvclkhdr_90_io_scan_mode)
  );
  rvclkhdr rvclkhdr_91 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_91_io_l1clk),
    .io_clk(rvclkhdr_91_io_clk),
    .io_en(rvclkhdr_91_io_en),
    .io_scan_mode(rvclkhdr_91_io_scan_mode)
  );
  rvclkhdr rvclkhdr_92 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_92_io_l1clk),
    .io_clk(rvclkhdr_92_io_clk),
    .io_en(rvclkhdr_92_io_en),
    .io_scan_mode(rvclkhdr_92_io_scan_mode)
  );
  rvclkhdr rvclkhdr_93 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_93_io_l1clk),
    .io_clk(rvclkhdr_93_io_clk),
    .io_en(rvclkhdr_93_io_en),
    .io_scan_mode(rvclkhdr_93_io_scan_mode)
  );
  assign io_dec_mem_ctrl_ifu_pmu_ic_miss = _T_9799; // @[ifu_mem_ctl.scala 752:35]
  assign io_dec_mem_ctrl_ifu_pmu_ic_hit = _T_9800; // @[ifu_mem_ctl.scala 753:34]
  assign io_dec_mem_ctrl_ifu_pmu_bus_error = _T_9801; // @[ifu_mem_ctl.scala 754:37]
  assign io_dec_mem_ctrl_ifu_pmu_bus_busy = _T_9805; // @[ifu_mem_ctl.scala 755:36]
  assign io_dec_mem_ctrl_ifu_pmu_bus_trxn = _T_9806; // @[ifu_mem_ctl.scala 756:36]
  assign io_dec_mem_ctrl_ifu_ic_error_start = _T_1200 | ic_rd_parity_final_err; // @[ifu_mem_ctl.scala 256:38]
  assign io_dec_mem_ctrl_ifu_iccm_rd_ecc_single_err = _T_3911 & ifc_fetch_req_f; // @[ifu_mem_ctl.scala 612:46]
  assign io_dec_mem_ctrl_ifu_ic_debug_rd_data = _T_1212; // @[ifu_mem_ctl.scala 263:40]
  assign io_dec_mem_ctrl_ifu_ic_debug_rd_data_valid = _T_9826; // @[ifu_mem_ctl.scala 770:46]
  assign io_dec_mem_ctrl_ifu_miss_state_idle = miss_state == 3'h0; // @[ifu_mem_ctl.scala 235:39]
  assign io_ifu_axi_ar_valid = ifu_bus_cmd_valid; // @[ifu_mem_ctl.scala 497:23]
  assign io_ifu_axi_ar_bits_id = bus_rd_addr_count & _T_2608; // @[ifu_mem_ctl.scala 498:25]
  assign io_ifu_axi_ar_bits_addr = _T_2610 & _T_2612; // @[ifu_mem_ctl.scala 499:27]
  assign io_ifu_axi_ar_bits_region = ifu_ic_req_addr_f[28:25]; // @[ifu_mem_ctl.scala 502:29]
  assign io_ifu_axi_r_ready = 1'h1; // @[ifu_mem_ctl.scala 504:22]
  assign io_iccm_rw_addr = _T_3110 ? io_dma_mem_ctl_dma_mem_addr[15:1] : _T_3117; // @[ifu_mem_ctl.scala 599:19]
  assign io_iccm_buf_correct_ecc = iccm_correct_ecc & _T_2497; // @[ifu_mem_ctl.scala 395:27]
  assign io_iccm_correction_state = _T_2526 ? 1'h0 : _GEN_42; // @[ifu_mem_ctl.scala 430:28 ifu_mem_ctl.scala 442:32 ifu_mem_ctl.scala 449:32 ifu_mem_ctl.scala 456:32]
  assign io_iccm_wren = _T_2710 | iccm_correct_ecc; // @[ifu_mem_ctl.scala 569:16]
  assign io_iccm_rden = _T_2714 | _T_2715; // @[ifu_mem_ctl.scala 570:16]
  assign io_iccm_wr_size = _T_2720 & io_dma_mem_ctl_dma_mem_sz; // @[ifu_mem_ctl.scala 572:19]
  assign io_iccm_wr_data = _T_3092 ? _T_3093 : _T_3100; // @[ifu_mem_ctl.scala 576:19]
  assign io_ic_rw_addr = _T_340 | _T_341; // @[ifu_mem_ctl.scala 244:17]
  assign io_ic_tag_valid = ic_tag_valid_unq & _T_9792; // @[ifu_mem_ctl.scala 747:19]
  assign io_ic_wr_en = bus_ic_wr_en & _T_3974; // @[ifu_mem_ctl.scala 635:15]
  assign io_ic_rd_en = _T_3966 | _T_3971; // @[ifu_mem_ctl.scala 626:15]
  assign io_ic_wr_data_0 = ic_wr_16bytes_data[70:0]; // @[ifu_mem_ctl.scala 253:17]
  assign io_ic_wr_data_1 = ic_wr_16bytes_data[141:71]; // @[ifu_mem_ctl.scala 253:17]
  assign io_ic_debug_wr_data = io_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_wrdata; // @[ifu_mem_ctl.scala 254:23]
  assign io_ic_debug_addr = io_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_dicawics[9:0]; // @[ifu_mem_ctl.scala 759:20]
  assign io_ic_debug_rd_en = io_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_rd_valid; // @[ifu_mem_ctl.scala 761:21]
  assign io_ic_debug_wr_en = io_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_wr_valid; // @[ifu_mem_ctl.scala 762:21]
  assign io_ic_debug_tag_array = io_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_dicawics[16]; // @[ifu_mem_ctl.scala 760:25]
  assign io_ic_debug_way = _T_9818[1:0]; // @[ifu_mem_ctl.scala 763:19]
  assign io_ic_premux_data = ic_premux_data_temp[63:0]; // @[ifu_mem_ctl.scala 295:21]
  assign io_ic_sel_premux_data = fetch_req_iccm_f | sel_byp_data; // @[ifu_mem_ctl.scala 296:25]
  assign io_ifu_ic_mb_empty = _T_328 | _T_231; // @[ifu_mem_ctl.scala 234:22]
  assign io_ic_dma_active = _T_11 | io_dec_mem_ctrl_dec_tlu_flush_err_wb; // @[ifu_mem_ctl.scala 97:20]
  assign io_ic_write_stall = write_ic_16_bytes & _T_3988; // @[ifu_mem_ctl.scala 636:21]
  assign io_iccm_dma_ecc_error = iccm_dma_ecc_error; // @[ifu_mem_ctl.scala 595:25]
  assign io_iccm_dma_rvalid = iccm_dma_rvalid_temp; // @[ifu_mem_ctl.scala 593:22]
  assign io_iccm_dma_rdata = iccm_dma_rdata_temp; // @[ifu_mem_ctl.scala 597:21]
  assign io_iccm_dma_rtag = iccm_dma_rtag_temp; // @[ifu_mem_ctl.scala 588:20]
  assign io_iccm_ready = _T_2706 & _T_2700; // @[ifu_mem_ctl.scala 567:17]
  assign io_iccm_rd_ecc_double_err = iccm_dma_ecc_error_in & ifc_iccm_access_f; // @[ifu_mem_ctl.scala 613:29]
  assign io_iccm_dma_sb_error = _T_3 & dma_iccm_req_f; // @[ifu_mem_ctl.scala 95:24]
  assign io_ic_hit_f = _T_263 | _T_264; // @[ifu_mem_ctl.scala 195:15]
  assign io_ic_access_fault_f = _T_2492 & _T_319; // @[ifu_mem_ctl.scala 301:24]
  assign io_ic_access_fault_type_f = io_iccm_rd_ecc_double_err ? 2'h1 : _T_1278; // @[ifu_mem_ctl.scala 302:29]
  assign io_ifu_async_error_start = io_dec_mem_ctrl_ifu_iccm_rd_ecc_single_err | io_dec_mem_ctrl_ifu_ic_error_start; // @[ifu_mem_ctl.scala 96:28]
  assign io_ic_fetch_val_f = {_T_1286,fetch_req_f_qual}; // @[ifu_mem_ctl.scala 305:21]
  assign io_ic_data_f = ic_final_data[31:0]; // @[ifu_mem_ctl.scala 298:16]
  assign rvclkhdr_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_io_en = ic_debug_rd_en_ff; // @[lib.scala 345:16]
  assign rvclkhdr_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_1_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_1_io_en = io_ic_debug_rd_en | io_ic_debug_wr_en; // @[lib.scala 345:16]
  assign rvclkhdr_1_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_2_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_2_io_en = _T_2 | scnd_miss_req; // @[lib.scala 345:16]
  assign rvclkhdr_2_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_3_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_3_io_en = _T_309 | io_dec_mem_ctrl_dec_tlu_force_halt; // @[lib.scala 345:16]
  assign rvclkhdr_3_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_4_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_4_io_en = bus_ifu_wr_en & _T_1289; // @[lib.scala 345:16]
  assign rvclkhdr_4_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_5_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_5_io_en = bus_ifu_wr_en & _T_1290; // @[lib.scala 345:16]
  assign rvclkhdr_5_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_6_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_6_io_en = bus_ifu_wr_en & _T_1291; // @[lib.scala 345:16]
  assign rvclkhdr_6_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_7_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_7_io_en = bus_ifu_wr_en & _T_1292; // @[lib.scala 345:16]
  assign rvclkhdr_7_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_8_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_8_io_en = bus_ifu_wr_en & _T_1293; // @[lib.scala 345:16]
  assign rvclkhdr_8_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_9_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_9_io_en = bus_ifu_wr_en & _T_1294; // @[lib.scala 345:16]
  assign rvclkhdr_9_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_10_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_10_io_en = bus_ifu_wr_en & _T_1295; // @[lib.scala 345:16]
  assign rvclkhdr_10_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_11_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_11_io_en = bus_ifu_wr_en & _T_1296; // @[lib.scala 345:16]
  assign rvclkhdr_11_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_12_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_12_io_en = bus_ifu_wr_en & _T_1289; // @[lib.scala 345:16]
  assign rvclkhdr_12_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_13_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_13_io_en = bus_ifu_wr_en & _T_1290; // @[lib.scala 345:16]
  assign rvclkhdr_13_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_14_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_14_io_en = bus_ifu_wr_en & _T_1291; // @[lib.scala 345:16]
  assign rvclkhdr_14_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_15_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_15_io_en = bus_ifu_wr_en & _T_1292; // @[lib.scala 345:16]
  assign rvclkhdr_15_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_16_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_16_io_en = bus_ifu_wr_en & _T_1293; // @[lib.scala 345:16]
  assign rvclkhdr_16_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_17_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_17_io_en = bus_ifu_wr_en & _T_1294; // @[lib.scala 345:16]
  assign rvclkhdr_17_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_18_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_18_io_en = bus_ifu_wr_en & _T_1295; // @[lib.scala 345:16]
  assign rvclkhdr_18_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_19_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_19_io_en = bus_ifu_wr_en & _T_1296; // @[lib.scala 345:16]
  assign rvclkhdr_19_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_20_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_20_io_en = bus_ifu_wr_en & _T_1289; // @[lib.scala 345:16]
  assign rvclkhdr_20_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_21_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_21_io_en = bus_ifu_wr_en & _T_1290; // @[lib.scala 345:16]
  assign rvclkhdr_21_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_22_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_22_io_en = bus_ifu_wr_en & _T_1291; // @[lib.scala 345:16]
  assign rvclkhdr_22_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_23_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_23_io_en = bus_ifu_wr_en & _T_1292; // @[lib.scala 345:16]
  assign rvclkhdr_23_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_24_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_24_io_en = bus_ifu_wr_en & _T_1293; // @[lib.scala 345:16]
  assign rvclkhdr_24_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_25_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_25_io_en = bus_ifu_wr_en & _T_1294; // @[lib.scala 345:16]
  assign rvclkhdr_25_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_26_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_26_io_en = bus_ifu_wr_en & _T_1295; // @[lib.scala 345:16]
  assign rvclkhdr_26_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_27_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_27_io_en = bus_ifu_wr_en & _T_1296; // @[lib.scala 345:16]
  assign rvclkhdr_27_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_28_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_28_io_en = bus_ifu_wr_en & _T_1289; // @[lib.scala 345:16]
  assign rvclkhdr_28_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_29_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_29_io_en = bus_ifu_wr_en & _T_1290; // @[lib.scala 345:16]
  assign rvclkhdr_29_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_30_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_30_io_en = bus_ifu_wr_en & _T_1291; // @[lib.scala 345:16]
  assign rvclkhdr_30_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_31_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_31_io_en = bus_ifu_wr_en & _T_1292; // @[lib.scala 345:16]
  assign rvclkhdr_31_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_32_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_32_io_en = bus_ifu_wr_en & _T_1293; // @[lib.scala 345:16]
  assign rvclkhdr_32_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_33_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_33_io_en = bus_ifu_wr_en & _T_1294; // @[lib.scala 345:16]
  assign rvclkhdr_33_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_34_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_34_io_en = bus_ifu_wr_en & _T_1295; // @[lib.scala 345:16]
  assign rvclkhdr_34_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_35_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_35_io_en = bus_ifu_wr_en & _T_1296; // @[lib.scala 345:16]
  assign rvclkhdr_35_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_36_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_36_io_en = bus_ifu_wr_en & _T_1289; // @[lib.scala 345:16]
  assign rvclkhdr_36_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_37_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_37_io_en = bus_ifu_wr_en & _T_1290; // @[lib.scala 345:16]
  assign rvclkhdr_37_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_38_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_38_io_en = bus_ifu_wr_en & _T_1291; // @[lib.scala 345:16]
  assign rvclkhdr_38_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_39_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_39_io_en = bus_ifu_wr_en & _T_1292; // @[lib.scala 345:16]
  assign rvclkhdr_39_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_40_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_40_io_en = bus_ifu_wr_en & _T_1293; // @[lib.scala 345:16]
  assign rvclkhdr_40_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_41_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_41_io_en = bus_ifu_wr_en & _T_1294; // @[lib.scala 345:16]
  assign rvclkhdr_41_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_42_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_42_io_en = bus_ifu_wr_en & _T_1295; // @[lib.scala 345:16]
  assign rvclkhdr_42_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_43_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_43_io_en = bus_ifu_wr_en & _T_1296; // @[lib.scala 345:16]
  assign rvclkhdr_43_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_44_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_44_io_en = bus_ifu_wr_en & _T_1289; // @[lib.scala 345:16]
  assign rvclkhdr_44_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_45_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_45_io_en = bus_ifu_wr_en & _T_1290; // @[lib.scala 345:16]
  assign rvclkhdr_45_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_46_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_46_io_en = bus_ifu_wr_en & _T_1291; // @[lib.scala 345:16]
  assign rvclkhdr_46_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_47_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_47_io_en = bus_ifu_wr_en & _T_1292; // @[lib.scala 345:16]
  assign rvclkhdr_47_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_48_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_48_io_en = bus_ifu_wr_en & _T_1293; // @[lib.scala 345:16]
  assign rvclkhdr_48_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_49_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_49_io_en = bus_ifu_wr_en & _T_1294; // @[lib.scala 345:16]
  assign rvclkhdr_49_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_50_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_50_io_en = bus_ifu_wr_en & _T_1295; // @[lib.scala 345:16]
  assign rvclkhdr_50_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_51_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_51_io_en = bus_ifu_wr_en & _T_1296; // @[lib.scala 345:16]
  assign rvclkhdr_51_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_52_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_52_io_en = bus_ifu_wr_en & _T_1289; // @[lib.scala 345:16]
  assign rvclkhdr_52_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_53_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_53_io_en = bus_ifu_wr_en & _T_1290; // @[lib.scala 345:16]
  assign rvclkhdr_53_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_54_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_54_io_en = bus_ifu_wr_en & _T_1291; // @[lib.scala 345:16]
  assign rvclkhdr_54_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_55_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_55_io_en = bus_ifu_wr_en & _T_1292; // @[lib.scala 345:16]
  assign rvclkhdr_55_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_56_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_56_io_en = bus_ifu_wr_en & _T_1293; // @[lib.scala 345:16]
  assign rvclkhdr_56_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_57_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_57_io_en = bus_ifu_wr_en & _T_1294; // @[lib.scala 345:16]
  assign rvclkhdr_57_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_58_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_58_io_en = bus_ifu_wr_en & _T_1295; // @[lib.scala 345:16]
  assign rvclkhdr_58_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_59_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_59_io_en = bus_ifu_wr_en & _T_1296; // @[lib.scala 345:16]
  assign rvclkhdr_59_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_60_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_60_io_en = bus_ifu_wr_en & _T_1289; // @[lib.scala 345:16]
  assign rvclkhdr_60_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_61_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_61_io_en = bus_ifu_wr_en & _T_1290; // @[lib.scala 345:16]
  assign rvclkhdr_61_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_62_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_62_io_en = bus_ifu_wr_en & _T_1291; // @[lib.scala 345:16]
  assign rvclkhdr_62_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_63_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_63_io_en = bus_ifu_wr_en & _T_1292; // @[lib.scala 345:16]
  assign rvclkhdr_63_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_64_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_64_io_en = bus_ifu_wr_en & _T_1293; // @[lib.scala 345:16]
  assign rvclkhdr_64_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_65_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_65_io_en = bus_ifu_wr_en & _T_1294; // @[lib.scala 345:16]
  assign rvclkhdr_65_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_66_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_66_io_en = bus_ifu_wr_en & _T_1295; // @[lib.scala 345:16]
  assign rvclkhdr_66_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_67_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_67_io_en = bus_ifu_wr_en & _T_1296; // @[lib.scala 345:16]
  assign rvclkhdr_67_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_68_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_68_io_en = io_ifu_bus_clk_en; // @[lib.scala 345:16]
  assign rvclkhdr_68_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_69_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_69_io_en = io_ifu_bus_clk_en | io_dec_mem_ctrl_dec_tlu_force_halt; // @[lib.scala 345:16]
  assign rvclkhdr_69_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_70_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_70_io_en = ifu_status_wr_addr_ff[6:3] == 4'h0; // @[lib.scala 345:16]
  assign rvclkhdr_70_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_71_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_71_io_en = ifu_status_wr_addr_ff[6:3] == 4'h1; // @[lib.scala 345:16]
  assign rvclkhdr_71_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_72_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_72_io_en = ifu_status_wr_addr_ff[6:3] == 4'h2; // @[lib.scala 345:16]
  assign rvclkhdr_72_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_73_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_73_io_en = ifu_status_wr_addr_ff[6:3] == 4'h3; // @[lib.scala 345:16]
  assign rvclkhdr_73_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_74_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_74_io_en = ifu_status_wr_addr_ff[6:3] == 4'h4; // @[lib.scala 345:16]
  assign rvclkhdr_74_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_75_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_75_io_en = ifu_status_wr_addr_ff[6:3] == 4'h5; // @[lib.scala 345:16]
  assign rvclkhdr_75_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_76_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_76_io_en = ifu_status_wr_addr_ff[6:3] == 4'h6; // @[lib.scala 345:16]
  assign rvclkhdr_76_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_77_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_77_io_en = ifu_status_wr_addr_ff[6:3] == 4'h7; // @[lib.scala 345:16]
  assign rvclkhdr_77_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_78_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_78_io_en = ifu_status_wr_addr_ff[6:3] == 4'h8; // @[lib.scala 345:16]
  assign rvclkhdr_78_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_79_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_79_io_en = ifu_status_wr_addr_ff[6:3] == 4'h9; // @[lib.scala 345:16]
  assign rvclkhdr_79_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_80_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_80_io_en = ifu_status_wr_addr_ff[6:3] == 4'ha; // @[lib.scala 345:16]
  assign rvclkhdr_80_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_81_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_81_io_en = ifu_status_wr_addr_ff[6:3] == 4'hb; // @[lib.scala 345:16]
  assign rvclkhdr_81_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_82_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_82_io_en = ifu_status_wr_addr_ff[6:3] == 4'hc; // @[lib.scala 345:16]
  assign rvclkhdr_82_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_83_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_83_io_en = ifu_status_wr_addr_ff[6:3] == 4'hd; // @[lib.scala 345:16]
  assign rvclkhdr_83_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_84_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_84_io_en = ifu_status_wr_addr_ff[6:3] == 4'he; // @[lib.scala 345:16]
  assign rvclkhdr_84_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_85_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_85_io_en = ifu_status_wr_addr_ff[6:3] == 4'hf; // @[lib.scala 345:16]
  assign rvclkhdr_85_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_86_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_86_io_en = tag_valid_clken_0[0]; // @[lib.scala 345:16]
  assign rvclkhdr_86_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_87_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_87_io_en = tag_valid_clken_0[1]; // @[lib.scala 345:16]
  assign rvclkhdr_87_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_88_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_88_io_en = tag_valid_clken_1[0]; // @[lib.scala 345:16]
  assign rvclkhdr_88_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_89_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_89_io_en = tag_valid_clken_1[1]; // @[lib.scala 345:16]
  assign rvclkhdr_89_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_90_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_90_io_en = tag_valid_clken_2[0]; // @[lib.scala 345:16]
  assign rvclkhdr_90_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_91_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_91_io_en = tag_valid_clken_2[1]; // @[lib.scala 345:16]
  assign rvclkhdr_91_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_92_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_92_io_en = tag_valid_clken_3[0]; // @[lib.scala 345:16]
  assign rvclkhdr_92_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_93_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_93_io_en = tag_valid_clken_3[1]; // @[lib.scala 345:16]
  assign rvclkhdr_93_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  flush_final_f = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  ifc_fetch_req_f_raw = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  miss_state = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  scnd_miss_req_q = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  ifu_fetch_addr_int_f = _RAND_4[30:0];
  _RAND_5 = {1{`RANDOM}};
  ifc_iccm_access_f = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  iccm_dma_rvalid_in = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  dma_iccm_req_f = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  perr_state = _RAND_8[2:0];
  _RAND_9 = {1{`RANDOM}};
  err_stop_state = _RAND_9[1:0];
  _RAND_10 = {1{`RANDOM}};
  reset_all_tags = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  ifc_region_acc_fault_final_f = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  ifu_bus_rvalid_unq_ff = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  bus_ifu_bus_clk_en_ff = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  uncacheable_miss_ff = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  bus_data_beat_count = _RAND_15[2:0];
  _RAND_16 = {1{`RANDOM}};
  ic_miss_buff_data_valid = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  imb_ff = _RAND_17[30:0];
  _RAND_18 = {1{`RANDOM}};
  last_data_recieved_ff = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  sel_mb_addr_ff = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  way_status_mb_scnd_ff = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  ifu_ic_rw_int_addr_ff = _RAND_21[6:0];
  _RAND_22 = {1{`RANDOM}};
  way_status_out_0 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  way_status_out_1 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  way_status_out_2 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  way_status_out_3 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  way_status_out_4 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  way_status_out_5 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  way_status_out_6 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  way_status_out_7 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  way_status_out_8 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  way_status_out_9 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  way_status_out_10 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  way_status_out_11 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  way_status_out_12 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  way_status_out_13 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  way_status_out_14 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  way_status_out_15 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  way_status_out_16 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  way_status_out_17 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  way_status_out_18 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  way_status_out_19 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  way_status_out_20 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  way_status_out_21 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  way_status_out_22 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  way_status_out_23 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  way_status_out_24 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  way_status_out_25 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  way_status_out_26 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  way_status_out_27 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  way_status_out_28 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  way_status_out_29 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  way_status_out_30 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  way_status_out_31 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  way_status_out_32 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  way_status_out_33 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  way_status_out_34 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  way_status_out_35 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  way_status_out_36 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  way_status_out_37 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  way_status_out_38 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  way_status_out_39 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  way_status_out_40 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  way_status_out_41 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  way_status_out_42 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  way_status_out_43 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  way_status_out_44 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  way_status_out_45 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  way_status_out_46 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  way_status_out_47 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  way_status_out_48 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  way_status_out_49 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  way_status_out_50 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  way_status_out_51 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  way_status_out_52 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  way_status_out_53 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  way_status_out_54 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  way_status_out_55 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  way_status_out_56 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  way_status_out_57 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  way_status_out_58 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  way_status_out_59 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  way_status_out_60 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  way_status_out_61 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  way_status_out_62 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  way_status_out_63 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  way_status_out_64 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  way_status_out_65 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  way_status_out_66 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  way_status_out_67 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  way_status_out_68 = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  way_status_out_69 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  way_status_out_70 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  way_status_out_71 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  way_status_out_72 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  way_status_out_73 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  way_status_out_74 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  way_status_out_75 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  way_status_out_76 = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  way_status_out_77 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  way_status_out_78 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  way_status_out_79 = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  way_status_out_80 = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  way_status_out_81 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  way_status_out_82 = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  way_status_out_83 = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  way_status_out_84 = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  way_status_out_85 = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  way_status_out_86 = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  way_status_out_87 = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  way_status_out_88 = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  way_status_out_89 = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  way_status_out_90 = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  way_status_out_91 = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  way_status_out_92 = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  way_status_out_93 = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  way_status_out_94 = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  way_status_out_95 = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  way_status_out_96 = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  way_status_out_97 = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  way_status_out_98 = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  way_status_out_99 = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  way_status_out_100 = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  way_status_out_101 = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  way_status_out_102 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  way_status_out_103 = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  way_status_out_104 = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  way_status_out_105 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  way_status_out_106 = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  way_status_out_107 = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  way_status_out_108 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  way_status_out_109 = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  way_status_out_110 = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  way_status_out_111 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  way_status_out_112 = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  way_status_out_113 = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  way_status_out_114 = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  way_status_out_115 = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  way_status_out_116 = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  way_status_out_117 = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  way_status_out_118 = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  way_status_out_119 = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  way_status_out_120 = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  way_status_out_121 = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  way_status_out_122 = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  way_status_out_123 = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  way_status_out_124 = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  way_status_out_125 = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  way_status_out_126 = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  way_status_out_127 = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  tagv_mb_scnd_ff = _RAND_150[1:0];
  _RAND_151 = {1{`RANDOM}};
  uncacheable_miss_scnd_ff = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  imb_scnd_ff = _RAND_152[30:0];
  _RAND_153 = {1{`RANDOM}};
  ifu_bus_rid_ff = _RAND_153[2:0];
  _RAND_154 = {1{`RANDOM}};
  ifu_bus_rresp_ff = _RAND_154[1:0];
  _RAND_155 = {1{`RANDOM}};
  ifu_wr_data_comb_err_ff = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  way_status_mb_ff = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  tagv_mb_ff = _RAND_157[1:0];
  _RAND_158 = {1{`RANDOM}};
  reset_ic_ff = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  fetch_uncacheable_ff = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  miss_addr = _RAND_160[25:0];
  _RAND_161 = {1{`RANDOM}};
  ifc_region_acc_fault_f = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  bus_rd_addr_count = _RAND_162[2:0];
  _RAND_163 = {1{`RANDOM}};
  ic_act_miss_f_delayed = _RAND_163[0:0];
  _RAND_164 = {2{`RANDOM}};
  ifu_bus_rdata_ff = _RAND_164[63:0];
  _RAND_165 = {1{`RANDOM}};
  ic_miss_buff_data_0 = _RAND_165[31:0];
  _RAND_166 = {1{`RANDOM}};
  ic_miss_buff_data_1 = _RAND_166[31:0];
  _RAND_167 = {1{`RANDOM}};
  ic_miss_buff_data_2 = _RAND_167[31:0];
  _RAND_168 = {1{`RANDOM}};
  ic_miss_buff_data_3 = _RAND_168[31:0];
  _RAND_169 = {1{`RANDOM}};
  ic_miss_buff_data_4 = _RAND_169[31:0];
  _RAND_170 = {1{`RANDOM}};
  ic_miss_buff_data_5 = _RAND_170[31:0];
  _RAND_171 = {1{`RANDOM}};
  ic_miss_buff_data_6 = _RAND_171[31:0];
  _RAND_172 = {1{`RANDOM}};
  ic_miss_buff_data_7 = _RAND_172[31:0];
  _RAND_173 = {1{`RANDOM}};
  ic_miss_buff_data_8 = _RAND_173[31:0];
  _RAND_174 = {1{`RANDOM}};
  ic_miss_buff_data_9 = _RAND_174[31:0];
  _RAND_175 = {1{`RANDOM}};
  ic_miss_buff_data_10 = _RAND_175[31:0];
  _RAND_176 = {1{`RANDOM}};
  ic_miss_buff_data_11 = _RAND_176[31:0];
  _RAND_177 = {1{`RANDOM}};
  ic_miss_buff_data_12 = _RAND_177[31:0];
  _RAND_178 = {1{`RANDOM}};
  ic_miss_buff_data_13 = _RAND_178[31:0];
  _RAND_179 = {1{`RANDOM}};
  ic_miss_buff_data_14 = _RAND_179[31:0];
  _RAND_180 = {1{`RANDOM}};
  ic_miss_buff_data_15 = _RAND_180[31:0];
  _RAND_181 = {1{`RANDOM}};
  ic_crit_wd_rdy_new_ff = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  ic_miss_buff_data_error = _RAND_182[7:0];
  _RAND_183 = {1{`RANDOM}};
  ic_debug_ict_array_sel_ff = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  ic_tag_valid_out_1_0 = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  ic_tag_valid_out_1_1 = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  ic_tag_valid_out_1_2 = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  ic_tag_valid_out_1_3 = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  ic_tag_valid_out_1_4 = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  ic_tag_valid_out_1_5 = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  ic_tag_valid_out_1_6 = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  ic_tag_valid_out_1_7 = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  ic_tag_valid_out_1_8 = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  ic_tag_valid_out_1_9 = _RAND_193[0:0];
  _RAND_194 = {1{`RANDOM}};
  ic_tag_valid_out_1_10 = _RAND_194[0:0];
  _RAND_195 = {1{`RANDOM}};
  ic_tag_valid_out_1_11 = _RAND_195[0:0];
  _RAND_196 = {1{`RANDOM}};
  ic_tag_valid_out_1_12 = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  ic_tag_valid_out_1_13 = _RAND_197[0:0];
  _RAND_198 = {1{`RANDOM}};
  ic_tag_valid_out_1_14 = _RAND_198[0:0];
  _RAND_199 = {1{`RANDOM}};
  ic_tag_valid_out_1_15 = _RAND_199[0:0];
  _RAND_200 = {1{`RANDOM}};
  ic_tag_valid_out_1_16 = _RAND_200[0:0];
  _RAND_201 = {1{`RANDOM}};
  ic_tag_valid_out_1_17 = _RAND_201[0:0];
  _RAND_202 = {1{`RANDOM}};
  ic_tag_valid_out_1_18 = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  ic_tag_valid_out_1_19 = _RAND_203[0:0];
  _RAND_204 = {1{`RANDOM}};
  ic_tag_valid_out_1_20 = _RAND_204[0:0];
  _RAND_205 = {1{`RANDOM}};
  ic_tag_valid_out_1_21 = _RAND_205[0:0];
  _RAND_206 = {1{`RANDOM}};
  ic_tag_valid_out_1_22 = _RAND_206[0:0];
  _RAND_207 = {1{`RANDOM}};
  ic_tag_valid_out_1_23 = _RAND_207[0:0];
  _RAND_208 = {1{`RANDOM}};
  ic_tag_valid_out_1_24 = _RAND_208[0:0];
  _RAND_209 = {1{`RANDOM}};
  ic_tag_valid_out_1_25 = _RAND_209[0:0];
  _RAND_210 = {1{`RANDOM}};
  ic_tag_valid_out_1_26 = _RAND_210[0:0];
  _RAND_211 = {1{`RANDOM}};
  ic_tag_valid_out_1_27 = _RAND_211[0:0];
  _RAND_212 = {1{`RANDOM}};
  ic_tag_valid_out_1_28 = _RAND_212[0:0];
  _RAND_213 = {1{`RANDOM}};
  ic_tag_valid_out_1_29 = _RAND_213[0:0];
  _RAND_214 = {1{`RANDOM}};
  ic_tag_valid_out_1_30 = _RAND_214[0:0];
  _RAND_215 = {1{`RANDOM}};
  ic_tag_valid_out_1_31 = _RAND_215[0:0];
  _RAND_216 = {1{`RANDOM}};
  ic_tag_valid_out_1_32 = _RAND_216[0:0];
  _RAND_217 = {1{`RANDOM}};
  ic_tag_valid_out_1_33 = _RAND_217[0:0];
  _RAND_218 = {1{`RANDOM}};
  ic_tag_valid_out_1_34 = _RAND_218[0:0];
  _RAND_219 = {1{`RANDOM}};
  ic_tag_valid_out_1_35 = _RAND_219[0:0];
  _RAND_220 = {1{`RANDOM}};
  ic_tag_valid_out_1_36 = _RAND_220[0:0];
  _RAND_221 = {1{`RANDOM}};
  ic_tag_valid_out_1_37 = _RAND_221[0:0];
  _RAND_222 = {1{`RANDOM}};
  ic_tag_valid_out_1_38 = _RAND_222[0:0];
  _RAND_223 = {1{`RANDOM}};
  ic_tag_valid_out_1_39 = _RAND_223[0:0];
  _RAND_224 = {1{`RANDOM}};
  ic_tag_valid_out_1_40 = _RAND_224[0:0];
  _RAND_225 = {1{`RANDOM}};
  ic_tag_valid_out_1_41 = _RAND_225[0:0];
  _RAND_226 = {1{`RANDOM}};
  ic_tag_valid_out_1_42 = _RAND_226[0:0];
  _RAND_227 = {1{`RANDOM}};
  ic_tag_valid_out_1_43 = _RAND_227[0:0];
  _RAND_228 = {1{`RANDOM}};
  ic_tag_valid_out_1_44 = _RAND_228[0:0];
  _RAND_229 = {1{`RANDOM}};
  ic_tag_valid_out_1_45 = _RAND_229[0:0];
  _RAND_230 = {1{`RANDOM}};
  ic_tag_valid_out_1_46 = _RAND_230[0:0];
  _RAND_231 = {1{`RANDOM}};
  ic_tag_valid_out_1_47 = _RAND_231[0:0];
  _RAND_232 = {1{`RANDOM}};
  ic_tag_valid_out_1_48 = _RAND_232[0:0];
  _RAND_233 = {1{`RANDOM}};
  ic_tag_valid_out_1_49 = _RAND_233[0:0];
  _RAND_234 = {1{`RANDOM}};
  ic_tag_valid_out_1_50 = _RAND_234[0:0];
  _RAND_235 = {1{`RANDOM}};
  ic_tag_valid_out_1_51 = _RAND_235[0:0];
  _RAND_236 = {1{`RANDOM}};
  ic_tag_valid_out_1_52 = _RAND_236[0:0];
  _RAND_237 = {1{`RANDOM}};
  ic_tag_valid_out_1_53 = _RAND_237[0:0];
  _RAND_238 = {1{`RANDOM}};
  ic_tag_valid_out_1_54 = _RAND_238[0:0];
  _RAND_239 = {1{`RANDOM}};
  ic_tag_valid_out_1_55 = _RAND_239[0:0];
  _RAND_240 = {1{`RANDOM}};
  ic_tag_valid_out_1_56 = _RAND_240[0:0];
  _RAND_241 = {1{`RANDOM}};
  ic_tag_valid_out_1_57 = _RAND_241[0:0];
  _RAND_242 = {1{`RANDOM}};
  ic_tag_valid_out_1_58 = _RAND_242[0:0];
  _RAND_243 = {1{`RANDOM}};
  ic_tag_valid_out_1_59 = _RAND_243[0:0];
  _RAND_244 = {1{`RANDOM}};
  ic_tag_valid_out_1_60 = _RAND_244[0:0];
  _RAND_245 = {1{`RANDOM}};
  ic_tag_valid_out_1_61 = _RAND_245[0:0];
  _RAND_246 = {1{`RANDOM}};
  ic_tag_valid_out_1_62 = _RAND_246[0:0];
  _RAND_247 = {1{`RANDOM}};
  ic_tag_valid_out_1_63 = _RAND_247[0:0];
  _RAND_248 = {1{`RANDOM}};
  ic_tag_valid_out_1_64 = _RAND_248[0:0];
  _RAND_249 = {1{`RANDOM}};
  ic_tag_valid_out_1_65 = _RAND_249[0:0];
  _RAND_250 = {1{`RANDOM}};
  ic_tag_valid_out_1_66 = _RAND_250[0:0];
  _RAND_251 = {1{`RANDOM}};
  ic_tag_valid_out_1_67 = _RAND_251[0:0];
  _RAND_252 = {1{`RANDOM}};
  ic_tag_valid_out_1_68 = _RAND_252[0:0];
  _RAND_253 = {1{`RANDOM}};
  ic_tag_valid_out_1_69 = _RAND_253[0:0];
  _RAND_254 = {1{`RANDOM}};
  ic_tag_valid_out_1_70 = _RAND_254[0:0];
  _RAND_255 = {1{`RANDOM}};
  ic_tag_valid_out_1_71 = _RAND_255[0:0];
  _RAND_256 = {1{`RANDOM}};
  ic_tag_valid_out_1_72 = _RAND_256[0:0];
  _RAND_257 = {1{`RANDOM}};
  ic_tag_valid_out_1_73 = _RAND_257[0:0];
  _RAND_258 = {1{`RANDOM}};
  ic_tag_valid_out_1_74 = _RAND_258[0:0];
  _RAND_259 = {1{`RANDOM}};
  ic_tag_valid_out_1_75 = _RAND_259[0:0];
  _RAND_260 = {1{`RANDOM}};
  ic_tag_valid_out_1_76 = _RAND_260[0:0];
  _RAND_261 = {1{`RANDOM}};
  ic_tag_valid_out_1_77 = _RAND_261[0:0];
  _RAND_262 = {1{`RANDOM}};
  ic_tag_valid_out_1_78 = _RAND_262[0:0];
  _RAND_263 = {1{`RANDOM}};
  ic_tag_valid_out_1_79 = _RAND_263[0:0];
  _RAND_264 = {1{`RANDOM}};
  ic_tag_valid_out_1_80 = _RAND_264[0:0];
  _RAND_265 = {1{`RANDOM}};
  ic_tag_valid_out_1_81 = _RAND_265[0:0];
  _RAND_266 = {1{`RANDOM}};
  ic_tag_valid_out_1_82 = _RAND_266[0:0];
  _RAND_267 = {1{`RANDOM}};
  ic_tag_valid_out_1_83 = _RAND_267[0:0];
  _RAND_268 = {1{`RANDOM}};
  ic_tag_valid_out_1_84 = _RAND_268[0:0];
  _RAND_269 = {1{`RANDOM}};
  ic_tag_valid_out_1_85 = _RAND_269[0:0];
  _RAND_270 = {1{`RANDOM}};
  ic_tag_valid_out_1_86 = _RAND_270[0:0];
  _RAND_271 = {1{`RANDOM}};
  ic_tag_valid_out_1_87 = _RAND_271[0:0];
  _RAND_272 = {1{`RANDOM}};
  ic_tag_valid_out_1_88 = _RAND_272[0:0];
  _RAND_273 = {1{`RANDOM}};
  ic_tag_valid_out_1_89 = _RAND_273[0:0];
  _RAND_274 = {1{`RANDOM}};
  ic_tag_valid_out_1_90 = _RAND_274[0:0];
  _RAND_275 = {1{`RANDOM}};
  ic_tag_valid_out_1_91 = _RAND_275[0:0];
  _RAND_276 = {1{`RANDOM}};
  ic_tag_valid_out_1_92 = _RAND_276[0:0];
  _RAND_277 = {1{`RANDOM}};
  ic_tag_valid_out_1_93 = _RAND_277[0:0];
  _RAND_278 = {1{`RANDOM}};
  ic_tag_valid_out_1_94 = _RAND_278[0:0];
  _RAND_279 = {1{`RANDOM}};
  ic_tag_valid_out_1_95 = _RAND_279[0:0];
  _RAND_280 = {1{`RANDOM}};
  ic_tag_valid_out_1_96 = _RAND_280[0:0];
  _RAND_281 = {1{`RANDOM}};
  ic_tag_valid_out_1_97 = _RAND_281[0:0];
  _RAND_282 = {1{`RANDOM}};
  ic_tag_valid_out_1_98 = _RAND_282[0:0];
  _RAND_283 = {1{`RANDOM}};
  ic_tag_valid_out_1_99 = _RAND_283[0:0];
  _RAND_284 = {1{`RANDOM}};
  ic_tag_valid_out_1_100 = _RAND_284[0:0];
  _RAND_285 = {1{`RANDOM}};
  ic_tag_valid_out_1_101 = _RAND_285[0:0];
  _RAND_286 = {1{`RANDOM}};
  ic_tag_valid_out_1_102 = _RAND_286[0:0];
  _RAND_287 = {1{`RANDOM}};
  ic_tag_valid_out_1_103 = _RAND_287[0:0];
  _RAND_288 = {1{`RANDOM}};
  ic_tag_valid_out_1_104 = _RAND_288[0:0];
  _RAND_289 = {1{`RANDOM}};
  ic_tag_valid_out_1_105 = _RAND_289[0:0];
  _RAND_290 = {1{`RANDOM}};
  ic_tag_valid_out_1_106 = _RAND_290[0:0];
  _RAND_291 = {1{`RANDOM}};
  ic_tag_valid_out_1_107 = _RAND_291[0:0];
  _RAND_292 = {1{`RANDOM}};
  ic_tag_valid_out_1_108 = _RAND_292[0:0];
  _RAND_293 = {1{`RANDOM}};
  ic_tag_valid_out_1_109 = _RAND_293[0:0];
  _RAND_294 = {1{`RANDOM}};
  ic_tag_valid_out_1_110 = _RAND_294[0:0];
  _RAND_295 = {1{`RANDOM}};
  ic_tag_valid_out_1_111 = _RAND_295[0:0];
  _RAND_296 = {1{`RANDOM}};
  ic_tag_valid_out_1_112 = _RAND_296[0:0];
  _RAND_297 = {1{`RANDOM}};
  ic_tag_valid_out_1_113 = _RAND_297[0:0];
  _RAND_298 = {1{`RANDOM}};
  ic_tag_valid_out_1_114 = _RAND_298[0:0];
  _RAND_299 = {1{`RANDOM}};
  ic_tag_valid_out_1_115 = _RAND_299[0:0];
  _RAND_300 = {1{`RANDOM}};
  ic_tag_valid_out_1_116 = _RAND_300[0:0];
  _RAND_301 = {1{`RANDOM}};
  ic_tag_valid_out_1_117 = _RAND_301[0:0];
  _RAND_302 = {1{`RANDOM}};
  ic_tag_valid_out_1_118 = _RAND_302[0:0];
  _RAND_303 = {1{`RANDOM}};
  ic_tag_valid_out_1_119 = _RAND_303[0:0];
  _RAND_304 = {1{`RANDOM}};
  ic_tag_valid_out_1_120 = _RAND_304[0:0];
  _RAND_305 = {1{`RANDOM}};
  ic_tag_valid_out_1_121 = _RAND_305[0:0];
  _RAND_306 = {1{`RANDOM}};
  ic_tag_valid_out_1_122 = _RAND_306[0:0];
  _RAND_307 = {1{`RANDOM}};
  ic_tag_valid_out_1_123 = _RAND_307[0:0];
  _RAND_308 = {1{`RANDOM}};
  ic_tag_valid_out_1_124 = _RAND_308[0:0];
  _RAND_309 = {1{`RANDOM}};
  ic_tag_valid_out_1_125 = _RAND_309[0:0];
  _RAND_310 = {1{`RANDOM}};
  ic_tag_valid_out_1_126 = _RAND_310[0:0];
  _RAND_311 = {1{`RANDOM}};
  ic_tag_valid_out_1_127 = _RAND_311[0:0];
  _RAND_312 = {1{`RANDOM}};
  ic_tag_valid_out_0_0 = _RAND_312[0:0];
  _RAND_313 = {1{`RANDOM}};
  ic_tag_valid_out_0_1 = _RAND_313[0:0];
  _RAND_314 = {1{`RANDOM}};
  ic_tag_valid_out_0_2 = _RAND_314[0:0];
  _RAND_315 = {1{`RANDOM}};
  ic_tag_valid_out_0_3 = _RAND_315[0:0];
  _RAND_316 = {1{`RANDOM}};
  ic_tag_valid_out_0_4 = _RAND_316[0:0];
  _RAND_317 = {1{`RANDOM}};
  ic_tag_valid_out_0_5 = _RAND_317[0:0];
  _RAND_318 = {1{`RANDOM}};
  ic_tag_valid_out_0_6 = _RAND_318[0:0];
  _RAND_319 = {1{`RANDOM}};
  ic_tag_valid_out_0_7 = _RAND_319[0:0];
  _RAND_320 = {1{`RANDOM}};
  ic_tag_valid_out_0_8 = _RAND_320[0:0];
  _RAND_321 = {1{`RANDOM}};
  ic_tag_valid_out_0_9 = _RAND_321[0:0];
  _RAND_322 = {1{`RANDOM}};
  ic_tag_valid_out_0_10 = _RAND_322[0:0];
  _RAND_323 = {1{`RANDOM}};
  ic_tag_valid_out_0_11 = _RAND_323[0:0];
  _RAND_324 = {1{`RANDOM}};
  ic_tag_valid_out_0_12 = _RAND_324[0:0];
  _RAND_325 = {1{`RANDOM}};
  ic_tag_valid_out_0_13 = _RAND_325[0:0];
  _RAND_326 = {1{`RANDOM}};
  ic_tag_valid_out_0_14 = _RAND_326[0:0];
  _RAND_327 = {1{`RANDOM}};
  ic_tag_valid_out_0_15 = _RAND_327[0:0];
  _RAND_328 = {1{`RANDOM}};
  ic_tag_valid_out_0_16 = _RAND_328[0:0];
  _RAND_329 = {1{`RANDOM}};
  ic_tag_valid_out_0_17 = _RAND_329[0:0];
  _RAND_330 = {1{`RANDOM}};
  ic_tag_valid_out_0_18 = _RAND_330[0:0];
  _RAND_331 = {1{`RANDOM}};
  ic_tag_valid_out_0_19 = _RAND_331[0:0];
  _RAND_332 = {1{`RANDOM}};
  ic_tag_valid_out_0_20 = _RAND_332[0:0];
  _RAND_333 = {1{`RANDOM}};
  ic_tag_valid_out_0_21 = _RAND_333[0:0];
  _RAND_334 = {1{`RANDOM}};
  ic_tag_valid_out_0_22 = _RAND_334[0:0];
  _RAND_335 = {1{`RANDOM}};
  ic_tag_valid_out_0_23 = _RAND_335[0:0];
  _RAND_336 = {1{`RANDOM}};
  ic_tag_valid_out_0_24 = _RAND_336[0:0];
  _RAND_337 = {1{`RANDOM}};
  ic_tag_valid_out_0_25 = _RAND_337[0:0];
  _RAND_338 = {1{`RANDOM}};
  ic_tag_valid_out_0_26 = _RAND_338[0:0];
  _RAND_339 = {1{`RANDOM}};
  ic_tag_valid_out_0_27 = _RAND_339[0:0];
  _RAND_340 = {1{`RANDOM}};
  ic_tag_valid_out_0_28 = _RAND_340[0:0];
  _RAND_341 = {1{`RANDOM}};
  ic_tag_valid_out_0_29 = _RAND_341[0:0];
  _RAND_342 = {1{`RANDOM}};
  ic_tag_valid_out_0_30 = _RAND_342[0:0];
  _RAND_343 = {1{`RANDOM}};
  ic_tag_valid_out_0_31 = _RAND_343[0:0];
  _RAND_344 = {1{`RANDOM}};
  ic_tag_valid_out_0_32 = _RAND_344[0:0];
  _RAND_345 = {1{`RANDOM}};
  ic_tag_valid_out_0_33 = _RAND_345[0:0];
  _RAND_346 = {1{`RANDOM}};
  ic_tag_valid_out_0_34 = _RAND_346[0:0];
  _RAND_347 = {1{`RANDOM}};
  ic_tag_valid_out_0_35 = _RAND_347[0:0];
  _RAND_348 = {1{`RANDOM}};
  ic_tag_valid_out_0_36 = _RAND_348[0:0];
  _RAND_349 = {1{`RANDOM}};
  ic_tag_valid_out_0_37 = _RAND_349[0:0];
  _RAND_350 = {1{`RANDOM}};
  ic_tag_valid_out_0_38 = _RAND_350[0:0];
  _RAND_351 = {1{`RANDOM}};
  ic_tag_valid_out_0_39 = _RAND_351[0:0];
  _RAND_352 = {1{`RANDOM}};
  ic_tag_valid_out_0_40 = _RAND_352[0:0];
  _RAND_353 = {1{`RANDOM}};
  ic_tag_valid_out_0_41 = _RAND_353[0:0];
  _RAND_354 = {1{`RANDOM}};
  ic_tag_valid_out_0_42 = _RAND_354[0:0];
  _RAND_355 = {1{`RANDOM}};
  ic_tag_valid_out_0_43 = _RAND_355[0:0];
  _RAND_356 = {1{`RANDOM}};
  ic_tag_valid_out_0_44 = _RAND_356[0:0];
  _RAND_357 = {1{`RANDOM}};
  ic_tag_valid_out_0_45 = _RAND_357[0:0];
  _RAND_358 = {1{`RANDOM}};
  ic_tag_valid_out_0_46 = _RAND_358[0:0];
  _RAND_359 = {1{`RANDOM}};
  ic_tag_valid_out_0_47 = _RAND_359[0:0];
  _RAND_360 = {1{`RANDOM}};
  ic_tag_valid_out_0_48 = _RAND_360[0:0];
  _RAND_361 = {1{`RANDOM}};
  ic_tag_valid_out_0_49 = _RAND_361[0:0];
  _RAND_362 = {1{`RANDOM}};
  ic_tag_valid_out_0_50 = _RAND_362[0:0];
  _RAND_363 = {1{`RANDOM}};
  ic_tag_valid_out_0_51 = _RAND_363[0:0];
  _RAND_364 = {1{`RANDOM}};
  ic_tag_valid_out_0_52 = _RAND_364[0:0];
  _RAND_365 = {1{`RANDOM}};
  ic_tag_valid_out_0_53 = _RAND_365[0:0];
  _RAND_366 = {1{`RANDOM}};
  ic_tag_valid_out_0_54 = _RAND_366[0:0];
  _RAND_367 = {1{`RANDOM}};
  ic_tag_valid_out_0_55 = _RAND_367[0:0];
  _RAND_368 = {1{`RANDOM}};
  ic_tag_valid_out_0_56 = _RAND_368[0:0];
  _RAND_369 = {1{`RANDOM}};
  ic_tag_valid_out_0_57 = _RAND_369[0:0];
  _RAND_370 = {1{`RANDOM}};
  ic_tag_valid_out_0_58 = _RAND_370[0:0];
  _RAND_371 = {1{`RANDOM}};
  ic_tag_valid_out_0_59 = _RAND_371[0:0];
  _RAND_372 = {1{`RANDOM}};
  ic_tag_valid_out_0_60 = _RAND_372[0:0];
  _RAND_373 = {1{`RANDOM}};
  ic_tag_valid_out_0_61 = _RAND_373[0:0];
  _RAND_374 = {1{`RANDOM}};
  ic_tag_valid_out_0_62 = _RAND_374[0:0];
  _RAND_375 = {1{`RANDOM}};
  ic_tag_valid_out_0_63 = _RAND_375[0:0];
  _RAND_376 = {1{`RANDOM}};
  ic_tag_valid_out_0_64 = _RAND_376[0:0];
  _RAND_377 = {1{`RANDOM}};
  ic_tag_valid_out_0_65 = _RAND_377[0:0];
  _RAND_378 = {1{`RANDOM}};
  ic_tag_valid_out_0_66 = _RAND_378[0:0];
  _RAND_379 = {1{`RANDOM}};
  ic_tag_valid_out_0_67 = _RAND_379[0:0];
  _RAND_380 = {1{`RANDOM}};
  ic_tag_valid_out_0_68 = _RAND_380[0:0];
  _RAND_381 = {1{`RANDOM}};
  ic_tag_valid_out_0_69 = _RAND_381[0:0];
  _RAND_382 = {1{`RANDOM}};
  ic_tag_valid_out_0_70 = _RAND_382[0:0];
  _RAND_383 = {1{`RANDOM}};
  ic_tag_valid_out_0_71 = _RAND_383[0:0];
  _RAND_384 = {1{`RANDOM}};
  ic_tag_valid_out_0_72 = _RAND_384[0:0];
  _RAND_385 = {1{`RANDOM}};
  ic_tag_valid_out_0_73 = _RAND_385[0:0];
  _RAND_386 = {1{`RANDOM}};
  ic_tag_valid_out_0_74 = _RAND_386[0:0];
  _RAND_387 = {1{`RANDOM}};
  ic_tag_valid_out_0_75 = _RAND_387[0:0];
  _RAND_388 = {1{`RANDOM}};
  ic_tag_valid_out_0_76 = _RAND_388[0:0];
  _RAND_389 = {1{`RANDOM}};
  ic_tag_valid_out_0_77 = _RAND_389[0:0];
  _RAND_390 = {1{`RANDOM}};
  ic_tag_valid_out_0_78 = _RAND_390[0:0];
  _RAND_391 = {1{`RANDOM}};
  ic_tag_valid_out_0_79 = _RAND_391[0:0];
  _RAND_392 = {1{`RANDOM}};
  ic_tag_valid_out_0_80 = _RAND_392[0:0];
  _RAND_393 = {1{`RANDOM}};
  ic_tag_valid_out_0_81 = _RAND_393[0:0];
  _RAND_394 = {1{`RANDOM}};
  ic_tag_valid_out_0_82 = _RAND_394[0:0];
  _RAND_395 = {1{`RANDOM}};
  ic_tag_valid_out_0_83 = _RAND_395[0:0];
  _RAND_396 = {1{`RANDOM}};
  ic_tag_valid_out_0_84 = _RAND_396[0:0];
  _RAND_397 = {1{`RANDOM}};
  ic_tag_valid_out_0_85 = _RAND_397[0:0];
  _RAND_398 = {1{`RANDOM}};
  ic_tag_valid_out_0_86 = _RAND_398[0:0];
  _RAND_399 = {1{`RANDOM}};
  ic_tag_valid_out_0_87 = _RAND_399[0:0];
  _RAND_400 = {1{`RANDOM}};
  ic_tag_valid_out_0_88 = _RAND_400[0:0];
  _RAND_401 = {1{`RANDOM}};
  ic_tag_valid_out_0_89 = _RAND_401[0:0];
  _RAND_402 = {1{`RANDOM}};
  ic_tag_valid_out_0_90 = _RAND_402[0:0];
  _RAND_403 = {1{`RANDOM}};
  ic_tag_valid_out_0_91 = _RAND_403[0:0];
  _RAND_404 = {1{`RANDOM}};
  ic_tag_valid_out_0_92 = _RAND_404[0:0];
  _RAND_405 = {1{`RANDOM}};
  ic_tag_valid_out_0_93 = _RAND_405[0:0];
  _RAND_406 = {1{`RANDOM}};
  ic_tag_valid_out_0_94 = _RAND_406[0:0];
  _RAND_407 = {1{`RANDOM}};
  ic_tag_valid_out_0_95 = _RAND_407[0:0];
  _RAND_408 = {1{`RANDOM}};
  ic_tag_valid_out_0_96 = _RAND_408[0:0];
  _RAND_409 = {1{`RANDOM}};
  ic_tag_valid_out_0_97 = _RAND_409[0:0];
  _RAND_410 = {1{`RANDOM}};
  ic_tag_valid_out_0_98 = _RAND_410[0:0];
  _RAND_411 = {1{`RANDOM}};
  ic_tag_valid_out_0_99 = _RAND_411[0:0];
  _RAND_412 = {1{`RANDOM}};
  ic_tag_valid_out_0_100 = _RAND_412[0:0];
  _RAND_413 = {1{`RANDOM}};
  ic_tag_valid_out_0_101 = _RAND_413[0:0];
  _RAND_414 = {1{`RANDOM}};
  ic_tag_valid_out_0_102 = _RAND_414[0:0];
  _RAND_415 = {1{`RANDOM}};
  ic_tag_valid_out_0_103 = _RAND_415[0:0];
  _RAND_416 = {1{`RANDOM}};
  ic_tag_valid_out_0_104 = _RAND_416[0:0];
  _RAND_417 = {1{`RANDOM}};
  ic_tag_valid_out_0_105 = _RAND_417[0:0];
  _RAND_418 = {1{`RANDOM}};
  ic_tag_valid_out_0_106 = _RAND_418[0:0];
  _RAND_419 = {1{`RANDOM}};
  ic_tag_valid_out_0_107 = _RAND_419[0:0];
  _RAND_420 = {1{`RANDOM}};
  ic_tag_valid_out_0_108 = _RAND_420[0:0];
  _RAND_421 = {1{`RANDOM}};
  ic_tag_valid_out_0_109 = _RAND_421[0:0];
  _RAND_422 = {1{`RANDOM}};
  ic_tag_valid_out_0_110 = _RAND_422[0:0];
  _RAND_423 = {1{`RANDOM}};
  ic_tag_valid_out_0_111 = _RAND_423[0:0];
  _RAND_424 = {1{`RANDOM}};
  ic_tag_valid_out_0_112 = _RAND_424[0:0];
  _RAND_425 = {1{`RANDOM}};
  ic_tag_valid_out_0_113 = _RAND_425[0:0];
  _RAND_426 = {1{`RANDOM}};
  ic_tag_valid_out_0_114 = _RAND_426[0:0];
  _RAND_427 = {1{`RANDOM}};
  ic_tag_valid_out_0_115 = _RAND_427[0:0];
  _RAND_428 = {1{`RANDOM}};
  ic_tag_valid_out_0_116 = _RAND_428[0:0];
  _RAND_429 = {1{`RANDOM}};
  ic_tag_valid_out_0_117 = _RAND_429[0:0];
  _RAND_430 = {1{`RANDOM}};
  ic_tag_valid_out_0_118 = _RAND_430[0:0];
  _RAND_431 = {1{`RANDOM}};
  ic_tag_valid_out_0_119 = _RAND_431[0:0];
  _RAND_432 = {1{`RANDOM}};
  ic_tag_valid_out_0_120 = _RAND_432[0:0];
  _RAND_433 = {1{`RANDOM}};
  ic_tag_valid_out_0_121 = _RAND_433[0:0];
  _RAND_434 = {1{`RANDOM}};
  ic_tag_valid_out_0_122 = _RAND_434[0:0];
  _RAND_435 = {1{`RANDOM}};
  ic_tag_valid_out_0_123 = _RAND_435[0:0];
  _RAND_436 = {1{`RANDOM}};
  ic_tag_valid_out_0_124 = _RAND_436[0:0];
  _RAND_437 = {1{`RANDOM}};
  ic_tag_valid_out_0_125 = _RAND_437[0:0];
  _RAND_438 = {1{`RANDOM}};
  ic_tag_valid_out_0_126 = _RAND_438[0:0];
  _RAND_439 = {1{`RANDOM}};
  ic_tag_valid_out_0_127 = _RAND_439[0:0];
  _RAND_440 = {1{`RANDOM}};
  ic_debug_way_ff = _RAND_440[1:0];
  _RAND_441 = {1{`RANDOM}};
  ic_debug_rd_en_ff = _RAND_441[0:0];
  _RAND_442 = {3{`RANDOM}};
  _T_1212 = _RAND_442[70:0];
  _RAND_443 = {1{`RANDOM}};
  ifc_region_acc_fault_memory_f = _RAND_443[0:0];
  _RAND_444 = {1{`RANDOM}};
  perr_ic_index_ff = _RAND_444[6:0];
  _RAND_445 = {1{`RANDOM}};
  dma_sb_err_state_ff = _RAND_445[0:0];
  _RAND_446 = {1{`RANDOM}};
  bus_cmd_req_hold = _RAND_446[0:0];
  _RAND_447 = {1{`RANDOM}};
  ifu_bus_cmd_valid = _RAND_447[0:0];
  _RAND_448 = {1{`RANDOM}};
  bus_cmd_beat_count = _RAND_448[2:0];
  _RAND_449 = {1{`RANDOM}};
  ifu_bus_arready_unq_ff = _RAND_449[0:0];
  _RAND_450 = {1{`RANDOM}};
  ifu_bus_arvalid_ff = _RAND_450[0:0];
  _RAND_451 = {1{`RANDOM}};
  ifc_dma_access_ok_prev = _RAND_451[0:0];
  _RAND_452 = {2{`RANDOM}};
  iccm_ecc_corr_data_ff = _RAND_452[38:0];
  _RAND_453 = {1{`RANDOM}};
  dma_mem_addr_ff = _RAND_453[1:0];
  _RAND_454 = {1{`RANDOM}};
  dma_mem_tag_ff = _RAND_454[2:0];
  _RAND_455 = {1{`RANDOM}};
  iccm_dma_rtag_temp = _RAND_455[2:0];
  _RAND_456 = {1{`RANDOM}};
  iccm_dma_rvalid_temp = _RAND_456[0:0];
  _RAND_457 = {1{`RANDOM}};
  iccm_dma_ecc_error = _RAND_457[0:0];
  _RAND_458 = {2{`RANDOM}};
  iccm_dma_rdata_temp = _RAND_458[63:0];
  _RAND_459 = {1{`RANDOM}};
  iccm_ecc_corr_index_ff = _RAND_459[13:0];
  _RAND_460 = {1{`RANDOM}};
  iccm_rd_ecc_single_err_ff = _RAND_460[0:0];
  _RAND_461 = {1{`RANDOM}};
  iccm_rw_addr_f = _RAND_461[13:0];
  _RAND_462 = {1{`RANDOM}};
  ifu_status_wr_addr_ff = _RAND_462[6:0];
  _RAND_463 = {1{`RANDOM}};
  way_status_wr_en_ff = _RAND_463[0:0];
  _RAND_464 = {1{`RANDOM}};
  way_status_new_ff = _RAND_464[0:0];
  _RAND_465 = {1{`RANDOM}};
  ifu_tag_wren_ff = _RAND_465[1:0];
  _RAND_466 = {1{`RANDOM}};
  ic_valid_ff = _RAND_466[0:0];
  _RAND_467 = {1{`RANDOM}};
  _T_9799 = _RAND_467[0:0];
  _RAND_468 = {1{`RANDOM}};
  _T_9800 = _RAND_468[0:0];
  _RAND_469 = {1{`RANDOM}};
  _T_9801 = _RAND_469[0:0];
  _RAND_470 = {1{`RANDOM}};
  _T_9805 = _RAND_470[0:0];
  _RAND_471 = {1{`RANDOM}};
  _T_9806 = _RAND_471[0:0];
  _RAND_472 = {1{`RANDOM}};
  _T_9826 = _RAND_472[0:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    flush_final_f = 1'h0;
  end
  if (reset) begin
    ifc_fetch_req_f_raw = 1'h0;
  end
  if (reset) begin
    miss_state = 3'h0;
  end
  if (reset) begin
    scnd_miss_req_q = 1'h0;
  end
  if (reset) begin
    ifu_fetch_addr_int_f = 31'h0;
  end
  if (reset) begin
    ifc_iccm_access_f = 1'h0;
  end
  if (reset) begin
    iccm_dma_rvalid_in = 1'h0;
  end
  if (reset) begin
    dma_iccm_req_f = 1'h0;
  end
  if (reset) begin
    perr_state = 3'h0;
  end
  if (reset) begin
    err_stop_state = 2'h0;
  end
  if (reset) begin
    reset_all_tags = 1'h0;
  end
  if (reset) begin
    ifc_region_acc_fault_final_f = 1'h0;
  end
  if (reset) begin
    ifu_bus_rvalid_unq_ff = 1'h0;
  end
  if (reset) begin
    bus_ifu_bus_clk_en_ff = 1'h0;
  end
  if (reset) begin
    uncacheable_miss_ff = 1'h0;
  end
  if (reset) begin
    bus_data_beat_count = 3'h0;
  end
  if (reset) begin
    ic_miss_buff_data_valid = 8'h0;
  end
  if (reset) begin
    imb_ff = 31'h0;
  end
  if (reset) begin
    last_data_recieved_ff = 1'h0;
  end
  if (reset) begin
    sel_mb_addr_ff = 1'h0;
  end
  if (reset) begin
    way_status_mb_scnd_ff = 1'h0;
  end
  if (reset) begin
    ifu_ic_rw_int_addr_ff = 7'h0;
  end
  if (reset) begin
    way_status_out_0 = 1'h0;
  end
  if (reset) begin
    way_status_out_1 = 1'h0;
  end
  if (reset) begin
    way_status_out_2 = 1'h0;
  end
  if (reset) begin
    way_status_out_3 = 1'h0;
  end
  if (reset) begin
    way_status_out_4 = 1'h0;
  end
  if (reset) begin
    way_status_out_5 = 1'h0;
  end
  if (reset) begin
    way_status_out_6 = 1'h0;
  end
  if (reset) begin
    way_status_out_7 = 1'h0;
  end
  if (reset) begin
    way_status_out_8 = 1'h0;
  end
  if (reset) begin
    way_status_out_9 = 1'h0;
  end
  if (reset) begin
    way_status_out_10 = 1'h0;
  end
  if (reset) begin
    way_status_out_11 = 1'h0;
  end
  if (reset) begin
    way_status_out_12 = 1'h0;
  end
  if (reset) begin
    way_status_out_13 = 1'h0;
  end
  if (reset) begin
    way_status_out_14 = 1'h0;
  end
  if (reset) begin
    way_status_out_15 = 1'h0;
  end
  if (reset) begin
    way_status_out_16 = 1'h0;
  end
  if (reset) begin
    way_status_out_17 = 1'h0;
  end
  if (reset) begin
    way_status_out_18 = 1'h0;
  end
  if (reset) begin
    way_status_out_19 = 1'h0;
  end
  if (reset) begin
    way_status_out_20 = 1'h0;
  end
  if (reset) begin
    way_status_out_21 = 1'h0;
  end
  if (reset) begin
    way_status_out_22 = 1'h0;
  end
  if (reset) begin
    way_status_out_23 = 1'h0;
  end
  if (reset) begin
    way_status_out_24 = 1'h0;
  end
  if (reset) begin
    way_status_out_25 = 1'h0;
  end
  if (reset) begin
    way_status_out_26 = 1'h0;
  end
  if (reset) begin
    way_status_out_27 = 1'h0;
  end
  if (reset) begin
    way_status_out_28 = 1'h0;
  end
  if (reset) begin
    way_status_out_29 = 1'h0;
  end
  if (reset) begin
    way_status_out_30 = 1'h0;
  end
  if (reset) begin
    way_status_out_31 = 1'h0;
  end
  if (reset) begin
    way_status_out_32 = 1'h0;
  end
  if (reset) begin
    way_status_out_33 = 1'h0;
  end
  if (reset) begin
    way_status_out_34 = 1'h0;
  end
  if (reset) begin
    way_status_out_35 = 1'h0;
  end
  if (reset) begin
    way_status_out_36 = 1'h0;
  end
  if (reset) begin
    way_status_out_37 = 1'h0;
  end
  if (reset) begin
    way_status_out_38 = 1'h0;
  end
  if (reset) begin
    way_status_out_39 = 1'h0;
  end
  if (reset) begin
    way_status_out_40 = 1'h0;
  end
  if (reset) begin
    way_status_out_41 = 1'h0;
  end
  if (reset) begin
    way_status_out_42 = 1'h0;
  end
  if (reset) begin
    way_status_out_43 = 1'h0;
  end
  if (reset) begin
    way_status_out_44 = 1'h0;
  end
  if (reset) begin
    way_status_out_45 = 1'h0;
  end
  if (reset) begin
    way_status_out_46 = 1'h0;
  end
  if (reset) begin
    way_status_out_47 = 1'h0;
  end
  if (reset) begin
    way_status_out_48 = 1'h0;
  end
  if (reset) begin
    way_status_out_49 = 1'h0;
  end
  if (reset) begin
    way_status_out_50 = 1'h0;
  end
  if (reset) begin
    way_status_out_51 = 1'h0;
  end
  if (reset) begin
    way_status_out_52 = 1'h0;
  end
  if (reset) begin
    way_status_out_53 = 1'h0;
  end
  if (reset) begin
    way_status_out_54 = 1'h0;
  end
  if (reset) begin
    way_status_out_55 = 1'h0;
  end
  if (reset) begin
    way_status_out_56 = 1'h0;
  end
  if (reset) begin
    way_status_out_57 = 1'h0;
  end
  if (reset) begin
    way_status_out_58 = 1'h0;
  end
  if (reset) begin
    way_status_out_59 = 1'h0;
  end
  if (reset) begin
    way_status_out_60 = 1'h0;
  end
  if (reset) begin
    way_status_out_61 = 1'h0;
  end
  if (reset) begin
    way_status_out_62 = 1'h0;
  end
  if (reset) begin
    way_status_out_63 = 1'h0;
  end
  if (reset) begin
    way_status_out_64 = 1'h0;
  end
  if (reset) begin
    way_status_out_65 = 1'h0;
  end
  if (reset) begin
    way_status_out_66 = 1'h0;
  end
  if (reset) begin
    way_status_out_67 = 1'h0;
  end
  if (reset) begin
    way_status_out_68 = 1'h0;
  end
  if (reset) begin
    way_status_out_69 = 1'h0;
  end
  if (reset) begin
    way_status_out_70 = 1'h0;
  end
  if (reset) begin
    way_status_out_71 = 1'h0;
  end
  if (reset) begin
    way_status_out_72 = 1'h0;
  end
  if (reset) begin
    way_status_out_73 = 1'h0;
  end
  if (reset) begin
    way_status_out_74 = 1'h0;
  end
  if (reset) begin
    way_status_out_75 = 1'h0;
  end
  if (reset) begin
    way_status_out_76 = 1'h0;
  end
  if (reset) begin
    way_status_out_77 = 1'h0;
  end
  if (reset) begin
    way_status_out_78 = 1'h0;
  end
  if (reset) begin
    way_status_out_79 = 1'h0;
  end
  if (reset) begin
    way_status_out_80 = 1'h0;
  end
  if (reset) begin
    way_status_out_81 = 1'h0;
  end
  if (reset) begin
    way_status_out_82 = 1'h0;
  end
  if (reset) begin
    way_status_out_83 = 1'h0;
  end
  if (reset) begin
    way_status_out_84 = 1'h0;
  end
  if (reset) begin
    way_status_out_85 = 1'h0;
  end
  if (reset) begin
    way_status_out_86 = 1'h0;
  end
  if (reset) begin
    way_status_out_87 = 1'h0;
  end
  if (reset) begin
    way_status_out_88 = 1'h0;
  end
  if (reset) begin
    way_status_out_89 = 1'h0;
  end
  if (reset) begin
    way_status_out_90 = 1'h0;
  end
  if (reset) begin
    way_status_out_91 = 1'h0;
  end
  if (reset) begin
    way_status_out_92 = 1'h0;
  end
  if (reset) begin
    way_status_out_93 = 1'h0;
  end
  if (reset) begin
    way_status_out_94 = 1'h0;
  end
  if (reset) begin
    way_status_out_95 = 1'h0;
  end
  if (reset) begin
    way_status_out_96 = 1'h0;
  end
  if (reset) begin
    way_status_out_97 = 1'h0;
  end
  if (reset) begin
    way_status_out_98 = 1'h0;
  end
  if (reset) begin
    way_status_out_99 = 1'h0;
  end
  if (reset) begin
    way_status_out_100 = 1'h0;
  end
  if (reset) begin
    way_status_out_101 = 1'h0;
  end
  if (reset) begin
    way_status_out_102 = 1'h0;
  end
  if (reset) begin
    way_status_out_103 = 1'h0;
  end
  if (reset) begin
    way_status_out_104 = 1'h0;
  end
  if (reset) begin
    way_status_out_105 = 1'h0;
  end
  if (reset) begin
    way_status_out_106 = 1'h0;
  end
  if (reset) begin
    way_status_out_107 = 1'h0;
  end
  if (reset) begin
    way_status_out_108 = 1'h0;
  end
  if (reset) begin
    way_status_out_109 = 1'h0;
  end
  if (reset) begin
    way_status_out_110 = 1'h0;
  end
  if (reset) begin
    way_status_out_111 = 1'h0;
  end
  if (reset) begin
    way_status_out_112 = 1'h0;
  end
  if (reset) begin
    way_status_out_113 = 1'h0;
  end
  if (reset) begin
    way_status_out_114 = 1'h0;
  end
  if (reset) begin
    way_status_out_115 = 1'h0;
  end
  if (reset) begin
    way_status_out_116 = 1'h0;
  end
  if (reset) begin
    way_status_out_117 = 1'h0;
  end
  if (reset) begin
    way_status_out_118 = 1'h0;
  end
  if (reset) begin
    way_status_out_119 = 1'h0;
  end
  if (reset) begin
    way_status_out_120 = 1'h0;
  end
  if (reset) begin
    way_status_out_121 = 1'h0;
  end
  if (reset) begin
    way_status_out_122 = 1'h0;
  end
  if (reset) begin
    way_status_out_123 = 1'h0;
  end
  if (reset) begin
    way_status_out_124 = 1'h0;
  end
  if (reset) begin
    way_status_out_125 = 1'h0;
  end
  if (reset) begin
    way_status_out_126 = 1'h0;
  end
  if (reset) begin
    way_status_out_127 = 1'h0;
  end
  if (reset) begin
    tagv_mb_scnd_ff = 2'h0;
  end
  if (reset) begin
    uncacheable_miss_scnd_ff = 1'h0;
  end
  if (reset) begin
    imb_scnd_ff = 31'h0;
  end
  if (reset) begin
    ifu_bus_rid_ff = 3'h0;
  end
  if (reset) begin
    ifu_bus_rresp_ff = 2'h0;
  end
  if (reset) begin
    ifu_wr_data_comb_err_ff = 1'h0;
  end
  if (reset) begin
    way_status_mb_ff = 1'h0;
  end
  if (reset) begin
    tagv_mb_ff = 2'h0;
  end
  if (reset) begin
    reset_ic_ff = 1'h0;
  end
  if (reset) begin
    fetch_uncacheable_ff = 1'h0;
  end
  if (reset) begin
    miss_addr = 26'h0;
  end
  if (reset) begin
    ifc_region_acc_fault_f = 1'h0;
  end
  if (reset) begin
    bus_rd_addr_count = 3'h0;
  end
  if (reset) begin
    ic_act_miss_f_delayed = 1'h0;
  end
  if (reset) begin
    ifu_bus_rdata_ff = 64'h0;
  end
  if (reset) begin
    ic_miss_buff_data_0 = 32'h0;
  end
  if (reset) begin
    ic_miss_buff_data_1 = 32'h0;
  end
  if (reset) begin
    ic_miss_buff_data_2 = 32'h0;
  end
  if (reset) begin
    ic_miss_buff_data_3 = 32'h0;
  end
  if (reset) begin
    ic_miss_buff_data_4 = 32'h0;
  end
  if (reset) begin
    ic_miss_buff_data_5 = 32'h0;
  end
  if (reset) begin
    ic_miss_buff_data_6 = 32'h0;
  end
  if (reset) begin
    ic_miss_buff_data_7 = 32'h0;
  end
  if (reset) begin
    ic_miss_buff_data_8 = 32'h0;
  end
  if (reset) begin
    ic_miss_buff_data_9 = 32'h0;
  end
  if (reset) begin
    ic_miss_buff_data_10 = 32'h0;
  end
  if (reset) begin
    ic_miss_buff_data_11 = 32'h0;
  end
  if (reset) begin
    ic_miss_buff_data_12 = 32'h0;
  end
  if (reset) begin
    ic_miss_buff_data_13 = 32'h0;
  end
  if (reset) begin
    ic_miss_buff_data_14 = 32'h0;
  end
  if (reset) begin
    ic_miss_buff_data_15 = 32'h0;
  end
  if (reset) begin
    ic_crit_wd_rdy_new_ff = 1'h0;
  end
  if (reset) begin
    ic_miss_buff_data_error = 8'h0;
  end
  if (reset) begin
    ic_debug_ict_array_sel_ff = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_0 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_1 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_2 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_3 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_4 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_5 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_6 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_7 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_8 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_9 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_10 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_11 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_12 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_13 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_14 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_15 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_16 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_17 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_18 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_19 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_20 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_21 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_22 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_23 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_24 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_25 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_26 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_27 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_28 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_29 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_30 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_31 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_32 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_33 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_34 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_35 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_36 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_37 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_38 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_39 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_40 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_41 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_42 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_43 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_44 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_45 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_46 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_47 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_48 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_49 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_50 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_51 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_52 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_53 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_54 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_55 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_56 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_57 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_58 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_59 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_60 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_61 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_62 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_63 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_64 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_65 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_66 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_67 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_68 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_69 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_70 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_71 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_72 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_73 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_74 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_75 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_76 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_77 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_78 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_79 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_80 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_81 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_82 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_83 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_84 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_85 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_86 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_87 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_88 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_89 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_90 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_91 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_92 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_93 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_94 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_95 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_96 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_97 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_98 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_99 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_100 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_101 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_102 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_103 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_104 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_105 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_106 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_107 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_108 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_109 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_110 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_111 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_112 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_113 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_114 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_115 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_116 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_117 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_118 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_119 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_120 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_121 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_122 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_123 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_124 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_125 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_126 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_127 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_0 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_1 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_2 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_3 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_4 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_5 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_6 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_7 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_8 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_9 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_10 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_11 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_12 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_13 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_14 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_15 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_16 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_17 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_18 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_19 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_20 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_21 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_22 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_23 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_24 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_25 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_26 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_27 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_28 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_29 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_30 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_31 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_32 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_33 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_34 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_35 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_36 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_37 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_38 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_39 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_40 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_41 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_42 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_43 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_44 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_45 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_46 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_47 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_48 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_49 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_50 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_51 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_52 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_53 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_54 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_55 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_56 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_57 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_58 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_59 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_60 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_61 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_62 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_63 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_64 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_65 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_66 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_67 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_68 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_69 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_70 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_71 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_72 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_73 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_74 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_75 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_76 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_77 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_78 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_79 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_80 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_81 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_82 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_83 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_84 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_85 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_86 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_87 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_88 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_89 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_90 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_91 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_92 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_93 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_94 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_95 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_96 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_97 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_98 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_99 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_100 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_101 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_102 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_103 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_104 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_105 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_106 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_107 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_108 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_109 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_110 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_111 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_112 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_113 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_114 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_115 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_116 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_117 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_118 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_119 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_120 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_121 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_122 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_123 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_124 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_125 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_126 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_127 = 1'h0;
  end
  if (reset) begin
    ic_debug_way_ff = 2'h0;
  end
  if (reset) begin
    ic_debug_rd_en_ff = 1'h0;
  end
  if (reset) begin
    _T_1212 = 71'h0;
  end
  if (reset) begin
    ifc_region_acc_fault_memory_f = 1'h0;
  end
  if (reset) begin
    perr_ic_index_ff = 7'h0;
  end
  if (reset) begin
    dma_sb_err_state_ff = 1'h0;
  end
  if (reset) begin
    bus_cmd_req_hold = 1'h0;
  end
  if (reset) begin
    ifu_bus_cmd_valid = 1'h0;
  end
  if (reset) begin
    bus_cmd_beat_count = 3'h0;
  end
  if (reset) begin
    ifu_bus_arready_unq_ff = 1'h0;
  end
  if (reset) begin
    ifu_bus_arvalid_ff = 1'h0;
  end
  if (reset) begin
    ifc_dma_access_ok_prev = 1'h0;
  end
  if (reset) begin
    iccm_ecc_corr_data_ff = 39'h0;
  end
  if (reset) begin
    dma_mem_addr_ff = 2'h0;
  end
  if (reset) begin
    dma_mem_tag_ff = 3'h0;
  end
  if (reset) begin
    iccm_dma_rtag_temp = 3'h0;
  end
  if (reset) begin
    iccm_dma_rvalid_temp = 1'h0;
  end
  if (reset) begin
    iccm_dma_ecc_error = 1'h0;
  end
  if (reset) begin
    iccm_dma_rdata_temp = 64'h0;
  end
  if (reset) begin
    iccm_ecc_corr_index_ff = 14'h0;
  end
  if (reset) begin
    iccm_rd_ecc_single_err_ff = 1'h0;
  end
  if (reset) begin
    iccm_rw_addr_f = 14'h0;
  end
  if (reset) begin
    ifu_status_wr_addr_ff = 7'h0;
  end
  if (reset) begin
    way_status_wr_en_ff = 1'h0;
  end
  if (reset) begin
    way_status_new_ff = 1'h0;
  end
  if (reset) begin
    ifu_tag_wren_ff = 2'h0;
  end
  if (reset) begin
    ic_valid_ff = 1'h0;
  end
  if (reset) begin
    _T_9799 = 1'h0;
  end
  if (reset) begin
    _T_9800 = 1'h0;
  end
  if (reset) begin
    _T_9801 = 1'h0;
  end
  if (reset) begin
    _T_9805 = 1'h0;
  end
  if (reset) begin
    _T_9806 = 1'h0;
  end
  if (reset) begin
    _T_9826 = 1'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      flush_final_f <= 1'h0;
    end else begin
      flush_final_f <= io_exu_flush_final;
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      ifc_fetch_req_f_raw <= 1'h0;
    end else begin
      ifc_fetch_req_f_raw <= _T_317 & _T_318;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      miss_state <= 3'h0;
    end else if (miss_state_en) begin
      if (_T_24) begin
        if (_T_26) begin
          miss_state <= 3'h1;
        end else begin
          miss_state <= 3'h2;
        end
      end else if (_T_31) begin
        if (_T_36) begin
          miss_state <= 3'h0;
        end else if (_T_40) begin
          miss_state <= 3'h3;
        end else if (_T_47) begin
          miss_state <= 3'h4;
        end else if (_T_51) begin
          miss_state <= 3'h0;
        end else if (_T_61) begin
          miss_state <= 3'h6;
        end else if (_T_71) begin
          miss_state <= 3'h6;
        end else if (_T_79) begin
          miss_state <= 3'h0;
        end else if (_T_84) begin
          miss_state <= 3'h2;
        end else begin
          miss_state <= 3'h0;
        end
      end else if (_T_102) begin
        miss_state <= 3'h0;
      end else if (_T_106) begin
        if (_T_113) begin
          miss_state <= 3'h2;
        end else begin
          miss_state <= 3'h0;
        end
      end else if (_T_121) begin
        if (_T_126) begin
          miss_state <= 3'h2;
        end else begin
          miss_state <= 3'h0;
        end
      end else if (_T_132) begin
        if (_T_137) begin
          miss_state <= 3'h5;
        end else if (_T_143) begin
          miss_state <= 3'h7;
        end else begin
          miss_state <= 3'h0;
        end
      end else if (_T_151) begin
        if (io_dec_mem_ctrl_dec_tlu_force_halt) begin
          miss_state <= 3'h0;
        end else if (io_exu_flush_final) begin
          if (_T_32) begin
            miss_state <= 3'h0;
          end else begin
            miss_state <= 3'h2;
          end
        end else begin
          miss_state <= 3'h1;
        end
      end else if (_T_160) begin
        if (io_dec_mem_ctrl_dec_tlu_force_halt) begin
          miss_state <= 3'h0;
        end else if (io_exu_flush_final) begin
          if (_T_32) begin
            miss_state <= 3'h0;
          end else begin
            miss_state <= 3'h2;
          end
        end else begin
          miss_state <= 3'h0;
        end
      end else begin
        miss_state <= 3'h0;
      end
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      scnd_miss_req_q <= 1'h0;
    end else begin
      scnd_miss_req_q <= _T_22 & _T_319;
    end
  end
  always @(posedge rvclkhdr_2_io_l1clk or posedge reset) begin
    if (reset) begin
      ifu_fetch_addr_int_f <= 31'h0;
    end else begin
      ifu_fetch_addr_int_f <= io_ifc_fetch_addr_bf;
    end
  end
  always @(posedge rvclkhdr_2_io_l1clk or posedge reset) begin
    if (reset) begin
      ifc_iccm_access_f <= 1'h0;
    end else begin
      ifc_iccm_access_f <= io_ifc_iccm_access_bf;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      iccm_dma_rvalid_in <= 1'h0;
    end else begin
      iccm_dma_rvalid_in <= _T_2709 & _T_2713;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      dma_iccm_req_f <= 1'h0;
    end else begin
      dma_iccm_req_f <= io_dma_mem_ctl_dma_iccm_req;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      perr_state <= 3'h0;
    end else if (perr_state_en) begin
      if (_T_2500) begin
        if (io_iccm_dma_sb_error) begin
          perr_state <= 3'h4;
        end else if (_T_2502) begin
          perr_state <= 3'h1;
        end else begin
          perr_state <= 3'h2;
        end
      end else if (_T_2512) begin
        perr_state <= 3'h0;
      end else if (_T_2515) begin
        if (_T_2518) begin
          perr_state <= 3'h0;
        end else begin
          perr_state <= 3'h3;
        end
      end else if (_T_2522) begin
        if (io_dec_mem_ctrl_dec_tlu_force_halt) begin
          perr_state <= 3'h0;
        end else begin
          perr_state <= 3'h3;
        end
      end else begin
        perr_state <= 3'h0;
      end
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      err_stop_state <= 2'h0;
    end else if (err_stop_state_en) begin
      if (_T_2526) begin
        err_stop_state <= 2'h1;
      end else if (_T_2531) begin
        if (_T_2533) begin
          err_stop_state <= 2'h0;
        end else if (_T_2554) begin
          err_stop_state <= 2'h3;
        end else if (io_ifu_fetch_val[0]) begin
          err_stop_state <= 2'h2;
        end else begin
          err_stop_state <= 2'h1;
        end
      end else if (_T_2558) begin
        if (_T_2533) begin
          err_stop_state <= 2'h0;
        end else if (io_ifu_fetch_val[0]) begin
          err_stop_state <= 2'h3;
        end else begin
          err_stop_state <= 2'h2;
        end
      end else if (_T_2575) begin
        if (_T_2579) begin
          err_stop_state <= 2'h0;
        end else if (io_dec_mem_ctrl_dec_tlu_flush_err_wb) begin
          err_stop_state <= 2'h1;
        end else begin
          err_stop_state <= 2'h3;
        end
      end else begin
        err_stop_state <= 2'h0;
      end
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      reset_all_tags <= 1'h0;
    end else begin
      reset_all_tags <= io_dec_mem_ctrl_dec_tlu_fence_i_wb;
    end
  end
  always @(posedge rvclkhdr_2_io_l1clk or posedge reset) begin
    if (reset) begin
      ifc_region_acc_fault_final_f <= 1'h0;
    end else begin
      ifc_region_acc_fault_final_f <= io_ifc_region_acc_fault_bf | ifc_region_acc_fault_memory_bf;
    end
  end
  always @(posedge rvclkhdr_68_io_l1clk or posedge reset) begin
    if (reset) begin
      ifu_bus_rvalid_unq_ff <= 1'h0;
    end else begin
      ifu_bus_rvalid_unq_ff <= io_ifu_axi_r_valid;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      bus_ifu_bus_clk_en_ff <= 1'h0;
    end else begin
      bus_ifu_bus_clk_en_ff <= io_ifu_bus_clk_en;
    end
  end
  always @(posedge rvclkhdr_2_io_l1clk or posedge reset) begin
    if (reset) begin
      uncacheable_miss_ff <= 1'h0;
    end else if (scnd_miss_req) begin
      uncacheable_miss_ff <= uncacheable_miss_scnd_ff;
    end else if (!(sel_hold_imb)) begin
      uncacheable_miss_ff <= io_ifc_fetch_uncacheable_bf;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      bus_data_beat_count <= 3'h0;
    end else begin
      bus_data_beat_count <= _T_2631 | _T_2632;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      ic_miss_buff_data_valid <= 8'h0;
    end else begin
      ic_miss_buff_data_valid <= {_T_1358,ic_miss_buff_data_valid_in_0};
    end
  end
  always @(posedge rvclkhdr_2_io_l1clk or posedge reset) begin
    if (reset) begin
      imb_ff <= 31'h0;
    end else if (scnd_miss_req) begin
      imb_ff <= imb_scnd_ff;
    end else if (!(sel_hold_imb)) begin
      imb_ff <= io_ifc_fetch_addr_bf;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      last_data_recieved_ff <= 1'h0;
    end else begin
      last_data_recieved_ff <= _T_2639 | _T_2641;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      sel_mb_addr_ff <= 1'h0;
    end else begin
      sel_mb_addr_ff <= _T_334 | reset_tag_valid_for_miss;
    end
  end
  always @(posedge rvclkhdr_2_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_mb_scnd_ff <= 1'h0;
    end else if (!(_T_19)) begin
      way_status_mb_scnd_ff <= way_status;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      ifu_ic_rw_int_addr_ff <= 7'h0;
    end else if (_T_3997) begin
      ifu_ic_rw_int_addr_ff <= io_ic_debug_addr[9:3];
    end else begin
      ifu_ic_rw_int_addr_ff <= ifu_ic_rw_int_addr[11:5];
    end
  end
  always @(posedge rvclkhdr_70_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_0 <= 1'h0;
    end else if (_T_4021) begin
      way_status_out_0 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_70_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_1 <= 1'h0;
    end else if (_T_4025) begin
      way_status_out_1 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_70_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_2 <= 1'h0;
    end else if (_T_4029) begin
      way_status_out_2 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_70_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_3 <= 1'h0;
    end else if (_T_4033) begin
      way_status_out_3 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_70_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_4 <= 1'h0;
    end else if (_T_4037) begin
      way_status_out_4 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_70_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_5 <= 1'h0;
    end else if (_T_4041) begin
      way_status_out_5 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_70_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_6 <= 1'h0;
    end else if (_T_4045) begin
      way_status_out_6 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_70_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_7 <= 1'h0;
    end else if (_T_4049) begin
      way_status_out_7 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_71_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_8 <= 1'h0;
    end else if (_T_4021) begin
      way_status_out_8 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_71_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_9 <= 1'h0;
    end else if (_T_4025) begin
      way_status_out_9 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_71_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_10 <= 1'h0;
    end else if (_T_4029) begin
      way_status_out_10 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_71_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_11 <= 1'h0;
    end else if (_T_4033) begin
      way_status_out_11 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_71_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_12 <= 1'h0;
    end else if (_T_4037) begin
      way_status_out_12 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_71_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_13 <= 1'h0;
    end else if (_T_4041) begin
      way_status_out_13 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_71_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_14 <= 1'h0;
    end else if (_T_4045) begin
      way_status_out_14 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_71_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_15 <= 1'h0;
    end else if (_T_4049) begin
      way_status_out_15 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_72_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_16 <= 1'h0;
    end else if (_T_4021) begin
      way_status_out_16 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_72_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_17 <= 1'h0;
    end else if (_T_4025) begin
      way_status_out_17 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_72_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_18 <= 1'h0;
    end else if (_T_4029) begin
      way_status_out_18 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_72_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_19 <= 1'h0;
    end else if (_T_4033) begin
      way_status_out_19 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_72_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_20 <= 1'h0;
    end else if (_T_4037) begin
      way_status_out_20 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_72_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_21 <= 1'h0;
    end else if (_T_4041) begin
      way_status_out_21 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_72_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_22 <= 1'h0;
    end else if (_T_4045) begin
      way_status_out_22 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_72_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_23 <= 1'h0;
    end else if (_T_4049) begin
      way_status_out_23 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_73_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_24 <= 1'h0;
    end else if (_T_4021) begin
      way_status_out_24 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_73_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_25 <= 1'h0;
    end else if (_T_4025) begin
      way_status_out_25 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_73_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_26 <= 1'h0;
    end else if (_T_4029) begin
      way_status_out_26 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_73_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_27 <= 1'h0;
    end else if (_T_4033) begin
      way_status_out_27 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_73_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_28 <= 1'h0;
    end else if (_T_4037) begin
      way_status_out_28 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_73_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_29 <= 1'h0;
    end else if (_T_4041) begin
      way_status_out_29 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_73_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_30 <= 1'h0;
    end else if (_T_4045) begin
      way_status_out_30 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_73_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_31 <= 1'h0;
    end else if (_T_4049) begin
      way_status_out_31 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_74_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_32 <= 1'h0;
    end else if (_T_4021) begin
      way_status_out_32 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_74_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_33 <= 1'h0;
    end else if (_T_4025) begin
      way_status_out_33 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_74_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_34 <= 1'h0;
    end else if (_T_4029) begin
      way_status_out_34 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_74_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_35 <= 1'h0;
    end else if (_T_4033) begin
      way_status_out_35 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_74_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_36 <= 1'h0;
    end else if (_T_4037) begin
      way_status_out_36 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_74_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_37 <= 1'h0;
    end else if (_T_4041) begin
      way_status_out_37 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_74_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_38 <= 1'h0;
    end else if (_T_4045) begin
      way_status_out_38 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_74_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_39 <= 1'h0;
    end else if (_T_4049) begin
      way_status_out_39 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_75_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_40 <= 1'h0;
    end else if (_T_4021) begin
      way_status_out_40 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_75_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_41 <= 1'h0;
    end else if (_T_4025) begin
      way_status_out_41 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_75_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_42 <= 1'h0;
    end else if (_T_4029) begin
      way_status_out_42 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_75_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_43 <= 1'h0;
    end else if (_T_4033) begin
      way_status_out_43 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_75_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_44 <= 1'h0;
    end else if (_T_4037) begin
      way_status_out_44 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_75_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_45 <= 1'h0;
    end else if (_T_4041) begin
      way_status_out_45 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_75_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_46 <= 1'h0;
    end else if (_T_4045) begin
      way_status_out_46 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_75_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_47 <= 1'h0;
    end else if (_T_4049) begin
      way_status_out_47 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_76_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_48 <= 1'h0;
    end else if (_T_4021) begin
      way_status_out_48 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_76_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_49 <= 1'h0;
    end else if (_T_4025) begin
      way_status_out_49 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_76_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_50 <= 1'h0;
    end else if (_T_4029) begin
      way_status_out_50 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_76_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_51 <= 1'h0;
    end else if (_T_4033) begin
      way_status_out_51 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_76_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_52 <= 1'h0;
    end else if (_T_4037) begin
      way_status_out_52 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_76_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_53 <= 1'h0;
    end else if (_T_4041) begin
      way_status_out_53 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_76_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_54 <= 1'h0;
    end else if (_T_4045) begin
      way_status_out_54 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_76_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_55 <= 1'h0;
    end else if (_T_4049) begin
      way_status_out_55 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_77_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_56 <= 1'h0;
    end else if (_T_4021) begin
      way_status_out_56 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_77_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_57 <= 1'h0;
    end else if (_T_4025) begin
      way_status_out_57 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_77_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_58 <= 1'h0;
    end else if (_T_4029) begin
      way_status_out_58 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_77_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_59 <= 1'h0;
    end else if (_T_4033) begin
      way_status_out_59 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_77_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_60 <= 1'h0;
    end else if (_T_4037) begin
      way_status_out_60 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_77_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_61 <= 1'h0;
    end else if (_T_4041) begin
      way_status_out_61 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_77_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_62 <= 1'h0;
    end else if (_T_4045) begin
      way_status_out_62 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_77_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_63 <= 1'h0;
    end else if (_T_4049) begin
      way_status_out_63 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_78_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_64 <= 1'h0;
    end else if (_T_4021) begin
      way_status_out_64 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_78_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_65 <= 1'h0;
    end else if (_T_4025) begin
      way_status_out_65 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_78_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_66 <= 1'h0;
    end else if (_T_4029) begin
      way_status_out_66 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_78_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_67 <= 1'h0;
    end else if (_T_4033) begin
      way_status_out_67 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_78_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_68 <= 1'h0;
    end else if (_T_4037) begin
      way_status_out_68 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_78_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_69 <= 1'h0;
    end else if (_T_4041) begin
      way_status_out_69 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_78_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_70 <= 1'h0;
    end else if (_T_4045) begin
      way_status_out_70 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_78_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_71 <= 1'h0;
    end else if (_T_4049) begin
      way_status_out_71 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_79_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_72 <= 1'h0;
    end else if (_T_4021) begin
      way_status_out_72 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_79_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_73 <= 1'h0;
    end else if (_T_4025) begin
      way_status_out_73 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_79_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_74 <= 1'h0;
    end else if (_T_4029) begin
      way_status_out_74 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_79_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_75 <= 1'h0;
    end else if (_T_4033) begin
      way_status_out_75 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_79_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_76 <= 1'h0;
    end else if (_T_4037) begin
      way_status_out_76 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_79_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_77 <= 1'h0;
    end else if (_T_4041) begin
      way_status_out_77 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_79_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_78 <= 1'h0;
    end else if (_T_4045) begin
      way_status_out_78 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_79_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_79 <= 1'h0;
    end else if (_T_4049) begin
      way_status_out_79 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_80_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_80 <= 1'h0;
    end else if (_T_4021) begin
      way_status_out_80 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_80_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_81 <= 1'h0;
    end else if (_T_4025) begin
      way_status_out_81 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_80_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_82 <= 1'h0;
    end else if (_T_4029) begin
      way_status_out_82 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_80_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_83 <= 1'h0;
    end else if (_T_4033) begin
      way_status_out_83 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_80_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_84 <= 1'h0;
    end else if (_T_4037) begin
      way_status_out_84 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_80_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_85 <= 1'h0;
    end else if (_T_4041) begin
      way_status_out_85 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_80_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_86 <= 1'h0;
    end else if (_T_4045) begin
      way_status_out_86 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_80_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_87 <= 1'h0;
    end else if (_T_4049) begin
      way_status_out_87 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_81_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_88 <= 1'h0;
    end else if (_T_4021) begin
      way_status_out_88 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_81_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_89 <= 1'h0;
    end else if (_T_4025) begin
      way_status_out_89 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_81_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_90 <= 1'h0;
    end else if (_T_4029) begin
      way_status_out_90 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_81_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_91 <= 1'h0;
    end else if (_T_4033) begin
      way_status_out_91 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_81_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_92 <= 1'h0;
    end else if (_T_4037) begin
      way_status_out_92 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_81_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_93 <= 1'h0;
    end else if (_T_4041) begin
      way_status_out_93 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_81_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_94 <= 1'h0;
    end else if (_T_4045) begin
      way_status_out_94 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_81_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_95 <= 1'h0;
    end else if (_T_4049) begin
      way_status_out_95 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_82_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_96 <= 1'h0;
    end else if (_T_4021) begin
      way_status_out_96 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_82_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_97 <= 1'h0;
    end else if (_T_4025) begin
      way_status_out_97 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_82_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_98 <= 1'h0;
    end else if (_T_4029) begin
      way_status_out_98 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_82_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_99 <= 1'h0;
    end else if (_T_4033) begin
      way_status_out_99 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_82_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_100 <= 1'h0;
    end else if (_T_4037) begin
      way_status_out_100 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_82_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_101 <= 1'h0;
    end else if (_T_4041) begin
      way_status_out_101 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_82_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_102 <= 1'h0;
    end else if (_T_4045) begin
      way_status_out_102 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_82_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_103 <= 1'h0;
    end else if (_T_4049) begin
      way_status_out_103 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_83_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_104 <= 1'h0;
    end else if (_T_4021) begin
      way_status_out_104 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_83_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_105 <= 1'h0;
    end else if (_T_4025) begin
      way_status_out_105 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_83_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_106 <= 1'h0;
    end else if (_T_4029) begin
      way_status_out_106 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_83_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_107 <= 1'h0;
    end else if (_T_4033) begin
      way_status_out_107 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_83_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_108 <= 1'h0;
    end else if (_T_4037) begin
      way_status_out_108 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_83_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_109 <= 1'h0;
    end else if (_T_4041) begin
      way_status_out_109 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_83_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_110 <= 1'h0;
    end else if (_T_4045) begin
      way_status_out_110 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_83_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_111 <= 1'h0;
    end else if (_T_4049) begin
      way_status_out_111 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_84_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_112 <= 1'h0;
    end else if (_T_4021) begin
      way_status_out_112 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_84_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_113 <= 1'h0;
    end else if (_T_4025) begin
      way_status_out_113 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_84_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_114 <= 1'h0;
    end else if (_T_4029) begin
      way_status_out_114 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_84_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_115 <= 1'h0;
    end else if (_T_4033) begin
      way_status_out_115 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_84_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_116 <= 1'h0;
    end else if (_T_4037) begin
      way_status_out_116 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_84_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_117 <= 1'h0;
    end else if (_T_4041) begin
      way_status_out_117 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_84_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_118 <= 1'h0;
    end else if (_T_4045) begin
      way_status_out_118 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_84_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_119 <= 1'h0;
    end else if (_T_4049) begin
      way_status_out_119 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_85_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_120 <= 1'h0;
    end else if (_T_4021) begin
      way_status_out_120 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_85_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_121 <= 1'h0;
    end else if (_T_4025) begin
      way_status_out_121 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_85_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_122 <= 1'h0;
    end else if (_T_4029) begin
      way_status_out_122 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_85_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_123 <= 1'h0;
    end else if (_T_4033) begin
      way_status_out_123 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_85_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_124 <= 1'h0;
    end else if (_T_4037) begin
      way_status_out_124 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_85_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_125 <= 1'h0;
    end else if (_T_4041) begin
      way_status_out_125 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_85_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_126 <= 1'h0;
    end else if (_T_4045) begin
      way_status_out_126 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_85_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_127 <= 1'h0;
    end else if (_T_4049) begin
      way_status_out_127 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_2_io_l1clk or posedge reset) begin
    if (reset) begin
      tagv_mb_scnd_ff <= 2'h0;
    end else if (!(_T_19)) begin
      tagv_mb_scnd_ff <= _T_198;
    end
  end
  always @(posedge rvclkhdr_2_io_l1clk or posedge reset) begin
    if (reset) begin
      uncacheable_miss_scnd_ff <= 1'h0;
    end else if (!(sel_hold_imb_scnd)) begin
      uncacheable_miss_scnd_ff <= io_ifc_fetch_uncacheable_bf;
    end
  end
  always @(posedge rvclkhdr_2_io_l1clk or posedge reset) begin
    if (reset) begin
      imb_scnd_ff <= 31'h0;
    end else if (!(sel_hold_imb_scnd)) begin
      imb_scnd_ff <= io_ifc_fetch_addr_bf;
    end
  end
  always @(posedge rvclkhdr_68_io_l1clk or posedge reset) begin
    if (reset) begin
      ifu_bus_rid_ff <= 3'h0;
    end else begin
      ifu_bus_rid_ff <= io_ifu_axi_r_bits_id;
    end
  end
  always @(posedge rvclkhdr_68_io_l1clk or posedge reset) begin
    if (reset) begin
      ifu_bus_rresp_ff <= 2'h0;
    end else begin
      ifu_bus_rresp_ff <= io_ifu_axi_r_bits_resp;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      ifu_wr_data_comb_err_ff <= 1'h0;
    end else begin
      ifu_wr_data_comb_err_ff <= ifu_wr_cumulative_err_data & _T_2627;
    end
  end
  always @(posedge rvclkhdr_2_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_mb_ff <= 1'h0;
    end else if (_T_278) begin
      way_status_mb_ff <= way_status_mb_scnd_ff;
    end else if (_T_280) begin
      way_status_mb_ff <= replace_way_mb_any_0;
    end else if (!(miss_pending)) begin
      way_status_mb_ff <= way_status;
    end
  end
  always @(posedge rvclkhdr_2_io_l1clk or posedge reset) begin
    if (reset) begin
      tagv_mb_ff <= 2'h0;
    end else if (scnd_miss_req) begin
      tagv_mb_ff <= _T_290;
    end else if (!(miss_pending)) begin
      tagv_mb_ff <= _T_295;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      reset_ic_ff <= 1'h0;
    end else begin
      reset_ic_ff <= _T_298 & _T_299;
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      fetch_uncacheable_ff <= 1'h0;
    end else begin
      fetch_uncacheable_ff <= io_ifc_fetch_uncacheable_bf;
    end
  end
  always @(posedge rvclkhdr_3_io_l1clk or posedge reset) begin
    if (reset) begin
      miss_addr <= 26'h0;
    end else if (_T_231) begin
      miss_addr <= imb_ff[30:5];
    end else if (scnd_miss_req_q) begin
      miss_addr <= imb_scnd_ff[30:5];
    end
  end
  always @(posedge rvclkhdr_2_io_l1clk or posedge reset) begin
    if (reset) begin
      ifc_region_acc_fault_f <= 1'h0;
    end else begin
      ifc_region_acc_fault_f <= io_ifc_region_acc_fault_bf;
    end
  end
  always @(posedge rvclkhdr_3_io_l1clk or posedge reset) begin
    if (reset) begin
      bus_rd_addr_count <= 3'h0;
    end else if (_T_231) begin
      bus_rd_addr_count <= imb_ff[4:2];
    end else if (scnd_miss_req_q) begin
      bus_rd_addr_count <= imb_scnd_ff[4:2];
    end else if (bus_cmd_sent) begin
      bus_rd_addr_count <= _T_2647;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      ic_act_miss_f_delayed <= 1'h0;
    end else begin
      ic_act_miss_f_delayed <= _T_233 & _T_209;
    end
  end
  always @(posedge rvclkhdr_68_io_l1clk or posedge reset) begin
    if (reset) begin
      ifu_bus_rdata_ff <= 64'h0;
    end else begin
      ifu_bus_rdata_ff <= io_ifu_axi_r_bits_data;
    end
  end
  always @(posedge rvclkhdr_4_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_miss_buff_data_0 <= 32'h0;
    end else begin
      ic_miss_buff_data_0 <= io_ifu_axi_r_bits_data[31:0];
    end
  end
  always @(posedge rvclkhdr_4_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_miss_buff_data_1 <= 32'h0;
    end else begin
      ic_miss_buff_data_1 <= io_ifu_axi_r_bits_data[63:32];
    end
  end
  always @(posedge rvclkhdr_13_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_miss_buff_data_2 <= 32'h0;
    end else begin
      ic_miss_buff_data_2 <= io_ifu_axi_r_bits_data[31:0];
    end
  end
  always @(posedge rvclkhdr_13_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_miss_buff_data_3 <= 32'h0;
    end else begin
      ic_miss_buff_data_3 <= io_ifu_axi_r_bits_data[63:32];
    end
  end
  always @(posedge rvclkhdr_22_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_miss_buff_data_4 <= 32'h0;
    end else begin
      ic_miss_buff_data_4 <= io_ifu_axi_r_bits_data[31:0];
    end
  end
  always @(posedge rvclkhdr_22_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_miss_buff_data_5 <= 32'h0;
    end else begin
      ic_miss_buff_data_5 <= io_ifu_axi_r_bits_data[63:32];
    end
  end
  always @(posedge rvclkhdr_31_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_miss_buff_data_6 <= 32'h0;
    end else begin
      ic_miss_buff_data_6 <= io_ifu_axi_r_bits_data[31:0];
    end
  end
  always @(posedge rvclkhdr_31_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_miss_buff_data_7 <= 32'h0;
    end else begin
      ic_miss_buff_data_7 <= io_ifu_axi_r_bits_data[63:32];
    end
  end
  always @(posedge rvclkhdr_40_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_miss_buff_data_8 <= 32'h0;
    end else begin
      ic_miss_buff_data_8 <= io_ifu_axi_r_bits_data[31:0];
    end
  end
  always @(posedge rvclkhdr_40_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_miss_buff_data_9 <= 32'h0;
    end else begin
      ic_miss_buff_data_9 <= io_ifu_axi_r_bits_data[63:32];
    end
  end
  always @(posedge rvclkhdr_49_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_miss_buff_data_10 <= 32'h0;
    end else begin
      ic_miss_buff_data_10 <= io_ifu_axi_r_bits_data[31:0];
    end
  end
  always @(posedge rvclkhdr_49_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_miss_buff_data_11 <= 32'h0;
    end else begin
      ic_miss_buff_data_11 <= io_ifu_axi_r_bits_data[63:32];
    end
  end
  always @(posedge rvclkhdr_58_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_miss_buff_data_12 <= 32'h0;
    end else begin
      ic_miss_buff_data_12 <= io_ifu_axi_r_bits_data[31:0];
    end
  end
  always @(posedge rvclkhdr_58_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_miss_buff_data_13 <= 32'h0;
    end else begin
      ic_miss_buff_data_13 <= io_ifu_axi_r_bits_data[63:32];
    end
  end
  always @(posedge rvclkhdr_67_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_miss_buff_data_14 <= 32'h0;
    end else begin
      ic_miss_buff_data_14 <= io_ifu_axi_r_bits_data[31:0];
    end
  end
  always @(posedge rvclkhdr_67_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_miss_buff_data_15 <= 32'h0;
    end else begin
      ic_miss_buff_data_15 <= io_ifu_axi_r_bits_data[63:32];
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      ic_crit_wd_rdy_new_ff <= 1'h0;
    end else begin
      ic_crit_wd_rdy_new_ff <= _T_1514 | _T_1519;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      ic_miss_buff_data_error <= 8'h0;
    end else begin
      ic_miss_buff_data_error <= {_T_1398,ic_miss_buff_data_error_in_0};
    end
  end
  always @(posedge rvclkhdr_1_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_debug_ict_array_sel_ff <= 1'h0;
    end else begin
      ic_debug_ict_array_sel_ff <= io_ic_debug_rd_en & io_ic_debug_tag_array;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_0 <= 1'h0;
    end else if (_T_5642) begin
      ic_tag_valid_out_1_0 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_1 <= 1'h0;
    end else if (_T_5657) begin
      ic_tag_valid_out_1_1 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_2 <= 1'h0;
    end else if (_T_5672) begin
      ic_tag_valid_out_1_2 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_3 <= 1'h0;
    end else if (_T_5687) begin
      ic_tag_valid_out_1_3 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_4 <= 1'h0;
    end else if (_T_5702) begin
      ic_tag_valid_out_1_4 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_5 <= 1'h0;
    end else if (_T_5717) begin
      ic_tag_valid_out_1_5 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_6 <= 1'h0;
    end else if (_T_5732) begin
      ic_tag_valid_out_1_6 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_7 <= 1'h0;
    end else if (_T_5747) begin
      ic_tag_valid_out_1_7 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_8 <= 1'h0;
    end else if (_T_5762) begin
      ic_tag_valid_out_1_8 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_9 <= 1'h0;
    end else if (_T_5777) begin
      ic_tag_valid_out_1_9 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_10 <= 1'h0;
    end else if (_T_5792) begin
      ic_tag_valid_out_1_10 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_11 <= 1'h0;
    end else if (_T_5807) begin
      ic_tag_valid_out_1_11 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_12 <= 1'h0;
    end else if (_T_5822) begin
      ic_tag_valid_out_1_12 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_13 <= 1'h0;
    end else if (_T_5837) begin
      ic_tag_valid_out_1_13 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_14 <= 1'h0;
    end else if (_T_5852) begin
      ic_tag_valid_out_1_14 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_15 <= 1'h0;
    end else if (_T_5867) begin
      ic_tag_valid_out_1_15 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_16 <= 1'h0;
    end else if (_T_5882) begin
      ic_tag_valid_out_1_16 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_17 <= 1'h0;
    end else if (_T_5897) begin
      ic_tag_valid_out_1_17 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_18 <= 1'h0;
    end else if (_T_5912) begin
      ic_tag_valid_out_1_18 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_19 <= 1'h0;
    end else if (_T_5927) begin
      ic_tag_valid_out_1_19 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_20 <= 1'h0;
    end else if (_T_5942) begin
      ic_tag_valid_out_1_20 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_21 <= 1'h0;
    end else if (_T_5957) begin
      ic_tag_valid_out_1_21 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_22 <= 1'h0;
    end else if (_T_5972) begin
      ic_tag_valid_out_1_22 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_23 <= 1'h0;
    end else if (_T_5987) begin
      ic_tag_valid_out_1_23 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_24 <= 1'h0;
    end else if (_T_6002) begin
      ic_tag_valid_out_1_24 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_25 <= 1'h0;
    end else if (_T_6017) begin
      ic_tag_valid_out_1_25 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_26 <= 1'h0;
    end else if (_T_6032) begin
      ic_tag_valid_out_1_26 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_27 <= 1'h0;
    end else if (_T_6047) begin
      ic_tag_valid_out_1_27 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_28 <= 1'h0;
    end else if (_T_6062) begin
      ic_tag_valid_out_1_28 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_29 <= 1'h0;
    end else if (_T_6077) begin
      ic_tag_valid_out_1_29 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_30 <= 1'h0;
    end else if (_T_6092) begin
      ic_tag_valid_out_1_30 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_31 <= 1'h0;
    end else if (_T_6107) begin
      ic_tag_valid_out_1_31 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_32 <= 1'h0;
    end else if (_T_6602) begin
      ic_tag_valid_out_1_32 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_33 <= 1'h0;
    end else if (_T_6617) begin
      ic_tag_valid_out_1_33 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_34 <= 1'h0;
    end else if (_T_6632) begin
      ic_tag_valid_out_1_34 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_35 <= 1'h0;
    end else if (_T_6647) begin
      ic_tag_valid_out_1_35 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_36 <= 1'h0;
    end else if (_T_6662) begin
      ic_tag_valid_out_1_36 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_37 <= 1'h0;
    end else if (_T_6677) begin
      ic_tag_valid_out_1_37 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_38 <= 1'h0;
    end else if (_T_6692) begin
      ic_tag_valid_out_1_38 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_39 <= 1'h0;
    end else if (_T_6707) begin
      ic_tag_valid_out_1_39 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_40 <= 1'h0;
    end else if (_T_6722) begin
      ic_tag_valid_out_1_40 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_41 <= 1'h0;
    end else if (_T_6737) begin
      ic_tag_valid_out_1_41 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_42 <= 1'h0;
    end else if (_T_6752) begin
      ic_tag_valid_out_1_42 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_43 <= 1'h0;
    end else if (_T_6767) begin
      ic_tag_valid_out_1_43 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_44 <= 1'h0;
    end else if (_T_6782) begin
      ic_tag_valid_out_1_44 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_45 <= 1'h0;
    end else if (_T_6797) begin
      ic_tag_valid_out_1_45 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_46 <= 1'h0;
    end else if (_T_6812) begin
      ic_tag_valid_out_1_46 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_47 <= 1'h0;
    end else if (_T_6827) begin
      ic_tag_valid_out_1_47 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_48 <= 1'h0;
    end else if (_T_6842) begin
      ic_tag_valid_out_1_48 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_49 <= 1'h0;
    end else if (_T_6857) begin
      ic_tag_valid_out_1_49 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_50 <= 1'h0;
    end else if (_T_6872) begin
      ic_tag_valid_out_1_50 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_51 <= 1'h0;
    end else if (_T_6887) begin
      ic_tag_valid_out_1_51 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_52 <= 1'h0;
    end else if (_T_6902) begin
      ic_tag_valid_out_1_52 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_53 <= 1'h0;
    end else if (_T_6917) begin
      ic_tag_valid_out_1_53 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_54 <= 1'h0;
    end else if (_T_6932) begin
      ic_tag_valid_out_1_54 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_55 <= 1'h0;
    end else if (_T_6947) begin
      ic_tag_valid_out_1_55 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_56 <= 1'h0;
    end else if (_T_6962) begin
      ic_tag_valid_out_1_56 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_57 <= 1'h0;
    end else if (_T_6977) begin
      ic_tag_valid_out_1_57 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_58 <= 1'h0;
    end else if (_T_6992) begin
      ic_tag_valid_out_1_58 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_59 <= 1'h0;
    end else if (_T_7007) begin
      ic_tag_valid_out_1_59 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_60 <= 1'h0;
    end else if (_T_7022) begin
      ic_tag_valid_out_1_60 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_61 <= 1'h0;
    end else if (_T_7037) begin
      ic_tag_valid_out_1_61 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_62 <= 1'h0;
    end else if (_T_7052) begin
      ic_tag_valid_out_1_62 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_63 <= 1'h0;
    end else if (_T_7067) begin
      ic_tag_valid_out_1_63 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_64 <= 1'h0;
    end else if (_T_7562) begin
      ic_tag_valid_out_1_64 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_65 <= 1'h0;
    end else if (_T_7577) begin
      ic_tag_valid_out_1_65 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_66 <= 1'h0;
    end else if (_T_7592) begin
      ic_tag_valid_out_1_66 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_67 <= 1'h0;
    end else if (_T_7607) begin
      ic_tag_valid_out_1_67 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_68 <= 1'h0;
    end else if (_T_7622) begin
      ic_tag_valid_out_1_68 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_69 <= 1'h0;
    end else if (_T_7637) begin
      ic_tag_valid_out_1_69 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_70 <= 1'h0;
    end else if (_T_7652) begin
      ic_tag_valid_out_1_70 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_71 <= 1'h0;
    end else if (_T_7667) begin
      ic_tag_valid_out_1_71 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_72 <= 1'h0;
    end else if (_T_7682) begin
      ic_tag_valid_out_1_72 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_73 <= 1'h0;
    end else if (_T_7697) begin
      ic_tag_valid_out_1_73 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_74 <= 1'h0;
    end else if (_T_7712) begin
      ic_tag_valid_out_1_74 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_75 <= 1'h0;
    end else if (_T_7727) begin
      ic_tag_valid_out_1_75 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_76 <= 1'h0;
    end else if (_T_7742) begin
      ic_tag_valid_out_1_76 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_77 <= 1'h0;
    end else if (_T_7757) begin
      ic_tag_valid_out_1_77 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_78 <= 1'h0;
    end else if (_T_7772) begin
      ic_tag_valid_out_1_78 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_79 <= 1'h0;
    end else if (_T_7787) begin
      ic_tag_valid_out_1_79 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_80 <= 1'h0;
    end else if (_T_7802) begin
      ic_tag_valid_out_1_80 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_81 <= 1'h0;
    end else if (_T_7817) begin
      ic_tag_valid_out_1_81 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_82 <= 1'h0;
    end else if (_T_7832) begin
      ic_tag_valid_out_1_82 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_83 <= 1'h0;
    end else if (_T_7847) begin
      ic_tag_valid_out_1_83 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_84 <= 1'h0;
    end else if (_T_7862) begin
      ic_tag_valid_out_1_84 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_85 <= 1'h0;
    end else if (_T_7877) begin
      ic_tag_valid_out_1_85 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_86 <= 1'h0;
    end else if (_T_7892) begin
      ic_tag_valid_out_1_86 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_87 <= 1'h0;
    end else if (_T_7907) begin
      ic_tag_valid_out_1_87 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_88 <= 1'h0;
    end else if (_T_7922) begin
      ic_tag_valid_out_1_88 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_89 <= 1'h0;
    end else if (_T_7937) begin
      ic_tag_valid_out_1_89 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_90 <= 1'h0;
    end else if (_T_7952) begin
      ic_tag_valid_out_1_90 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_91 <= 1'h0;
    end else if (_T_7967) begin
      ic_tag_valid_out_1_91 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_92 <= 1'h0;
    end else if (_T_7982) begin
      ic_tag_valid_out_1_92 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_93 <= 1'h0;
    end else if (_T_7997) begin
      ic_tag_valid_out_1_93 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_94 <= 1'h0;
    end else if (_T_8012) begin
      ic_tag_valid_out_1_94 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_95 <= 1'h0;
    end else if (_T_8027) begin
      ic_tag_valid_out_1_95 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_96 <= 1'h0;
    end else if (_T_8522) begin
      ic_tag_valid_out_1_96 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_97 <= 1'h0;
    end else if (_T_8537) begin
      ic_tag_valid_out_1_97 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_98 <= 1'h0;
    end else if (_T_8552) begin
      ic_tag_valid_out_1_98 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_99 <= 1'h0;
    end else if (_T_8567) begin
      ic_tag_valid_out_1_99 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_100 <= 1'h0;
    end else if (_T_8582) begin
      ic_tag_valid_out_1_100 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_101 <= 1'h0;
    end else if (_T_8597) begin
      ic_tag_valid_out_1_101 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_102 <= 1'h0;
    end else if (_T_8612) begin
      ic_tag_valid_out_1_102 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_103 <= 1'h0;
    end else if (_T_8627) begin
      ic_tag_valid_out_1_103 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_104 <= 1'h0;
    end else if (_T_8642) begin
      ic_tag_valid_out_1_104 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_105 <= 1'h0;
    end else if (_T_8657) begin
      ic_tag_valid_out_1_105 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_106 <= 1'h0;
    end else if (_T_8672) begin
      ic_tag_valid_out_1_106 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_107 <= 1'h0;
    end else if (_T_8687) begin
      ic_tag_valid_out_1_107 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_108 <= 1'h0;
    end else if (_T_8702) begin
      ic_tag_valid_out_1_108 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_109 <= 1'h0;
    end else if (_T_8717) begin
      ic_tag_valid_out_1_109 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_110 <= 1'h0;
    end else if (_T_8732) begin
      ic_tag_valid_out_1_110 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_111 <= 1'h0;
    end else if (_T_8747) begin
      ic_tag_valid_out_1_111 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_112 <= 1'h0;
    end else if (_T_8762) begin
      ic_tag_valid_out_1_112 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_113 <= 1'h0;
    end else if (_T_8777) begin
      ic_tag_valid_out_1_113 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_114 <= 1'h0;
    end else if (_T_8792) begin
      ic_tag_valid_out_1_114 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_115 <= 1'h0;
    end else if (_T_8807) begin
      ic_tag_valid_out_1_115 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_116 <= 1'h0;
    end else if (_T_8822) begin
      ic_tag_valid_out_1_116 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_117 <= 1'h0;
    end else if (_T_8837) begin
      ic_tag_valid_out_1_117 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_118 <= 1'h0;
    end else if (_T_8852) begin
      ic_tag_valid_out_1_118 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_119 <= 1'h0;
    end else if (_T_8867) begin
      ic_tag_valid_out_1_119 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_120 <= 1'h0;
    end else if (_T_8882) begin
      ic_tag_valid_out_1_120 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_121 <= 1'h0;
    end else if (_T_8897) begin
      ic_tag_valid_out_1_121 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_122 <= 1'h0;
    end else if (_T_8912) begin
      ic_tag_valid_out_1_122 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_123 <= 1'h0;
    end else if (_T_8927) begin
      ic_tag_valid_out_1_123 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_124 <= 1'h0;
    end else if (_T_8942) begin
      ic_tag_valid_out_1_124 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_125 <= 1'h0;
    end else if (_T_8957) begin
      ic_tag_valid_out_1_125 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_126 <= 1'h0;
    end else if (_T_8972) begin
      ic_tag_valid_out_1_126 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_127 <= 1'h0;
    end else if (_T_8987) begin
      ic_tag_valid_out_1_127 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_0 <= 1'h0;
    end else if (_T_5162) begin
      ic_tag_valid_out_0_0 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_1 <= 1'h0;
    end else if (_T_5177) begin
      ic_tag_valid_out_0_1 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_2 <= 1'h0;
    end else if (_T_5192) begin
      ic_tag_valid_out_0_2 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_3 <= 1'h0;
    end else if (_T_5207) begin
      ic_tag_valid_out_0_3 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_4 <= 1'h0;
    end else if (_T_5222) begin
      ic_tag_valid_out_0_4 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_5 <= 1'h0;
    end else if (_T_5237) begin
      ic_tag_valid_out_0_5 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_6 <= 1'h0;
    end else if (_T_5252) begin
      ic_tag_valid_out_0_6 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_7 <= 1'h0;
    end else if (_T_5267) begin
      ic_tag_valid_out_0_7 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_8 <= 1'h0;
    end else if (_T_5282) begin
      ic_tag_valid_out_0_8 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_9 <= 1'h0;
    end else if (_T_5297) begin
      ic_tag_valid_out_0_9 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_10 <= 1'h0;
    end else if (_T_5312) begin
      ic_tag_valid_out_0_10 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_11 <= 1'h0;
    end else if (_T_5327) begin
      ic_tag_valid_out_0_11 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_12 <= 1'h0;
    end else if (_T_5342) begin
      ic_tag_valid_out_0_12 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_13 <= 1'h0;
    end else if (_T_5357) begin
      ic_tag_valid_out_0_13 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_14 <= 1'h0;
    end else if (_T_5372) begin
      ic_tag_valid_out_0_14 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_15 <= 1'h0;
    end else if (_T_5387) begin
      ic_tag_valid_out_0_15 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_16 <= 1'h0;
    end else if (_T_5402) begin
      ic_tag_valid_out_0_16 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_17 <= 1'h0;
    end else if (_T_5417) begin
      ic_tag_valid_out_0_17 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_18 <= 1'h0;
    end else if (_T_5432) begin
      ic_tag_valid_out_0_18 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_19 <= 1'h0;
    end else if (_T_5447) begin
      ic_tag_valid_out_0_19 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_20 <= 1'h0;
    end else if (_T_5462) begin
      ic_tag_valid_out_0_20 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_21 <= 1'h0;
    end else if (_T_5477) begin
      ic_tag_valid_out_0_21 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_22 <= 1'h0;
    end else if (_T_5492) begin
      ic_tag_valid_out_0_22 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_23 <= 1'h0;
    end else if (_T_5507) begin
      ic_tag_valid_out_0_23 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_24 <= 1'h0;
    end else if (_T_5522) begin
      ic_tag_valid_out_0_24 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_25 <= 1'h0;
    end else if (_T_5537) begin
      ic_tag_valid_out_0_25 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_26 <= 1'h0;
    end else if (_T_5552) begin
      ic_tag_valid_out_0_26 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_27 <= 1'h0;
    end else if (_T_5567) begin
      ic_tag_valid_out_0_27 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_28 <= 1'h0;
    end else if (_T_5582) begin
      ic_tag_valid_out_0_28 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_29 <= 1'h0;
    end else if (_T_5597) begin
      ic_tag_valid_out_0_29 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_30 <= 1'h0;
    end else if (_T_5612) begin
      ic_tag_valid_out_0_30 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_31 <= 1'h0;
    end else if (_T_5627) begin
      ic_tag_valid_out_0_31 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_32 <= 1'h0;
    end else if (_T_6122) begin
      ic_tag_valid_out_0_32 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_33 <= 1'h0;
    end else if (_T_6137) begin
      ic_tag_valid_out_0_33 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_34 <= 1'h0;
    end else if (_T_6152) begin
      ic_tag_valid_out_0_34 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_35 <= 1'h0;
    end else if (_T_6167) begin
      ic_tag_valid_out_0_35 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_36 <= 1'h0;
    end else if (_T_6182) begin
      ic_tag_valid_out_0_36 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_37 <= 1'h0;
    end else if (_T_6197) begin
      ic_tag_valid_out_0_37 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_38 <= 1'h0;
    end else if (_T_6212) begin
      ic_tag_valid_out_0_38 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_39 <= 1'h0;
    end else if (_T_6227) begin
      ic_tag_valid_out_0_39 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_40 <= 1'h0;
    end else if (_T_6242) begin
      ic_tag_valid_out_0_40 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_41 <= 1'h0;
    end else if (_T_6257) begin
      ic_tag_valid_out_0_41 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_42 <= 1'h0;
    end else if (_T_6272) begin
      ic_tag_valid_out_0_42 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_43 <= 1'h0;
    end else if (_T_6287) begin
      ic_tag_valid_out_0_43 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_44 <= 1'h0;
    end else if (_T_6302) begin
      ic_tag_valid_out_0_44 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_45 <= 1'h0;
    end else if (_T_6317) begin
      ic_tag_valid_out_0_45 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_46 <= 1'h0;
    end else if (_T_6332) begin
      ic_tag_valid_out_0_46 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_47 <= 1'h0;
    end else if (_T_6347) begin
      ic_tag_valid_out_0_47 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_48 <= 1'h0;
    end else if (_T_6362) begin
      ic_tag_valid_out_0_48 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_49 <= 1'h0;
    end else if (_T_6377) begin
      ic_tag_valid_out_0_49 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_50 <= 1'h0;
    end else if (_T_6392) begin
      ic_tag_valid_out_0_50 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_51 <= 1'h0;
    end else if (_T_6407) begin
      ic_tag_valid_out_0_51 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_52 <= 1'h0;
    end else if (_T_6422) begin
      ic_tag_valid_out_0_52 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_53 <= 1'h0;
    end else if (_T_6437) begin
      ic_tag_valid_out_0_53 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_54 <= 1'h0;
    end else if (_T_6452) begin
      ic_tag_valid_out_0_54 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_55 <= 1'h0;
    end else if (_T_6467) begin
      ic_tag_valid_out_0_55 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_56 <= 1'h0;
    end else if (_T_6482) begin
      ic_tag_valid_out_0_56 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_57 <= 1'h0;
    end else if (_T_6497) begin
      ic_tag_valid_out_0_57 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_58 <= 1'h0;
    end else if (_T_6512) begin
      ic_tag_valid_out_0_58 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_59 <= 1'h0;
    end else if (_T_6527) begin
      ic_tag_valid_out_0_59 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_60 <= 1'h0;
    end else if (_T_6542) begin
      ic_tag_valid_out_0_60 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_61 <= 1'h0;
    end else if (_T_6557) begin
      ic_tag_valid_out_0_61 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_62 <= 1'h0;
    end else if (_T_6572) begin
      ic_tag_valid_out_0_62 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_63 <= 1'h0;
    end else if (_T_6587) begin
      ic_tag_valid_out_0_63 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_64 <= 1'h0;
    end else if (_T_7082) begin
      ic_tag_valid_out_0_64 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_65 <= 1'h0;
    end else if (_T_7097) begin
      ic_tag_valid_out_0_65 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_66 <= 1'h0;
    end else if (_T_7112) begin
      ic_tag_valid_out_0_66 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_67 <= 1'h0;
    end else if (_T_7127) begin
      ic_tag_valid_out_0_67 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_68 <= 1'h0;
    end else if (_T_7142) begin
      ic_tag_valid_out_0_68 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_69 <= 1'h0;
    end else if (_T_7157) begin
      ic_tag_valid_out_0_69 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_70 <= 1'h0;
    end else if (_T_7172) begin
      ic_tag_valid_out_0_70 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_71 <= 1'h0;
    end else if (_T_7187) begin
      ic_tag_valid_out_0_71 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_72 <= 1'h0;
    end else if (_T_7202) begin
      ic_tag_valid_out_0_72 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_73 <= 1'h0;
    end else if (_T_7217) begin
      ic_tag_valid_out_0_73 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_74 <= 1'h0;
    end else if (_T_7232) begin
      ic_tag_valid_out_0_74 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_75 <= 1'h0;
    end else if (_T_7247) begin
      ic_tag_valid_out_0_75 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_76 <= 1'h0;
    end else if (_T_7262) begin
      ic_tag_valid_out_0_76 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_77 <= 1'h0;
    end else if (_T_7277) begin
      ic_tag_valid_out_0_77 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_78 <= 1'h0;
    end else if (_T_7292) begin
      ic_tag_valid_out_0_78 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_79 <= 1'h0;
    end else if (_T_7307) begin
      ic_tag_valid_out_0_79 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_80 <= 1'h0;
    end else if (_T_7322) begin
      ic_tag_valid_out_0_80 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_81 <= 1'h0;
    end else if (_T_7337) begin
      ic_tag_valid_out_0_81 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_82 <= 1'h0;
    end else if (_T_7352) begin
      ic_tag_valid_out_0_82 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_83 <= 1'h0;
    end else if (_T_7367) begin
      ic_tag_valid_out_0_83 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_84 <= 1'h0;
    end else if (_T_7382) begin
      ic_tag_valid_out_0_84 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_85 <= 1'h0;
    end else if (_T_7397) begin
      ic_tag_valid_out_0_85 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_86 <= 1'h0;
    end else if (_T_7412) begin
      ic_tag_valid_out_0_86 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_87 <= 1'h0;
    end else if (_T_7427) begin
      ic_tag_valid_out_0_87 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_88 <= 1'h0;
    end else if (_T_7442) begin
      ic_tag_valid_out_0_88 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_89 <= 1'h0;
    end else if (_T_7457) begin
      ic_tag_valid_out_0_89 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_90 <= 1'h0;
    end else if (_T_7472) begin
      ic_tag_valid_out_0_90 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_91 <= 1'h0;
    end else if (_T_7487) begin
      ic_tag_valid_out_0_91 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_92 <= 1'h0;
    end else if (_T_7502) begin
      ic_tag_valid_out_0_92 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_93 <= 1'h0;
    end else if (_T_7517) begin
      ic_tag_valid_out_0_93 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_94 <= 1'h0;
    end else if (_T_7532) begin
      ic_tag_valid_out_0_94 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_95 <= 1'h0;
    end else if (_T_7547) begin
      ic_tag_valid_out_0_95 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_96 <= 1'h0;
    end else if (_T_8042) begin
      ic_tag_valid_out_0_96 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_97 <= 1'h0;
    end else if (_T_8057) begin
      ic_tag_valid_out_0_97 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_98 <= 1'h0;
    end else if (_T_8072) begin
      ic_tag_valid_out_0_98 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_99 <= 1'h0;
    end else if (_T_8087) begin
      ic_tag_valid_out_0_99 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_100 <= 1'h0;
    end else if (_T_8102) begin
      ic_tag_valid_out_0_100 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_101 <= 1'h0;
    end else if (_T_8117) begin
      ic_tag_valid_out_0_101 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_102 <= 1'h0;
    end else if (_T_8132) begin
      ic_tag_valid_out_0_102 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_103 <= 1'h0;
    end else if (_T_8147) begin
      ic_tag_valid_out_0_103 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_104 <= 1'h0;
    end else if (_T_8162) begin
      ic_tag_valid_out_0_104 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_105 <= 1'h0;
    end else if (_T_8177) begin
      ic_tag_valid_out_0_105 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_106 <= 1'h0;
    end else if (_T_8192) begin
      ic_tag_valid_out_0_106 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_107 <= 1'h0;
    end else if (_T_8207) begin
      ic_tag_valid_out_0_107 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_108 <= 1'h0;
    end else if (_T_8222) begin
      ic_tag_valid_out_0_108 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_109 <= 1'h0;
    end else if (_T_8237) begin
      ic_tag_valid_out_0_109 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_110 <= 1'h0;
    end else if (_T_8252) begin
      ic_tag_valid_out_0_110 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_111 <= 1'h0;
    end else if (_T_8267) begin
      ic_tag_valid_out_0_111 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_112 <= 1'h0;
    end else if (_T_8282) begin
      ic_tag_valid_out_0_112 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_113 <= 1'h0;
    end else if (_T_8297) begin
      ic_tag_valid_out_0_113 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_114 <= 1'h0;
    end else if (_T_8312) begin
      ic_tag_valid_out_0_114 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_115 <= 1'h0;
    end else if (_T_8327) begin
      ic_tag_valid_out_0_115 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_116 <= 1'h0;
    end else if (_T_8342) begin
      ic_tag_valid_out_0_116 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_117 <= 1'h0;
    end else if (_T_8357) begin
      ic_tag_valid_out_0_117 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_118 <= 1'h0;
    end else if (_T_8372) begin
      ic_tag_valid_out_0_118 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_119 <= 1'h0;
    end else if (_T_8387) begin
      ic_tag_valid_out_0_119 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_120 <= 1'h0;
    end else if (_T_8402) begin
      ic_tag_valid_out_0_120 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_121 <= 1'h0;
    end else if (_T_8417) begin
      ic_tag_valid_out_0_121 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_122 <= 1'h0;
    end else if (_T_8432) begin
      ic_tag_valid_out_0_122 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_123 <= 1'h0;
    end else if (_T_8447) begin
      ic_tag_valid_out_0_123 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_124 <= 1'h0;
    end else if (_T_8462) begin
      ic_tag_valid_out_0_124 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_125 <= 1'h0;
    end else if (_T_8477) begin
      ic_tag_valid_out_0_125 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_126 <= 1'h0;
    end else if (_T_8492) begin
      ic_tag_valid_out_0_126 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_127 <= 1'h0;
    end else if (_T_8507) begin
      ic_tag_valid_out_0_127 <= _T_5154;
    end
  end
  always @(posedge rvclkhdr_1_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_debug_way_ff <= 2'h0;
    end else begin
      ic_debug_way_ff <= io_ic_debug_way;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      ic_debug_rd_en_ff <= 1'h0;
    end else begin
      ic_debug_rd_en_ff <= io_ic_debug_rd_en;
    end
  end
  always @(posedge rvclkhdr_io_l1clk or posedge reset) begin
    if (reset) begin
      _T_1212 <= 71'h0;
    end else if (ic_debug_ict_array_sel_ff) begin
      _T_1212 <= _T_1211;
    end else begin
      _T_1212 <= io_ic_debug_rd_data;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      ifc_region_acc_fault_memory_f <= 1'h0;
    end else begin
      ifc_region_acc_fault_memory_f <= _T_9885 & io_ifc_fetch_req_bf;
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      perr_ic_index_ff <= 7'h0;
    end else if (perr_sb_write_status) begin
      perr_ic_index_ff <= ifu_ic_rw_int_addr_ff;
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      dma_sb_err_state_ff <= 1'h0;
    end else begin
      dma_sb_err_state_ff <= perr_state == 3'h4;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      bus_cmd_req_hold <= 1'h0;
    end else begin
      bus_cmd_req_hold <= _T_2604 & _T_2623;
    end
  end
  always @(posedge rvclkhdr_69_io_l1clk or posedge reset) begin
    if (reset) begin
      ifu_bus_cmd_valid <= 1'h0;
    end else begin
      ifu_bus_cmd_valid <= _T_2594 & _T_2600;
    end
  end
  always @(posedge rvclkhdr_3_io_l1clk or posedge reset) begin
    if (reset) begin
      bus_cmd_beat_count <= 3'h0;
    end else if (bus_cmd_beat_en) begin
      bus_cmd_beat_count <= bus_new_cmd_beat_count;
    end
  end
  always @(posedge rvclkhdr_68_io_l1clk or posedge reset) begin
    if (reset) begin
      ifu_bus_arready_unq_ff <= 1'h0;
    end else begin
      ifu_bus_arready_unq_ff <= io_ifu_axi_ar_ready;
    end
  end
  always @(posedge rvclkhdr_68_io_l1clk or posedge reset) begin
    if (reset) begin
      ifu_bus_arvalid_ff <= 1'h0;
    end else begin
      ifu_bus_arvalid_ff <= io_ifu_axi_ar_valid;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      ifc_dma_access_ok_prev <= 1'h0;
    end else begin
      ifc_dma_access_ok_prev <= _T_2699 & _T_2700;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      iccm_ecc_corr_data_ff <= 39'h0;
    end else if (iccm_ecc_write_status) begin
      iccm_ecc_corr_data_ff <= _T_3932;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      dma_mem_addr_ff <= 2'h0;
    end else begin
      dma_mem_addr_ff <= io_dma_mem_ctl_dma_mem_addr[3:2];
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      dma_mem_tag_ff <= 3'h0;
    end else begin
      dma_mem_tag_ff <= io_dma_mem_ctl_dma_mem_tag;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      iccm_dma_rtag_temp <= 3'h0;
    end else begin
      iccm_dma_rtag_temp <= dma_mem_tag_ff;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      iccm_dma_rvalid_temp <= 1'h0;
    end else begin
      iccm_dma_rvalid_temp <= iccm_dma_rvalid_in;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      iccm_dma_ecc_error <= 1'h0;
    end else begin
      iccm_dma_ecc_error <= |iccm_double_ecc_error;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      iccm_dma_rdata_temp <= 64'h0;
    end else if (iccm_dma_ecc_error_in) begin
      iccm_dma_rdata_temp <= _T_3104;
    end else begin
      iccm_dma_rdata_temp <= _T_3105;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      iccm_ecc_corr_index_ff <= 14'h0;
    end else if (iccm_ecc_write_status) begin
      if (iccm_single_ecc_error[0]) begin
        iccm_ecc_corr_index_ff <= iccm_rw_addr_f;
      end else begin
        iccm_ecc_corr_index_ff <= _T_3928;
      end
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      iccm_rd_ecc_single_err_ff <= 1'h0;
    end else begin
      iccm_rd_ecc_single_err_ff <= _T_3923 & _T_319;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      iccm_rw_addr_f <= 14'h0;
    end else begin
      iccm_rw_addr_f <= io_iccm_rw_addr[14:1];
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      ifu_status_wr_addr_ff <= 7'h0;
    end else if (_T_3997) begin
      ifu_status_wr_addr_ff <= io_ic_debug_addr[9:3];
    end else begin
      ifu_status_wr_addr_ff <= ifu_status_wr_addr[11:5];
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      way_status_wr_en_ff <= 1'h0;
    end else begin
      way_status_wr_en_ff <= way_status_wr_en | _T_4000;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      way_status_new_ff <= 1'h0;
    end else if (_T_4000) begin
      way_status_new_ff <= io_ic_debug_wr_data[4];
    end else if (_T_9777) begin
      way_status_new_ff <= replace_way_mb_any_0;
    end else begin
      way_status_new_ff <= way_status_hit_new;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      ifu_tag_wren_ff <= 2'h0;
    end else begin
      ifu_tag_wren_ff <= ifu_tag_wren | ic_debug_tag_wr_en;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      ic_valid_ff <= 1'h0;
    end else if (_T_4000) begin
      ic_valid_ff <= io_ic_debug_wr_data[0];
    end else begin
      ic_valid_ff <= ic_valid;
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      _T_9799 <= 1'h0;
    end else begin
      _T_9799 <= _T_233 & _T_209;
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      _T_9800 <= 1'h0;
    end else begin
      _T_9800 <= _T_225 & _T_247;
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      _T_9801 <= 1'h0;
    end else begin
      _T_9801 <= ic_byp_hit_f & ifu_byp_data_err_new;
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      _T_9805 <= 1'h0;
    end else begin
      _T_9805 <= _T_9803 & miss_pending;
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      _T_9806 <= 1'h0;
    end else begin
      _T_9806 <= _T_2618 & _T_2623;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      _T_9826 <= 1'h0;
    end else begin
      _T_9826 <= ic_debug_rd_en_ff;
    end
  end
endmodule
module ifu_bp_ctl(
  input         clock,
  input         reset,
  input         io_active_clk,
  input         io_ic_hit_f,
  input         io_exu_flush_final,
  input  [30:0] io_ifc_fetch_addr_f,
  input         io_ifc_fetch_req_f,
  input         io_dec_bp_dec_tlu_br0_r_pkt_valid,
  input  [1:0]  io_dec_bp_dec_tlu_br0_r_pkt_bits_hist,
  input         io_dec_bp_dec_tlu_br0_r_pkt_bits_br_error,
  input         io_dec_bp_dec_tlu_br0_r_pkt_bits_br_start_error,
  input         io_dec_bp_dec_tlu_br0_r_pkt_bits_way,
  input         io_dec_bp_dec_tlu_br0_r_pkt_bits_middle,
  input         io_dec_bp_dec_tlu_flush_leak_one_wb,
  input         io_dec_bp_dec_tlu_bpred_disable,
  input         io_dec_tlu_flush_lower_wb,
  input  [7:0]  io_exu_bp_exu_i0_br_index_r,
  input  [7:0]  io_exu_bp_exu_i0_br_fghr_r,
  input         io_exu_bp_exu_mp_pkt_bits_misp,
  input         io_exu_bp_exu_mp_pkt_bits_ataken,
  input         io_exu_bp_exu_mp_pkt_bits_boffset,
  input         io_exu_bp_exu_mp_pkt_bits_pc4,
  input  [1:0]  io_exu_bp_exu_mp_pkt_bits_hist,
  input  [11:0] io_exu_bp_exu_mp_pkt_bits_toffset,
  input         io_exu_bp_exu_mp_pkt_bits_pcall,
  input         io_exu_bp_exu_mp_pkt_bits_pret,
  input         io_exu_bp_exu_mp_pkt_bits_pja,
  input         io_exu_bp_exu_mp_pkt_bits_way,
  input  [7:0]  io_exu_bp_exu_mp_eghr,
  input  [7:0]  io_exu_bp_exu_mp_fghr,
  input  [7:0]  io_exu_bp_exu_mp_index,
  input  [4:0]  io_exu_bp_exu_mp_btag,
  output        io_ifu_bp_hit_taken_f,
  output [30:0] io_ifu_bp_btb_target_f,
  output        io_ifu_bp_inst_mask_f,
  output [7:0]  io_ifu_bp_fghr_f,
  output [1:0]  io_ifu_bp_way_f,
  output [1:0]  io_ifu_bp_ret_f,
  output [1:0]  io_ifu_bp_hist1_f,
  output [1:0]  io_ifu_bp_hist0_f,
  output [1:0]  io_ifu_bp_pc4_f,
  output [1:0]  io_ifu_bp_valid_f,
  output [11:0] io_ifu_bp_poffset_f,
  input         io_scan_mode
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_576;
  reg [31:0] _RAND_577;
  reg [31:0] _RAND_578;
  reg [31:0] _RAND_579;
  reg [31:0] _RAND_580;
  reg [31:0] _RAND_581;
  reg [31:0] _RAND_582;
  reg [31:0] _RAND_583;
  reg [31:0] _RAND_584;
  reg [31:0] _RAND_585;
  reg [31:0] _RAND_586;
  reg [31:0] _RAND_587;
  reg [31:0] _RAND_588;
  reg [31:0] _RAND_589;
  reg [31:0] _RAND_590;
  reg [31:0] _RAND_591;
  reg [31:0] _RAND_592;
  reg [31:0] _RAND_593;
  reg [31:0] _RAND_594;
  reg [31:0] _RAND_595;
  reg [31:0] _RAND_596;
  reg [31:0] _RAND_597;
  reg [31:0] _RAND_598;
  reg [31:0] _RAND_599;
  reg [31:0] _RAND_600;
  reg [31:0] _RAND_601;
  reg [31:0] _RAND_602;
  reg [31:0] _RAND_603;
  reg [31:0] _RAND_604;
  reg [31:0] _RAND_605;
  reg [31:0] _RAND_606;
  reg [31:0] _RAND_607;
  reg [31:0] _RAND_608;
  reg [31:0] _RAND_609;
  reg [31:0] _RAND_610;
  reg [31:0] _RAND_611;
  reg [31:0] _RAND_612;
  reg [31:0] _RAND_613;
  reg [31:0] _RAND_614;
  reg [31:0] _RAND_615;
  reg [31:0] _RAND_616;
  reg [31:0] _RAND_617;
  reg [31:0] _RAND_618;
  reg [31:0] _RAND_619;
  reg [31:0] _RAND_620;
  reg [31:0] _RAND_621;
  reg [31:0] _RAND_622;
  reg [31:0] _RAND_623;
  reg [31:0] _RAND_624;
  reg [31:0] _RAND_625;
  reg [31:0] _RAND_626;
  reg [31:0] _RAND_627;
  reg [31:0] _RAND_628;
  reg [31:0] _RAND_629;
  reg [31:0] _RAND_630;
  reg [31:0] _RAND_631;
  reg [31:0] _RAND_632;
  reg [31:0] _RAND_633;
  reg [31:0] _RAND_634;
  reg [31:0] _RAND_635;
  reg [31:0] _RAND_636;
  reg [31:0] _RAND_637;
  reg [31:0] _RAND_638;
  reg [31:0] _RAND_639;
  reg [31:0] _RAND_640;
  reg [31:0] _RAND_641;
  reg [31:0] _RAND_642;
  reg [31:0] _RAND_643;
  reg [31:0] _RAND_644;
  reg [31:0] _RAND_645;
  reg [31:0] _RAND_646;
  reg [31:0] _RAND_647;
  reg [31:0] _RAND_648;
  reg [31:0] _RAND_649;
  reg [31:0] _RAND_650;
  reg [31:0] _RAND_651;
  reg [31:0] _RAND_652;
  reg [31:0] _RAND_653;
  reg [31:0] _RAND_654;
  reg [31:0] _RAND_655;
  reg [31:0] _RAND_656;
  reg [31:0] _RAND_657;
  reg [31:0] _RAND_658;
  reg [31:0] _RAND_659;
  reg [31:0] _RAND_660;
  reg [31:0] _RAND_661;
  reg [31:0] _RAND_662;
  reg [31:0] _RAND_663;
  reg [31:0] _RAND_664;
  reg [31:0] _RAND_665;
  reg [31:0] _RAND_666;
  reg [31:0] _RAND_667;
  reg [31:0] _RAND_668;
  reg [31:0] _RAND_669;
  reg [31:0] _RAND_670;
  reg [31:0] _RAND_671;
  reg [31:0] _RAND_672;
  reg [31:0] _RAND_673;
  reg [31:0] _RAND_674;
  reg [31:0] _RAND_675;
  reg [31:0] _RAND_676;
  reg [31:0] _RAND_677;
  reg [31:0] _RAND_678;
  reg [31:0] _RAND_679;
  reg [31:0] _RAND_680;
  reg [31:0] _RAND_681;
  reg [31:0] _RAND_682;
  reg [31:0] _RAND_683;
  reg [31:0] _RAND_684;
  reg [31:0] _RAND_685;
  reg [31:0] _RAND_686;
  reg [31:0] _RAND_687;
  reg [31:0] _RAND_688;
  reg [31:0] _RAND_689;
  reg [31:0] _RAND_690;
  reg [31:0] _RAND_691;
  reg [31:0] _RAND_692;
  reg [31:0] _RAND_693;
  reg [31:0] _RAND_694;
  reg [31:0] _RAND_695;
  reg [31:0] _RAND_696;
  reg [31:0] _RAND_697;
  reg [31:0] _RAND_698;
  reg [31:0] _RAND_699;
  reg [31:0] _RAND_700;
  reg [31:0] _RAND_701;
  reg [31:0] _RAND_702;
  reg [31:0] _RAND_703;
  reg [31:0] _RAND_704;
  reg [31:0] _RAND_705;
  reg [31:0] _RAND_706;
  reg [31:0] _RAND_707;
  reg [31:0] _RAND_708;
  reg [31:0] _RAND_709;
  reg [31:0] _RAND_710;
  reg [31:0] _RAND_711;
  reg [31:0] _RAND_712;
  reg [31:0] _RAND_713;
  reg [31:0] _RAND_714;
  reg [31:0] _RAND_715;
  reg [31:0] _RAND_716;
  reg [31:0] _RAND_717;
  reg [31:0] _RAND_718;
  reg [31:0] _RAND_719;
  reg [31:0] _RAND_720;
  reg [31:0] _RAND_721;
  reg [31:0] _RAND_722;
  reg [31:0] _RAND_723;
  reg [31:0] _RAND_724;
  reg [31:0] _RAND_725;
  reg [31:0] _RAND_726;
  reg [31:0] _RAND_727;
  reg [31:0] _RAND_728;
  reg [31:0] _RAND_729;
  reg [31:0] _RAND_730;
  reg [31:0] _RAND_731;
  reg [31:0] _RAND_732;
  reg [31:0] _RAND_733;
  reg [31:0] _RAND_734;
  reg [31:0] _RAND_735;
  reg [31:0] _RAND_736;
  reg [31:0] _RAND_737;
  reg [31:0] _RAND_738;
  reg [31:0] _RAND_739;
  reg [31:0] _RAND_740;
  reg [31:0] _RAND_741;
  reg [31:0] _RAND_742;
  reg [31:0] _RAND_743;
  reg [31:0] _RAND_744;
  reg [31:0] _RAND_745;
  reg [31:0] _RAND_746;
  reg [31:0] _RAND_747;
  reg [31:0] _RAND_748;
  reg [31:0] _RAND_749;
  reg [31:0] _RAND_750;
  reg [31:0] _RAND_751;
  reg [31:0] _RAND_752;
  reg [31:0] _RAND_753;
  reg [31:0] _RAND_754;
  reg [31:0] _RAND_755;
  reg [31:0] _RAND_756;
  reg [31:0] _RAND_757;
  reg [31:0] _RAND_758;
  reg [31:0] _RAND_759;
  reg [31:0] _RAND_760;
  reg [31:0] _RAND_761;
  reg [31:0] _RAND_762;
  reg [31:0] _RAND_763;
  reg [31:0] _RAND_764;
  reg [31:0] _RAND_765;
  reg [31:0] _RAND_766;
  reg [31:0] _RAND_767;
  reg [31:0] _RAND_768;
  reg [31:0] _RAND_769;
  reg [31:0] _RAND_770;
  reg [31:0] _RAND_771;
  reg [31:0] _RAND_772;
  reg [31:0] _RAND_773;
  reg [31:0] _RAND_774;
  reg [31:0] _RAND_775;
  reg [31:0] _RAND_776;
  reg [31:0] _RAND_777;
  reg [31:0] _RAND_778;
  reg [31:0] _RAND_779;
  reg [31:0] _RAND_780;
  reg [31:0] _RAND_781;
  reg [31:0] _RAND_782;
  reg [31:0] _RAND_783;
  reg [31:0] _RAND_784;
  reg [31:0] _RAND_785;
  reg [31:0] _RAND_786;
  reg [31:0] _RAND_787;
  reg [31:0] _RAND_788;
  reg [31:0] _RAND_789;
  reg [31:0] _RAND_790;
  reg [31:0] _RAND_791;
  reg [31:0] _RAND_792;
  reg [31:0] _RAND_793;
  reg [31:0] _RAND_794;
  reg [31:0] _RAND_795;
  reg [31:0] _RAND_796;
  reg [31:0] _RAND_797;
  reg [31:0] _RAND_798;
  reg [31:0] _RAND_799;
  reg [31:0] _RAND_800;
  reg [31:0] _RAND_801;
  reg [31:0] _RAND_802;
  reg [31:0] _RAND_803;
  reg [31:0] _RAND_804;
  reg [31:0] _RAND_805;
  reg [31:0] _RAND_806;
  reg [31:0] _RAND_807;
  reg [31:0] _RAND_808;
  reg [31:0] _RAND_809;
  reg [31:0] _RAND_810;
  reg [31:0] _RAND_811;
  reg [31:0] _RAND_812;
  reg [31:0] _RAND_813;
  reg [31:0] _RAND_814;
  reg [31:0] _RAND_815;
  reg [31:0] _RAND_816;
  reg [31:0] _RAND_817;
  reg [31:0] _RAND_818;
  reg [31:0] _RAND_819;
  reg [31:0] _RAND_820;
  reg [31:0] _RAND_821;
  reg [31:0] _RAND_822;
  reg [31:0] _RAND_823;
  reg [31:0] _RAND_824;
  reg [31:0] _RAND_825;
  reg [31:0] _RAND_826;
  reg [31:0] _RAND_827;
  reg [31:0] _RAND_828;
  reg [31:0] _RAND_829;
  reg [31:0] _RAND_830;
  reg [31:0] _RAND_831;
  reg [31:0] _RAND_832;
  reg [31:0] _RAND_833;
  reg [31:0] _RAND_834;
  reg [31:0] _RAND_835;
  reg [31:0] _RAND_836;
  reg [31:0] _RAND_837;
  reg [31:0] _RAND_838;
  reg [31:0] _RAND_839;
  reg [31:0] _RAND_840;
  reg [31:0] _RAND_841;
  reg [31:0] _RAND_842;
  reg [31:0] _RAND_843;
  reg [31:0] _RAND_844;
  reg [31:0] _RAND_845;
  reg [31:0] _RAND_846;
  reg [31:0] _RAND_847;
  reg [31:0] _RAND_848;
  reg [31:0] _RAND_849;
  reg [31:0] _RAND_850;
  reg [31:0] _RAND_851;
  reg [31:0] _RAND_852;
  reg [31:0] _RAND_853;
  reg [31:0] _RAND_854;
  reg [31:0] _RAND_855;
  reg [31:0] _RAND_856;
  reg [31:0] _RAND_857;
  reg [31:0] _RAND_858;
  reg [31:0] _RAND_859;
  reg [31:0] _RAND_860;
  reg [31:0] _RAND_861;
  reg [31:0] _RAND_862;
  reg [31:0] _RAND_863;
  reg [31:0] _RAND_864;
  reg [31:0] _RAND_865;
  reg [31:0] _RAND_866;
  reg [31:0] _RAND_867;
  reg [31:0] _RAND_868;
  reg [31:0] _RAND_869;
  reg [31:0] _RAND_870;
  reg [31:0] _RAND_871;
  reg [31:0] _RAND_872;
  reg [31:0] _RAND_873;
  reg [31:0] _RAND_874;
  reg [31:0] _RAND_875;
  reg [31:0] _RAND_876;
  reg [31:0] _RAND_877;
  reg [31:0] _RAND_878;
  reg [31:0] _RAND_879;
  reg [31:0] _RAND_880;
  reg [31:0] _RAND_881;
  reg [31:0] _RAND_882;
  reg [31:0] _RAND_883;
  reg [31:0] _RAND_884;
  reg [31:0] _RAND_885;
  reg [31:0] _RAND_886;
  reg [31:0] _RAND_887;
  reg [31:0] _RAND_888;
  reg [31:0] _RAND_889;
  reg [31:0] _RAND_890;
  reg [31:0] _RAND_891;
  reg [31:0] _RAND_892;
  reg [31:0] _RAND_893;
  reg [31:0] _RAND_894;
  reg [31:0] _RAND_895;
  reg [31:0] _RAND_896;
  reg [31:0] _RAND_897;
  reg [31:0] _RAND_898;
  reg [31:0] _RAND_899;
  reg [31:0] _RAND_900;
  reg [31:0] _RAND_901;
  reg [31:0] _RAND_902;
  reg [31:0] _RAND_903;
  reg [31:0] _RAND_904;
  reg [31:0] _RAND_905;
  reg [31:0] _RAND_906;
  reg [31:0] _RAND_907;
  reg [31:0] _RAND_908;
  reg [31:0] _RAND_909;
  reg [31:0] _RAND_910;
  reg [31:0] _RAND_911;
  reg [31:0] _RAND_912;
  reg [31:0] _RAND_913;
  reg [31:0] _RAND_914;
  reg [31:0] _RAND_915;
  reg [31:0] _RAND_916;
  reg [31:0] _RAND_917;
  reg [31:0] _RAND_918;
  reg [31:0] _RAND_919;
  reg [31:0] _RAND_920;
  reg [31:0] _RAND_921;
  reg [31:0] _RAND_922;
  reg [31:0] _RAND_923;
  reg [31:0] _RAND_924;
  reg [31:0] _RAND_925;
  reg [31:0] _RAND_926;
  reg [31:0] _RAND_927;
  reg [31:0] _RAND_928;
  reg [31:0] _RAND_929;
  reg [31:0] _RAND_930;
  reg [31:0] _RAND_931;
  reg [31:0] _RAND_932;
  reg [31:0] _RAND_933;
  reg [31:0] _RAND_934;
  reg [31:0] _RAND_935;
  reg [31:0] _RAND_936;
  reg [31:0] _RAND_937;
  reg [31:0] _RAND_938;
  reg [31:0] _RAND_939;
  reg [31:0] _RAND_940;
  reg [31:0] _RAND_941;
  reg [31:0] _RAND_942;
  reg [31:0] _RAND_943;
  reg [31:0] _RAND_944;
  reg [31:0] _RAND_945;
  reg [31:0] _RAND_946;
  reg [31:0] _RAND_947;
  reg [31:0] _RAND_948;
  reg [31:0] _RAND_949;
  reg [31:0] _RAND_950;
  reg [31:0] _RAND_951;
  reg [31:0] _RAND_952;
  reg [31:0] _RAND_953;
  reg [31:0] _RAND_954;
  reg [31:0] _RAND_955;
  reg [31:0] _RAND_956;
  reg [31:0] _RAND_957;
  reg [31:0] _RAND_958;
  reg [31:0] _RAND_959;
  reg [31:0] _RAND_960;
  reg [31:0] _RAND_961;
  reg [31:0] _RAND_962;
  reg [31:0] _RAND_963;
  reg [31:0] _RAND_964;
  reg [31:0] _RAND_965;
  reg [31:0] _RAND_966;
  reg [31:0] _RAND_967;
  reg [31:0] _RAND_968;
  reg [31:0] _RAND_969;
  reg [31:0] _RAND_970;
  reg [31:0] _RAND_971;
  reg [31:0] _RAND_972;
  reg [31:0] _RAND_973;
  reg [31:0] _RAND_974;
  reg [31:0] _RAND_975;
  reg [31:0] _RAND_976;
  reg [31:0] _RAND_977;
  reg [31:0] _RAND_978;
  reg [31:0] _RAND_979;
  reg [31:0] _RAND_980;
  reg [31:0] _RAND_981;
  reg [31:0] _RAND_982;
  reg [31:0] _RAND_983;
  reg [31:0] _RAND_984;
  reg [31:0] _RAND_985;
  reg [31:0] _RAND_986;
  reg [31:0] _RAND_987;
  reg [31:0] _RAND_988;
  reg [31:0] _RAND_989;
  reg [31:0] _RAND_990;
  reg [31:0] _RAND_991;
  reg [31:0] _RAND_992;
  reg [31:0] _RAND_993;
  reg [31:0] _RAND_994;
  reg [31:0] _RAND_995;
  reg [31:0] _RAND_996;
  reg [31:0] _RAND_997;
  reg [31:0] _RAND_998;
  reg [31:0] _RAND_999;
  reg [31:0] _RAND_1000;
  reg [31:0] _RAND_1001;
  reg [31:0] _RAND_1002;
  reg [31:0] _RAND_1003;
  reg [31:0] _RAND_1004;
  reg [31:0] _RAND_1005;
  reg [31:0] _RAND_1006;
  reg [31:0] _RAND_1007;
  reg [31:0] _RAND_1008;
  reg [31:0] _RAND_1009;
  reg [31:0] _RAND_1010;
  reg [31:0] _RAND_1011;
  reg [31:0] _RAND_1012;
  reg [31:0] _RAND_1013;
  reg [31:0] _RAND_1014;
  reg [31:0] _RAND_1015;
  reg [31:0] _RAND_1016;
  reg [31:0] _RAND_1017;
  reg [31:0] _RAND_1018;
  reg [31:0] _RAND_1019;
  reg [31:0] _RAND_1020;
  reg [31:0] _RAND_1021;
  reg [31:0] _RAND_1022;
  reg [31:0] _RAND_1023;
  reg [31:0] _RAND_1024;
  reg [31:0] _RAND_1025;
  reg [31:0] _RAND_1026;
  reg [31:0] _RAND_1027;
  reg [31:0] _RAND_1028;
  reg [255:0] _RAND_1029;
  reg [31:0] _RAND_1030;
  reg [31:0] _RAND_1031;
  reg [31:0] _RAND_1032;
  reg [31:0] _RAND_1033;
  reg [31:0] _RAND_1034;
  reg [31:0] _RAND_1035;
  reg [31:0] _RAND_1036;
  reg [31:0] _RAND_1037;
  reg [31:0] _RAND_1038;
`endif // RANDOMIZE_REG_INIT
  wire  rvclkhdr_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_1_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_1_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_1_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_1_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_2_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_2_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_2_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_2_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_3_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_3_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_3_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_3_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_4_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_4_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_4_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_4_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_5_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_5_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_5_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_5_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_6_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_6_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_6_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_6_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_7_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_7_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_7_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_7_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_8_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_8_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_8_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_8_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_9_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_9_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_9_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_9_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_10_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_10_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_10_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_10_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_11_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_11_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_11_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_11_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_12_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_12_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_12_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_12_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_13_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_13_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_13_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_13_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_14_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_14_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_14_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_14_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_15_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_15_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_15_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_15_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_16_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_16_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_16_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_16_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_17_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_17_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_17_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_17_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_18_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_18_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_18_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_18_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_19_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_19_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_19_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_19_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_20_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_20_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_20_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_20_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_21_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_21_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_21_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_21_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_22_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_22_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_22_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_22_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_23_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_23_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_23_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_23_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_24_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_24_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_24_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_24_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_25_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_25_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_25_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_25_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_26_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_26_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_26_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_26_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_27_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_27_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_27_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_27_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_28_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_28_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_28_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_28_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_29_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_29_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_29_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_29_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_30_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_30_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_30_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_30_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_31_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_31_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_31_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_31_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_32_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_32_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_32_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_32_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_33_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_33_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_33_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_33_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_34_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_34_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_34_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_34_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_35_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_35_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_35_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_35_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_36_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_36_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_36_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_36_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_37_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_37_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_37_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_37_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_38_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_38_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_38_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_38_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_39_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_39_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_39_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_39_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_40_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_40_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_40_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_40_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_41_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_41_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_41_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_41_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_42_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_42_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_42_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_42_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_43_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_43_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_43_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_43_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_44_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_44_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_44_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_44_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_45_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_45_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_45_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_45_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_46_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_46_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_46_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_46_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_47_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_47_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_47_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_47_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_48_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_48_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_48_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_48_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_49_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_49_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_49_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_49_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_50_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_50_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_50_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_50_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_51_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_51_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_51_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_51_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_52_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_52_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_52_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_52_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_53_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_53_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_53_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_53_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_54_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_54_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_54_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_54_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_55_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_55_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_55_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_55_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_56_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_56_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_56_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_56_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_57_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_57_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_57_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_57_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_58_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_58_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_58_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_58_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_59_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_59_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_59_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_59_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_60_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_60_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_60_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_60_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_61_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_61_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_61_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_61_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_62_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_62_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_62_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_62_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_63_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_63_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_63_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_63_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_64_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_64_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_64_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_64_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_65_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_65_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_65_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_65_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_66_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_66_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_66_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_66_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_67_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_67_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_67_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_67_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_68_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_68_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_68_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_68_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_69_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_69_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_69_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_69_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_70_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_70_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_70_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_70_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_71_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_71_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_71_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_71_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_72_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_72_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_72_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_72_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_73_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_73_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_73_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_73_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_74_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_74_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_74_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_74_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_75_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_75_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_75_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_75_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_76_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_76_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_76_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_76_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_77_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_77_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_77_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_77_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_78_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_78_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_78_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_78_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_79_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_79_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_79_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_79_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_80_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_80_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_80_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_80_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_81_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_81_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_81_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_81_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_82_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_82_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_82_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_82_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_83_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_83_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_83_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_83_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_84_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_84_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_84_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_84_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_85_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_85_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_85_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_85_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_86_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_86_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_86_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_86_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_87_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_87_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_87_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_87_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_88_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_88_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_88_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_88_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_89_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_89_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_89_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_89_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_90_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_90_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_90_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_90_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_91_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_91_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_91_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_91_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_92_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_92_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_92_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_92_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_93_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_93_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_93_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_93_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_94_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_94_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_94_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_94_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_95_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_95_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_95_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_95_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_96_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_96_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_96_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_96_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_97_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_97_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_97_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_97_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_98_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_98_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_98_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_98_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_99_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_99_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_99_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_99_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_100_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_100_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_100_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_100_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_101_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_101_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_101_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_101_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_102_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_102_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_102_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_102_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_103_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_103_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_103_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_103_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_104_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_104_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_104_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_104_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_105_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_105_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_105_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_105_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_106_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_106_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_106_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_106_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_107_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_107_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_107_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_107_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_108_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_108_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_108_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_108_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_109_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_109_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_109_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_109_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_110_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_110_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_110_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_110_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_111_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_111_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_111_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_111_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_112_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_112_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_112_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_112_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_113_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_113_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_113_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_113_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_114_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_114_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_114_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_114_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_115_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_115_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_115_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_115_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_116_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_116_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_116_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_116_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_117_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_117_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_117_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_117_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_118_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_118_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_118_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_118_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_119_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_119_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_119_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_119_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_120_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_120_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_120_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_120_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_121_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_121_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_121_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_121_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_122_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_122_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_122_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_122_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_123_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_123_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_123_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_123_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_124_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_124_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_124_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_124_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_125_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_125_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_125_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_125_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_126_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_126_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_126_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_126_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_127_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_127_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_127_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_127_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_128_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_128_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_128_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_128_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_129_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_129_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_129_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_129_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_130_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_130_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_130_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_130_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_131_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_131_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_131_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_131_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_132_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_132_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_132_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_132_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_133_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_133_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_133_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_133_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_134_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_134_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_134_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_134_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_135_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_135_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_135_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_135_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_136_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_136_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_136_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_136_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_137_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_137_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_137_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_137_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_138_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_138_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_138_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_138_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_139_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_139_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_139_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_139_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_140_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_140_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_140_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_140_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_141_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_141_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_141_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_141_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_142_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_142_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_142_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_142_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_143_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_143_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_143_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_143_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_144_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_144_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_144_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_144_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_145_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_145_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_145_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_145_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_146_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_146_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_146_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_146_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_147_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_147_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_147_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_147_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_148_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_148_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_148_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_148_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_149_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_149_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_149_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_149_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_150_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_150_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_150_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_150_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_151_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_151_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_151_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_151_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_152_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_152_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_152_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_152_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_153_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_153_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_153_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_153_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_154_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_154_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_154_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_154_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_155_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_155_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_155_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_155_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_156_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_156_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_156_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_156_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_157_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_157_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_157_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_157_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_158_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_158_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_158_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_158_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_159_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_159_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_159_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_159_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_160_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_160_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_160_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_160_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_161_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_161_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_161_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_161_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_162_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_162_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_162_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_162_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_163_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_163_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_163_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_163_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_164_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_164_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_164_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_164_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_165_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_165_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_165_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_165_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_166_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_166_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_166_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_166_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_167_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_167_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_167_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_167_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_168_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_168_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_168_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_168_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_169_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_169_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_169_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_169_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_170_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_170_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_170_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_170_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_171_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_171_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_171_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_171_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_172_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_172_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_172_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_172_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_173_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_173_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_173_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_173_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_174_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_174_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_174_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_174_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_175_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_175_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_175_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_175_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_176_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_176_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_176_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_176_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_177_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_177_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_177_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_177_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_178_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_178_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_178_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_178_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_179_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_179_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_179_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_179_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_180_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_180_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_180_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_180_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_181_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_181_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_181_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_181_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_182_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_182_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_182_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_182_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_183_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_183_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_183_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_183_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_184_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_184_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_184_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_184_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_185_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_185_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_185_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_185_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_186_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_186_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_186_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_186_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_187_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_187_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_187_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_187_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_188_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_188_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_188_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_188_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_189_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_189_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_189_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_189_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_190_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_190_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_190_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_190_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_191_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_191_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_191_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_191_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_192_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_192_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_192_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_192_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_193_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_193_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_193_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_193_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_194_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_194_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_194_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_194_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_195_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_195_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_195_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_195_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_196_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_196_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_196_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_196_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_197_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_197_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_197_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_197_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_198_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_198_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_198_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_198_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_199_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_199_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_199_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_199_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_200_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_200_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_200_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_200_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_201_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_201_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_201_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_201_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_202_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_202_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_202_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_202_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_203_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_203_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_203_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_203_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_204_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_204_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_204_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_204_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_205_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_205_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_205_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_205_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_206_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_206_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_206_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_206_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_207_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_207_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_207_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_207_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_208_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_208_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_208_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_208_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_209_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_209_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_209_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_209_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_210_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_210_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_210_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_210_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_211_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_211_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_211_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_211_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_212_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_212_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_212_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_212_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_213_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_213_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_213_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_213_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_214_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_214_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_214_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_214_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_215_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_215_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_215_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_215_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_216_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_216_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_216_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_216_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_217_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_217_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_217_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_217_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_218_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_218_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_218_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_218_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_219_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_219_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_219_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_219_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_220_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_220_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_220_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_220_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_221_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_221_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_221_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_221_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_222_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_222_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_222_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_222_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_223_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_223_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_223_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_223_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_224_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_224_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_224_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_224_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_225_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_225_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_225_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_225_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_226_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_226_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_226_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_226_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_227_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_227_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_227_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_227_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_228_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_228_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_228_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_228_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_229_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_229_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_229_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_229_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_230_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_230_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_230_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_230_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_231_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_231_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_231_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_231_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_232_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_232_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_232_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_232_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_233_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_233_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_233_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_233_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_234_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_234_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_234_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_234_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_235_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_235_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_235_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_235_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_236_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_236_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_236_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_236_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_237_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_237_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_237_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_237_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_238_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_238_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_238_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_238_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_239_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_239_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_239_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_239_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_240_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_240_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_240_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_240_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_241_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_241_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_241_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_241_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_242_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_242_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_242_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_242_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_243_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_243_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_243_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_243_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_244_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_244_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_244_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_244_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_245_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_245_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_245_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_245_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_246_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_246_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_246_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_246_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_247_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_247_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_247_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_247_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_248_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_248_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_248_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_248_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_249_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_249_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_249_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_249_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_250_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_250_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_250_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_250_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_251_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_251_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_251_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_251_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_252_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_252_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_252_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_252_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_253_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_253_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_253_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_253_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_254_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_254_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_254_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_254_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_255_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_255_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_255_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_255_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_256_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_256_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_256_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_256_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_257_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_257_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_257_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_257_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_258_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_258_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_258_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_258_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_259_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_259_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_259_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_259_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_260_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_260_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_260_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_260_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_261_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_261_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_261_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_261_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_262_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_262_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_262_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_262_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_263_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_263_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_263_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_263_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_264_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_264_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_264_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_264_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_265_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_265_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_265_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_265_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_266_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_266_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_266_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_266_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_267_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_267_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_267_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_267_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_268_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_268_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_268_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_268_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_269_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_269_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_269_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_269_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_270_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_270_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_270_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_270_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_271_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_271_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_271_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_271_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_272_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_272_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_272_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_272_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_273_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_273_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_273_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_273_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_274_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_274_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_274_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_274_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_275_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_275_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_275_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_275_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_276_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_276_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_276_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_276_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_277_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_277_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_277_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_277_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_278_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_278_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_278_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_278_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_279_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_279_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_279_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_279_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_280_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_280_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_280_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_280_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_281_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_281_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_281_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_281_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_282_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_282_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_282_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_282_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_283_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_283_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_283_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_283_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_284_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_284_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_284_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_284_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_285_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_285_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_285_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_285_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_286_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_286_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_286_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_286_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_287_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_287_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_287_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_287_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_288_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_288_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_288_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_288_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_289_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_289_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_289_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_289_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_290_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_290_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_290_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_290_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_291_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_291_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_291_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_291_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_292_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_292_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_292_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_292_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_293_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_293_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_293_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_293_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_294_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_294_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_294_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_294_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_295_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_295_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_295_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_295_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_296_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_296_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_296_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_296_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_297_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_297_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_297_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_297_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_298_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_298_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_298_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_298_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_299_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_299_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_299_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_299_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_300_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_300_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_300_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_300_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_301_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_301_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_301_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_301_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_302_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_302_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_302_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_302_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_303_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_303_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_303_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_303_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_304_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_304_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_304_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_304_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_305_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_305_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_305_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_305_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_306_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_306_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_306_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_306_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_307_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_307_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_307_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_307_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_308_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_308_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_308_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_308_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_309_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_309_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_309_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_309_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_310_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_310_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_310_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_310_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_311_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_311_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_311_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_311_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_312_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_312_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_312_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_312_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_313_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_313_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_313_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_313_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_314_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_314_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_314_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_314_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_315_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_315_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_315_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_315_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_316_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_316_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_316_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_316_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_317_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_317_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_317_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_317_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_318_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_318_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_318_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_318_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_319_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_319_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_319_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_319_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_320_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_320_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_320_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_320_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_321_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_321_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_321_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_321_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_322_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_322_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_322_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_322_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_323_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_323_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_323_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_323_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_324_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_324_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_324_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_324_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_325_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_325_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_325_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_325_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_326_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_326_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_326_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_326_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_327_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_327_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_327_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_327_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_328_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_328_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_328_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_328_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_329_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_329_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_329_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_329_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_330_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_330_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_330_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_330_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_331_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_331_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_331_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_331_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_332_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_332_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_332_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_332_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_333_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_333_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_333_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_333_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_334_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_334_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_334_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_334_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_335_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_335_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_335_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_335_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_336_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_336_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_336_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_336_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_337_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_337_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_337_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_337_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_338_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_338_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_338_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_338_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_339_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_339_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_339_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_339_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_340_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_340_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_340_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_340_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_341_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_341_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_341_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_341_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_342_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_342_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_342_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_342_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_343_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_343_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_343_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_343_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_344_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_344_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_344_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_344_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_345_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_345_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_345_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_345_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_346_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_346_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_346_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_346_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_347_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_347_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_347_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_347_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_348_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_348_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_348_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_348_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_349_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_349_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_349_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_349_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_350_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_350_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_350_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_350_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_351_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_351_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_351_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_351_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_352_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_352_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_352_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_352_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_353_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_353_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_353_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_353_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_354_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_354_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_354_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_354_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_355_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_355_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_355_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_355_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_356_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_356_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_356_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_356_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_357_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_357_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_357_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_357_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_358_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_358_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_358_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_358_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_359_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_359_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_359_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_359_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_360_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_360_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_360_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_360_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_361_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_361_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_361_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_361_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_362_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_362_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_362_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_362_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_363_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_363_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_363_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_363_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_364_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_364_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_364_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_364_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_365_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_365_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_365_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_365_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_366_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_366_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_366_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_366_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_367_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_367_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_367_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_367_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_368_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_368_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_368_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_368_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_369_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_369_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_369_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_369_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_370_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_370_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_370_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_370_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_371_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_371_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_371_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_371_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_372_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_372_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_372_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_372_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_373_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_373_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_373_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_373_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_374_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_374_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_374_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_374_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_375_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_375_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_375_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_375_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_376_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_376_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_376_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_376_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_377_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_377_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_377_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_377_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_378_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_378_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_378_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_378_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_379_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_379_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_379_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_379_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_380_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_380_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_380_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_380_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_381_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_381_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_381_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_381_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_382_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_382_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_382_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_382_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_383_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_383_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_383_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_383_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_384_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_384_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_384_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_384_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_385_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_385_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_385_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_385_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_386_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_386_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_386_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_386_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_387_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_387_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_387_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_387_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_388_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_388_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_388_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_388_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_389_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_389_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_389_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_389_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_390_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_390_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_390_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_390_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_391_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_391_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_391_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_391_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_392_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_392_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_392_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_392_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_393_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_393_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_393_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_393_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_394_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_394_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_394_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_394_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_395_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_395_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_395_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_395_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_396_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_396_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_396_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_396_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_397_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_397_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_397_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_397_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_398_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_398_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_398_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_398_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_399_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_399_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_399_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_399_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_400_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_400_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_400_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_400_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_401_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_401_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_401_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_401_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_402_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_402_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_402_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_402_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_403_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_403_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_403_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_403_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_404_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_404_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_404_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_404_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_405_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_405_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_405_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_405_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_406_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_406_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_406_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_406_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_407_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_407_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_407_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_407_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_408_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_408_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_408_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_408_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_409_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_409_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_409_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_409_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_410_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_410_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_410_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_410_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_411_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_411_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_411_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_411_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_412_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_412_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_412_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_412_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_413_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_413_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_413_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_413_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_414_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_414_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_414_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_414_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_415_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_415_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_415_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_415_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_416_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_416_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_416_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_416_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_417_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_417_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_417_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_417_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_418_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_418_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_418_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_418_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_419_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_419_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_419_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_419_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_420_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_420_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_420_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_420_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_421_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_421_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_421_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_421_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_422_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_422_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_422_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_422_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_423_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_423_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_423_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_423_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_424_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_424_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_424_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_424_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_425_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_425_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_425_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_425_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_426_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_426_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_426_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_426_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_427_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_427_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_427_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_427_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_428_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_428_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_428_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_428_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_429_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_429_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_429_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_429_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_430_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_430_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_430_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_430_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_431_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_431_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_431_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_431_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_432_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_432_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_432_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_432_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_433_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_433_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_433_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_433_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_434_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_434_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_434_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_434_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_435_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_435_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_435_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_435_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_436_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_436_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_436_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_436_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_437_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_437_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_437_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_437_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_438_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_438_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_438_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_438_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_439_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_439_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_439_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_439_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_440_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_440_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_440_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_440_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_441_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_441_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_441_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_441_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_442_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_442_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_442_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_442_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_443_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_443_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_443_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_443_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_444_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_444_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_444_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_444_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_445_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_445_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_445_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_445_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_446_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_446_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_446_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_446_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_447_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_447_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_447_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_447_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_448_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_448_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_448_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_448_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_449_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_449_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_449_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_449_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_450_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_450_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_450_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_450_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_451_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_451_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_451_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_451_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_452_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_452_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_452_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_452_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_453_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_453_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_453_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_453_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_454_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_454_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_454_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_454_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_455_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_455_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_455_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_455_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_456_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_456_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_456_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_456_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_457_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_457_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_457_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_457_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_458_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_458_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_458_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_458_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_459_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_459_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_459_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_459_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_460_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_460_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_460_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_460_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_461_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_461_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_461_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_461_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_462_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_462_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_462_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_462_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_463_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_463_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_463_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_463_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_464_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_464_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_464_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_464_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_465_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_465_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_465_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_465_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_466_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_466_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_466_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_466_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_467_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_467_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_467_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_467_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_468_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_468_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_468_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_468_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_469_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_469_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_469_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_469_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_470_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_470_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_470_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_470_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_471_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_471_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_471_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_471_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_472_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_472_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_472_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_472_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_473_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_473_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_473_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_473_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_474_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_474_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_474_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_474_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_475_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_475_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_475_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_475_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_476_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_476_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_476_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_476_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_477_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_477_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_477_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_477_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_478_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_478_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_478_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_478_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_479_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_479_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_479_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_479_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_480_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_480_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_480_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_480_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_481_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_481_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_481_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_481_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_482_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_482_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_482_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_482_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_483_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_483_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_483_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_483_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_484_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_484_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_484_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_484_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_485_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_485_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_485_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_485_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_486_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_486_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_486_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_486_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_487_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_487_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_487_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_487_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_488_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_488_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_488_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_488_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_489_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_489_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_489_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_489_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_490_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_490_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_490_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_490_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_491_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_491_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_491_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_491_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_492_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_492_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_492_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_492_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_493_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_493_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_493_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_493_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_494_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_494_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_494_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_494_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_495_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_495_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_495_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_495_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_496_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_496_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_496_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_496_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_497_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_497_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_497_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_497_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_498_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_498_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_498_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_498_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_499_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_499_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_499_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_499_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_500_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_500_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_500_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_500_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_501_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_501_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_501_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_501_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_502_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_502_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_502_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_502_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_503_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_503_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_503_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_503_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_504_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_504_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_504_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_504_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_505_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_505_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_505_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_505_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_506_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_506_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_506_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_506_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_507_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_507_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_507_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_507_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_508_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_508_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_508_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_508_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_509_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_509_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_509_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_509_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_510_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_510_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_510_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_510_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_511_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_511_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_511_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_511_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_512_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_512_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_512_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_512_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_513_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_513_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_513_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_513_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_514_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_514_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_514_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_514_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_515_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_515_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_515_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_515_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_516_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_516_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_516_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_516_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_517_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_517_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_517_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_517_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_518_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_518_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_518_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_518_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_519_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_519_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_519_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_519_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_520_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_520_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_520_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_520_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_521_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_521_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_521_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_521_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_522_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_522_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_522_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_522_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_523_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_523_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_523_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_523_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_524_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_524_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_524_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_524_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_525_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_525_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_525_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_525_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_526_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_526_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_526_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_526_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_527_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_527_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_527_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_527_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_528_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_528_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_528_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_528_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_529_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_529_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_529_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_529_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_530_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_530_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_530_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_530_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_531_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_531_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_531_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_531_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_532_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_532_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_532_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_532_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_533_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_533_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_533_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_533_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_534_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_534_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_534_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_534_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_535_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_535_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_535_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_535_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_536_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_536_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_536_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_536_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_537_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_537_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_537_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_537_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_538_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_538_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_538_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_538_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_539_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_539_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_539_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_539_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_540_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_540_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_540_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_540_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_541_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_541_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_541_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_541_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_542_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_542_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_542_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_542_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_543_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_543_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_543_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_543_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_544_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_544_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_544_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_544_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_545_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_545_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_545_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_545_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_546_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_546_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_546_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_546_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_547_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_547_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_547_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_547_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_548_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_548_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_548_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_548_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_549_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_549_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_549_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_549_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_550_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_550_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_550_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_550_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_551_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_551_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_551_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_551_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_552_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_552_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_552_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_552_io_scan_mode; // @[lib.scala 343:22]
  wire  rvclkhdr_553_io_l1clk; // @[lib.scala 343:22]
  wire  rvclkhdr_553_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_553_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_553_io_scan_mode; // @[lib.scala 343:22]
  wire  _T_40 = io_dec_bp_dec_tlu_flush_leak_one_wb & io_dec_tlu_flush_lower_wb; // @[ifu_bp_ctl.scala 123:54]
  reg  leak_one_f_d1; // @[ifu_bp_ctl.scala 117:56]
  wire  _T_41 = ~io_dec_tlu_flush_lower_wb; // @[ifu_bp_ctl.scala 123:102]
  wire  _T_42 = leak_one_f_d1 & _T_41; // @[ifu_bp_ctl.scala 123:100]
  wire  leak_one_f = _T_40 | _T_42; // @[ifu_bp_ctl.scala 123:83]
  wire  _T = ~leak_one_f; // @[ifu_bp_ctl.scala 60:58]
  wire  exu_mp_valid = io_exu_bp_exu_mp_pkt_bits_misp & _T; // @[ifu_bp_ctl.scala 60:56]
  wire  dec_tlu_error_wb = io_dec_bp_dec_tlu_br0_r_pkt_bits_br_start_error | io_dec_bp_dec_tlu_br0_r_pkt_bits_br_error; // @[ifu_bp_ctl.scala 82:50]
  wire [7:0] _T_4 = io_ifc_fetch_addr_f[8:1] ^ io_ifc_fetch_addr_f[16:9]; // @[lib.scala 51:47]
  wire [7:0] btb_rd_addr_f = _T_4 ^ io_ifc_fetch_addr_f[24:17]; // @[lib.scala 51:85]
  wire [29:0] fetch_addr_p1_f = io_ifc_fetch_addr_f[30:1] + 30'h1; // @[ifu_bp_ctl.scala 90:51]
  wire [30:0] _T_8 = {fetch_addr_p1_f,1'h0}; // @[Cat.scala 29:58]
  wire [7:0] _T_11 = _T_8[8:1] ^ _T_8[16:9]; // @[lib.scala 51:47]
  wire [7:0] btb_rd_addr_p1_f = _T_11 ^ _T_8[24:17]; // @[lib.scala 51:85]
  wire  _T_144 = ~io_ifc_fetch_addr_f[0]; // @[ifu_bp_ctl.scala 174:40]
  wire  _T_2112 = btb_rd_addr_f == 8'h0; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_0; // @[lib.scala 374:16]
  wire [21:0] _T_2624 = _T_2112 ? btb_bank0_rd_data_way0_out_0 : 22'h0; // @[Mux.scala 27:72]
  wire  _T_2114 = btb_rd_addr_f == 8'h1; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_1; // @[lib.scala 374:16]
  wire [21:0] _T_2625 = _T_2114 ? btb_bank0_rd_data_way0_out_1 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2880 = _T_2624 | _T_2625; // @[Mux.scala 27:72]
  wire  _T_2116 = btb_rd_addr_f == 8'h2; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_2; // @[lib.scala 374:16]
  wire [21:0] _T_2626 = _T_2116 ? btb_bank0_rd_data_way0_out_2 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2881 = _T_2880 | _T_2626; // @[Mux.scala 27:72]
  wire  _T_2118 = btb_rd_addr_f == 8'h3; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_3; // @[lib.scala 374:16]
  wire [21:0] _T_2627 = _T_2118 ? btb_bank0_rd_data_way0_out_3 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2882 = _T_2881 | _T_2627; // @[Mux.scala 27:72]
  wire  _T_2120 = btb_rd_addr_f == 8'h4; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_4; // @[lib.scala 374:16]
  wire [21:0] _T_2628 = _T_2120 ? btb_bank0_rd_data_way0_out_4 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2883 = _T_2882 | _T_2628; // @[Mux.scala 27:72]
  wire  _T_2122 = btb_rd_addr_f == 8'h5; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_5; // @[lib.scala 374:16]
  wire [21:0] _T_2629 = _T_2122 ? btb_bank0_rd_data_way0_out_5 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2884 = _T_2883 | _T_2629; // @[Mux.scala 27:72]
  wire  _T_2124 = btb_rd_addr_f == 8'h6; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_6; // @[lib.scala 374:16]
  wire [21:0] _T_2630 = _T_2124 ? btb_bank0_rd_data_way0_out_6 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2885 = _T_2884 | _T_2630; // @[Mux.scala 27:72]
  wire  _T_2126 = btb_rd_addr_f == 8'h7; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_7; // @[lib.scala 374:16]
  wire [21:0] _T_2631 = _T_2126 ? btb_bank0_rd_data_way0_out_7 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2886 = _T_2885 | _T_2631; // @[Mux.scala 27:72]
  wire  _T_2128 = btb_rd_addr_f == 8'h8; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_8; // @[lib.scala 374:16]
  wire [21:0] _T_2632 = _T_2128 ? btb_bank0_rd_data_way0_out_8 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2887 = _T_2886 | _T_2632; // @[Mux.scala 27:72]
  wire  _T_2130 = btb_rd_addr_f == 8'h9; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_9; // @[lib.scala 374:16]
  wire [21:0] _T_2633 = _T_2130 ? btb_bank0_rd_data_way0_out_9 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2888 = _T_2887 | _T_2633; // @[Mux.scala 27:72]
  wire  _T_2132 = btb_rd_addr_f == 8'ha; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_10; // @[lib.scala 374:16]
  wire [21:0] _T_2634 = _T_2132 ? btb_bank0_rd_data_way0_out_10 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2889 = _T_2888 | _T_2634; // @[Mux.scala 27:72]
  wire  _T_2134 = btb_rd_addr_f == 8'hb; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_11; // @[lib.scala 374:16]
  wire [21:0] _T_2635 = _T_2134 ? btb_bank0_rd_data_way0_out_11 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2890 = _T_2889 | _T_2635; // @[Mux.scala 27:72]
  wire  _T_2136 = btb_rd_addr_f == 8'hc; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_12; // @[lib.scala 374:16]
  wire [21:0] _T_2636 = _T_2136 ? btb_bank0_rd_data_way0_out_12 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2891 = _T_2890 | _T_2636; // @[Mux.scala 27:72]
  wire  _T_2138 = btb_rd_addr_f == 8'hd; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_13; // @[lib.scala 374:16]
  wire [21:0] _T_2637 = _T_2138 ? btb_bank0_rd_data_way0_out_13 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2892 = _T_2891 | _T_2637; // @[Mux.scala 27:72]
  wire  _T_2140 = btb_rd_addr_f == 8'he; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_14; // @[lib.scala 374:16]
  wire [21:0] _T_2638 = _T_2140 ? btb_bank0_rd_data_way0_out_14 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2893 = _T_2892 | _T_2638; // @[Mux.scala 27:72]
  wire  _T_2142 = btb_rd_addr_f == 8'hf; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_15; // @[lib.scala 374:16]
  wire [21:0] _T_2639 = _T_2142 ? btb_bank0_rd_data_way0_out_15 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2894 = _T_2893 | _T_2639; // @[Mux.scala 27:72]
  wire  _T_2144 = btb_rd_addr_f == 8'h10; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_16; // @[lib.scala 374:16]
  wire [21:0] _T_2640 = _T_2144 ? btb_bank0_rd_data_way0_out_16 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2895 = _T_2894 | _T_2640; // @[Mux.scala 27:72]
  wire  _T_2146 = btb_rd_addr_f == 8'h11; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_17; // @[lib.scala 374:16]
  wire [21:0] _T_2641 = _T_2146 ? btb_bank0_rd_data_way0_out_17 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2896 = _T_2895 | _T_2641; // @[Mux.scala 27:72]
  wire  _T_2148 = btb_rd_addr_f == 8'h12; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_18; // @[lib.scala 374:16]
  wire [21:0] _T_2642 = _T_2148 ? btb_bank0_rd_data_way0_out_18 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2897 = _T_2896 | _T_2642; // @[Mux.scala 27:72]
  wire  _T_2150 = btb_rd_addr_f == 8'h13; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_19; // @[lib.scala 374:16]
  wire [21:0] _T_2643 = _T_2150 ? btb_bank0_rd_data_way0_out_19 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2898 = _T_2897 | _T_2643; // @[Mux.scala 27:72]
  wire  _T_2152 = btb_rd_addr_f == 8'h14; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_20; // @[lib.scala 374:16]
  wire [21:0] _T_2644 = _T_2152 ? btb_bank0_rd_data_way0_out_20 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2899 = _T_2898 | _T_2644; // @[Mux.scala 27:72]
  wire  _T_2154 = btb_rd_addr_f == 8'h15; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_21; // @[lib.scala 374:16]
  wire [21:0] _T_2645 = _T_2154 ? btb_bank0_rd_data_way0_out_21 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2900 = _T_2899 | _T_2645; // @[Mux.scala 27:72]
  wire  _T_2156 = btb_rd_addr_f == 8'h16; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_22; // @[lib.scala 374:16]
  wire [21:0] _T_2646 = _T_2156 ? btb_bank0_rd_data_way0_out_22 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2901 = _T_2900 | _T_2646; // @[Mux.scala 27:72]
  wire  _T_2158 = btb_rd_addr_f == 8'h17; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_23; // @[lib.scala 374:16]
  wire [21:0] _T_2647 = _T_2158 ? btb_bank0_rd_data_way0_out_23 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2902 = _T_2901 | _T_2647; // @[Mux.scala 27:72]
  wire  _T_2160 = btb_rd_addr_f == 8'h18; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_24; // @[lib.scala 374:16]
  wire [21:0] _T_2648 = _T_2160 ? btb_bank0_rd_data_way0_out_24 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2903 = _T_2902 | _T_2648; // @[Mux.scala 27:72]
  wire  _T_2162 = btb_rd_addr_f == 8'h19; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_25; // @[lib.scala 374:16]
  wire [21:0] _T_2649 = _T_2162 ? btb_bank0_rd_data_way0_out_25 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2904 = _T_2903 | _T_2649; // @[Mux.scala 27:72]
  wire  _T_2164 = btb_rd_addr_f == 8'h1a; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_26; // @[lib.scala 374:16]
  wire [21:0] _T_2650 = _T_2164 ? btb_bank0_rd_data_way0_out_26 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2905 = _T_2904 | _T_2650; // @[Mux.scala 27:72]
  wire  _T_2166 = btb_rd_addr_f == 8'h1b; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_27; // @[lib.scala 374:16]
  wire [21:0] _T_2651 = _T_2166 ? btb_bank0_rd_data_way0_out_27 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2906 = _T_2905 | _T_2651; // @[Mux.scala 27:72]
  wire  _T_2168 = btb_rd_addr_f == 8'h1c; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_28; // @[lib.scala 374:16]
  wire [21:0] _T_2652 = _T_2168 ? btb_bank0_rd_data_way0_out_28 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2907 = _T_2906 | _T_2652; // @[Mux.scala 27:72]
  wire  _T_2170 = btb_rd_addr_f == 8'h1d; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_29; // @[lib.scala 374:16]
  wire [21:0] _T_2653 = _T_2170 ? btb_bank0_rd_data_way0_out_29 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2908 = _T_2907 | _T_2653; // @[Mux.scala 27:72]
  wire  _T_2172 = btb_rd_addr_f == 8'h1e; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_30; // @[lib.scala 374:16]
  wire [21:0] _T_2654 = _T_2172 ? btb_bank0_rd_data_way0_out_30 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2909 = _T_2908 | _T_2654; // @[Mux.scala 27:72]
  wire  _T_2174 = btb_rd_addr_f == 8'h1f; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_31; // @[lib.scala 374:16]
  wire [21:0] _T_2655 = _T_2174 ? btb_bank0_rd_data_way0_out_31 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2910 = _T_2909 | _T_2655; // @[Mux.scala 27:72]
  wire  _T_2176 = btb_rd_addr_f == 8'h20; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_32; // @[lib.scala 374:16]
  wire [21:0] _T_2656 = _T_2176 ? btb_bank0_rd_data_way0_out_32 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2911 = _T_2910 | _T_2656; // @[Mux.scala 27:72]
  wire  _T_2178 = btb_rd_addr_f == 8'h21; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_33; // @[lib.scala 374:16]
  wire [21:0] _T_2657 = _T_2178 ? btb_bank0_rd_data_way0_out_33 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2912 = _T_2911 | _T_2657; // @[Mux.scala 27:72]
  wire  _T_2180 = btb_rd_addr_f == 8'h22; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_34; // @[lib.scala 374:16]
  wire [21:0] _T_2658 = _T_2180 ? btb_bank0_rd_data_way0_out_34 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2913 = _T_2912 | _T_2658; // @[Mux.scala 27:72]
  wire  _T_2182 = btb_rd_addr_f == 8'h23; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_35; // @[lib.scala 374:16]
  wire [21:0] _T_2659 = _T_2182 ? btb_bank0_rd_data_way0_out_35 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2914 = _T_2913 | _T_2659; // @[Mux.scala 27:72]
  wire  _T_2184 = btb_rd_addr_f == 8'h24; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_36; // @[lib.scala 374:16]
  wire [21:0] _T_2660 = _T_2184 ? btb_bank0_rd_data_way0_out_36 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2915 = _T_2914 | _T_2660; // @[Mux.scala 27:72]
  wire  _T_2186 = btb_rd_addr_f == 8'h25; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_37; // @[lib.scala 374:16]
  wire [21:0] _T_2661 = _T_2186 ? btb_bank0_rd_data_way0_out_37 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2916 = _T_2915 | _T_2661; // @[Mux.scala 27:72]
  wire  _T_2188 = btb_rd_addr_f == 8'h26; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_38; // @[lib.scala 374:16]
  wire [21:0] _T_2662 = _T_2188 ? btb_bank0_rd_data_way0_out_38 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2917 = _T_2916 | _T_2662; // @[Mux.scala 27:72]
  wire  _T_2190 = btb_rd_addr_f == 8'h27; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_39; // @[lib.scala 374:16]
  wire [21:0] _T_2663 = _T_2190 ? btb_bank0_rd_data_way0_out_39 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2918 = _T_2917 | _T_2663; // @[Mux.scala 27:72]
  wire  _T_2192 = btb_rd_addr_f == 8'h28; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_40; // @[lib.scala 374:16]
  wire [21:0] _T_2664 = _T_2192 ? btb_bank0_rd_data_way0_out_40 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2919 = _T_2918 | _T_2664; // @[Mux.scala 27:72]
  wire  _T_2194 = btb_rd_addr_f == 8'h29; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_41; // @[lib.scala 374:16]
  wire [21:0] _T_2665 = _T_2194 ? btb_bank0_rd_data_way0_out_41 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2920 = _T_2919 | _T_2665; // @[Mux.scala 27:72]
  wire  _T_2196 = btb_rd_addr_f == 8'h2a; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_42; // @[lib.scala 374:16]
  wire [21:0] _T_2666 = _T_2196 ? btb_bank0_rd_data_way0_out_42 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2921 = _T_2920 | _T_2666; // @[Mux.scala 27:72]
  wire  _T_2198 = btb_rd_addr_f == 8'h2b; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_43; // @[lib.scala 374:16]
  wire [21:0] _T_2667 = _T_2198 ? btb_bank0_rd_data_way0_out_43 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2922 = _T_2921 | _T_2667; // @[Mux.scala 27:72]
  wire  _T_2200 = btb_rd_addr_f == 8'h2c; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_44; // @[lib.scala 374:16]
  wire [21:0] _T_2668 = _T_2200 ? btb_bank0_rd_data_way0_out_44 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2923 = _T_2922 | _T_2668; // @[Mux.scala 27:72]
  wire  _T_2202 = btb_rd_addr_f == 8'h2d; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_45; // @[lib.scala 374:16]
  wire [21:0] _T_2669 = _T_2202 ? btb_bank0_rd_data_way0_out_45 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2924 = _T_2923 | _T_2669; // @[Mux.scala 27:72]
  wire  _T_2204 = btb_rd_addr_f == 8'h2e; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_46; // @[lib.scala 374:16]
  wire [21:0] _T_2670 = _T_2204 ? btb_bank0_rd_data_way0_out_46 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2925 = _T_2924 | _T_2670; // @[Mux.scala 27:72]
  wire  _T_2206 = btb_rd_addr_f == 8'h2f; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_47; // @[lib.scala 374:16]
  wire [21:0] _T_2671 = _T_2206 ? btb_bank0_rd_data_way0_out_47 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2926 = _T_2925 | _T_2671; // @[Mux.scala 27:72]
  wire  _T_2208 = btb_rd_addr_f == 8'h30; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_48; // @[lib.scala 374:16]
  wire [21:0] _T_2672 = _T_2208 ? btb_bank0_rd_data_way0_out_48 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2927 = _T_2926 | _T_2672; // @[Mux.scala 27:72]
  wire  _T_2210 = btb_rd_addr_f == 8'h31; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_49; // @[lib.scala 374:16]
  wire [21:0] _T_2673 = _T_2210 ? btb_bank0_rd_data_way0_out_49 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2928 = _T_2927 | _T_2673; // @[Mux.scala 27:72]
  wire  _T_2212 = btb_rd_addr_f == 8'h32; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_50; // @[lib.scala 374:16]
  wire [21:0] _T_2674 = _T_2212 ? btb_bank0_rd_data_way0_out_50 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2929 = _T_2928 | _T_2674; // @[Mux.scala 27:72]
  wire  _T_2214 = btb_rd_addr_f == 8'h33; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_51; // @[lib.scala 374:16]
  wire [21:0] _T_2675 = _T_2214 ? btb_bank0_rd_data_way0_out_51 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2930 = _T_2929 | _T_2675; // @[Mux.scala 27:72]
  wire  _T_2216 = btb_rd_addr_f == 8'h34; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_52; // @[lib.scala 374:16]
  wire [21:0] _T_2676 = _T_2216 ? btb_bank0_rd_data_way0_out_52 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2931 = _T_2930 | _T_2676; // @[Mux.scala 27:72]
  wire  _T_2218 = btb_rd_addr_f == 8'h35; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_53; // @[lib.scala 374:16]
  wire [21:0] _T_2677 = _T_2218 ? btb_bank0_rd_data_way0_out_53 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2932 = _T_2931 | _T_2677; // @[Mux.scala 27:72]
  wire  _T_2220 = btb_rd_addr_f == 8'h36; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_54; // @[lib.scala 374:16]
  wire [21:0] _T_2678 = _T_2220 ? btb_bank0_rd_data_way0_out_54 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2933 = _T_2932 | _T_2678; // @[Mux.scala 27:72]
  wire  _T_2222 = btb_rd_addr_f == 8'h37; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_55; // @[lib.scala 374:16]
  wire [21:0] _T_2679 = _T_2222 ? btb_bank0_rd_data_way0_out_55 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2934 = _T_2933 | _T_2679; // @[Mux.scala 27:72]
  wire  _T_2224 = btb_rd_addr_f == 8'h38; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_56; // @[lib.scala 374:16]
  wire [21:0] _T_2680 = _T_2224 ? btb_bank0_rd_data_way0_out_56 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2935 = _T_2934 | _T_2680; // @[Mux.scala 27:72]
  wire  _T_2226 = btb_rd_addr_f == 8'h39; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_57; // @[lib.scala 374:16]
  wire [21:0] _T_2681 = _T_2226 ? btb_bank0_rd_data_way0_out_57 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2936 = _T_2935 | _T_2681; // @[Mux.scala 27:72]
  wire  _T_2228 = btb_rd_addr_f == 8'h3a; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_58; // @[lib.scala 374:16]
  wire [21:0] _T_2682 = _T_2228 ? btb_bank0_rd_data_way0_out_58 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2937 = _T_2936 | _T_2682; // @[Mux.scala 27:72]
  wire  _T_2230 = btb_rd_addr_f == 8'h3b; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_59; // @[lib.scala 374:16]
  wire [21:0] _T_2683 = _T_2230 ? btb_bank0_rd_data_way0_out_59 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2938 = _T_2937 | _T_2683; // @[Mux.scala 27:72]
  wire  _T_2232 = btb_rd_addr_f == 8'h3c; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_60; // @[lib.scala 374:16]
  wire [21:0] _T_2684 = _T_2232 ? btb_bank0_rd_data_way0_out_60 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2939 = _T_2938 | _T_2684; // @[Mux.scala 27:72]
  wire  _T_2234 = btb_rd_addr_f == 8'h3d; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_61; // @[lib.scala 374:16]
  wire [21:0] _T_2685 = _T_2234 ? btb_bank0_rd_data_way0_out_61 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2940 = _T_2939 | _T_2685; // @[Mux.scala 27:72]
  wire  _T_2236 = btb_rd_addr_f == 8'h3e; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_62; // @[lib.scala 374:16]
  wire [21:0] _T_2686 = _T_2236 ? btb_bank0_rd_data_way0_out_62 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2941 = _T_2940 | _T_2686; // @[Mux.scala 27:72]
  wire  _T_2238 = btb_rd_addr_f == 8'h3f; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_63; // @[lib.scala 374:16]
  wire [21:0] _T_2687 = _T_2238 ? btb_bank0_rd_data_way0_out_63 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2942 = _T_2941 | _T_2687; // @[Mux.scala 27:72]
  wire  _T_2240 = btb_rd_addr_f == 8'h40; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_64; // @[lib.scala 374:16]
  wire [21:0] _T_2688 = _T_2240 ? btb_bank0_rd_data_way0_out_64 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2943 = _T_2942 | _T_2688; // @[Mux.scala 27:72]
  wire  _T_2242 = btb_rd_addr_f == 8'h41; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_65; // @[lib.scala 374:16]
  wire [21:0] _T_2689 = _T_2242 ? btb_bank0_rd_data_way0_out_65 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2944 = _T_2943 | _T_2689; // @[Mux.scala 27:72]
  wire  _T_2244 = btb_rd_addr_f == 8'h42; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_66; // @[lib.scala 374:16]
  wire [21:0] _T_2690 = _T_2244 ? btb_bank0_rd_data_way0_out_66 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2945 = _T_2944 | _T_2690; // @[Mux.scala 27:72]
  wire  _T_2246 = btb_rd_addr_f == 8'h43; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_67; // @[lib.scala 374:16]
  wire [21:0] _T_2691 = _T_2246 ? btb_bank0_rd_data_way0_out_67 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2946 = _T_2945 | _T_2691; // @[Mux.scala 27:72]
  wire  _T_2248 = btb_rd_addr_f == 8'h44; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_68; // @[lib.scala 374:16]
  wire [21:0] _T_2692 = _T_2248 ? btb_bank0_rd_data_way0_out_68 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2947 = _T_2946 | _T_2692; // @[Mux.scala 27:72]
  wire  _T_2250 = btb_rd_addr_f == 8'h45; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_69; // @[lib.scala 374:16]
  wire [21:0] _T_2693 = _T_2250 ? btb_bank0_rd_data_way0_out_69 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2948 = _T_2947 | _T_2693; // @[Mux.scala 27:72]
  wire  _T_2252 = btb_rd_addr_f == 8'h46; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_70; // @[lib.scala 374:16]
  wire [21:0] _T_2694 = _T_2252 ? btb_bank0_rd_data_way0_out_70 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2949 = _T_2948 | _T_2694; // @[Mux.scala 27:72]
  wire  _T_2254 = btb_rd_addr_f == 8'h47; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_71; // @[lib.scala 374:16]
  wire [21:0] _T_2695 = _T_2254 ? btb_bank0_rd_data_way0_out_71 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2950 = _T_2949 | _T_2695; // @[Mux.scala 27:72]
  wire  _T_2256 = btb_rd_addr_f == 8'h48; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_72; // @[lib.scala 374:16]
  wire [21:0] _T_2696 = _T_2256 ? btb_bank0_rd_data_way0_out_72 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2951 = _T_2950 | _T_2696; // @[Mux.scala 27:72]
  wire  _T_2258 = btb_rd_addr_f == 8'h49; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_73; // @[lib.scala 374:16]
  wire [21:0] _T_2697 = _T_2258 ? btb_bank0_rd_data_way0_out_73 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2952 = _T_2951 | _T_2697; // @[Mux.scala 27:72]
  wire  _T_2260 = btb_rd_addr_f == 8'h4a; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_74; // @[lib.scala 374:16]
  wire [21:0] _T_2698 = _T_2260 ? btb_bank0_rd_data_way0_out_74 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2953 = _T_2952 | _T_2698; // @[Mux.scala 27:72]
  wire  _T_2262 = btb_rd_addr_f == 8'h4b; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_75; // @[lib.scala 374:16]
  wire [21:0] _T_2699 = _T_2262 ? btb_bank0_rd_data_way0_out_75 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2954 = _T_2953 | _T_2699; // @[Mux.scala 27:72]
  wire  _T_2264 = btb_rd_addr_f == 8'h4c; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_76; // @[lib.scala 374:16]
  wire [21:0] _T_2700 = _T_2264 ? btb_bank0_rd_data_way0_out_76 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2955 = _T_2954 | _T_2700; // @[Mux.scala 27:72]
  wire  _T_2266 = btb_rd_addr_f == 8'h4d; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_77; // @[lib.scala 374:16]
  wire [21:0] _T_2701 = _T_2266 ? btb_bank0_rd_data_way0_out_77 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2956 = _T_2955 | _T_2701; // @[Mux.scala 27:72]
  wire  _T_2268 = btb_rd_addr_f == 8'h4e; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_78; // @[lib.scala 374:16]
  wire [21:0] _T_2702 = _T_2268 ? btb_bank0_rd_data_way0_out_78 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2957 = _T_2956 | _T_2702; // @[Mux.scala 27:72]
  wire  _T_2270 = btb_rd_addr_f == 8'h4f; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_79; // @[lib.scala 374:16]
  wire [21:0] _T_2703 = _T_2270 ? btb_bank0_rd_data_way0_out_79 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2958 = _T_2957 | _T_2703; // @[Mux.scala 27:72]
  wire  _T_2272 = btb_rd_addr_f == 8'h50; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_80; // @[lib.scala 374:16]
  wire [21:0] _T_2704 = _T_2272 ? btb_bank0_rd_data_way0_out_80 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2959 = _T_2958 | _T_2704; // @[Mux.scala 27:72]
  wire  _T_2274 = btb_rd_addr_f == 8'h51; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_81; // @[lib.scala 374:16]
  wire [21:0] _T_2705 = _T_2274 ? btb_bank0_rd_data_way0_out_81 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2960 = _T_2959 | _T_2705; // @[Mux.scala 27:72]
  wire  _T_2276 = btb_rd_addr_f == 8'h52; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_82; // @[lib.scala 374:16]
  wire [21:0] _T_2706 = _T_2276 ? btb_bank0_rd_data_way0_out_82 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2961 = _T_2960 | _T_2706; // @[Mux.scala 27:72]
  wire  _T_2278 = btb_rd_addr_f == 8'h53; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_83; // @[lib.scala 374:16]
  wire [21:0] _T_2707 = _T_2278 ? btb_bank0_rd_data_way0_out_83 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2962 = _T_2961 | _T_2707; // @[Mux.scala 27:72]
  wire  _T_2280 = btb_rd_addr_f == 8'h54; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_84; // @[lib.scala 374:16]
  wire [21:0] _T_2708 = _T_2280 ? btb_bank0_rd_data_way0_out_84 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2963 = _T_2962 | _T_2708; // @[Mux.scala 27:72]
  wire  _T_2282 = btb_rd_addr_f == 8'h55; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_85; // @[lib.scala 374:16]
  wire [21:0] _T_2709 = _T_2282 ? btb_bank0_rd_data_way0_out_85 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2964 = _T_2963 | _T_2709; // @[Mux.scala 27:72]
  wire  _T_2284 = btb_rd_addr_f == 8'h56; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_86; // @[lib.scala 374:16]
  wire [21:0] _T_2710 = _T_2284 ? btb_bank0_rd_data_way0_out_86 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2965 = _T_2964 | _T_2710; // @[Mux.scala 27:72]
  wire  _T_2286 = btb_rd_addr_f == 8'h57; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_87; // @[lib.scala 374:16]
  wire [21:0] _T_2711 = _T_2286 ? btb_bank0_rd_data_way0_out_87 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2966 = _T_2965 | _T_2711; // @[Mux.scala 27:72]
  wire  _T_2288 = btb_rd_addr_f == 8'h58; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_88; // @[lib.scala 374:16]
  wire [21:0] _T_2712 = _T_2288 ? btb_bank0_rd_data_way0_out_88 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2967 = _T_2966 | _T_2712; // @[Mux.scala 27:72]
  wire  _T_2290 = btb_rd_addr_f == 8'h59; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_89; // @[lib.scala 374:16]
  wire [21:0] _T_2713 = _T_2290 ? btb_bank0_rd_data_way0_out_89 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2968 = _T_2967 | _T_2713; // @[Mux.scala 27:72]
  wire  _T_2292 = btb_rd_addr_f == 8'h5a; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_90; // @[lib.scala 374:16]
  wire [21:0] _T_2714 = _T_2292 ? btb_bank0_rd_data_way0_out_90 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2969 = _T_2968 | _T_2714; // @[Mux.scala 27:72]
  wire  _T_2294 = btb_rd_addr_f == 8'h5b; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_91; // @[lib.scala 374:16]
  wire [21:0] _T_2715 = _T_2294 ? btb_bank0_rd_data_way0_out_91 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2970 = _T_2969 | _T_2715; // @[Mux.scala 27:72]
  wire  _T_2296 = btb_rd_addr_f == 8'h5c; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_92; // @[lib.scala 374:16]
  wire [21:0] _T_2716 = _T_2296 ? btb_bank0_rd_data_way0_out_92 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2971 = _T_2970 | _T_2716; // @[Mux.scala 27:72]
  wire  _T_2298 = btb_rd_addr_f == 8'h5d; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_93; // @[lib.scala 374:16]
  wire [21:0] _T_2717 = _T_2298 ? btb_bank0_rd_data_way0_out_93 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2972 = _T_2971 | _T_2717; // @[Mux.scala 27:72]
  wire  _T_2300 = btb_rd_addr_f == 8'h5e; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_94; // @[lib.scala 374:16]
  wire [21:0] _T_2718 = _T_2300 ? btb_bank0_rd_data_way0_out_94 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2973 = _T_2972 | _T_2718; // @[Mux.scala 27:72]
  wire  _T_2302 = btb_rd_addr_f == 8'h5f; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_95; // @[lib.scala 374:16]
  wire [21:0] _T_2719 = _T_2302 ? btb_bank0_rd_data_way0_out_95 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2974 = _T_2973 | _T_2719; // @[Mux.scala 27:72]
  wire  _T_2304 = btb_rd_addr_f == 8'h60; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_96; // @[lib.scala 374:16]
  wire [21:0] _T_2720 = _T_2304 ? btb_bank0_rd_data_way0_out_96 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2975 = _T_2974 | _T_2720; // @[Mux.scala 27:72]
  wire  _T_2306 = btb_rd_addr_f == 8'h61; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_97; // @[lib.scala 374:16]
  wire [21:0] _T_2721 = _T_2306 ? btb_bank0_rd_data_way0_out_97 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2976 = _T_2975 | _T_2721; // @[Mux.scala 27:72]
  wire  _T_2308 = btb_rd_addr_f == 8'h62; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_98; // @[lib.scala 374:16]
  wire [21:0] _T_2722 = _T_2308 ? btb_bank0_rd_data_way0_out_98 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2977 = _T_2976 | _T_2722; // @[Mux.scala 27:72]
  wire  _T_2310 = btb_rd_addr_f == 8'h63; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_99; // @[lib.scala 374:16]
  wire [21:0] _T_2723 = _T_2310 ? btb_bank0_rd_data_way0_out_99 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2978 = _T_2977 | _T_2723; // @[Mux.scala 27:72]
  wire  _T_2312 = btb_rd_addr_f == 8'h64; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_100; // @[lib.scala 374:16]
  wire [21:0] _T_2724 = _T_2312 ? btb_bank0_rd_data_way0_out_100 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2979 = _T_2978 | _T_2724; // @[Mux.scala 27:72]
  wire  _T_2314 = btb_rd_addr_f == 8'h65; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_101; // @[lib.scala 374:16]
  wire [21:0] _T_2725 = _T_2314 ? btb_bank0_rd_data_way0_out_101 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2980 = _T_2979 | _T_2725; // @[Mux.scala 27:72]
  wire  _T_2316 = btb_rd_addr_f == 8'h66; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_102; // @[lib.scala 374:16]
  wire [21:0] _T_2726 = _T_2316 ? btb_bank0_rd_data_way0_out_102 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2981 = _T_2980 | _T_2726; // @[Mux.scala 27:72]
  wire  _T_2318 = btb_rd_addr_f == 8'h67; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_103; // @[lib.scala 374:16]
  wire [21:0] _T_2727 = _T_2318 ? btb_bank0_rd_data_way0_out_103 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2982 = _T_2981 | _T_2727; // @[Mux.scala 27:72]
  wire  _T_2320 = btb_rd_addr_f == 8'h68; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_104; // @[lib.scala 374:16]
  wire [21:0] _T_2728 = _T_2320 ? btb_bank0_rd_data_way0_out_104 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2983 = _T_2982 | _T_2728; // @[Mux.scala 27:72]
  wire  _T_2322 = btb_rd_addr_f == 8'h69; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_105; // @[lib.scala 374:16]
  wire [21:0] _T_2729 = _T_2322 ? btb_bank0_rd_data_way0_out_105 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2984 = _T_2983 | _T_2729; // @[Mux.scala 27:72]
  wire  _T_2324 = btb_rd_addr_f == 8'h6a; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_106; // @[lib.scala 374:16]
  wire [21:0] _T_2730 = _T_2324 ? btb_bank0_rd_data_way0_out_106 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2985 = _T_2984 | _T_2730; // @[Mux.scala 27:72]
  wire  _T_2326 = btb_rd_addr_f == 8'h6b; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_107; // @[lib.scala 374:16]
  wire [21:0] _T_2731 = _T_2326 ? btb_bank0_rd_data_way0_out_107 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2986 = _T_2985 | _T_2731; // @[Mux.scala 27:72]
  wire  _T_2328 = btb_rd_addr_f == 8'h6c; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_108; // @[lib.scala 374:16]
  wire [21:0] _T_2732 = _T_2328 ? btb_bank0_rd_data_way0_out_108 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2987 = _T_2986 | _T_2732; // @[Mux.scala 27:72]
  wire  _T_2330 = btb_rd_addr_f == 8'h6d; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_109; // @[lib.scala 374:16]
  wire [21:0] _T_2733 = _T_2330 ? btb_bank0_rd_data_way0_out_109 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2988 = _T_2987 | _T_2733; // @[Mux.scala 27:72]
  wire  _T_2332 = btb_rd_addr_f == 8'h6e; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_110; // @[lib.scala 374:16]
  wire [21:0] _T_2734 = _T_2332 ? btb_bank0_rd_data_way0_out_110 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2989 = _T_2988 | _T_2734; // @[Mux.scala 27:72]
  wire  _T_2334 = btb_rd_addr_f == 8'h6f; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_111; // @[lib.scala 374:16]
  wire [21:0] _T_2735 = _T_2334 ? btb_bank0_rd_data_way0_out_111 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2990 = _T_2989 | _T_2735; // @[Mux.scala 27:72]
  wire  _T_2336 = btb_rd_addr_f == 8'h70; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_112; // @[lib.scala 374:16]
  wire [21:0] _T_2736 = _T_2336 ? btb_bank0_rd_data_way0_out_112 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2991 = _T_2990 | _T_2736; // @[Mux.scala 27:72]
  wire  _T_2338 = btb_rd_addr_f == 8'h71; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_113; // @[lib.scala 374:16]
  wire [21:0] _T_2737 = _T_2338 ? btb_bank0_rd_data_way0_out_113 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2992 = _T_2991 | _T_2737; // @[Mux.scala 27:72]
  wire  _T_2340 = btb_rd_addr_f == 8'h72; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_114; // @[lib.scala 374:16]
  wire [21:0] _T_2738 = _T_2340 ? btb_bank0_rd_data_way0_out_114 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2993 = _T_2992 | _T_2738; // @[Mux.scala 27:72]
  wire  _T_2342 = btb_rd_addr_f == 8'h73; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_115; // @[lib.scala 374:16]
  wire [21:0] _T_2739 = _T_2342 ? btb_bank0_rd_data_way0_out_115 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2994 = _T_2993 | _T_2739; // @[Mux.scala 27:72]
  wire  _T_2344 = btb_rd_addr_f == 8'h74; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_116; // @[lib.scala 374:16]
  wire [21:0] _T_2740 = _T_2344 ? btb_bank0_rd_data_way0_out_116 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2995 = _T_2994 | _T_2740; // @[Mux.scala 27:72]
  wire  _T_2346 = btb_rd_addr_f == 8'h75; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_117; // @[lib.scala 374:16]
  wire [21:0] _T_2741 = _T_2346 ? btb_bank0_rd_data_way0_out_117 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2996 = _T_2995 | _T_2741; // @[Mux.scala 27:72]
  wire  _T_2348 = btb_rd_addr_f == 8'h76; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_118; // @[lib.scala 374:16]
  wire [21:0] _T_2742 = _T_2348 ? btb_bank0_rd_data_way0_out_118 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2997 = _T_2996 | _T_2742; // @[Mux.scala 27:72]
  wire  _T_2350 = btb_rd_addr_f == 8'h77; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_119; // @[lib.scala 374:16]
  wire [21:0] _T_2743 = _T_2350 ? btb_bank0_rd_data_way0_out_119 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2998 = _T_2997 | _T_2743; // @[Mux.scala 27:72]
  wire  _T_2352 = btb_rd_addr_f == 8'h78; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_120; // @[lib.scala 374:16]
  wire [21:0] _T_2744 = _T_2352 ? btb_bank0_rd_data_way0_out_120 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2999 = _T_2998 | _T_2744; // @[Mux.scala 27:72]
  wire  _T_2354 = btb_rd_addr_f == 8'h79; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_121; // @[lib.scala 374:16]
  wire [21:0] _T_2745 = _T_2354 ? btb_bank0_rd_data_way0_out_121 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3000 = _T_2999 | _T_2745; // @[Mux.scala 27:72]
  wire  _T_2356 = btb_rd_addr_f == 8'h7a; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_122; // @[lib.scala 374:16]
  wire [21:0] _T_2746 = _T_2356 ? btb_bank0_rd_data_way0_out_122 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3001 = _T_3000 | _T_2746; // @[Mux.scala 27:72]
  wire  _T_2358 = btb_rd_addr_f == 8'h7b; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_123; // @[lib.scala 374:16]
  wire [21:0] _T_2747 = _T_2358 ? btb_bank0_rd_data_way0_out_123 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3002 = _T_3001 | _T_2747; // @[Mux.scala 27:72]
  wire  _T_2360 = btb_rd_addr_f == 8'h7c; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_124; // @[lib.scala 374:16]
  wire [21:0] _T_2748 = _T_2360 ? btb_bank0_rd_data_way0_out_124 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3003 = _T_3002 | _T_2748; // @[Mux.scala 27:72]
  wire  _T_2362 = btb_rd_addr_f == 8'h7d; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_125; // @[lib.scala 374:16]
  wire [21:0] _T_2749 = _T_2362 ? btb_bank0_rd_data_way0_out_125 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3004 = _T_3003 | _T_2749; // @[Mux.scala 27:72]
  wire  _T_2364 = btb_rd_addr_f == 8'h7e; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_126; // @[lib.scala 374:16]
  wire [21:0] _T_2750 = _T_2364 ? btb_bank0_rd_data_way0_out_126 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3005 = _T_3004 | _T_2750; // @[Mux.scala 27:72]
  wire  _T_2366 = btb_rd_addr_f == 8'h7f; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_127; // @[lib.scala 374:16]
  wire [21:0] _T_2751 = _T_2366 ? btb_bank0_rd_data_way0_out_127 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3006 = _T_3005 | _T_2751; // @[Mux.scala 27:72]
  wire  _T_2368 = btb_rd_addr_f == 8'h80; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_128; // @[lib.scala 374:16]
  wire [21:0] _T_2752 = _T_2368 ? btb_bank0_rd_data_way0_out_128 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3007 = _T_3006 | _T_2752; // @[Mux.scala 27:72]
  wire  _T_2370 = btb_rd_addr_f == 8'h81; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_129; // @[lib.scala 374:16]
  wire [21:0] _T_2753 = _T_2370 ? btb_bank0_rd_data_way0_out_129 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3008 = _T_3007 | _T_2753; // @[Mux.scala 27:72]
  wire  _T_2372 = btb_rd_addr_f == 8'h82; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_130; // @[lib.scala 374:16]
  wire [21:0] _T_2754 = _T_2372 ? btb_bank0_rd_data_way0_out_130 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3009 = _T_3008 | _T_2754; // @[Mux.scala 27:72]
  wire  _T_2374 = btb_rd_addr_f == 8'h83; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_131; // @[lib.scala 374:16]
  wire [21:0] _T_2755 = _T_2374 ? btb_bank0_rd_data_way0_out_131 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3010 = _T_3009 | _T_2755; // @[Mux.scala 27:72]
  wire  _T_2376 = btb_rd_addr_f == 8'h84; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_132; // @[lib.scala 374:16]
  wire [21:0] _T_2756 = _T_2376 ? btb_bank0_rd_data_way0_out_132 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3011 = _T_3010 | _T_2756; // @[Mux.scala 27:72]
  wire  _T_2378 = btb_rd_addr_f == 8'h85; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_133; // @[lib.scala 374:16]
  wire [21:0] _T_2757 = _T_2378 ? btb_bank0_rd_data_way0_out_133 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3012 = _T_3011 | _T_2757; // @[Mux.scala 27:72]
  wire  _T_2380 = btb_rd_addr_f == 8'h86; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_134; // @[lib.scala 374:16]
  wire [21:0] _T_2758 = _T_2380 ? btb_bank0_rd_data_way0_out_134 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3013 = _T_3012 | _T_2758; // @[Mux.scala 27:72]
  wire  _T_2382 = btb_rd_addr_f == 8'h87; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_135; // @[lib.scala 374:16]
  wire [21:0] _T_2759 = _T_2382 ? btb_bank0_rd_data_way0_out_135 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3014 = _T_3013 | _T_2759; // @[Mux.scala 27:72]
  wire  _T_2384 = btb_rd_addr_f == 8'h88; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_136; // @[lib.scala 374:16]
  wire [21:0] _T_2760 = _T_2384 ? btb_bank0_rd_data_way0_out_136 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3015 = _T_3014 | _T_2760; // @[Mux.scala 27:72]
  wire  _T_2386 = btb_rd_addr_f == 8'h89; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_137; // @[lib.scala 374:16]
  wire [21:0] _T_2761 = _T_2386 ? btb_bank0_rd_data_way0_out_137 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3016 = _T_3015 | _T_2761; // @[Mux.scala 27:72]
  wire  _T_2388 = btb_rd_addr_f == 8'h8a; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_138; // @[lib.scala 374:16]
  wire [21:0] _T_2762 = _T_2388 ? btb_bank0_rd_data_way0_out_138 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3017 = _T_3016 | _T_2762; // @[Mux.scala 27:72]
  wire  _T_2390 = btb_rd_addr_f == 8'h8b; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_139; // @[lib.scala 374:16]
  wire [21:0] _T_2763 = _T_2390 ? btb_bank0_rd_data_way0_out_139 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3018 = _T_3017 | _T_2763; // @[Mux.scala 27:72]
  wire  _T_2392 = btb_rd_addr_f == 8'h8c; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_140; // @[lib.scala 374:16]
  wire [21:0] _T_2764 = _T_2392 ? btb_bank0_rd_data_way0_out_140 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3019 = _T_3018 | _T_2764; // @[Mux.scala 27:72]
  wire  _T_2394 = btb_rd_addr_f == 8'h8d; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_141; // @[lib.scala 374:16]
  wire [21:0] _T_2765 = _T_2394 ? btb_bank0_rd_data_way0_out_141 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3020 = _T_3019 | _T_2765; // @[Mux.scala 27:72]
  wire  _T_2396 = btb_rd_addr_f == 8'h8e; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_142; // @[lib.scala 374:16]
  wire [21:0] _T_2766 = _T_2396 ? btb_bank0_rd_data_way0_out_142 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3021 = _T_3020 | _T_2766; // @[Mux.scala 27:72]
  wire  _T_2398 = btb_rd_addr_f == 8'h8f; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_143; // @[lib.scala 374:16]
  wire [21:0] _T_2767 = _T_2398 ? btb_bank0_rd_data_way0_out_143 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3022 = _T_3021 | _T_2767; // @[Mux.scala 27:72]
  wire  _T_2400 = btb_rd_addr_f == 8'h90; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_144; // @[lib.scala 374:16]
  wire [21:0] _T_2768 = _T_2400 ? btb_bank0_rd_data_way0_out_144 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3023 = _T_3022 | _T_2768; // @[Mux.scala 27:72]
  wire  _T_2402 = btb_rd_addr_f == 8'h91; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_145; // @[lib.scala 374:16]
  wire [21:0] _T_2769 = _T_2402 ? btb_bank0_rd_data_way0_out_145 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3024 = _T_3023 | _T_2769; // @[Mux.scala 27:72]
  wire  _T_2404 = btb_rd_addr_f == 8'h92; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_146; // @[lib.scala 374:16]
  wire [21:0] _T_2770 = _T_2404 ? btb_bank0_rd_data_way0_out_146 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3025 = _T_3024 | _T_2770; // @[Mux.scala 27:72]
  wire  _T_2406 = btb_rd_addr_f == 8'h93; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_147; // @[lib.scala 374:16]
  wire [21:0] _T_2771 = _T_2406 ? btb_bank0_rd_data_way0_out_147 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3026 = _T_3025 | _T_2771; // @[Mux.scala 27:72]
  wire  _T_2408 = btb_rd_addr_f == 8'h94; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_148; // @[lib.scala 374:16]
  wire [21:0] _T_2772 = _T_2408 ? btb_bank0_rd_data_way0_out_148 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3027 = _T_3026 | _T_2772; // @[Mux.scala 27:72]
  wire  _T_2410 = btb_rd_addr_f == 8'h95; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_149; // @[lib.scala 374:16]
  wire [21:0] _T_2773 = _T_2410 ? btb_bank0_rd_data_way0_out_149 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3028 = _T_3027 | _T_2773; // @[Mux.scala 27:72]
  wire  _T_2412 = btb_rd_addr_f == 8'h96; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_150; // @[lib.scala 374:16]
  wire [21:0] _T_2774 = _T_2412 ? btb_bank0_rd_data_way0_out_150 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3029 = _T_3028 | _T_2774; // @[Mux.scala 27:72]
  wire  _T_2414 = btb_rd_addr_f == 8'h97; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_151; // @[lib.scala 374:16]
  wire [21:0] _T_2775 = _T_2414 ? btb_bank0_rd_data_way0_out_151 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3030 = _T_3029 | _T_2775; // @[Mux.scala 27:72]
  wire  _T_2416 = btb_rd_addr_f == 8'h98; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_152; // @[lib.scala 374:16]
  wire [21:0] _T_2776 = _T_2416 ? btb_bank0_rd_data_way0_out_152 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3031 = _T_3030 | _T_2776; // @[Mux.scala 27:72]
  wire  _T_2418 = btb_rd_addr_f == 8'h99; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_153; // @[lib.scala 374:16]
  wire [21:0] _T_2777 = _T_2418 ? btb_bank0_rd_data_way0_out_153 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3032 = _T_3031 | _T_2777; // @[Mux.scala 27:72]
  wire  _T_2420 = btb_rd_addr_f == 8'h9a; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_154; // @[lib.scala 374:16]
  wire [21:0] _T_2778 = _T_2420 ? btb_bank0_rd_data_way0_out_154 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3033 = _T_3032 | _T_2778; // @[Mux.scala 27:72]
  wire  _T_2422 = btb_rd_addr_f == 8'h9b; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_155; // @[lib.scala 374:16]
  wire [21:0] _T_2779 = _T_2422 ? btb_bank0_rd_data_way0_out_155 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3034 = _T_3033 | _T_2779; // @[Mux.scala 27:72]
  wire  _T_2424 = btb_rd_addr_f == 8'h9c; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_156; // @[lib.scala 374:16]
  wire [21:0] _T_2780 = _T_2424 ? btb_bank0_rd_data_way0_out_156 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3035 = _T_3034 | _T_2780; // @[Mux.scala 27:72]
  wire  _T_2426 = btb_rd_addr_f == 8'h9d; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_157; // @[lib.scala 374:16]
  wire [21:0] _T_2781 = _T_2426 ? btb_bank0_rd_data_way0_out_157 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3036 = _T_3035 | _T_2781; // @[Mux.scala 27:72]
  wire  _T_2428 = btb_rd_addr_f == 8'h9e; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_158; // @[lib.scala 374:16]
  wire [21:0] _T_2782 = _T_2428 ? btb_bank0_rd_data_way0_out_158 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3037 = _T_3036 | _T_2782; // @[Mux.scala 27:72]
  wire  _T_2430 = btb_rd_addr_f == 8'h9f; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_159; // @[lib.scala 374:16]
  wire [21:0] _T_2783 = _T_2430 ? btb_bank0_rd_data_way0_out_159 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3038 = _T_3037 | _T_2783; // @[Mux.scala 27:72]
  wire  _T_2432 = btb_rd_addr_f == 8'ha0; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_160; // @[lib.scala 374:16]
  wire [21:0] _T_2784 = _T_2432 ? btb_bank0_rd_data_way0_out_160 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3039 = _T_3038 | _T_2784; // @[Mux.scala 27:72]
  wire  _T_2434 = btb_rd_addr_f == 8'ha1; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_161; // @[lib.scala 374:16]
  wire [21:0] _T_2785 = _T_2434 ? btb_bank0_rd_data_way0_out_161 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3040 = _T_3039 | _T_2785; // @[Mux.scala 27:72]
  wire  _T_2436 = btb_rd_addr_f == 8'ha2; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_162; // @[lib.scala 374:16]
  wire [21:0] _T_2786 = _T_2436 ? btb_bank0_rd_data_way0_out_162 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3041 = _T_3040 | _T_2786; // @[Mux.scala 27:72]
  wire  _T_2438 = btb_rd_addr_f == 8'ha3; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_163; // @[lib.scala 374:16]
  wire [21:0] _T_2787 = _T_2438 ? btb_bank0_rd_data_way0_out_163 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3042 = _T_3041 | _T_2787; // @[Mux.scala 27:72]
  wire  _T_2440 = btb_rd_addr_f == 8'ha4; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_164; // @[lib.scala 374:16]
  wire [21:0] _T_2788 = _T_2440 ? btb_bank0_rd_data_way0_out_164 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3043 = _T_3042 | _T_2788; // @[Mux.scala 27:72]
  wire  _T_2442 = btb_rd_addr_f == 8'ha5; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_165; // @[lib.scala 374:16]
  wire [21:0] _T_2789 = _T_2442 ? btb_bank0_rd_data_way0_out_165 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3044 = _T_3043 | _T_2789; // @[Mux.scala 27:72]
  wire  _T_2444 = btb_rd_addr_f == 8'ha6; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_166; // @[lib.scala 374:16]
  wire [21:0] _T_2790 = _T_2444 ? btb_bank0_rd_data_way0_out_166 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3045 = _T_3044 | _T_2790; // @[Mux.scala 27:72]
  wire  _T_2446 = btb_rd_addr_f == 8'ha7; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_167; // @[lib.scala 374:16]
  wire [21:0] _T_2791 = _T_2446 ? btb_bank0_rd_data_way0_out_167 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3046 = _T_3045 | _T_2791; // @[Mux.scala 27:72]
  wire  _T_2448 = btb_rd_addr_f == 8'ha8; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_168; // @[lib.scala 374:16]
  wire [21:0] _T_2792 = _T_2448 ? btb_bank0_rd_data_way0_out_168 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3047 = _T_3046 | _T_2792; // @[Mux.scala 27:72]
  wire  _T_2450 = btb_rd_addr_f == 8'ha9; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_169; // @[lib.scala 374:16]
  wire [21:0] _T_2793 = _T_2450 ? btb_bank0_rd_data_way0_out_169 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3048 = _T_3047 | _T_2793; // @[Mux.scala 27:72]
  wire  _T_2452 = btb_rd_addr_f == 8'haa; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_170; // @[lib.scala 374:16]
  wire [21:0] _T_2794 = _T_2452 ? btb_bank0_rd_data_way0_out_170 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3049 = _T_3048 | _T_2794; // @[Mux.scala 27:72]
  wire  _T_2454 = btb_rd_addr_f == 8'hab; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_171; // @[lib.scala 374:16]
  wire [21:0] _T_2795 = _T_2454 ? btb_bank0_rd_data_way0_out_171 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3050 = _T_3049 | _T_2795; // @[Mux.scala 27:72]
  wire  _T_2456 = btb_rd_addr_f == 8'hac; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_172; // @[lib.scala 374:16]
  wire [21:0] _T_2796 = _T_2456 ? btb_bank0_rd_data_way0_out_172 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3051 = _T_3050 | _T_2796; // @[Mux.scala 27:72]
  wire  _T_2458 = btb_rd_addr_f == 8'had; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_173; // @[lib.scala 374:16]
  wire [21:0] _T_2797 = _T_2458 ? btb_bank0_rd_data_way0_out_173 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3052 = _T_3051 | _T_2797; // @[Mux.scala 27:72]
  wire  _T_2460 = btb_rd_addr_f == 8'hae; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_174; // @[lib.scala 374:16]
  wire [21:0] _T_2798 = _T_2460 ? btb_bank0_rd_data_way0_out_174 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3053 = _T_3052 | _T_2798; // @[Mux.scala 27:72]
  wire  _T_2462 = btb_rd_addr_f == 8'haf; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_175; // @[lib.scala 374:16]
  wire [21:0] _T_2799 = _T_2462 ? btb_bank0_rd_data_way0_out_175 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3054 = _T_3053 | _T_2799; // @[Mux.scala 27:72]
  wire  _T_2464 = btb_rd_addr_f == 8'hb0; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_176; // @[lib.scala 374:16]
  wire [21:0] _T_2800 = _T_2464 ? btb_bank0_rd_data_way0_out_176 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3055 = _T_3054 | _T_2800; // @[Mux.scala 27:72]
  wire  _T_2466 = btb_rd_addr_f == 8'hb1; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_177; // @[lib.scala 374:16]
  wire [21:0] _T_2801 = _T_2466 ? btb_bank0_rd_data_way0_out_177 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3056 = _T_3055 | _T_2801; // @[Mux.scala 27:72]
  wire  _T_2468 = btb_rd_addr_f == 8'hb2; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_178; // @[lib.scala 374:16]
  wire [21:0] _T_2802 = _T_2468 ? btb_bank0_rd_data_way0_out_178 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3057 = _T_3056 | _T_2802; // @[Mux.scala 27:72]
  wire  _T_2470 = btb_rd_addr_f == 8'hb3; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_179; // @[lib.scala 374:16]
  wire [21:0] _T_2803 = _T_2470 ? btb_bank0_rd_data_way0_out_179 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3058 = _T_3057 | _T_2803; // @[Mux.scala 27:72]
  wire  _T_2472 = btb_rd_addr_f == 8'hb4; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_180; // @[lib.scala 374:16]
  wire [21:0] _T_2804 = _T_2472 ? btb_bank0_rd_data_way0_out_180 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3059 = _T_3058 | _T_2804; // @[Mux.scala 27:72]
  wire  _T_2474 = btb_rd_addr_f == 8'hb5; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_181; // @[lib.scala 374:16]
  wire [21:0] _T_2805 = _T_2474 ? btb_bank0_rd_data_way0_out_181 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3060 = _T_3059 | _T_2805; // @[Mux.scala 27:72]
  wire  _T_2476 = btb_rd_addr_f == 8'hb6; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_182; // @[lib.scala 374:16]
  wire [21:0] _T_2806 = _T_2476 ? btb_bank0_rd_data_way0_out_182 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3061 = _T_3060 | _T_2806; // @[Mux.scala 27:72]
  wire  _T_2478 = btb_rd_addr_f == 8'hb7; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_183; // @[lib.scala 374:16]
  wire [21:0] _T_2807 = _T_2478 ? btb_bank0_rd_data_way0_out_183 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3062 = _T_3061 | _T_2807; // @[Mux.scala 27:72]
  wire  _T_2480 = btb_rd_addr_f == 8'hb8; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_184; // @[lib.scala 374:16]
  wire [21:0] _T_2808 = _T_2480 ? btb_bank0_rd_data_way0_out_184 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3063 = _T_3062 | _T_2808; // @[Mux.scala 27:72]
  wire  _T_2482 = btb_rd_addr_f == 8'hb9; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_185; // @[lib.scala 374:16]
  wire [21:0] _T_2809 = _T_2482 ? btb_bank0_rd_data_way0_out_185 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3064 = _T_3063 | _T_2809; // @[Mux.scala 27:72]
  wire  _T_2484 = btb_rd_addr_f == 8'hba; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_186; // @[lib.scala 374:16]
  wire [21:0] _T_2810 = _T_2484 ? btb_bank0_rd_data_way0_out_186 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3065 = _T_3064 | _T_2810; // @[Mux.scala 27:72]
  wire  _T_2486 = btb_rd_addr_f == 8'hbb; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_187; // @[lib.scala 374:16]
  wire [21:0] _T_2811 = _T_2486 ? btb_bank0_rd_data_way0_out_187 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3066 = _T_3065 | _T_2811; // @[Mux.scala 27:72]
  wire  _T_2488 = btb_rd_addr_f == 8'hbc; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_188; // @[lib.scala 374:16]
  wire [21:0] _T_2812 = _T_2488 ? btb_bank0_rd_data_way0_out_188 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3067 = _T_3066 | _T_2812; // @[Mux.scala 27:72]
  wire  _T_2490 = btb_rd_addr_f == 8'hbd; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_189; // @[lib.scala 374:16]
  wire [21:0] _T_2813 = _T_2490 ? btb_bank0_rd_data_way0_out_189 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3068 = _T_3067 | _T_2813; // @[Mux.scala 27:72]
  wire  _T_2492 = btb_rd_addr_f == 8'hbe; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_190; // @[lib.scala 374:16]
  wire [21:0] _T_2814 = _T_2492 ? btb_bank0_rd_data_way0_out_190 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3069 = _T_3068 | _T_2814; // @[Mux.scala 27:72]
  wire  _T_2494 = btb_rd_addr_f == 8'hbf; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_191; // @[lib.scala 374:16]
  wire [21:0] _T_2815 = _T_2494 ? btb_bank0_rd_data_way0_out_191 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3070 = _T_3069 | _T_2815; // @[Mux.scala 27:72]
  wire  _T_2496 = btb_rd_addr_f == 8'hc0; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_192; // @[lib.scala 374:16]
  wire [21:0] _T_2816 = _T_2496 ? btb_bank0_rd_data_way0_out_192 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3071 = _T_3070 | _T_2816; // @[Mux.scala 27:72]
  wire  _T_2498 = btb_rd_addr_f == 8'hc1; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_193; // @[lib.scala 374:16]
  wire [21:0] _T_2817 = _T_2498 ? btb_bank0_rd_data_way0_out_193 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3072 = _T_3071 | _T_2817; // @[Mux.scala 27:72]
  wire  _T_2500 = btb_rd_addr_f == 8'hc2; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_194; // @[lib.scala 374:16]
  wire [21:0] _T_2818 = _T_2500 ? btb_bank0_rd_data_way0_out_194 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3073 = _T_3072 | _T_2818; // @[Mux.scala 27:72]
  wire  _T_2502 = btb_rd_addr_f == 8'hc3; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_195; // @[lib.scala 374:16]
  wire [21:0] _T_2819 = _T_2502 ? btb_bank0_rd_data_way0_out_195 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3074 = _T_3073 | _T_2819; // @[Mux.scala 27:72]
  wire  _T_2504 = btb_rd_addr_f == 8'hc4; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_196; // @[lib.scala 374:16]
  wire [21:0] _T_2820 = _T_2504 ? btb_bank0_rd_data_way0_out_196 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3075 = _T_3074 | _T_2820; // @[Mux.scala 27:72]
  wire  _T_2506 = btb_rd_addr_f == 8'hc5; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_197; // @[lib.scala 374:16]
  wire [21:0] _T_2821 = _T_2506 ? btb_bank0_rd_data_way0_out_197 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3076 = _T_3075 | _T_2821; // @[Mux.scala 27:72]
  wire  _T_2508 = btb_rd_addr_f == 8'hc6; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_198; // @[lib.scala 374:16]
  wire [21:0] _T_2822 = _T_2508 ? btb_bank0_rd_data_way0_out_198 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3077 = _T_3076 | _T_2822; // @[Mux.scala 27:72]
  wire  _T_2510 = btb_rd_addr_f == 8'hc7; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_199; // @[lib.scala 374:16]
  wire [21:0] _T_2823 = _T_2510 ? btb_bank0_rd_data_way0_out_199 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3078 = _T_3077 | _T_2823; // @[Mux.scala 27:72]
  wire  _T_2512 = btb_rd_addr_f == 8'hc8; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_200; // @[lib.scala 374:16]
  wire [21:0] _T_2824 = _T_2512 ? btb_bank0_rd_data_way0_out_200 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3079 = _T_3078 | _T_2824; // @[Mux.scala 27:72]
  wire  _T_2514 = btb_rd_addr_f == 8'hc9; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_201; // @[lib.scala 374:16]
  wire [21:0] _T_2825 = _T_2514 ? btb_bank0_rd_data_way0_out_201 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3080 = _T_3079 | _T_2825; // @[Mux.scala 27:72]
  wire  _T_2516 = btb_rd_addr_f == 8'hca; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_202; // @[lib.scala 374:16]
  wire [21:0] _T_2826 = _T_2516 ? btb_bank0_rd_data_way0_out_202 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3081 = _T_3080 | _T_2826; // @[Mux.scala 27:72]
  wire  _T_2518 = btb_rd_addr_f == 8'hcb; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_203; // @[lib.scala 374:16]
  wire [21:0] _T_2827 = _T_2518 ? btb_bank0_rd_data_way0_out_203 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3082 = _T_3081 | _T_2827; // @[Mux.scala 27:72]
  wire  _T_2520 = btb_rd_addr_f == 8'hcc; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_204; // @[lib.scala 374:16]
  wire [21:0] _T_2828 = _T_2520 ? btb_bank0_rd_data_way0_out_204 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3083 = _T_3082 | _T_2828; // @[Mux.scala 27:72]
  wire  _T_2522 = btb_rd_addr_f == 8'hcd; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_205; // @[lib.scala 374:16]
  wire [21:0] _T_2829 = _T_2522 ? btb_bank0_rd_data_way0_out_205 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3084 = _T_3083 | _T_2829; // @[Mux.scala 27:72]
  wire  _T_2524 = btb_rd_addr_f == 8'hce; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_206; // @[lib.scala 374:16]
  wire [21:0] _T_2830 = _T_2524 ? btb_bank0_rd_data_way0_out_206 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3085 = _T_3084 | _T_2830; // @[Mux.scala 27:72]
  wire  _T_2526 = btb_rd_addr_f == 8'hcf; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_207; // @[lib.scala 374:16]
  wire [21:0] _T_2831 = _T_2526 ? btb_bank0_rd_data_way0_out_207 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3086 = _T_3085 | _T_2831; // @[Mux.scala 27:72]
  wire  _T_2528 = btb_rd_addr_f == 8'hd0; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_208; // @[lib.scala 374:16]
  wire [21:0] _T_2832 = _T_2528 ? btb_bank0_rd_data_way0_out_208 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3087 = _T_3086 | _T_2832; // @[Mux.scala 27:72]
  wire  _T_2530 = btb_rd_addr_f == 8'hd1; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_209; // @[lib.scala 374:16]
  wire [21:0] _T_2833 = _T_2530 ? btb_bank0_rd_data_way0_out_209 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3088 = _T_3087 | _T_2833; // @[Mux.scala 27:72]
  wire  _T_2532 = btb_rd_addr_f == 8'hd2; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_210; // @[lib.scala 374:16]
  wire [21:0] _T_2834 = _T_2532 ? btb_bank0_rd_data_way0_out_210 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3089 = _T_3088 | _T_2834; // @[Mux.scala 27:72]
  wire  _T_2534 = btb_rd_addr_f == 8'hd3; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_211; // @[lib.scala 374:16]
  wire [21:0] _T_2835 = _T_2534 ? btb_bank0_rd_data_way0_out_211 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3090 = _T_3089 | _T_2835; // @[Mux.scala 27:72]
  wire  _T_2536 = btb_rd_addr_f == 8'hd4; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_212; // @[lib.scala 374:16]
  wire [21:0] _T_2836 = _T_2536 ? btb_bank0_rd_data_way0_out_212 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3091 = _T_3090 | _T_2836; // @[Mux.scala 27:72]
  wire  _T_2538 = btb_rd_addr_f == 8'hd5; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_213; // @[lib.scala 374:16]
  wire [21:0] _T_2837 = _T_2538 ? btb_bank0_rd_data_way0_out_213 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3092 = _T_3091 | _T_2837; // @[Mux.scala 27:72]
  wire  _T_2540 = btb_rd_addr_f == 8'hd6; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_214; // @[lib.scala 374:16]
  wire [21:0] _T_2838 = _T_2540 ? btb_bank0_rd_data_way0_out_214 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3093 = _T_3092 | _T_2838; // @[Mux.scala 27:72]
  wire  _T_2542 = btb_rd_addr_f == 8'hd7; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_215; // @[lib.scala 374:16]
  wire [21:0] _T_2839 = _T_2542 ? btb_bank0_rd_data_way0_out_215 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3094 = _T_3093 | _T_2839; // @[Mux.scala 27:72]
  wire  _T_2544 = btb_rd_addr_f == 8'hd8; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_216; // @[lib.scala 374:16]
  wire [21:0] _T_2840 = _T_2544 ? btb_bank0_rd_data_way0_out_216 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3095 = _T_3094 | _T_2840; // @[Mux.scala 27:72]
  wire  _T_2546 = btb_rd_addr_f == 8'hd9; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_217; // @[lib.scala 374:16]
  wire [21:0] _T_2841 = _T_2546 ? btb_bank0_rd_data_way0_out_217 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3096 = _T_3095 | _T_2841; // @[Mux.scala 27:72]
  wire  _T_2548 = btb_rd_addr_f == 8'hda; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_218; // @[lib.scala 374:16]
  wire [21:0] _T_2842 = _T_2548 ? btb_bank0_rd_data_way0_out_218 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3097 = _T_3096 | _T_2842; // @[Mux.scala 27:72]
  wire  _T_2550 = btb_rd_addr_f == 8'hdb; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_219; // @[lib.scala 374:16]
  wire [21:0] _T_2843 = _T_2550 ? btb_bank0_rd_data_way0_out_219 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3098 = _T_3097 | _T_2843; // @[Mux.scala 27:72]
  wire  _T_2552 = btb_rd_addr_f == 8'hdc; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_220; // @[lib.scala 374:16]
  wire [21:0] _T_2844 = _T_2552 ? btb_bank0_rd_data_way0_out_220 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3099 = _T_3098 | _T_2844; // @[Mux.scala 27:72]
  wire  _T_2554 = btb_rd_addr_f == 8'hdd; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_221; // @[lib.scala 374:16]
  wire [21:0] _T_2845 = _T_2554 ? btb_bank0_rd_data_way0_out_221 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3100 = _T_3099 | _T_2845; // @[Mux.scala 27:72]
  wire  _T_2556 = btb_rd_addr_f == 8'hde; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_222; // @[lib.scala 374:16]
  wire [21:0] _T_2846 = _T_2556 ? btb_bank0_rd_data_way0_out_222 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3101 = _T_3100 | _T_2846; // @[Mux.scala 27:72]
  wire  _T_2558 = btb_rd_addr_f == 8'hdf; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_223; // @[lib.scala 374:16]
  wire [21:0] _T_2847 = _T_2558 ? btb_bank0_rd_data_way0_out_223 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3102 = _T_3101 | _T_2847; // @[Mux.scala 27:72]
  wire  _T_2560 = btb_rd_addr_f == 8'he0; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_224; // @[lib.scala 374:16]
  wire [21:0] _T_2848 = _T_2560 ? btb_bank0_rd_data_way0_out_224 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3103 = _T_3102 | _T_2848; // @[Mux.scala 27:72]
  wire  _T_2562 = btb_rd_addr_f == 8'he1; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_225; // @[lib.scala 374:16]
  wire [21:0] _T_2849 = _T_2562 ? btb_bank0_rd_data_way0_out_225 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3104 = _T_3103 | _T_2849; // @[Mux.scala 27:72]
  wire  _T_2564 = btb_rd_addr_f == 8'he2; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_226; // @[lib.scala 374:16]
  wire [21:0] _T_2850 = _T_2564 ? btb_bank0_rd_data_way0_out_226 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3105 = _T_3104 | _T_2850; // @[Mux.scala 27:72]
  wire  _T_2566 = btb_rd_addr_f == 8'he3; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_227; // @[lib.scala 374:16]
  wire [21:0] _T_2851 = _T_2566 ? btb_bank0_rd_data_way0_out_227 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3106 = _T_3105 | _T_2851; // @[Mux.scala 27:72]
  wire  _T_2568 = btb_rd_addr_f == 8'he4; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_228; // @[lib.scala 374:16]
  wire [21:0] _T_2852 = _T_2568 ? btb_bank0_rd_data_way0_out_228 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3107 = _T_3106 | _T_2852; // @[Mux.scala 27:72]
  wire  _T_2570 = btb_rd_addr_f == 8'he5; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_229; // @[lib.scala 374:16]
  wire [21:0] _T_2853 = _T_2570 ? btb_bank0_rd_data_way0_out_229 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3108 = _T_3107 | _T_2853; // @[Mux.scala 27:72]
  wire  _T_2572 = btb_rd_addr_f == 8'he6; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_230; // @[lib.scala 374:16]
  wire [21:0] _T_2854 = _T_2572 ? btb_bank0_rd_data_way0_out_230 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3109 = _T_3108 | _T_2854; // @[Mux.scala 27:72]
  wire  _T_2574 = btb_rd_addr_f == 8'he7; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_231; // @[lib.scala 374:16]
  wire [21:0] _T_2855 = _T_2574 ? btb_bank0_rd_data_way0_out_231 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3110 = _T_3109 | _T_2855; // @[Mux.scala 27:72]
  wire  _T_2576 = btb_rd_addr_f == 8'he8; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_232; // @[lib.scala 374:16]
  wire [21:0] _T_2856 = _T_2576 ? btb_bank0_rd_data_way0_out_232 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3111 = _T_3110 | _T_2856; // @[Mux.scala 27:72]
  wire  _T_2578 = btb_rd_addr_f == 8'he9; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_233; // @[lib.scala 374:16]
  wire [21:0] _T_2857 = _T_2578 ? btb_bank0_rd_data_way0_out_233 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3112 = _T_3111 | _T_2857; // @[Mux.scala 27:72]
  wire  _T_2580 = btb_rd_addr_f == 8'hea; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_234; // @[lib.scala 374:16]
  wire [21:0] _T_2858 = _T_2580 ? btb_bank0_rd_data_way0_out_234 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3113 = _T_3112 | _T_2858; // @[Mux.scala 27:72]
  wire  _T_2582 = btb_rd_addr_f == 8'heb; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_235; // @[lib.scala 374:16]
  wire [21:0] _T_2859 = _T_2582 ? btb_bank0_rd_data_way0_out_235 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3114 = _T_3113 | _T_2859; // @[Mux.scala 27:72]
  wire  _T_2584 = btb_rd_addr_f == 8'hec; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_236; // @[lib.scala 374:16]
  wire [21:0] _T_2860 = _T_2584 ? btb_bank0_rd_data_way0_out_236 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3115 = _T_3114 | _T_2860; // @[Mux.scala 27:72]
  wire  _T_2586 = btb_rd_addr_f == 8'hed; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_237; // @[lib.scala 374:16]
  wire [21:0] _T_2861 = _T_2586 ? btb_bank0_rd_data_way0_out_237 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3116 = _T_3115 | _T_2861; // @[Mux.scala 27:72]
  wire  _T_2588 = btb_rd_addr_f == 8'hee; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_238; // @[lib.scala 374:16]
  wire [21:0] _T_2862 = _T_2588 ? btb_bank0_rd_data_way0_out_238 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3117 = _T_3116 | _T_2862; // @[Mux.scala 27:72]
  wire  _T_2590 = btb_rd_addr_f == 8'hef; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_239; // @[lib.scala 374:16]
  wire [21:0] _T_2863 = _T_2590 ? btb_bank0_rd_data_way0_out_239 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3118 = _T_3117 | _T_2863; // @[Mux.scala 27:72]
  wire  _T_2592 = btb_rd_addr_f == 8'hf0; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_240; // @[lib.scala 374:16]
  wire [21:0] _T_2864 = _T_2592 ? btb_bank0_rd_data_way0_out_240 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3119 = _T_3118 | _T_2864; // @[Mux.scala 27:72]
  wire  _T_2594 = btb_rd_addr_f == 8'hf1; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_241; // @[lib.scala 374:16]
  wire [21:0] _T_2865 = _T_2594 ? btb_bank0_rd_data_way0_out_241 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3120 = _T_3119 | _T_2865; // @[Mux.scala 27:72]
  wire  _T_2596 = btb_rd_addr_f == 8'hf2; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_242; // @[lib.scala 374:16]
  wire [21:0] _T_2866 = _T_2596 ? btb_bank0_rd_data_way0_out_242 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3121 = _T_3120 | _T_2866; // @[Mux.scala 27:72]
  wire  _T_2598 = btb_rd_addr_f == 8'hf3; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_243; // @[lib.scala 374:16]
  wire [21:0] _T_2867 = _T_2598 ? btb_bank0_rd_data_way0_out_243 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3122 = _T_3121 | _T_2867; // @[Mux.scala 27:72]
  wire  _T_2600 = btb_rd_addr_f == 8'hf4; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_244; // @[lib.scala 374:16]
  wire [21:0] _T_2868 = _T_2600 ? btb_bank0_rd_data_way0_out_244 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3123 = _T_3122 | _T_2868; // @[Mux.scala 27:72]
  wire  _T_2602 = btb_rd_addr_f == 8'hf5; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_245; // @[lib.scala 374:16]
  wire [21:0] _T_2869 = _T_2602 ? btb_bank0_rd_data_way0_out_245 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3124 = _T_3123 | _T_2869; // @[Mux.scala 27:72]
  wire  _T_2604 = btb_rd_addr_f == 8'hf6; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_246; // @[lib.scala 374:16]
  wire [21:0] _T_2870 = _T_2604 ? btb_bank0_rd_data_way0_out_246 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3125 = _T_3124 | _T_2870; // @[Mux.scala 27:72]
  wire  _T_2606 = btb_rd_addr_f == 8'hf7; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_247; // @[lib.scala 374:16]
  wire [21:0] _T_2871 = _T_2606 ? btb_bank0_rd_data_way0_out_247 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3126 = _T_3125 | _T_2871; // @[Mux.scala 27:72]
  wire  _T_2608 = btb_rd_addr_f == 8'hf8; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_248; // @[lib.scala 374:16]
  wire [21:0] _T_2872 = _T_2608 ? btb_bank0_rd_data_way0_out_248 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3127 = _T_3126 | _T_2872; // @[Mux.scala 27:72]
  wire  _T_2610 = btb_rd_addr_f == 8'hf9; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_249; // @[lib.scala 374:16]
  wire [21:0] _T_2873 = _T_2610 ? btb_bank0_rd_data_way0_out_249 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3128 = _T_3127 | _T_2873; // @[Mux.scala 27:72]
  wire  _T_2612 = btb_rd_addr_f == 8'hfa; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_250; // @[lib.scala 374:16]
  wire [21:0] _T_2874 = _T_2612 ? btb_bank0_rd_data_way0_out_250 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3129 = _T_3128 | _T_2874; // @[Mux.scala 27:72]
  wire  _T_2614 = btb_rd_addr_f == 8'hfb; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_251; // @[lib.scala 374:16]
  wire [21:0] _T_2875 = _T_2614 ? btb_bank0_rd_data_way0_out_251 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3130 = _T_3129 | _T_2875; // @[Mux.scala 27:72]
  wire  _T_2616 = btb_rd_addr_f == 8'hfc; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_252; // @[lib.scala 374:16]
  wire [21:0] _T_2876 = _T_2616 ? btb_bank0_rd_data_way0_out_252 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3131 = _T_3130 | _T_2876; // @[Mux.scala 27:72]
  wire  _T_2618 = btb_rd_addr_f == 8'hfd; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_253; // @[lib.scala 374:16]
  wire [21:0] _T_2877 = _T_2618 ? btb_bank0_rd_data_way0_out_253 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3132 = _T_3131 | _T_2877; // @[Mux.scala 27:72]
  wire  _T_2620 = btb_rd_addr_f == 8'hfe; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_254; // @[lib.scala 374:16]
  wire [21:0] _T_2878 = _T_2620 ? btb_bank0_rd_data_way0_out_254 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3133 = _T_3132 | _T_2878; // @[Mux.scala 27:72]
  wire  _T_2622 = btb_rd_addr_f == 8'hff; // @[ifu_bp_ctl.scala 418:77]
  reg [21:0] btb_bank0_rd_data_way0_out_255; // @[lib.scala 374:16]
  wire [21:0] _T_2879 = _T_2622 ? btb_bank0_rd_data_way0_out_255 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] btb_bank0_rd_data_way0_f = _T_3133 | _T_2879; // @[Mux.scala 27:72]
  wire [4:0] _T_25 = io_ifc_fetch_addr_f[13:9] ^ io_ifc_fetch_addr_f[18:14]; // @[lib.scala 42:111]
  wire [4:0] fetch_rd_tag_f = _T_25 ^ io_ifc_fetch_addr_f[23:19]; // @[lib.scala 42:111]
  wire  _T_46 = btb_bank0_rd_data_way0_f[21:17] == fetch_rd_tag_f; // @[ifu_bp_ctl.scala 127:97]
  wire  _T_47 = btb_bank0_rd_data_way0_f[0] & _T_46; // @[ifu_bp_ctl.scala 127:55]
  reg  dec_tlu_way_wb_f; // @[ifu_bp_ctl.scala 118:59]
  wire  _T_19 = io_exu_bp_exu_i0_br_index_r == btb_rd_addr_f; // @[ifu_bp_ctl.scala 102:72]
  wire  branch_error_collision_f = dec_tlu_error_wb & _T_19; // @[ifu_bp_ctl.scala 102:51]
  wire  branch_error_bank_conflict_f = branch_error_collision_f & dec_tlu_error_wb; // @[ifu_bp_ctl.scala 106:63]
  wire  _T_48 = dec_tlu_way_wb_f & branch_error_bank_conflict_f; // @[ifu_bp_ctl.scala 128:44]
  wire  _T_49 = ~_T_48; // @[ifu_bp_ctl.scala 128:25]
  wire  _T_50 = _T_47 & _T_49; // @[ifu_bp_ctl.scala 127:117]
  wire  _T_51 = _T_50 & io_ifc_fetch_req_f; // @[ifu_bp_ctl.scala 128:76]
  wire  tag_match_way0_f = _T_51 & _T; // @[ifu_bp_ctl.scala 128:97]
  wire  _T_82 = btb_bank0_rd_data_way0_f[3] ^ btb_bank0_rd_data_way0_f[4]; // @[ifu_bp_ctl.scala 142:91]
  wire  _T_83 = tag_match_way0_f & _T_82; // @[ifu_bp_ctl.scala 142:56]
  wire  _T_87 = ~_T_82; // @[ifu_bp_ctl.scala 143:58]
  wire  _T_88 = tag_match_way0_f & _T_87; // @[ifu_bp_ctl.scala 143:56]
  wire [1:0] tag_match_way0_expanded_f = {_T_83,_T_88}; // @[Cat.scala 29:58]
  wire [21:0] _T_127 = tag_match_way0_expanded_f[1] ? btb_bank0_rd_data_way0_f : 22'h0; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_0; // @[lib.scala 374:16]
  wire [21:0] _T_3648 = _T_2112 ? btb_bank0_rd_data_way1_out_0 : 22'h0; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_1; // @[lib.scala 374:16]
  wire [21:0] _T_3649 = _T_2114 ? btb_bank0_rd_data_way1_out_1 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3904 = _T_3648 | _T_3649; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_2; // @[lib.scala 374:16]
  wire [21:0] _T_3650 = _T_2116 ? btb_bank0_rd_data_way1_out_2 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3905 = _T_3904 | _T_3650; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_3; // @[lib.scala 374:16]
  wire [21:0] _T_3651 = _T_2118 ? btb_bank0_rd_data_way1_out_3 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3906 = _T_3905 | _T_3651; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_4; // @[lib.scala 374:16]
  wire [21:0] _T_3652 = _T_2120 ? btb_bank0_rd_data_way1_out_4 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3907 = _T_3906 | _T_3652; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_5; // @[lib.scala 374:16]
  wire [21:0] _T_3653 = _T_2122 ? btb_bank0_rd_data_way1_out_5 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3908 = _T_3907 | _T_3653; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_6; // @[lib.scala 374:16]
  wire [21:0] _T_3654 = _T_2124 ? btb_bank0_rd_data_way1_out_6 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3909 = _T_3908 | _T_3654; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_7; // @[lib.scala 374:16]
  wire [21:0] _T_3655 = _T_2126 ? btb_bank0_rd_data_way1_out_7 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3910 = _T_3909 | _T_3655; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_8; // @[lib.scala 374:16]
  wire [21:0] _T_3656 = _T_2128 ? btb_bank0_rd_data_way1_out_8 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3911 = _T_3910 | _T_3656; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_9; // @[lib.scala 374:16]
  wire [21:0] _T_3657 = _T_2130 ? btb_bank0_rd_data_way1_out_9 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3912 = _T_3911 | _T_3657; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_10; // @[lib.scala 374:16]
  wire [21:0] _T_3658 = _T_2132 ? btb_bank0_rd_data_way1_out_10 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3913 = _T_3912 | _T_3658; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_11; // @[lib.scala 374:16]
  wire [21:0] _T_3659 = _T_2134 ? btb_bank0_rd_data_way1_out_11 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3914 = _T_3913 | _T_3659; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_12; // @[lib.scala 374:16]
  wire [21:0] _T_3660 = _T_2136 ? btb_bank0_rd_data_way1_out_12 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3915 = _T_3914 | _T_3660; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_13; // @[lib.scala 374:16]
  wire [21:0] _T_3661 = _T_2138 ? btb_bank0_rd_data_way1_out_13 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3916 = _T_3915 | _T_3661; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_14; // @[lib.scala 374:16]
  wire [21:0] _T_3662 = _T_2140 ? btb_bank0_rd_data_way1_out_14 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3917 = _T_3916 | _T_3662; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_15; // @[lib.scala 374:16]
  wire [21:0] _T_3663 = _T_2142 ? btb_bank0_rd_data_way1_out_15 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3918 = _T_3917 | _T_3663; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_16; // @[lib.scala 374:16]
  wire [21:0] _T_3664 = _T_2144 ? btb_bank0_rd_data_way1_out_16 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3919 = _T_3918 | _T_3664; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_17; // @[lib.scala 374:16]
  wire [21:0] _T_3665 = _T_2146 ? btb_bank0_rd_data_way1_out_17 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3920 = _T_3919 | _T_3665; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_18; // @[lib.scala 374:16]
  wire [21:0] _T_3666 = _T_2148 ? btb_bank0_rd_data_way1_out_18 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3921 = _T_3920 | _T_3666; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_19; // @[lib.scala 374:16]
  wire [21:0] _T_3667 = _T_2150 ? btb_bank0_rd_data_way1_out_19 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3922 = _T_3921 | _T_3667; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_20; // @[lib.scala 374:16]
  wire [21:0] _T_3668 = _T_2152 ? btb_bank0_rd_data_way1_out_20 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3923 = _T_3922 | _T_3668; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_21; // @[lib.scala 374:16]
  wire [21:0] _T_3669 = _T_2154 ? btb_bank0_rd_data_way1_out_21 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3924 = _T_3923 | _T_3669; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_22; // @[lib.scala 374:16]
  wire [21:0] _T_3670 = _T_2156 ? btb_bank0_rd_data_way1_out_22 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3925 = _T_3924 | _T_3670; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_23; // @[lib.scala 374:16]
  wire [21:0] _T_3671 = _T_2158 ? btb_bank0_rd_data_way1_out_23 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3926 = _T_3925 | _T_3671; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_24; // @[lib.scala 374:16]
  wire [21:0] _T_3672 = _T_2160 ? btb_bank0_rd_data_way1_out_24 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3927 = _T_3926 | _T_3672; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_25; // @[lib.scala 374:16]
  wire [21:0] _T_3673 = _T_2162 ? btb_bank0_rd_data_way1_out_25 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3928 = _T_3927 | _T_3673; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_26; // @[lib.scala 374:16]
  wire [21:0] _T_3674 = _T_2164 ? btb_bank0_rd_data_way1_out_26 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3929 = _T_3928 | _T_3674; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_27; // @[lib.scala 374:16]
  wire [21:0] _T_3675 = _T_2166 ? btb_bank0_rd_data_way1_out_27 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3930 = _T_3929 | _T_3675; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_28; // @[lib.scala 374:16]
  wire [21:0] _T_3676 = _T_2168 ? btb_bank0_rd_data_way1_out_28 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3931 = _T_3930 | _T_3676; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_29; // @[lib.scala 374:16]
  wire [21:0] _T_3677 = _T_2170 ? btb_bank0_rd_data_way1_out_29 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3932 = _T_3931 | _T_3677; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_30; // @[lib.scala 374:16]
  wire [21:0] _T_3678 = _T_2172 ? btb_bank0_rd_data_way1_out_30 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3933 = _T_3932 | _T_3678; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_31; // @[lib.scala 374:16]
  wire [21:0] _T_3679 = _T_2174 ? btb_bank0_rd_data_way1_out_31 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3934 = _T_3933 | _T_3679; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_32; // @[lib.scala 374:16]
  wire [21:0] _T_3680 = _T_2176 ? btb_bank0_rd_data_way1_out_32 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3935 = _T_3934 | _T_3680; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_33; // @[lib.scala 374:16]
  wire [21:0] _T_3681 = _T_2178 ? btb_bank0_rd_data_way1_out_33 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3936 = _T_3935 | _T_3681; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_34; // @[lib.scala 374:16]
  wire [21:0] _T_3682 = _T_2180 ? btb_bank0_rd_data_way1_out_34 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3937 = _T_3936 | _T_3682; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_35; // @[lib.scala 374:16]
  wire [21:0] _T_3683 = _T_2182 ? btb_bank0_rd_data_way1_out_35 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3938 = _T_3937 | _T_3683; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_36; // @[lib.scala 374:16]
  wire [21:0] _T_3684 = _T_2184 ? btb_bank0_rd_data_way1_out_36 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3939 = _T_3938 | _T_3684; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_37; // @[lib.scala 374:16]
  wire [21:0] _T_3685 = _T_2186 ? btb_bank0_rd_data_way1_out_37 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3940 = _T_3939 | _T_3685; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_38; // @[lib.scala 374:16]
  wire [21:0] _T_3686 = _T_2188 ? btb_bank0_rd_data_way1_out_38 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3941 = _T_3940 | _T_3686; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_39; // @[lib.scala 374:16]
  wire [21:0] _T_3687 = _T_2190 ? btb_bank0_rd_data_way1_out_39 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3942 = _T_3941 | _T_3687; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_40; // @[lib.scala 374:16]
  wire [21:0] _T_3688 = _T_2192 ? btb_bank0_rd_data_way1_out_40 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3943 = _T_3942 | _T_3688; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_41; // @[lib.scala 374:16]
  wire [21:0] _T_3689 = _T_2194 ? btb_bank0_rd_data_way1_out_41 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3944 = _T_3943 | _T_3689; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_42; // @[lib.scala 374:16]
  wire [21:0] _T_3690 = _T_2196 ? btb_bank0_rd_data_way1_out_42 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3945 = _T_3944 | _T_3690; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_43; // @[lib.scala 374:16]
  wire [21:0] _T_3691 = _T_2198 ? btb_bank0_rd_data_way1_out_43 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3946 = _T_3945 | _T_3691; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_44; // @[lib.scala 374:16]
  wire [21:0] _T_3692 = _T_2200 ? btb_bank0_rd_data_way1_out_44 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3947 = _T_3946 | _T_3692; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_45; // @[lib.scala 374:16]
  wire [21:0] _T_3693 = _T_2202 ? btb_bank0_rd_data_way1_out_45 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3948 = _T_3947 | _T_3693; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_46; // @[lib.scala 374:16]
  wire [21:0] _T_3694 = _T_2204 ? btb_bank0_rd_data_way1_out_46 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3949 = _T_3948 | _T_3694; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_47; // @[lib.scala 374:16]
  wire [21:0] _T_3695 = _T_2206 ? btb_bank0_rd_data_way1_out_47 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3950 = _T_3949 | _T_3695; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_48; // @[lib.scala 374:16]
  wire [21:0] _T_3696 = _T_2208 ? btb_bank0_rd_data_way1_out_48 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3951 = _T_3950 | _T_3696; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_49; // @[lib.scala 374:16]
  wire [21:0] _T_3697 = _T_2210 ? btb_bank0_rd_data_way1_out_49 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3952 = _T_3951 | _T_3697; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_50; // @[lib.scala 374:16]
  wire [21:0] _T_3698 = _T_2212 ? btb_bank0_rd_data_way1_out_50 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3953 = _T_3952 | _T_3698; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_51; // @[lib.scala 374:16]
  wire [21:0] _T_3699 = _T_2214 ? btb_bank0_rd_data_way1_out_51 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3954 = _T_3953 | _T_3699; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_52; // @[lib.scala 374:16]
  wire [21:0] _T_3700 = _T_2216 ? btb_bank0_rd_data_way1_out_52 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3955 = _T_3954 | _T_3700; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_53; // @[lib.scala 374:16]
  wire [21:0] _T_3701 = _T_2218 ? btb_bank0_rd_data_way1_out_53 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3956 = _T_3955 | _T_3701; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_54; // @[lib.scala 374:16]
  wire [21:0] _T_3702 = _T_2220 ? btb_bank0_rd_data_way1_out_54 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3957 = _T_3956 | _T_3702; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_55; // @[lib.scala 374:16]
  wire [21:0] _T_3703 = _T_2222 ? btb_bank0_rd_data_way1_out_55 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3958 = _T_3957 | _T_3703; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_56; // @[lib.scala 374:16]
  wire [21:0] _T_3704 = _T_2224 ? btb_bank0_rd_data_way1_out_56 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3959 = _T_3958 | _T_3704; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_57; // @[lib.scala 374:16]
  wire [21:0] _T_3705 = _T_2226 ? btb_bank0_rd_data_way1_out_57 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3960 = _T_3959 | _T_3705; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_58; // @[lib.scala 374:16]
  wire [21:0] _T_3706 = _T_2228 ? btb_bank0_rd_data_way1_out_58 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3961 = _T_3960 | _T_3706; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_59; // @[lib.scala 374:16]
  wire [21:0] _T_3707 = _T_2230 ? btb_bank0_rd_data_way1_out_59 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3962 = _T_3961 | _T_3707; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_60; // @[lib.scala 374:16]
  wire [21:0] _T_3708 = _T_2232 ? btb_bank0_rd_data_way1_out_60 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3963 = _T_3962 | _T_3708; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_61; // @[lib.scala 374:16]
  wire [21:0] _T_3709 = _T_2234 ? btb_bank0_rd_data_way1_out_61 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3964 = _T_3963 | _T_3709; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_62; // @[lib.scala 374:16]
  wire [21:0] _T_3710 = _T_2236 ? btb_bank0_rd_data_way1_out_62 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3965 = _T_3964 | _T_3710; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_63; // @[lib.scala 374:16]
  wire [21:0] _T_3711 = _T_2238 ? btb_bank0_rd_data_way1_out_63 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3966 = _T_3965 | _T_3711; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_64; // @[lib.scala 374:16]
  wire [21:0] _T_3712 = _T_2240 ? btb_bank0_rd_data_way1_out_64 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3967 = _T_3966 | _T_3712; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_65; // @[lib.scala 374:16]
  wire [21:0] _T_3713 = _T_2242 ? btb_bank0_rd_data_way1_out_65 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3968 = _T_3967 | _T_3713; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_66; // @[lib.scala 374:16]
  wire [21:0] _T_3714 = _T_2244 ? btb_bank0_rd_data_way1_out_66 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3969 = _T_3968 | _T_3714; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_67; // @[lib.scala 374:16]
  wire [21:0] _T_3715 = _T_2246 ? btb_bank0_rd_data_way1_out_67 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3970 = _T_3969 | _T_3715; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_68; // @[lib.scala 374:16]
  wire [21:0] _T_3716 = _T_2248 ? btb_bank0_rd_data_way1_out_68 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3971 = _T_3970 | _T_3716; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_69; // @[lib.scala 374:16]
  wire [21:0] _T_3717 = _T_2250 ? btb_bank0_rd_data_way1_out_69 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3972 = _T_3971 | _T_3717; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_70; // @[lib.scala 374:16]
  wire [21:0] _T_3718 = _T_2252 ? btb_bank0_rd_data_way1_out_70 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3973 = _T_3972 | _T_3718; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_71; // @[lib.scala 374:16]
  wire [21:0] _T_3719 = _T_2254 ? btb_bank0_rd_data_way1_out_71 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3974 = _T_3973 | _T_3719; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_72; // @[lib.scala 374:16]
  wire [21:0] _T_3720 = _T_2256 ? btb_bank0_rd_data_way1_out_72 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3975 = _T_3974 | _T_3720; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_73; // @[lib.scala 374:16]
  wire [21:0] _T_3721 = _T_2258 ? btb_bank0_rd_data_way1_out_73 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3976 = _T_3975 | _T_3721; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_74; // @[lib.scala 374:16]
  wire [21:0] _T_3722 = _T_2260 ? btb_bank0_rd_data_way1_out_74 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3977 = _T_3976 | _T_3722; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_75; // @[lib.scala 374:16]
  wire [21:0] _T_3723 = _T_2262 ? btb_bank0_rd_data_way1_out_75 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3978 = _T_3977 | _T_3723; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_76; // @[lib.scala 374:16]
  wire [21:0] _T_3724 = _T_2264 ? btb_bank0_rd_data_way1_out_76 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3979 = _T_3978 | _T_3724; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_77; // @[lib.scala 374:16]
  wire [21:0] _T_3725 = _T_2266 ? btb_bank0_rd_data_way1_out_77 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3980 = _T_3979 | _T_3725; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_78; // @[lib.scala 374:16]
  wire [21:0] _T_3726 = _T_2268 ? btb_bank0_rd_data_way1_out_78 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3981 = _T_3980 | _T_3726; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_79; // @[lib.scala 374:16]
  wire [21:0] _T_3727 = _T_2270 ? btb_bank0_rd_data_way1_out_79 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3982 = _T_3981 | _T_3727; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_80; // @[lib.scala 374:16]
  wire [21:0] _T_3728 = _T_2272 ? btb_bank0_rd_data_way1_out_80 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3983 = _T_3982 | _T_3728; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_81; // @[lib.scala 374:16]
  wire [21:0] _T_3729 = _T_2274 ? btb_bank0_rd_data_way1_out_81 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3984 = _T_3983 | _T_3729; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_82; // @[lib.scala 374:16]
  wire [21:0] _T_3730 = _T_2276 ? btb_bank0_rd_data_way1_out_82 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3985 = _T_3984 | _T_3730; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_83; // @[lib.scala 374:16]
  wire [21:0] _T_3731 = _T_2278 ? btb_bank0_rd_data_way1_out_83 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3986 = _T_3985 | _T_3731; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_84; // @[lib.scala 374:16]
  wire [21:0] _T_3732 = _T_2280 ? btb_bank0_rd_data_way1_out_84 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3987 = _T_3986 | _T_3732; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_85; // @[lib.scala 374:16]
  wire [21:0] _T_3733 = _T_2282 ? btb_bank0_rd_data_way1_out_85 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3988 = _T_3987 | _T_3733; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_86; // @[lib.scala 374:16]
  wire [21:0] _T_3734 = _T_2284 ? btb_bank0_rd_data_way1_out_86 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3989 = _T_3988 | _T_3734; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_87; // @[lib.scala 374:16]
  wire [21:0] _T_3735 = _T_2286 ? btb_bank0_rd_data_way1_out_87 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3990 = _T_3989 | _T_3735; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_88; // @[lib.scala 374:16]
  wire [21:0] _T_3736 = _T_2288 ? btb_bank0_rd_data_way1_out_88 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3991 = _T_3990 | _T_3736; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_89; // @[lib.scala 374:16]
  wire [21:0] _T_3737 = _T_2290 ? btb_bank0_rd_data_way1_out_89 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3992 = _T_3991 | _T_3737; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_90; // @[lib.scala 374:16]
  wire [21:0] _T_3738 = _T_2292 ? btb_bank0_rd_data_way1_out_90 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3993 = _T_3992 | _T_3738; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_91; // @[lib.scala 374:16]
  wire [21:0] _T_3739 = _T_2294 ? btb_bank0_rd_data_way1_out_91 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3994 = _T_3993 | _T_3739; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_92; // @[lib.scala 374:16]
  wire [21:0] _T_3740 = _T_2296 ? btb_bank0_rd_data_way1_out_92 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3995 = _T_3994 | _T_3740; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_93; // @[lib.scala 374:16]
  wire [21:0] _T_3741 = _T_2298 ? btb_bank0_rd_data_way1_out_93 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3996 = _T_3995 | _T_3741; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_94; // @[lib.scala 374:16]
  wire [21:0] _T_3742 = _T_2300 ? btb_bank0_rd_data_way1_out_94 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3997 = _T_3996 | _T_3742; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_95; // @[lib.scala 374:16]
  wire [21:0] _T_3743 = _T_2302 ? btb_bank0_rd_data_way1_out_95 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3998 = _T_3997 | _T_3743; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_96; // @[lib.scala 374:16]
  wire [21:0] _T_3744 = _T_2304 ? btb_bank0_rd_data_way1_out_96 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3999 = _T_3998 | _T_3744; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_97; // @[lib.scala 374:16]
  wire [21:0] _T_3745 = _T_2306 ? btb_bank0_rd_data_way1_out_97 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4000 = _T_3999 | _T_3745; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_98; // @[lib.scala 374:16]
  wire [21:0] _T_3746 = _T_2308 ? btb_bank0_rd_data_way1_out_98 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4001 = _T_4000 | _T_3746; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_99; // @[lib.scala 374:16]
  wire [21:0] _T_3747 = _T_2310 ? btb_bank0_rd_data_way1_out_99 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4002 = _T_4001 | _T_3747; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_100; // @[lib.scala 374:16]
  wire [21:0] _T_3748 = _T_2312 ? btb_bank0_rd_data_way1_out_100 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4003 = _T_4002 | _T_3748; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_101; // @[lib.scala 374:16]
  wire [21:0] _T_3749 = _T_2314 ? btb_bank0_rd_data_way1_out_101 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4004 = _T_4003 | _T_3749; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_102; // @[lib.scala 374:16]
  wire [21:0] _T_3750 = _T_2316 ? btb_bank0_rd_data_way1_out_102 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4005 = _T_4004 | _T_3750; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_103; // @[lib.scala 374:16]
  wire [21:0] _T_3751 = _T_2318 ? btb_bank0_rd_data_way1_out_103 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4006 = _T_4005 | _T_3751; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_104; // @[lib.scala 374:16]
  wire [21:0] _T_3752 = _T_2320 ? btb_bank0_rd_data_way1_out_104 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4007 = _T_4006 | _T_3752; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_105; // @[lib.scala 374:16]
  wire [21:0] _T_3753 = _T_2322 ? btb_bank0_rd_data_way1_out_105 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4008 = _T_4007 | _T_3753; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_106; // @[lib.scala 374:16]
  wire [21:0] _T_3754 = _T_2324 ? btb_bank0_rd_data_way1_out_106 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4009 = _T_4008 | _T_3754; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_107; // @[lib.scala 374:16]
  wire [21:0] _T_3755 = _T_2326 ? btb_bank0_rd_data_way1_out_107 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4010 = _T_4009 | _T_3755; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_108; // @[lib.scala 374:16]
  wire [21:0] _T_3756 = _T_2328 ? btb_bank0_rd_data_way1_out_108 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4011 = _T_4010 | _T_3756; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_109; // @[lib.scala 374:16]
  wire [21:0] _T_3757 = _T_2330 ? btb_bank0_rd_data_way1_out_109 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4012 = _T_4011 | _T_3757; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_110; // @[lib.scala 374:16]
  wire [21:0] _T_3758 = _T_2332 ? btb_bank0_rd_data_way1_out_110 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4013 = _T_4012 | _T_3758; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_111; // @[lib.scala 374:16]
  wire [21:0] _T_3759 = _T_2334 ? btb_bank0_rd_data_way1_out_111 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4014 = _T_4013 | _T_3759; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_112; // @[lib.scala 374:16]
  wire [21:0] _T_3760 = _T_2336 ? btb_bank0_rd_data_way1_out_112 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4015 = _T_4014 | _T_3760; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_113; // @[lib.scala 374:16]
  wire [21:0] _T_3761 = _T_2338 ? btb_bank0_rd_data_way1_out_113 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4016 = _T_4015 | _T_3761; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_114; // @[lib.scala 374:16]
  wire [21:0] _T_3762 = _T_2340 ? btb_bank0_rd_data_way1_out_114 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4017 = _T_4016 | _T_3762; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_115; // @[lib.scala 374:16]
  wire [21:0] _T_3763 = _T_2342 ? btb_bank0_rd_data_way1_out_115 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4018 = _T_4017 | _T_3763; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_116; // @[lib.scala 374:16]
  wire [21:0] _T_3764 = _T_2344 ? btb_bank0_rd_data_way1_out_116 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4019 = _T_4018 | _T_3764; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_117; // @[lib.scala 374:16]
  wire [21:0] _T_3765 = _T_2346 ? btb_bank0_rd_data_way1_out_117 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4020 = _T_4019 | _T_3765; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_118; // @[lib.scala 374:16]
  wire [21:0] _T_3766 = _T_2348 ? btb_bank0_rd_data_way1_out_118 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4021 = _T_4020 | _T_3766; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_119; // @[lib.scala 374:16]
  wire [21:0] _T_3767 = _T_2350 ? btb_bank0_rd_data_way1_out_119 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4022 = _T_4021 | _T_3767; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_120; // @[lib.scala 374:16]
  wire [21:0] _T_3768 = _T_2352 ? btb_bank0_rd_data_way1_out_120 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4023 = _T_4022 | _T_3768; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_121; // @[lib.scala 374:16]
  wire [21:0] _T_3769 = _T_2354 ? btb_bank0_rd_data_way1_out_121 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4024 = _T_4023 | _T_3769; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_122; // @[lib.scala 374:16]
  wire [21:0] _T_3770 = _T_2356 ? btb_bank0_rd_data_way1_out_122 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4025 = _T_4024 | _T_3770; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_123; // @[lib.scala 374:16]
  wire [21:0] _T_3771 = _T_2358 ? btb_bank0_rd_data_way1_out_123 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4026 = _T_4025 | _T_3771; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_124; // @[lib.scala 374:16]
  wire [21:0] _T_3772 = _T_2360 ? btb_bank0_rd_data_way1_out_124 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4027 = _T_4026 | _T_3772; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_125; // @[lib.scala 374:16]
  wire [21:0] _T_3773 = _T_2362 ? btb_bank0_rd_data_way1_out_125 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4028 = _T_4027 | _T_3773; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_126; // @[lib.scala 374:16]
  wire [21:0] _T_3774 = _T_2364 ? btb_bank0_rd_data_way1_out_126 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4029 = _T_4028 | _T_3774; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_127; // @[lib.scala 374:16]
  wire [21:0] _T_3775 = _T_2366 ? btb_bank0_rd_data_way1_out_127 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4030 = _T_4029 | _T_3775; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_128; // @[lib.scala 374:16]
  wire [21:0] _T_3776 = _T_2368 ? btb_bank0_rd_data_way1_out_128 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4031 = _T_4030 | _T_3776; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_129; // @[lib.scala 374:16]
  wire [21:0] _T_3777 = _T_2370 ? btb_bank0_rd_data_way1_out_129 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4032 = _T_4031 | _T_3777; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_130; // @[lib.scala 374:16]
  wire [21:0] _T_3778 = _T_2372 ? btb_bank0_rd_data_way1_out_130 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4033 = _T_4032 | _T_3778; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_131; // @[lib.scala 374:16]
  wire [21:0] _T_3779 = _T_2374 ? btb_bank0_rd_data_way1_out_131 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4034 = _T_4033 | _T_3779; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_132; // @[lib.scala 374:16]
  wire [21:0] _T_3780 = _T_2376 ? btb_bank0_rd_data_way1_out_132 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4035 = _T_4034 | _T_3780; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_133; // @[lib.scala 374:16]
  wire [21:0] _T_3781 = _T_2378 ? btb_bank0_rd_data_way1_out_133 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4036 = _T_4035 | _T_3781; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_134; // @[lib.scala 374:16]
  wire [21:0] _T_3782 = _T_2380 ? btb_bank0_rd_data_way1_out_134 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4037 = _T_4036 | _T_3782; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_135; // @[lib.scala 374:16]
  wire [21:0] _T_3783 = _T_2382 ? btb_bank0_rd_data_way1_out_135 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4038 = _T_4037 | _T_3783; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_136; // @[lib.scala 374:16]
  wire [21:0] _T_3784 = _T_2384 ? btb_bank0_rd_data_way1_out_136 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4039 = _T_4038 | _T_3784; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_137; // @[lib.scala 374:16]
  wire [21:0] _T_3785 = _T_2386 ? btb_bank0_rd_data_way1_out_137 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4040 = _T_4039 | _T_3785; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_138; // @[lib.scala 374:16]
  wire [21:0] _T_3786 = _T_2388 ? btb_bank0_rd_data_way1_out_138 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4041 = _T_4040 | _T_3786; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_139; // @[lib.scala 374:16]
  wire [21:0] _T_3787 = _T_2390 ? btb_bank0_rd_data_way1_out_139 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4042 = _T_4041 | _T_3787; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_140; // @[lib.scala 374:16]
  wire [21:0] _T_3788 = _T_2392 ? btb_bank0_rd_data_way1_out_140 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4043 = _T_4042 | _T_3788; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_141; // @[lib.scala 374:16]
  wire [21:0] _T_3789 = _T_2394 ? btb_bank0_rd_data_way1_out_141 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4044 = _T_4043 | _T_3789; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_142; // @[lib.scala 374:16]
  wire [21:0] _T_3790 = _T_2396 ? btb_bank0_rd_data_way1_out_142 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4045 = _T_4044 | _T_3790; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_143; // @[lib.scala 374:16]
  wire [21:0] _T_3791 = _T_2398 ? btb_bank0_rd_data_way1_out_143 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4046 = _T_4045 | _T_3791; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_144; // @[lib.scala 374:16]
  wire [21:0] _T_3792 = _T_2400 ? btb_bank0_rd_data_way1_out_144 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4047 = _T_4046 | _T_3792; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_145; // @[lib.scala 374:16]
  wire [21:0] _T_3793 = _T_2402 ? btb_bank0_rd_data_way1_out_145 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4048 = _T_4047 | _T_3793; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_146; // @[lib.scala 374:16]
  wire [21:0] _T_3794 = _T_2404 ? btb_bank0_rd_data_way1_out_146 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4049 = _T_4048 | _T_3794; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_147; // @[lib.scala 374:16]
  wire [21:0] _T_3795 = _T_2406 ? btb_bank0_rd_data_way1_out_147 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4050 = _T_4049 | _T_3795; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_148; // @[lib.scala 374:16]
  wire [21:0] _T_3796 = _T_2408 ? btb_bank0_rd_data_way1_out_148 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4051 = _T_4050 | _T_3796; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_149; // @[lib.scala 374:16]
  wire [21:0] _T_3797 = _T_2410 ? btb_bank0_rd_data_way1_out_149 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4052 = _T_4051 | _T_3797; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_150; // @[lib.scala 374:16]
  wire [21:0] _T_3798 = _T_2412 ? btb_bank0_rd_data_way1_out_150 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4053 = _T_4052 | _T_3798; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_151; // @[lib.scala 374:16]
  wire [21:0] _T_3799 = _T_2414 ? btb_bank0_rd_data_way1_out_151 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4054 = _T_4053 | _T_3799; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_152; // @[lib.scala 374:16]
  wire [21:0] _T_3800 = _T_2416 ? btb_bank0_rd_data_way1_out_152 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4055 = _T_4054 | _T_3800; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_153; // @[lib.scala 374:16]
  wire [21:0] _T_3801 = _T_2418 ? btb_bank0_rd_data_way1_out_153 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4056 = _T_4055 | _T_3801; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_154; // @[lib.scala 374:16]
  wire [21:0] _T_3802 = _T_2420 ? btb_bank0_rd_data_way1_out_154 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4057 = _T_4056 | _T_3802; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_155; // @[lib.scala 374:16]
  wire [21:0] _T_3803 = _T_2422 ? btb_bank0_rd_data_way1_out_155 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4058 = _T_4057 | _T_3803; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_156; // @[lib.scala 374:16]
  wire [21:0] _T_3804 = _T_2424 ? btb_bank0_rd_data_way1_out_156 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4059 = _T_4058 | _T_3804; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_157; // @[lib.scala 374:16]
  wire [21:0] _T_3805 = _T_2426 ? btb_bank0_rd_data_way1_out_157 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4060 = _T_4059 | _T_3805; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_158; // @[lib.scala 374:16]
  wire [21:0] _T_3806 = _T_2428 ? btb_bank0_rd_data_way1_out_158 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4061 = _T_4060 | _T_3806; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_159; // @[lib.scala 374:16]
  wire [21:0] _T_3807 = _T_2430 ? btb_bank0_rd_data_way1_out_159 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4062 = _T_4061 | _T_3807; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_160; // @[lib.scala 374:16]
  wire [21:0] _T_3808 = _T_2432 ? btb_bank0_rd_data_way1_out_160 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4063 = _T_4062 | _T_3808; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_161; // @[lib.scala 374:16]
  wire [21:0] _T_3809 = _T_2434 ? btb_bank0_rd_data_way1_out_161 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4064 = _T_4063 | _T_3809; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_162; // @[lib.scala 374:16]
  wire [21:0] _T_3810 = _T_2436 ? btb_bank0_rd_data_way1_out_162 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4065 = _T_4064 | _T_3810; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_163; // @[lib.scala 374:16]
  wire [21:0] _T_3811 = _T_2438 ? btb_bank0_rd_data_way1_out_163 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4066 = _T_4065 | _T_3811; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_164; // @[lib.scala 374:16]
  wire [21:0] _T_3812 = _T_2440 ? btb_bank0_rd_data_way1_out_164 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4067 = _T_4066 | _T_3812; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_165; // @[lib.scala 374:16]
  wire [21:0] _T_3813 = _T_2442 ? btb_bank0_rd_data_way1_out_165 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4068 = _T_4067 | _T_3813; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_166; // @[lib.scala 374:16]
  wire [21:0] _T_3814 = _T_2444 ? btb_bank0_rd_data_way1_out_166 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4069 = _T_4068 | _T_3814; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_167; // @[lib.scala 374:16]
  wire [21:0] _T_3815 = _T_2446 ? btb_bank0_rd_data_way1_out_167 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4070 = _T_4069 | _T_3815; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_168; // @[lib.scala 374:16]
  wire [21:0] _T_3816 = _T_2448 ? btb_bank0_rd_data_way1_out_168 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4071 = _T_4070 | _T_3816; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_169; // @[lib.scala 374:16]
  wire [21:0] _T_3817 = _T_2450 ? btb_bank0_rd_data_way1_out_169 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4072 = _T_4071 | _T_3817; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_170; // @[lib.scala 374:16]
  wire [21:0] _T_3818 = _T_2452 ? btb_bank0_rd_data_way1_out_170 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4073 = _T_4072 | _T_3818; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_171; // @[lib.scala 374:16]
  wire [21:0] _T_3819 = _T_2454 ? btb_bank0_rd_data_way1_out_171 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4074 = _T_4073 | _T_3819; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_172; // @[lib.scala 374:16]
  wire [21:0] _T_3820 = _T_2456 ? btb_bank0_rd_data_way1_out_172 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4075 = _T_4074 | _T_3820; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_173; // @[lib.scala 374:16]
  wire [21:0] _T_3821 = _T_2458 ? btb_bank0_rd_data_way1_out_173 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4076 = _T_4075 | _T_3821; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_174; // @[lib.scala 374:16]
  wire [21:0] _T_3822 = _T_2460 ? btb_bank0_rd_data_way1_out_174 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4077 = _T_4076 | _T_3822; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_175; // @[lib.scala 374:16]
  wire [21:0] _T_3823 = _T_2462 ? btb_bank0_rd_data_way1_out_175 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4078 = _T_4077 | _T_3823; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_176; // @[lib.scala 374:16]
  wire [21:0] _T_3824 = _T_2464 ? btb_bank0_rd_data_way1_out_176 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4079 = _T_4078 | _T_3824; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_177; // @[lib.scala 374:16]
  wire [21:0] _T_3825 = _T_2466 ? btb_bank0_rd_data_way1_out_177 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4080 = _T_4079 | _T_3825; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_178; // @[lib.scala 374:16]
  wire [21:0] _T_3826 = _T_2468 ? btb_bank0_rd_data_way1_out_178 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4081 = _T_4080 | _T_3826; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_179; // @[lib.scala 374:16]
  wire [21:0] _T_3827 = _T_2470 ? btb_bank0_rd_data_way1_out_179 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4082 = _T_4081 | _T_3827; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_180; // @[lib.scala 374:16]
  wire [21:0] _T_3828 = _T_2472 ? btb_bank0_rd_data_way1_out_180 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4083 = _T_4082 | _T_3828; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_181; // @[lib.scala 374:16]
  wire [21:0] _T_3829 = _T_2474 ? btb_bank0_rd_data_way1_out_181 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4084 = _T_4083 | _T_3829; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_182; // @[lib.scala 374:16]
  wire [21:0] _T_3830 = _T_2476 ? btb_bank0_rd_data_way1_out_182 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4085 = _T_4084 | _T_3830; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_183; // @[lib.scala 374:16]
  wire [21:0] _T_3831 = _T_2478 ? btb_bank0_rd_data_way1_out_183 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4086 = _T_4085 | _T_3831; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_184; // @[lib.scala 374:16]
  wire [21:0] _T_3832 = _T_2480 ? btb_bank0_rd_data_way1_out_184 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4087 = _T_4086 | _T_3832; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_185; // @[lib.scala 374:16]
  wire [21:0] _T_3833 = _T_2482 ? btb_bank0_rd_data_way1_out_185 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4088 = _T_4087 | _T_3833; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_186; // @[lib.scala 374:16]
  wire [21:0] _T_3834 = _T_2484 ? btb_bank0_rd_data_way1_out_186 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4089 = _T_4088 | _T_3834; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_187; // @[lib.scala 374:16]
  wire [21:0] _T_3835 = _T_2486 ? btb_bank0_rd_data_way1_out_187 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4090 = _T_4089 | _T_3835; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_188; // @[lib.scala 374:16]
  wire [21:0] _T_3836 = _T_2488 ? btb_bank0_rd_data_way1_out_188 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4091 = _T_4090 | _T_3836; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_189; // @[lib.scala 374:16]
  wire [21:0] _T_3837 = _T_2490 ? btb_bank0_rd_data_way1_out_189 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4092 = _T_4091 | _T_3837; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_190; // @[lib.scala 374:16]
  wire [21:0] _T_3838 = _T_2492 ? btb_bank0_rd_data_way1_out_190 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4093 = _T_4092 | _T_3838; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_191; // @[lib.scala 374:16]
  wire [21:0] _T_3839 = _T_2494 ? btb_bank0_rd_data_way1_out_191 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4094 = _T_4093 | _T_3839; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_192; // @[lib.scala 374:16]
  wire [21:0] _T_3840 = _T_2496 ? btb_bank0_rd_data_way1_out_192 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4095 = _T_4094 | _T_3840; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_193; // @[lib.scala 374:16]
  wire [21:0] _T_3841 = _T_2498 ? btb_bank0_rd_data_way1_out_193 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4096 = _T_4095 | _T_3841; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_194; // @[lib.scala 374:16]
  wire [21:0] _T_3842 = _T_2500 ? btb_bank0_rd_data_way1_out_194 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4097 = _T_4096 | _T_3842; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_195; // @[lib.scala 374:16]
  wire [21:0] _T_3843 = _T_2502 ? btb_bank0_rd_data_way1_out_195 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4098 = _T_4097 | _T_3843; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_196; // @[lib.scala 374:16]
  wire [21:0] _T_3844 = _T_2504 ? btb_bank0_rd_data_way1_out_196 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4099 = _T_4098 | _T_3844; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_197; // @[lib.scala 374:16]
  wire [21:0] _T_3845 = _T_2506 ? btb_bank0_rd_data_way1_out_197 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4100 = _T_4099 | _T_3845; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_198; // @[lib.scala 374:16]
  wire [21:0] _T_3846 = _T_2508 ? btb_bank0_rd_data_way1_out_198 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4101 = _T_4100 | _T_3846; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_199; // @[lib.scala 374:16]
  wire [21:0] _T_3847 = _T_2510 ? btb_bank0_rd_data_way1_out_199 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4102 = _T_4101 | _T_3847; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_200; // @[lib.scala 374:16]
  wire [21:0] _T_3848 = _T_2512 ? btb_bank0_rd_data_way1_out_200 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4103 = _T_4102 | _T_3848; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_201; // @[lib.scala 374:16]
  wire [21:0] _T_3849 = _T_2514 ? btb_bank0_rd_data_way1_out_201 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4104 = _T_4103 | _T_3849; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_202; // @[lib.scala 374:16]
  wire [21:0] _T_3850 = _T_2516 ? btb_bank0_rd_data_way1_out_202 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4105 = _T_4104 | _T_3850; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_203; // @[lib.scala 374:16]
  wire [21:0] _T_3851 = _T_2518 ? btb_bank0_rd_data_way1_out_203 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4106 = _T_4105 | _T_3851; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_204; // @[lib.scala 374:16]
  wire [21:0] _T_3852 = _T_2520 ? btb_bank0_rd_data_way1_out_204 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4107 = _T_4106 | _T_3852; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_205; // @[lib.scala 374:16]
  wire [21:0] _T_3853 = _T_2522 ? btb_bank0_rd_data_way1_out_205 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4108 = _T_4107 | _T_3853; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_206; // @[lib.scala 374:16]
  wire [21:0] _T_3854 = _T_2524 ? btb_bank0_rd_data_way1_out_206 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4109 = _T_4108 | _T_3854; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_207; // @[lib.scala 374:16]
  wire [21:0] _T_3855 = _T_2526 ? btb_bank0_rd_data_way1_out_207 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4110 = _T_4109 | _T_3855; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_208; // @[lib.scala 374:16]
  wire [21:0] _T_3856 = _T_2528 ? btb_bank0_rd_data_way1_out_208 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4111 = _T_4110 | _T_3856; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_209; // @[lib.scala 374:16]
  wire [21:0] _T_3857 = _T_2530 ? btb_bank0_rd_data_way1_out_209 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4112 = _T_4111 | _T_3857; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_210; // @[lib.scala 374:16]
  wire [21:0] _T_3858 = _T_2532 ? btb_bank0_rd_data_way1_out_210 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4113 = _T_4112 | _T_3858; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_211; // @[lib.scala 374:16]
  wire [21:0] _T_3859 = _T_2534 ? btb_bank0_rd_data_way1_out_211 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4114 = _T_4113 | _T_3859; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_212; // @[lib.scala 374:16]
  wire [21:0] _T_3860 = _T_2536 ? btb_bank0_rd_data_way1_out_212 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4115 = _T_4114 | _T_3860; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_213; // @[lib.scala 374:16]
  wire [21:0] _T_3861 = _T_2538 ? btb_bank0_rd_data_way1_out_213 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4116 = _T_4115 | _T_3861; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_214; // @[lib.scala 374:16]
  wire [21:0] _T_3862 = _T_2540 ? btb_bank0_rd_data_way1_out_214 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4117 = _T_4116 | _T_3862; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_215; // @[lib.scala 374:16]
  wire [21:0] _T_3863 = _T_2542 ? btb_bank0_rd_data_way1_out_215 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4118 = _T_4117 | _T_3863; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_216; // @[lib.scala 374:16]
  wire [21:0] _T_3864 = _T_2544 ? btb_bank0_rd_data_way1_out_216 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4119 = _T_4118 | _T_3864; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_217; // @[lib.scala 374:16]
  wire [21:0] _T_3865 = _T_2546 ? btb_bank0_rd_data_way1_out_217 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4120 = _T_4119 | _T_3865; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_218; // @[lib.scala 374:16]
  wire [21:0] _T_3866 = _T_2548 ? btb_bank0_rd_data_way1_out_218 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4121 = _T_4120 | _T_3866; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_219; // @[lib.scala 374:16]
  wire [21:0] _T_3867 = _T_2550 ? btb_bank0_rd_data_way1_out_219 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4122 = _T_4121 | _T_3867; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_220; // @[lib.scala 374:16]
  wire [21:0] _T_3868 = _T_2552 ? btb_bank0_rd_data_way1_out_220 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4123 = _T_4122 | _T_3868; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_221; // @[lib.scala 374:16]
  wire [21:0] _T_3869 = _T_2554 ? btb_bank0_rd_data_way1_out_221 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4124 = _T_4123 | _T_3869; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_222; // @[lib.scala 374:16]
  wire [21:0] _T_3870 = _T_2556 ? btb_bank0_rd_data_way1_out_222 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4125 = _T_4124 | _T_3870; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_223; // @[lib.scala 374:16]
  wire [21:0] _T_3871 = _T_2558 ? btb_bank0_rd_data_way1_out_223 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4126 = _T_4125 | _T_3871; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_224; // @[lib.scala 374:16]
  wire [21:0] _T_3872 = _T_2560 ? btb_bank0_rd_data_way1_out_224 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4127 = _T_4126 | _T_3872; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_225; // @[lib.scala 374:16]
  wire [21:0] _T_3873 = _T_2562 ? btb_bank0_rd_data_way1_out_225 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4128 = _T_4127 | _T_3873; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_226; // @[lib.scala 374:16]
  wire [21:0] _T_3874 = _T_2564 ? btb_bank0_rd_data_way1_out_226 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4129 = _T_4128 | _T_3874; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_227; // @[lib.scala 374:16]
  wire [21:0] _T_3875 = _T_2566 ? btb_bank0_rd_data_way1_out_227 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4130 = _T_4129 | _T_3875; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_228; // @[lib.scala 374:16]
  wire [21:0] _T_3876 = _T_2568 ? btb_bank0_rd_data_way1_out_228 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4131 = _T_4130 | _T_3876; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_229; // @[lib.scala 374:16]
  wire [21:0] _T_3877 = _T_2570 ? btb_bank0_rd_data_way1_out_229 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4132 = _T_4131 | _T_3877; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_230; // @[lib.scala 374:16]
  wire [21:0] _T_3878 = _T_2572 ? btb_bank0_rd_data_way1_out_230 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4133 = _T_4132 | _T_3878; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_231; // @[lib.scala 374:16]
  wire [21:0] _T_3879 = _T_2574 ? btb_bank0_rd_data_way1_out_231 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4134 = _T_4133 | _T_3879; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_232; // @[lib.scala 374:16]
  wire [21:0] _T_3880 = _T_2576 ? btb_bank0_rd_data_way1_out_232 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4135 = _T_4134 | _T_3880; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_233; // @[lib.scala 374:16]
  wire [21:0] _T_3881 = _T_2578 ? btb_bank0_rd_data_way1_out_233 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4136 = _T_4135 | _T_3881; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_234; // @[lib.scala 374:16]
  wire [21:0] _T_3882 = _T_2580 ? btb_bank0_rd_data_way1_out_234 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4137 = _T_4136 | _T_3882; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_235; // @[lib.scala 374:16]
  wire [21:0] _T_3883 = _T_2582 ? btb_bank0_rd_data_way1_out_235 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4138 = _T_4137 | _T_3883; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_236; // @[lib.scala 374:16]
  wire [21:0] _T_3884 = _T_2584 ? btb_bank0_rd_data_way1_out_236 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4139 = _T_4138 | _T_3884; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_237; // @[lib.scala 374:16]
  wire [21:0] _T_3885 = _T_2586 ? btb_bank0_rd_data_way1_out_237 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4140 = _T_4139 | _T_3885; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_238; // @[lib.scala 374:16]
  wire [21:0] _T_3886 = _T_2588 ? btb_bank0_rd_data_way1_out_238 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4141 = _T_4140 | _T_3886; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_239; // @[lib.scala 374:16]
  wire [21:0] _T_3887 = _T_2590 ? btb_bank0_rd_data_way1_out_239 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4142 = _T_4141 | _T_3887; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_240; // @[lib.scala 374:16]
  wire [21:0] _T_3888 = _T_2592 ? btb_bank0_rd_data_way1_out_240 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4143 = _T_4142 | _T_3888; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_241; // @[lib.scala 374:16]
  wire [21:0] _T_3889 = _T_2594 ? btb_bank0_rd_data_way1_out_241 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4144 = _T_4143 | _T_3889; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_242; // @[lib.scala 374:16]
  wire [21:0] _T_3890 = _T_2596 ? btb_bank0_rd_data_way1_out_242 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4145 = _T_4144 | _T_3890; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_243; // @[lib.scala 374:16]
  wire [21:0] _T_3891 = _T_2598 ? btb_bank0_rd_data_way1_out_243 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4146 = _T_4145 | _T_3891; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_244; // @[lib.scala 374:16]
  wire [21:0] _T_3892 = _T_2600 ? btb_bank0_rd_data_way1_out_244 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4147 = _T_4146 | _T_3892; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_245; // @[lib.scala 374:16]
  wire [21:0] _T_3893 = _T_2602 ? btb_bank0_rd_data_way1_out_245 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4148 = _T_4147 | _T_3893; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_246; // @[lib.scala 374:16]
  wire [21:0] _T_3894 = _T_2604 ? btb_bank0_rd_data_way1_out_246 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4149 = _T_4148 | _T_3894; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_247; // @[lib.scala 374:16]
  wire [21:0] _T_3895 = _T_2606 ? btb_bank0_rd_data_way1_out_247 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4150 = _T_4149 | _T_3895; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_248; // @[lib.scala 374:16]
  wire [21:0] _T_3896 = _T_2608 ? btb_bank0_rd_data_way1_out_248 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4151 = _T_4150 | _T_3896; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_249; // @[lib.scala 374:16]
  wire [21:0] _T_3897 = _T_2610 ? btb_bank0_rd_data_way1_out_249 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4152 = _T_4151 | _T_3897; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_250; // @[lib.scala 374:16]
  wire [21:0] _T_3898 = _T_2612 ? btb_bank0_rd_data_way1_out_250 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4153 = _T_4152 | _T_3898; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_251; // @[lib.scala 374:16]
  wire [21:0] _T_3899 = _T_2614 ? btb_bank0_rd_data_way1_out_251 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4154 = _T_4153 | _T_3899; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_252; // @[lib.scala 374:16]
  wire [21:0] _T_3900 = _T_2616 ? btb_bank0_rd_data_way1_out_252 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4155 = _T_4154 | _T_3900; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_253; // @[lib.scala 374:16]
  wire [21:0] _T_3901 = _T_2618 ? btb_bank0_rd_data_way1_out_253 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4156 = _T_4155 | _T_3901; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_254; // @[lib.scala 374:16]
  wire [21:0] _T_3902 = _T_2620 ? btb_bank0_rd_data_way1_out_254 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4157 = _T_4156 | _T_3902; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_255; // @[lib.scala 374:16]
  wire [21:0] _T_3903 = _T_2622 ? btb_bank0_rd_data_way1_out_255 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] btb_bank0_rd_data_way1_f = _T_4157 | _T_3903; // @[Mux.scala 27:72]
  wire  _T_55 = btb_bank0_rd_data_way1_f[21:17] == fetch_rd_tag_f; // @[ifu_bp_ctl.scala 131:97]
  wire  _T_56 = btb_bank0_rd_data_way1_f[0] & _T_55; // @[ifu_bp_ctl.scala 131:55]
  wire  _T_59 = _T_56 & _T_49; // @[ifu_bp_ctl.scala 131:117]
  wire  _T_60 = _T_59 & io_ifc_fetch_req_f; // @[ifu_bp_ctl.scala 132:76]
  wire  tag_match_way1_f = _T_60 & _T; // @[ifu_bp_ctl.scala 132:97]
  wire  _T_91 = btb_bank0_rd_data_way1_f[3] ^ btb_bank0_rd_data_way1_f[4]; // @[ifu_bp_ctl.scala 145:91]
  wire  _T_92 = tag_match_way1_f & _T_91; // @[ifu_bp_ctl.scala 145:56]
  wire  _T_96 = ~_T_91; // @[ifu_bp_ctl.scala 146:58]
  wire  _T_97 = tag_match_way1_f & _T_96; // @[ifu_bp_ctl.scala 146:56]
  wire [1:0] tag_match_way1_expanded_f = {_T_92,_T_97}; // @[Cat.scala 29:58]
  wire [21:0] _T_128 = tag_match_way1_expanded_f[1] ? btb_bank0_rd_data_way1_f : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] btb_bank0o_rd_data_f = _T_127 | _T_128; // @[Mux.scala 27:72]
  wire [21:0] _T_146 = _T_144 ? btb_bank0o_rd_data_f : 22'h0; // @[Mux.scala 27:72]
  wire  _T_4160 = btb_rd_addr_p1_f == 8'h0; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4672 = _T_4160 ? btb_bank0_rd_data_way0_out_0 : 22'h0; // @[Mux.scala 27:72]
  wire  _T_4162 = btb_rd_addr_p1_f == 8'h1; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4673 = _T_4162 ? btb_bank0_rd_data_way0_out_1 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4928 = _T_4672 | _T_4673; // @[Mux.scala 27:72]
  wire  _T_4164 = btb_rd_addr_p1_f == 8'h2; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4674 = _T_4164 ? btb_bank0_rd_data_way0_out_2 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4929 = _T_4928 | _T_4674; // @[Mux.scala 27:72]
  wire  _T_4166 = btb_rd_addr_p1_f == 8'h3; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4675 = _T_4166 ? btb_bank0_rd_data_way0_out_3 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4930 = _T_4929 | _T_4675; // @[Mux.scala 27:72]
  wire  _T_4168 = btb_rd_addr_p1_f == 8'h4; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4676 = _T_4168 ? btb_bank0_rd_data_way0_out_4 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4931 = _T_4930 | _T_4676; // @[Mux.scala 27:72]
  wire  _T_4170 = btb_rd_addr_p1_f == 8'h5; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4677 = _T_4170 ? btb_bank0_rd_data_way0_out_5 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4932 = _T_4931 | _T_4677; // @[Mux.scala 27:72]
  wire  _T_4172 = btb_rd_addr_p1_f == 8'h6; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4678 = _T_4172 ? btb_bank0_rd_data_way0_out_6 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4933 = _T_4932 | _T_4678; // @[Mux.scala 27:72]
  wire  _T_4174 = btb_rd_addr_p1_f == 8'h7; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4679 = _T_4174 ? btb_bank0_rd_data_way0_out_7 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4934 = _T_4933 | _T_4679; // @[Mux.scala 27:72]
  wire  _T_4176 = btb_rd_addr_p1_f == 8'h8; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4680 = _T_4176 ? btb_bank0_rd_data_way0_out_8 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4935 = _T_4934 | _T_4680; // @[Mux.scala 27:72]
  wire  _T_4178 = btb_rd_addr_p1_f == 8'h9; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4681 = _T_4178 ? btb_bank0_rd_data_way0_out_9 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4936 = _T_4935 | _T_4681; // @[Mux.scala 27:72]
  wire  _T_4180 = btb_rd_addr_p1_f == 8'ha; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4682 = _T_4180 ? btb_bank0_rd_data_way0_out_10 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4937 = _T_4936 | _T_4682; // @[Mux.scala 27:72]
  wire  _T_4182 = btb_rd_addr_p1_f == 8'hb; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4683 = _T_4182 ? btb_bank0_rd_data_way0_out_11 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4938 = _T_4937 | _T_4683; // @[Mux.scala 27:72]
  wire  _T_4184 = btb_rd_addr_p1_f == 8'hc; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4684 = _T_4184 ? btb_bank0_rd_data_way0_out_12 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4939 = _T_4938 | _T_4684; // @[Mux.scala 27:72]
  wire  _T_4186 = btb_rd_addr_p1_f == 8'hd; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4685 = _T_4186 ? btb_bank0_rd_data_way0_out_13 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4940 = _T_4939 | _T_4685; // @[Mux.scala 27:72]
  wire  _T_4188 = btb_rd_addr_p1_f == 8'he; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4686 = _T_4188 ? btb_bank0_rd_data_way0_out_14 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4941 = _T_4940 | _T_4686; // @[Mux.scala 27:72]
  wire  _T_4190 = btb_rd_addr_p1_f == 8'hf; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4687 = _T_4190 ? btb_bank0_rd_data_way0_out_15 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4942 = _T_4941 | _T_4687; // @[Mux.scala 27:72]
  wire  _T_4192 = btb_rd_addr_p1_f == 8'h10; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4688 = _T_4192 ? btb_bank0_rd_data_way0_out_16 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4943 = _T_4942 | _T_4688; // @[Mux.scala 27:72]
  wire  _T_4194 = btb_rd_addr_p1_f == 8'h11; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4689 = _T_4194 ? btb_bank0_rd_data_way0_out_17 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4944 = _T_4943 | _T_4689; // @[Mux.scala 27:72]
  wire  _T_4196 = btb_rd_addr_p1_f == 8'h12; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4690 = _T_4196 ? btb_bank0_rd_data_way0_out_18 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4945 = _T_4944 | _T_4690; // @[Mux.scala 27:72]
  wire  _T_4198 = btb_rd_addr_p1_f == 8'h13; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4691 = _T_4198 ? btb_bank0_rd_data_way0_out_19 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4946 = _T_4945 | _T_4691; // @[Mux.scala 27:72]
  wire  _T_4200 = btb_rd_addr_p1_f == 8'h14; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4692 = _T_4200 ? btb_bank0_rd_data_way0_out_20 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4947 = _T_4946 | _T_4692; // @[Mux.scala 27:72]
  wire  _T_4202 = btb_rd_addr_p1_f == 8'h15; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4693 = _T_4202 ? btb_bank0_rd_data_way0_out_21 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4948 = _T_4947 | _T_4693; // @[Mux.scala 27:72]
  wire  _T_4204 = btb_rd_addr_p1_f == 8'h16; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4694 = _T_4204 ? btb_bank0_rd_data_way0_out_22 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4949 = _T_4948 | _T_4694; // @[Mux.scala 27:72]
  wire  _T_4206 = btb_rd_addr_p1_f == 8'h17; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4695 = _T_4206 ? btb_bank0_rd_data_way0_out_23 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4950 = _T_4949 | _T_4695; // @[Mux.scala 27:72]
  wire  _T_4208 = btb_rd_addr_p1_f == 8'h18; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4696 = _T_4208 ? btb_bank0_rd_data_way0_out_24 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4951 = _T_4950 | _T_4696; // @[Mux.scala 27:72]
  wire  _T_4210 = btb_rd_addr_p1_f == 8'h19; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4697 = _T_4210 ? btb_bank0_rd_data_way0_out_25 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4952 = _T_4951 | _T_4697; // @[Mux.scala 27:72]
  wire  _T_4212 = btb_rd_addr_p1_f == 8'h1a; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4698 = _T_4212 ? btb_bank0_rd_data_way0_out_26 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4953 = _T_4952 | _T_4698; // @[Mux.scala 27:72]
  wire  _T_4214 = btb_rd_addr_p1_f == 8'h1b; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4699 = _T_4214 ? btb_bank0_rd_data_way0_out_27 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4954 = _T_4953 | _T_4699; // @[Mux.scala 27:72]
  wire  _T_4216 = btb_rd_addr_p1_f == 8'h1c; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4700 = _T_4216 ? btb_bank0_rd_data_way0_out_28 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4955 = _T_4954 | _T_4700; // @[Mux.scala 27:72]
  wire  _T_4218 = btb_rd_addr_p1_f == 8'h1d; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4701 = _T_4218 ? btb_bank0_rd_data_way0_out_29 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4956 = _T_4955 | _T_4701; // @[Mux.scala 27:72]
  wire  _T_4220 = btb_rd_addr_p1_f == 8'h1e; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4702 = _T_4220 ? btb_bank0_rd_data_way0_out_30 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4957 = _T_4956 | _T_4702; // @[Mux.scala 27:72]
  wire  _T_4222 = btb_rd_addr_p1_f == 8'h1f; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4703 = _T_4222 ? btb_bank0_rd_data_way0_out_31 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4958 = _T_4957 | _T_4703; // @[Mux.scala 27:72]
  wire  _T_4224 = btb_rd_addr_p1_f == 8'h20; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4704 = _T_4224 ? btb_bank0_rd_data_way0_out_32 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4959 = _T_4958 | _T_4704; // @[Mux.scala 27:72]
  wire  _T_4226 = btb_rd_addr_p1_f == 8'h21; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4705 = _T_4226 ? btb_bank0_rd_data_way0_out_33 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4960 = _T_4959 | _T_4705; // @[Mux.scala 27:72]
  wire  _T_4228 = btb_rd_addr_p1_f == 8'h22; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4706 = _T_4228 ? btb_bank0_rd_data_way0_out_34 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4961 = _T_4960 | _T_4706; // @[Mux.scala 27:72]
  wire  _T_4230 = btb_rd_addr_p1_f == 8'h23; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4707 = _T_4230 ? btb_bank0_rd_data_way0_out_35 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4962 = _T_4961 | _T_4707; // @[Mux.scala 27:72]
  wire  _T_4232 = btb_rd_addr_p1_f == 8'h24; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4708 = _T_4232 ? btb_bank0_rd_data_way0_out_36 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4963 = _T_4962 | _T_4708; // @[Mux.scala 27:72]
  wire  _T_4234 = btb_rd_addr_p1_f == 8'h25; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4709 = _T_4234 ? btb_bank0_rd_data_way0_out_37 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4964 = _T_4963 | _T_4709; // @[Mux.scala 27:72]
  wire  _T_4236 = btb_rd_addr_p1_f == 8'h26; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4710 = _T_4236 ? btb_bank0_rd_data_way0_out_38 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4965 = _T_4964 | _T_4710; // @[Mux.scala 27:72]
  wire  _T_4238 = btb_rd_addr_p1_f == 8'h27; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4711 = _T_4238 ? btb_bank0_rd_data_way0_out_39 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4966 = _T_4965 | _T_4711; // @[Mux.scala 27:72]
  wire  _T_4240 = btb_rd_addr_p1_f == 8'h28; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4712 = _T_4240 ? btb_bank0_rd_data_way0_out_40 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4967 = _T_4966 | _T_4712; // @[Mux.scala 27:72]
  wire  _T_4242 = btb_rd_addr_p1_f == 8'h29; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4713 = _T_4242 ? btb_bank0_rd_data_way0_out_41 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4968 = _T_4967 | _T_4713; // @[Mux.scala 27:72]
  wire  _T_4244 = btb_rd_addr_p1_f == 8'h2a; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4714 = _T_4244 ? btb_bank0_rd_data_way0_out_42 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4969 = _T_4968 | _T_4714; // @[Mux.scala 27:72]
  wire  _T_4246 = btb_rd_addr_p1_f == 8'h2b; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4715 = _T_4246 ? btb_bank0_rd_data_way0_out_43 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4970 = _T_4969 | _T_4715; // @[Mux.scala 27:72]
  wire  _T_4248 = btb_rd_addr_p1_f == 8'h2c; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4716 = _T_4248 ? btb_bank0_rd_data_way0_out_44 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4971 = _T_4970 | _T_4716; // @[Mux.scala 27:72]
  wire  _T_4250 = btb_rd_addr_p1_f == 8'h2d; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4717 = _T_4250 ? btb_bank0_rd_data_way0_out_45 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4972 = _T_4971 | _T_4717; // @[Mux.scala 27:72]
  wire  _T_4252 = btb_rd_addr_p1_f == 8'h2e; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4718 = _T_4252 ? btb_bank0_rd_data_way0_out_46 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4973 = _T_4972 | _T_4718; // @[Mux.scala 27:72]
  wire  _T_4254 = btb_rd_addr_p1_f == 8'h2f; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4719 = _T_4254 ? btb_bank0_rd_data_way0_out_47 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4974 = _T_4973 | _T_4719; // @[Mux.scala 27:72]
  wire  _T_4256 = btb_rd_addr_p1_f == 8'h30; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4720 = _T_4256 ? btb_bank0_rd_data_way0_out_48 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4975 = _T_4974 | _T_4720; // @[Mux.scala 27:72]
  wire  _T_4258 = btb_rd_addr_p1_f == 8'h31; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4721 = _T_4258 ? btb_bank0_rd_data_way0_out_49 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4976 = _T_4975 | _T_4721; // @[Mux.scala 27:72]
  wire  _T_4260 = btb_rd_addr_p1_f == 8'h32; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4722 = _T_4260 ? btb_bank0_rd_data_way0_out_50 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4977 = _T_4976 | _T_4722; // @[Mux.scala 27:72]
  wire  _T_4262 = btb_rd_addr_p1_f == 8'h33; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4723 = _T_4262 ? btb_bank0_rd_data_way0_out_51 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4978 = _T_4977 | _T_4723; // @[Mux.scala 27:72]
  wire  _T_4264 = btb_rd_addr_p1_f == 8'h34; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4724 = _T_4264 ? btb_bank0_rd_data_way0_out_52 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4979 = _T_4978 | _T_4724; // @[Mux.scala 27:72]
  wire  _T_4266 = btb_rd_addr_p1_f == 8'h35; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4725 = _T_4266 ? btb_bank0_rd_data_way0_out_53 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4980 = _T_4979 | _T_4725; // @[Mux.scala 27:72]
  wire  _T_4268 = btb_rd_addr_p1_f == 8'h36; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4726 = _T_4268 ? btb_bank0_rd_data_way0_out_54 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4981 = _T_4980 | _T_4726; // @[Mux.scala 27:72]
  wire  _T_4270 = btb_rd_addr_p1_f == 8'h37; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4727 = _T_4270 ? btb_bank0_rd_data_way0_out_55 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4982 = _T_4981 | _T_4727; // @[Mux.scala 27:72]
  wire  _T_4272 = btb_rd_addr_p1_f == 8'h38; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4728 = _T_4272 ? btb_bank0_rd_data_way0_out_56 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4983 = _T_4982 | _T_4728; // @[Mux.scala 27:72]
  wire  _T_4274 = btb_rd_addr_p1_f == 8'h39; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4729 = _T_4274 ? btb_bank0_rd_data_way0_out_57 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4984 = _T_4983 | _T_4729; // @[Mux.scala 27:72]
  wire  _T_4276 = btb_rd_addr_p1_f == 8'h3a; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4730 = _T_4276 ? btb_bank0_rd_data_way0_out_58 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4985 = _T_4984 | _T_4730; // @[Mux.scala 27:72]
  wire  _T_4278 = btb_rd_addr_p1_f == 8'h3b; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4731 = _T_4278 ? btb_bank0_rd_data_way0_out_59 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4986 = _T_4985 | _T_4731; // @[Mux.scala 27:72]
  wire  _T_4280 = btb_rd_addr_p1_f == 8'h3c; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4732 = _T_4280 ? btb_bank0_rd_data_way0_out_60 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4987 = _T_4986 | _T_4732; // @[Mux.scala 27:72]
  wire  _T_4282 = btb_rd_addr_p1_f == 8'h3d; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4733 = _T_4282 ? btb_bank0_rd_data_way0_out_61 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4988 = _T_4987 | _T_4733; // @[Mux.scala 27:72]
  wire  _T_4284 = btb_rd_addr_p1_f == 8'h3e; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4734 = _T_4284 ? btb_bank0_rd_data_way0_out_62 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4989 = _T_4988 | _T_4734; // @[Mux.scala 27:72]
  wire  _T_4286 = btb_rd_addr_p1_f == 8'h3f; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4735 = _T_4286 ? btb_bank0_rd_data_way0_out_63 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4990 = _T_4989 | _T_4735; // @[Mux.scala 27:72]
  wire  _T_4288 = btb_rd_addr_p1_f == 8'h40; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4736 = _T_4288 ? btb_bank0_rd_data_way0_out_64 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4991 = _T_4990 | _T_4736; // @[Mux.scala 27:72]
  wire  _T_4290 = btb_rd_addr_p1_f == 8'h41; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4737 = _T_4290 ? btb_bank0_rd_data_way0_out_65 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4992 = _T_4991 | _T_4737; // @[Mux.scala 27:72]
  wire  _T_4292 = btb_rd_addr_p1_f == 8'h42; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4738 = _T_4292 ? btb_bank0_rd_data_way0_out_66 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4993 = _T_4992 | _T_4738; // @[Mux.scala 27:72]
  wire  _T_4294 = btb_rd_addr_p1_f == 8'h43; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4739 = _T_4294 ? btb_bank0_rd_data_way0_out_67 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4994 = _T_4993 | _T_4739; // @[Mux.scala 27:72]
  wire  _T_4296 = btb_rd_addr_p1_f == 8'h44; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4740 = _T_4296 ? btb_bank0_rd_data_way0_out_68 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4995 = _T_4994 | _T_4740; // @[Mux.scala 27:72]
  wire  _T_4298 = btb_rd_addr_p1_f == 8'h45; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4741 = _T_4298 ? btb_bank0_rd_data_way0_out_69 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4996 = _T_4995 | _T_4741; // @[Mux.scala 27:72]
  wire  _T_4300 = btb_rd_addr_p1_f == 8'h46; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4742 = _T_4300 ? btb_bank0_rd_data_way0_out_70 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4997 = _T_4996 | _T_4742; // @[Mux.scala 27:72]
  wire  _T_4302 = btb_rd_addr_p1_f == 8'h47; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4743 = _T_4302 ? btb_bank0_rd_data_way0_out_71 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4998 = _T_4997 | _T_4743; // @[Mux.scala 27:72]
  wire  _T_4304 = btb_rd_addr_p1_f == 8'h48; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4744 = _T_4304 ? btb_bank0_rd_data_way0_out_72 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4999 = _T_4998 | _T_4744; // @[Mux.scala 27:72]
  wire  _T_4306 = btb_rd_addr_p1_f == 8'h49; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4745 = _T_4306 ? btb_bank0_rd_data_way0_out_73 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5000 = _T_4999 | _T_4745; // @[Mux.scala 27:72]
  wire  _T_4308 = btb_rd_addr_p1_f == 8'h4a; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4746 = _T_4308 ? btb_bank0_rd_data_way0_out_74 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5001 = _T_5000 | _T_4746; // @[Mux.scala 27:72]
  wire  _T_4310 = btb_rd_addr_p1_f == 8'h4b; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4747 = _T_4310 ? btb_bank0_rd_data_way0_out_75 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5002 = _T_5001 | _T_4747; // @[Mux.scala 27:72]
  wire  _T_4312 = btb_rd_addr_p1_f == 8'h4c; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4748 = _T_4312 ? btb_bank0_rd_data_way0_out_76 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5003 = _T_5002 | _T_4748; // @[Mux.scala 27:72]
  wire  _T_4314 = btb_rd_addr_p1_f == 8'h4d; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4749 = _T_4314 ? btb_bank0_rd_data_way0_out_77 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5004 = _T_5003 | _T_4749; // @[Mux.scala 27:72]
  wire  _T_4316 = btb_rd_addr_p1_f == 8'h4e; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4750 = _T_4316 ? btb_bank0_rd_data_way0_out_78 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5005 = _T_5004 | _T_4750; // @[Mux.scala 27:72]
  wire  _T_4318 = btb_rd_addr_p1_f == 8'h4f; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4751 = _T_4318 ? btb_bank0_rd_data_way0_out_79 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5006 = _T_5005 | _T_4751; // @[Mux.scala 27:72]
  wire  _T_4320 = btb_rd_addr_p1_f == 8'h50; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4752 = _T_4320 ? btb_bank0_rd_data_way0_out_80 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5007 = _T_5006 | _T_4752; // @[Mux.scala 27:72]
  wire  _T_4322 = btb_rd_addr_p1_f == 8'h51; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4753 = _T_4322 ? btb_bank0_rd_data_way0_out_81 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5008 = _T_5007 | _T_4753; // @[Mux.scala 27:72]
  wire  _T_4324 = btb_rd_addr_p1_f == 8'h52; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4754 = _T_4324 ? btb_bank0_rd_data_way0_out_82 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5009 = _T_5008 | _T_4754; // @[Mux.scala 27:72]
  wire  _T_4326 = btb_rd_addr_p1_f == 8'h53; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4755 = _T_4326 ? btb_bank0_rd_data_way0_out_83 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5010 = _T_5009 | _T_4755; // @[Mux.scala 27:72]
  wire  _T_4328 = btb_rd_addr_p1_f == 8'h54; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4756 = _T_4328 ? btb_bank0_rd_data_way0_out_84 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5011 = _T_5010 | _T_4756; // @[Mux.scala 27:72]
  wire  _T_4330 = btb_rd_addr_p1_f == 8'h55; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4757 = _T_4330 ? btb_bank0_rd_data_way0_out_85 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5012 = _T_5011 | _T_4757; // @[Mux.scala 27:72]
  wire  _T_4332 = btb_rd_addr_p1_f == 8'h56; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4758 = _T_4332 ? btb_bank0_rd_data_way0_out_86 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5013 = _T_5012 | _T_4758; // @[Mux.scala 27:72]
  wire  _T_4334 = btb_rd_addr_p1_f == 8'h57; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4759 = _T_4334 ? btb_bank0_rd_data_way0_out_87 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5014 = _T_5013 | _T_4759; // @[Mux.scala 27:72]
  wire  _T_4336 = btb_rd_addr_p1_f == 8'h58; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4760 = _T_4336 ? btb_bank0_rd_data_way0_out_88 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5015 = _T_5014 | _T_4760; // @[Mux.scala 27:72]
  wire  _T_4338 = btb_rd_addr_p1_f == 8'h59; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4761 = _T_4338 ? btb_bank0_rd_data_way0_out_89 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5016 = _T_5015 | _T_4761; // @[Mux.scala 27:72]
  wire  _T_4340 = btb_rd_addr_p1_f == 8'h5a; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4762 = _T_4340 ? btb_bank0_rd_data_way0_out_90 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5017 = _T_5016 | _T_4762; // @[Mux.scala 27:72]
  wire  _T_4342 = btb_rd_addr_p1_f == 8'h5b; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4763 = _T_4342 ? btb_bank0_rd_data_way0_out_91 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5018 = _T_5017 | _T_4763; // @[Mux.scala 27:72]
  wire  _T_4344 = btb_rd_addr_p1_f == 8'h5c; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4764 = _T_4344 ? btb_bank0_rd_data_way0_out_92 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5019 = _T_5018 | _T_4764; // @[Mux.scala 27:72]
  wire  _T_4346 = btb_rd_addr_p1_f == 8'h5d; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4765 = _T_4346 ? btb_bank0_rd_data_way0_out_93 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5020 = _T_5019 | _T_4765; // @[Mux.scala 27:72]
  wire  _T_4348 = btb_rd_addr_p1_f == 8'h5e; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4766 = _T_4348 ? btb_bank0_rd_data_way0_out_94 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5021 = _T_5020 | _T_4766; // @[Mux.scala 27:72]
  wire  _T_4350 = btb_rd_addr_p1_f == 8'h5f; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4767 = _T_4350 ? btb_bank0_rd_data_way0_out_95 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5022 = _T_5021 | _T_4767; // @[Mux.scala 27:72]
  wire  _T_4352 = btb_rd_addr_p1_f == 8'h60; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4768 = _T_4352 ? btb_bank0_rd_data_way0_out_96 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5023 = _T_5022 | _T_4768; // @[Mux.scala 27:72]
  wire  _T_4354 = btb_rd_addr_p1_f == 8'h61; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4769 = _T_4354 ? btb_bank0_rd_data_way0_out_97 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5024 = _T_5023 | _T_4769; // @[Mux.scala 27:72]
  wire  _T_4356 = btb_rd_addr_p1_f == 8'h62; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4770 = _T_4356 ? btb_bank0_rd_data_way0_out_98 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5025 = _T_5024 | _T_4770; // @[Mux.scala 27:72]
  wire  _T_4358 = btb_rd_addr_p1_f == 8'h63; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4771 = _T_4358 ? btb_bank0_rd_data_way0_out_99 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5026 = _T_5025 | _T_4771; // @[Mux.scala 27:72]
  wire  _T_4360 = btb_rd_addr_p1_f == 8'h64; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4772 = _T_4360 ? btb_bank0_rd_data_way0_out_100 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5027 = _T_5026 | _T_4772; // @[Mux.scala 27:72]
  wire  _T_4362 = btb_rd_addr_p1_f == 8'h65; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4773 = _T_4362 ? btb_bank0_rd_data_way0_out_101 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5028 = _T_5027 | _T_4773; // @[Mux.scala 27:72]
  wire  _T_4364 = btb_rd_addr_p1_f == 8'h66; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4774 = _T_4364 ? btb_bank0_rd_data_way0_out_102 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5029 = _T_5028 | _T_4774; // @[Mux.scala 27:72]
  wire  _T_4366 = btb_rd_addr_p1_f == 8'h67; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4775 = _T_4366 ? btb_bank0_rd_data_way0_out_103 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5030 = _T_5029 | _T_4775; // @[Mux.scala 27:72]
  wire  _T_4368 = btb_rd_addr_p1_f == 8'h68; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4776 = _T_4368 ? btb_bank0_rd_data_way0_out_104 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5031 = _T_5030 | _T_4776; // @[Mux.scala 27:72]
  wire  _T_4370 = btb_rd_addr_p1_f == 8'h69; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4777 = _T_4370 ? btb_bank0_rd_data_way0_out_105 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5032 = _T_5031 | _T_4777; // @[Mux.scala 27:72]
  wire  _T_4372 = btb_rd_addr_p1_f == 8'h6a; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4778 = _T_4372 ? btb_bank0_rd_data_way0_out_106 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5033 = _T_5032 | _T_4778; // @[Mux.scala 27:72]
  wire  _T_4374 = btb_rd_addr_p1_f == 8'h6b; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4779 = _T_4374 ? btb_bank0_rd_data_way0_out_107 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5034 = _T_5033 | _T_4779; // @[Mux.scala 27:72]
  wire  _T_4376 = btb_rd_addr_p1_f == 8'h6c; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4780 = _T_4376 ? btb_bank0_rd_data_way0_out_108 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5035 = _T_5034 | _T_4780; // @[Mux.scala 27:72]
  wire  _T_4378 = btb_rd_addr_p1_f == 8'h6d; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4781 = _T_4378 ? btb_bank0_rd_data_way0_out_109 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5036 = _T_5035 | _T_4781; // @[Mux.scala 27:72]
  wire  _T_4380 = btb_rd_addr_p1_f == 8'h6e; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4782 = _T_4380 ? btb_bank0_rd_data_way0_out_110 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5037 = _T_5036 | _T_4782; // @[Mux.scala 27:72]
  wire  _T_4382 = btb_rd_addr_p1_f == 8'h6f; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4783 = _T_4382 ? btb_bank0_rd_data_way0_out_111 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5038 = _T_5037 | _T_4783; // @[Mux.scala 27:72]
  wire  _T_4384 = btb_rd_addr_p1_f == 8'h70; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4784 = _T_4384 ? btb_bank0_rd_data_way0_out_112 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5039 = _T_5038 | _T_4784; // @[Mux.scala 27:72]
  wire  _T_4386 = btb_rd_addr_p1_f == 8'h71; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4785 = _T_4386 ? btb_bank0_rd_data_way0_out_113 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5040 = _T_5039 | _T_4785; // @[Mux.scala 27:72]
  wire  _T_4388 = btb_rd_addr_p1_f == 8'h72; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4786 = _T_4388 ? btb_bank0_rd_data_way0_out_114 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5041 = _T_5040 | _T_4786; // @[Mux.scala 27:72]
  wire  _T_4390 = btb_rd_addr_p1_f == 8'h73; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4787 = _T_4390 ? btb_bank0_rd_data_way0_out_115 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5042 = _T_5041 | _T_4787; // @[Mux.scala 27:72]
  wire  _T_4392 = btb_rd_addr_p1_f == 8'h74; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4788 = _T_4392 ? btb_bank0_rd_data_way0_out_116 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5043 = _T_5042 | _T_4788; // @[Mux.scala 27:72]
  wire  _T_4394 = btb_rd_addr_p1_f == 8'h75; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4789 = _T_4394 ? btb_bank0_rd_data_way0_out_117 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5044 = _T_5043 | _T_4789; // @[Mux.scala 27:72]
  wire  _T_4396 = btb_rd_addr_p1_f == 8'h76; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4790 = _T_4396 ? btb_bank0_rd_data_way0_out_118 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5045 = _T_5044 | _T_4790; // @[Mux.scala 27:72]
  wire  _T_4398 = btb_rd_addr_p1_f == 8'h77; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4791 = _T_4398 ? btb_bank0_rd_data_way0_out_119 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5046 = _T_5045 | _T_4791; // @[Mux.scala 27:72]
  wire  _T_4400 = btb_rd_addr_p1_f == 8'h78; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4792 = _T_4400 ? btb_bank0_rd_data_way0_out_120 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5047 = _T_5046 | _T_4792; // @[Mux.scala 27:72]
  wire  _T_4402 = btb_rd_addr_p1_f == 8'h79; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4793 = _T_4402 ? btb_bank0_rd_data_way0_out_121 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5048 = _T_5047 | _T_4793; // @[Mux.scala 27:72]
  wire  _T_4404 = btb_rd_addr_p1_f == 8'h7a; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4794 = _T_4404 ? btb_bank0_rd_data_way0_out_122 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5049 = _T_5048 | _T_4794; // @[Mux.scala 27:72]
  wire  _T_4406 = btb_rd_addr_p1_f == 8'h7b; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4795 = _T_4406 ? btb_bank0_rd_data_way0_out_123 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5050 = _T_5049 | _T_4795; // @[Mux.scala 27:72]
  wire  _T_4408 = btb_rd_addr_p1_f == 8'h7c; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4796 = _T_4408 ? btb_bank0_rd_data_way0_out_124 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5051 = _T_5050 | _T_4796; // @[Mux.scala 27:72]
  wire  _T_4410 = btb_rd_addr_p1_f == 8'h7d; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4797 = _T_4410 ? btb_bank0_rd_data_way0_out_125 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5052 = _T_5051 | _T_4797; // @[Mux.scala 27:72]
  wire  _T_4412 = btb_rd_addr_p1_f == 8'h7e; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4798 = _T_4412 ? btb_bank0_rd_data_way0_out_126 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5053 = _T_5052 | _T_4798; // @[Mux.scala 27:72]
  wire  _T_4414 = btb_rd_addr_p1_f == 8'h7f; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4799 = _T_4414 ? btb_bank0_rd_data_way0_out_127 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5054 = _T_5053 | _T_4799; // @[Mux.scala 27:72]
  wire  _T_4416 = btb_rd_addr_p1_f == 8'h80; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4800 = _T_4416 ? btb_bank0_rd_data_way0_out_128 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5055 = _T_5054 | _T_4800; // @[Mux.scala 27:72]
  wire  _T_4418 = btb_rd_addr_p1_f == 8'h81; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4801 = _T_4418 ? btb_bank0_rd_data_way0_out_129 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5056 = _T_5055 | _T_4801; // @[Mux.scala 27:72]
  wire  _T_4420 = btb_rd_addr_p1_f == 8'h82; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4802 = _T_4420 ? btb_bank0_rd_data_way0_out_130 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5057 = _T_5056 | _T_4802; // @[Mux.scala 27:72]
  wire  _T_4422 = btb_rd_addr_p1_f == 8'h83; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4803 = _T_4422 ? btb_bank0_rd_data_way0_out_131 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5058 = _T_5057 | _T_4803; // @[Mux.scala 27:72]
  wire  _T_4424 = btb_rd_addr_p1_f == 8'h84; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4804 = _T_4424 ? btb_bank0_rd_data_way0_out_132 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5059 = _T_5058 | _T_4804; // @[Mux.scala 27:72]
  wire  _T_4426 = btb_rd_addr_p1_f == 8'h85; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4805 = _T_4426 ? btb_bank0_rd_data_way0_out_133 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5060 = _T_5059 | _T_4805; // @[Mux.scala 27:72]
  wire  _T_4428 = btb_rd_addr_p1_f == 8'h86; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4806 = _T_4428 ? btb_bank0_rd_data_way0_out_134 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5061 = _T_5060 | _T_4806; // @[Mux.scala 27:72]
  wire  _T_4430 = btb_rd_addr_p1_f == 8'h87; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4807 = _T_4430 ? btb_bank0_rd_data_way0_out_135 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5062 = _T_5061 | _T_4807; // @[Mux.scala 27:72]
  wire  _T_4432 = btb_rd_addr_p1_f == 8'h88; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4808 = _T_4432 ? btb_bank0_rd_data_way0_out_136 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5063 = _T_5062 | _T_4808; // @[Mux.scala 27:72]
  wire  _T_4434 = btb_rd_addr_p1_f == 8'h89; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4809 = _T_4434 ? btb_bank0_rd_data_way0_out_137 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5064 = _T_5063 | _T_4809; // @[Mux.scala 27:72]
  wire  _T_4436 = btb_rd_addr_p1_f == 8'h8a; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4810 = _T_4436 ? btb_bank0_rd_data_way0_out_138 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5065 = _T_5064 | _T_4810; // @[Mux.scala 27:72]
  wire  _T_4438 = btb_rd_addr_p1_f == 8'h8b; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4811 = _T_4438 ? btb_bank0_rd_data_way0_out_139 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5066 = _T_5065 | _T_4811; // @[Mux.scala 27:72]
  wire  _T_4440 = btb_rd_addr_p1_f == 8'h8c; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4812 = _T_4440 ? btb_bank0_rd_data_way0_out_140 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5067 = _T_5066 | _T_4812; // @[Mux.scala 27:72]
  wire  _T_4442 = btb_rd_addr_p1_f == 8'h8d; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4813 = _T_4442 ? btb_bank0_rd_data_way0_out_141 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5068 = _T_5067 | _T_4813; // @[Mux.scala 27:72]
  wire  _T_4444 = btb_rd_addr_p1_f == 8'h8e; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4814 = _T_4444 ? btb_bank0_rd_data_way0_out_142 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5069 = _T_5068 | _T_4814; // @[Mux.scala 27:72]
  wire  _T_4446 = btb_rd_addr_p1_f == 8'h8f; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4815 = _T_4446 ? btb_bank0_rd_data_way0_out_143 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5070 = _T_5069 | _T_4815; // @[Mux.scala 27:72]
  wire  _T_4448 = btb_rd_addr_p1_f == 8'h90; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4816 = _T_4448 ? btb_bank0_rd_data_way0_out_144 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5071 = _T_5070 | _T_4816; // @[Mux.scala 27:72]
  wire  _T_4450 = btb_rd_addr_p1_f == 8'h91; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4817 = _T_4450 ? btb_bank0_rd_data_way0_out_145 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5072 = _T_5071 | _T_4817; // @[Mux.scala 27:72]
  wire  _T_4452 = btb_rd_addr_p1_f == 8'h92; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4818 = _T_4452 ? btb_bank0_rd_data_way0_out_146 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5073 = _T_5072 | _T_4818; // @[Mux.scala 27:72]
  wire  _T_4454 = btb_rd_addr_p1_f == 8'h93; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4819 = _T_4454 ? btb_bank0_rd_data_way0_out_147 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5074 = _T_5073 | _T_4819; // @[Mux.scala 27:72]
  wire  _T_4456 = btb_rd_addr_p1_f == 8'h94; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4820 = _T_4456 ? btb_bank0_rd_data_way0_out_148 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5075 = _T_5074 | _T_4820; // @[Mux.scala 27:72]
  wire  _T_4458 = btb_rd_addr_p1_f == 8'h95; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4821 = _T_4458 ? btb_bank0_rd_data_way0_out_149 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5076 = _T_5075 | _T_4821; // @[Mux.scala 27:72]
  wire  _T_4460 = btb_rd_addr_p1_f == 8'h96; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4822 = _T_4460 ? btb_bank0_rd_data_way0_out_150 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5077 = _T_5076 | _T_4822; // @[Mux.scala 27:72]
  wire  _T_4462 = btb_rd_addr_p1_f == 8'h97; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4823 = _T_4462 ? btb_bank0_rd_data_way0_out_151 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5078 = _T_5077 | _T_4823; // @[Mux.scala 27:72]
  wire  _T_4464 = btb_rd_addr_p1_f == 8'h98; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4824 = _T_4464 ? btb_bank0_rd_data_way0_out_152 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5079 = _T_5078 | _T_4824; // @[Mux.scala 27:72]
  wire  _T_4466 = btb_rd_addr_p1_f == 8'h99; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4825 = _T_4466 ? btb_bank0_rd_data_way0_out_153 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5080 = _T_5079 | _T_4825; // @[Mux.scala 27:72]
  wire  _T_4468 = btb_rd_addr_p1_f == 8'h9a; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4826 = _T_4468 ? btb_bank0_rd_data_way0_out_154 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5081 = _T_5080 | _T_4826; // @[Mux.scala 27:72]
  wire  _T_4470 = btb_rd_addr_p1_f == 8'h9b; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4827 = _T_4470 ? btb_bank0_rd_data_way0_out_155 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5082 = _T_5081 | _T_4827; // @[Mux.scala 27:72]
  wire  _T_4472 = btb_rd_addr_p1_f == 8'h9c; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4828 = _T_4472 ? btb_bank0_rd_data_way0_out_156 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5083 = _T_5082 | _T_4828; // @[Mux.scala 27:72]
  wire  _T_4474 = btb_rd_addr_p1_f == 8'h9d; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4829 = _T_4474 ? btb_bank0_rd_data_way0_out_157 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5084 = _T_5083 | _T_4829; // @[Mux.scala 27:72]
  wire  _T_4476 = btb_rd_addr_p1_f == 8'h9e; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4830 = _T_4476 ? btb_bank0_rd_data_way0_out_158 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5085 = _T_5084 | _T_4830; // @[Mux.scala 27:72]
  wire  _T_4478 = btb_rd_addr_p1_f == 8'h9f; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4831 = _T_4478 ? btb_bank0_rd_data_way0_out_159 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5086 = _T_5085 | _T_4831; // @[Mux.scala 27:72]
  wire  _T_4480 = btb_rd_addr_p1_f == 8'ha0; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4832 = _T_4480 ? btb_bank0_rd_data_way0_out_160 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5087 = _T_5086 | _T_4832; // @[Mux.scala 27:72]
  wire  _T_4482 = btb_rd_addr_p1_f == 8'ha1; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4833 = _T_4482 ? btb_bank0_rd_data_way0_out_161 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5088 = _T_5087 | _T_4833; // @[Mux.scala 27:72]
  wire  _T_4484 = btb_rd_addr_p1_f == 8'ha2; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4834 = _T_4484 ? btb_bank0_rd_data_way0_out_162 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5089 = _T_5088 | _T_4834; // @[Mux.scala 27:72]
  wire  _T_4486 = btb_rd_addr_p1_f == 8'ha3; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4835 = _T_4486 ? btb_bank0_rd_data_way0_out_163 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5090 = _T_5089 | _T_4835; // @[Mux.scala 27:72]
  wire  _T_4488 = btb_rd_addr_p1_f == 8'ha4; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4836 = _T_4488 ? btb_bank0_rd_data_way0_out_164 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5091 = _T_5090 | _T_4836; // @[Mux.scala 27:72]
  wire  _T_4490 = btb_rd_addr_p1_f == 8'ha5; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4837 = _T_4490 ? btb_bank0_rd_data_way0_out_165 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5092 = _T_5091 | _T_4837; // @[Mux.scala 27:72]
  wire  _T_4492 = btb_rd_addr_p1_f == 8'ha6; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4838 = _T_4492 ? btb_bank0_rd_data_way0_out_166 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5093 = _T_5092 | _T_4838; // @[Mux.scala 27:72]
  wire  _T_4494 = btb_rd_addr_p1_f == 8'ha7; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4839 = _T_4494 ? btb_bank0_rd_data_way0_out_167 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5094 = _T_5093 | _T_4839; // @[Mux.scala 27:72]
  wire  _T_4496 = btb_rd_addr_p1_f == 8'ha8; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4840 = _T_4496 ? btb_bank0_rd_data_way0_out_168 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5095 = _T_5094 | _T_4840; // @[Mux.scala 27:72]
  wire  _T_4498 = btb_rd_addr_p1_f == 8'ha9; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4841 = _T_4498 ? btb_bank0_rd_data_way0_out_169 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5096 = _T_5095 | _T_4841; // @[Mux.scala 27:72]
  wire  _T_4500 = btb_rd_addr_p1_f == 8'haa; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4842 = _T_4500 ? btb_bank0_rd_data_way0_out_170 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5097 = _T_5096 | _T_4842; // @[Mux.scala 27:72]
  wire  _T_4502 = btb_rd_addr_p1_f == 8'hab; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4843 = _T_4502 ? btb_bank0_rd_data_way0_out_171 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5098 = _T_5097 | _T_4843; // @[Mux.scala 27:72]
  wire  _T_4504 = btb_rd_addr_p1_f == 8'hac; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4844 = _T_4504 ? btb_bank0_rd_data_way0_out_172 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5099 = _T_5098 | _T_4844; // @[Mux.scala 27:72]
  wire  _T_4506 = btb_rd_addr_p1_f == 8'had; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4845 = _T_4506 ? btb_bank0_rd_data_way0_out_173 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5100 = _T_5099 | _T_4845; // @[Mux.scala 27:72]
  wire  _T_4508 = btb_rd_addr_p1_f == 8'hae; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4846 = _T_4508 ? btb_bank0_rd_data_way0_out_174 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5101 = _T_5100 | _T_4846; // @[Mux.scala 27:72]
  wire  _T_4510 = btb_rd_addr_p1_f == 8'haf; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4847 = _T_4510 ? btb_bank0_rd_data_way0_out_175 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5102 = _T_5101 | _T_4847; // @[Mux.scala 27:72]
  wire  _T_4512 = btb_rd_addr_p1_f == 8'hb0; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4848 = _T_4512 ? btb_bank0_rd_data_way0_out_176 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5103 = _T_5102 | _T_4848; // @[Mux.scala 27:72]
  wire  _T_4514 = btb_rd_addr_p1_f == 8'hb1; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4849 = _T_4514 ? btb_bank0_rd_data_way0_out_177 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5104 = _T_5103 | _T_4849; // @[Mux.scala 27:72]
  wire  _T_4516 = btb_rd_addr_p1_f == 8'hb2; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4850 = _T_4516 ? btb_bank0_rd_data_way0_out_178 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5105 = _T_5104 | _T_4850; // @[Mux.scala 27:72]
  wire  _T_4518 = btb_rd_addr_p1_f == 8'hb3; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4851 = _T_4518 ? btb_bank0_rd_data_way0_out_179 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5106 = _T_5105 | _T_4851; // @[Mux.scala 27:72]
  wire  _T_4520 = btb_rd_addr_p1_f == 8'hb4; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4852 = _T_4520 ? btb_bank0_rd_data_way0_out_180 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5107 = _T_5106 | _T_4852; // @[Mux.scala 27:72]
  wire  _T_4522 = btb_rd_addr_p1_f == 8'hb5; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4853 = _T_4522 ? btb_bank0_rd_data_way0_out_181 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5108 = _T_5107 | _T_4853; // @[Mux.scala 27:72]
  wire  _T_4524 = btb_rd_addr_p1_f == 8'hb6; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4854 = _T_4524 ? btb_bank0_rd_data_way0_out_182 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5109 = _T_5108 | _T_4854; // @[Mux.scala 27:72]
  wire  _T_4526 = btb_rd_addr_p1_f == 8'hb7; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4855 = _T_4526 ? btb_bank0_rd_data_way0_out_183 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5110 = _T_5109 | _T_4855; // @[Mux.scala 27:72]
  wire  _T_4528 = btb_rd_addr_p1_f == 8'hb8; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4856 = _T_4528 ? btb_bank0_rd_data_way0_out_184 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5111 = _T_5110 | _T_4856; // @[Mux.scala 27:72]
  wire  _T_4530 = btb_rd_addr_p1_f == 8'hb9; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4857 = _T_4530 ? btb_bank0_rd_data_way0_out_185 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5112 = _T_5111 | _T_4857; // @[Mux.scala 27:72]
  wire  _T_4532 = btb_rd_addr_p1_f == 8'hba; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4858 = _T_4532 ? btb_bank0_rd_data_way0_out_186 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5113 = _T_5112 | _T_4858; // @[Mux.scala 27:72]
  wire  _T_4534 = btb_rd_addr_p1_f == 8'hbb; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4859 = _T_4534 ? btb_bank0_rd_data_way0_out_187 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5114 = _T_5113 | _T_4859; // @[Mux.scala 27:72]
  wire  _T_4536 = btb_rd_addr_p1_f == 8'hbc; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4860 = _T_4536 ? btb_bank0_rd_data_way0_out_188 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5115 = _T_5114 | _T_4860; // @[Mux.scala 27:72]
  wire  _T_4538 = btb_rd_addr_p1_f == 8'hbd; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4861 = _T_4538 ? btb_bank0_rd_data_way0_out_189 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5116 = _T_5115 | _T_4861; // @[Mux.scala 27:72]
  wire  _T_4540 = btb_rd_addr_p1_f == 8'hbe; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4862 = _T_4540 ? btb_bank0_rd_data_way0_out_190 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5117 = _T_5116 | _T_4862; // @[Mux.scala 27:72]
  wire  _T_4542 = btb_rd_addr_p1_f == 8'hbf; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4863 = _T_4542 ? btb_bank0_rd_data_way0_out_191 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5118 = _T_5117 | _T_4863; // @[Mux.scala 27:72]
  wire  _T_4544 = btb_rd_addr_p1_f == 8'hc0; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4864 = _T_4544 ? btb_bank0_rd_data_way0_out_192 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5119 = _T_5118 | _T_4864; // @[Mux.scala 27:72]
  wire  _T_4546 = btb_rd_addr_p1_f == 8'hc1; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4865 = _T_4546 ? btb_bank0_rd_data_way0_out_193 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5120 = _T_5119 | _T_4865; // @[Mux.scala 27:72]
  wire  _T_4548 = btb_rd_addr_p1_f == 8'hc2; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4866 = _T_4548 ? btb_bank0_rd_data_way0_out_194 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5121 = _T_5120 | _T_4866; // @[Mux.scala 27:72]
  wire  _T_4550 = btb_rd_addr_p1_f == 8'hc3; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4867 = _T_4550 ? btb_bank0_rd_data_way0_out_195 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5122 = _T_5121 | _T_4867; // @[Mux.scala 27:72]
  wire  _T_4552 = btb_rd_addr_p1_f == 8'hc4; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4868 = _T_4552 ? btb_bank0_rd_data_way0_out_196 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5123 = _T_5122 | _T_4868; // @[Mux.scala 27:72]
  wire  _T_4554 = btb_rd_addr_p1_f == 8'hc5; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4869 = _T_4554 ? btb_bank0_rd_data_way0_out_197 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5124 = _T_5123 | _T_4869; // @[Mux.scala 27:72]
  wire  _T_4556 = btb_rd_addr_p1_f == 8'hc6; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4870 = _T_4556 ? btb_bank0_rd_data_way0_out_198 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5125 = _T_5124 | _T_4870; // @[Mux.scala 27:72]
  wire  _T_4558 = btb_rd_addr_p1_f == 8'hc7; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4871 = _T_4558 ? btb_bank0_rd_data_way0_out_199 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5126 = _T_5125 | _T_4871; // @[Mux.scala 27:72]
  wire  _T_4560 = btb_rd_addr_p1_f == 8'hc8; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4872 = _T_4560 ? btb_bank0_rd_data_way0_out_200 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5127 = _T_5126 | _T_4872; // @[Mux.scala 27:72]
  wire  _T_4562 = btb_rd_addr_p1_f == 8'hc9; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4873 = _T_4562 ? btb_bank0_rd_data_way0_out_201 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5128 = _T_5127 | _T_4873; // @[Mux.scala 27:72]
  wire  _T_4564 = btb_rd_addr_p1_f == 8'hca; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4874 = _T_4564 ? btb_bank0_rd_data_way0_out_202 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5129 = _T_5128 | _T_4874; // @[Mux.scala 27:72]
  wire  _T_4566 = btb_rd_addr_p1_f == 8'hcb; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4875 = _T_4566 ? btb_bank0_rd_data_way0_out_203 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5130 = _T_5129 | _T_4875; // @[Mux.scala 27:72]
  wire  _T_4568 = btb_rd_addr_p1_f == 8'hcc; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4876 = _T_4568 ? btb_bank0_rd_data_way0_out_204 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5131 = _T_5130 | _T_4876; // @[Mux.scala 27:72]
  wire  _T_4570 = btb_rd_addr_p1_f == 8'hcd; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4877 = _T_4570 ? btb_bank0_rd_data_way0_out_205 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5132 = _T_5131 | _T_4877; // @[Mux.scala 27:72]
  wire  _T_4572 = btb_rd_addr_p1_f == 8'hce; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4878 = _T_4572 ? btb_bank0_rd_data_way0_out_206 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5133 = _T_5132 | _T_4878; // @[Mux.scala 27:72]
  wire  _T_4574 = btb_rd_addr_p1_f == 8'hcf; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4879 = _T_4574 ? btb_bank0_rd_data_way0_out_207 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5134 = _T_5133 | _T_4879; // @[Mux.scala 27:72]
  wire  _T_4576 = btb_rd_addr_p1_f == 8'hd0; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4880 = _T_4576 ? btb_bank0_rd_data_way0_out_208 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5135 = _T_5134 | _T_4880; // @[Mux.scala 27:72]
  wire  _T_4578 = btb_rd_addr_p1_f == 8'hd1; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4881 = _T_4578 ? btb_bank0_rd_data_way0_out_209 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5136 = _T_5135 | _T_4881; // @[Mux.scala 27:72]
  wire  _T_4580 = btb_rd_addr_p1_f == 8'hd2; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4882 = _T_4580 ? btb_bank0_rd_data_way0_out_210 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5137 = _T_5136 | _T_4882; // @[Mux.scala 27:72]
  wire  _T_4582 = btb_rd_addr_p1_f == 8'hd3; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4883 = _T_4582 ? btb_bank0_rd_data_way0_out_211 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5138 = _T_5137 | _T_4883; // @[Mux.scala 27:72]
  wire  _T_4584 = btb_rd_addr_p1_f == 8'hd4; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4884 = _T_4584 ? btb_bank0_rd_data_way0_out_212 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5139 = _T_5138 | _T_4884; // @[Mux.scala 27:72]
  wire  _T_4586 = btb_rd_addr_p1_f == 8'hd5; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4885 = _T_4586 ? btb_bank0_rd_data_way0_out_213 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5140 = _T_5139 | _T_4885; // @[Mux.scala 27:72]
  wire  _T_4588 = btb_rd_addr_p1_f == 8'hd6; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4886 = _T_4588 ? btb_bank0_rd_data_way0_out_214 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5141 = _T_5140 | _T_4886; // @[Mux.scala 27:72]
  wire  _T_4590 = btb_rd_addr_p1_f == 8'hd7; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4887 = _T_4590 ? btb_bank0_rd_data_way0_out_215 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5142 = _T_5141 | _T_4887; // @[Mux.scala 27:72]
  wire  _T_4592 = btb_rd_addr_p1_f == 8'hd8; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4888 = _T_4592 ? btb_bank0_rd_data_way0_out_216 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5143 = _T_5142 | _T_4888; // @[Mux.scala 27:72]
  wire  _T_4594 = btb_rd_addr_p1_f == 8'hd9; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4889 = _T_4594 ? btb_bank0_rd_data_way0_out_217 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5144 = _T_5143 | _T_4889; // @[Mux.scala 27:72]
  wire  _T_4596 = btb_rd_addr_p1_f == 8'hda; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4890 = _T_4596 ? btb_bank0_rd_data_way0_out_218 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5145 = _T_5144 | _T_4890; // @[Mux.scala 27:72]
  wire  _T_4598 = btb_rd_addr_p1_f == 8'hdb; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4891 = _T_4598 ? btb_bank0_rd_data_way0_out_219 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5146 = _T_5145 | _T_4891; // @[Mux.scala 27:72]
  wire  _T_4600 = btb_rd_addr_p1_f == 8'hdc; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4892 = _T_4600 ? btb_bank0_rd_data_way0_out_220 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5147 = _T_5146 | _T_4892; // @[Mux.scala 27:72]
  wire  _T_4602 = btb_rd_addr_p1_f == 8'hdd; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4893 = _T_4602 ? btb_bank0_rd_data_way0_out_221 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5148 = _T_5147 | _T_4893; // @[Mux.scala 27:72]
  wire  _T_4604 = btb_rd_addr_p1_f == 8'hde; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4894 = _T_4604 ? btb_bank0_rd_data_way0_out_222 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5149 = _T_5148 | _T_4894; // @[Mux.scala 27:72]
  wire  _T_4606 = btb_rd_addr_p1_f == 8'hdf; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4895 = _T_4606 ? btb_bank0_rd_data_way0_out_223 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5150 = _T_5149 | _T_4895; // @[Mux.scala 27:72]
  wire  _T_4608 = btb_rd_addr_p1_f == 8'he0; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4896 = _T_4608 ? btb_bank0_rd_data_way0_out_224 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5151 = _T_5150 | _T_4896; // @[Mux.scala 27:72]
  wire  _T_4610 = btb_rd_addr_p1_f == 8'he1; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4897 = _T_4610 ? btb_bank0_rd_data_way0_out_225 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5152 = _T_5151 | _T_4897; // @[Mux.scala 27:72]
  wire  _T_4612 = btb_rd_addr_p1_f == 8'he2; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4898 = _T_4612 ? btb_bank0_rd_data_way0_out_226 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5153 = _T_5152 | _T_4898; // @[Mux.scala 27:72]
  wire  _T_4614 = btb_rd_addr_p1_f == 8'he3; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4899 = _T_4614 ? btb_bank0_rd_data_way0_out_227 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5154 = _T_5153 | _T_4899; // @[Mux.scala 27:72]
  wire  _T_4616 = btb_rd_addr_p1_f == 8'he4; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4900 = _T_4616 ? btb_bank0_rd_data_way0_out_228 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5155 = _T_5154 | _T_4900; // @[Mux.scala 27:72]
  wire  _T_4618 = btb_rd_addr_p1_f == 8'he5; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4901 = _T_4618 ? btb_bank0_rd_data_way0_out_229 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5156 = _T_5155 | _T_4901; // @[Mux.scala 27:72]
  wire  _T_4620 = btb_rd_addr_p1_f == 8'he6; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4902 = _T_4620 ? btb_bank0_rd_data_way0_out_230 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5157 = _T_5156 | _T_4902; // @[Mux.scala 27:72]
  wire  _T_4622 = btb_rd_addr_p1_f == 8'he7; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4903 = _T_4622 ? btb_bank0_rd_data_way0_out_231 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5158 = _T_5157 | _T_4903; // @[Mux.scala 27:72]
  wire  _T_4624 = btb_rd_addr_p1_f == 8'he8; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4904 = _T_4624 ? btb_bank0_rd_data_way0_out_232 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5159 = _T_5158 | _T_4904; // @[Mux.scala 27:72]
  wire  _T_4626 = btb_rd_addr_p1_f == 8'he9; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4905 = _T_4626 ? btb_bank0_rd_data_way0_out_233 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5160 = _T_5159 | _T_4905; // @[Mux.scala 27:72]
  wire  _T_4628 = btb_rd_addr_p1_f == 8'hea; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4906 = _T_4628 ? btb_bank0_rd_data_way0_out_234 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5161 = _T_5160 | _T_4906; // @[Mux.scala 27:72]
  wire  _T_4630 = btb_rd_addr_p1_f == 8'heb; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4907 = _T_4630 ? btb_bank0_rd_data_way0_out_235 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5162 = _T_5161 | _T_4907; // @[Mux.scala 27:72]
  wire  _T_4632 = btb_rd_addr_p1_f == 8'hec; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4908 = _T_4632 ? btb_bank0_rd_data_way0_out_236 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5163 = _T_5162 | _T_4908; // @[Mux.scala 27:72]
  wire  _T_4634 = btb_rd_addr_p1_f == 8'hed; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4909 = _T_4634 ? btb_bank0_rd_data_way0_out_237 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5164 = _T_5163 | _T_4909; // @[Mux.scala 27:72]
  wire  _T_4636 = btb_rd_addr_p1_f == 8'hee; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4910 = _T_4636 ? btb_bank0_rd_data_way0_out_238 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5165 = _T_5164 | _T_4910; // @[Mux.scala 27:72]
  wire  _T_4638 = btb_rd_addr_p1_f == 8'hef; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4911 = _T_4638 ? btb_bank0_rd_data_way0_out_239 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5166 = _T_5165 | _T_4911; // @[Mux.scala 27:72]
  wire  _T_4640 = btb_rd_addr_p1_f == 8'hf0; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4912 = _T_4640 ? btb_bank0_rd_data_way0_out_240 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5167 = _T_5166 | _T_4912; // @[Mux.scala 27:72]
  wire  _T_4642 = btb_rd_addr_p1_f == 8'hf1; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4913 = _T_4642 ? btb_bank0_rd_data_way0_out_241 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5168 = _T_5167 | _T_4913; // @[Mux.scala 27:72]
  wire  _T_4644 = btb_rd_addr_p1_f == 8'hf2; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4914 = _T_4644 ? btb_bank0_rd_data_way0_out_242 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5169 = _T_5168 | _T_4914; // @[Mux.scala 27:72]
  wire  _T_4646 = btb_rd_addr_p1_f == 8'hf3; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4915 = _T_4646 ? btb_bank0_rd_data_way0_out_243 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5170 = _T_5169 | _T_4915; // @[Mux.scala 27:72]
  wire  _T_4648 = btb_rd_addr_p1_f == 8'hf4; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4916 = _T_4648 ? btb_bank0_rd_data_way0_out_244 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5171 = _T_5170 | _T_4916; // @[Mux.scala 27:72]
  wire  _T_4650 = btb_rd_addr_p1_f == 8'hf5; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4917 = _T_4650 ? btb_bank0_rd_data_way0_out_245 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5172 = _T_5171 | _T_4917; // @[Mux.scala 27:72]
  wire  _T_4652 = btb_rd_addr_p1_f == 8'hf6; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4918 = _T_4652 ? btb_bank0_rd_data_way0_out_246 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5173 = _T_5172 | _T_4918; // @[Mux.scala 27:72]
  wire  _T_4654 = btb_rd_addr_p1_f == 8'hf7; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4919 = _T_4654 ? btb_bank0_rd_data_way0_out_247 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5174 = _T_5173 | _T_4919; // @[Mux.scala 27:72]
  wire  _T_4656 = btb_rd_addr_p1_f == 8'hf8; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4920 = _T_4656 ? btb_bank0_rd_data_way0_out_248 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5175 = _T_5174 | _T_4920; // @[Mux.scala 27:72]
  wire  _T_4658 = btb_rd_addr_p1_f == 8'hf9; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4921 = _T_4658 ? btb_bank0_rd_data_way0_out_249 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5176 = _T_5175 | _T_4921; // @[Mux.scala 27:72]
  wire  _T_4660 = btb_rd_addr_p1_f == 8'hfa; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4922 = _T_4660 ? btb_bank0_rd_data_way0_out_250 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5177 = _T_5176 | _T_4922; // @[Mux.scala 27:72]
  wire  _T_4662 = btb_rd_addr_p1_f == 8'hfb; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4923 = _T_4662 ? btb_bank0_rd_data_way0_out_251 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5178 = _T_5177 | _T_4923; // @[Mux.scala 27:72]
  wire  _T_4664 = btb_rd_addr_p1_f == 8'hfc; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4924 = _T_4664 ? btb_bank0_rd_data_way0_out_252 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5179 = _T_5178 | _T_4924; // @[Mux.scala 27:72]
  wire  _T_4666 = btb_rd_addr_p1_f == 8'hfd; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4925 = _T_4666 ? btb_bank0_rd_data_way0_out_253 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5180 = _T_5179 | _T_4925; // @[Mux.scala 27:72]
  wire  _T_4668 = btb_rd_addr_p1_f == 8'hfe; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4926 = _T_4668 ? btb_bank0_rd_data_way0_out_254 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5181 = _T_5180 | _T_4926; // @[Mux.scala 27:72]
  wire  _T_4670 = btb_rd_addr_p1_f == 8'hff; // @[ifu_bp_ctl.scala 422:83]
  wire [21:0] _T_4927 = _T_4670 ? btb_bank0_rd_data_way0_out_255 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] btb_bank0_rd_data_way0_p1_f = _T_5181 | _T_4927; // @[Mux.scala 27:72]
  wire [4:0] _T_31 = _T_8[13:9] ^ _T_8[18:14]; // @[lib.scala 42:111]
  wire [4:0] fetch_rd_tag_p1_f = _T_31 ^ _T_8[23:19]; // @[lib.scala 42:111]
  wire  _T_64 = btb_bank0_rd_data_way0_p1_f[21:17] == fetch_rd_tag_p1_f; // @[ifu_bp_ctl.scala 135:106]
  wire  _T_65 = btb_bank0_rd_data_way0_p1_f[0] & _T_64; // @[ifu_bp_ctl.scala 135:61]
  wire  _T_20 = io_exu_bp_exu_i0_br_index_r == btb_rd_addr_p1_f; // @[ifu_bp_ctl.scala 103:75]
  wire  branch_error_collision_p1_f = dec_tlu_error_wb & _T_20; // @[ifu_bp_ctl.scala 103:54]
  wire  branch_error_bank_conflict_p1_f = branch_error_collision_p1_f & dec_tlu_error_wb; // @[ifu_bp_ctl.scala 107:69]
  wire  _T_66 = dec_tlu_way_wb_f & branch_error_bank_conflict_p1_f; // @[ifu_bp_ctl.scala 136:24]
  wire  _T_67 = ~_T_66; // @[ifu_bp_ctl.scala 136:5]
  wire  _T_68 = _T_65 & _T_67; // @[ifu_bp_ctl.scala 135:129]
  wire  _T_69 = _T_68 & io_ifc_fetch_req_f; // @[ifu_bp_ctl.scala 136:59]
  wire  tag_match_way0_p1_f = _T_69 & _T; // @[ifu_bp_ctl.scala 136:80]
  wire  _T_100 = btb_bank0_rd_data_way0_p1_f[3] ^ btb_bank0_rd_data_way0_p1_f[4]; // @[ifu_bp_ctl.scala 148:100]
  wire  _T_101 = tag_match_way0_p1_f & _T_100; // @[ifu_bp_ctl.scala 148:62]
  wire  _T_105 = ~_T_100; // @[ifu_bp_ctl.scala 149:64]
  wire  _T_106 = tag_match_way0_p1_f & _T_105; // @[ifu_bp_ctl.scala 149:62]
  wire [1:0] tag_match_way0_expanded_p1_f = {_T_101,_T_106}; // @[Cat.scala 29:58]
  wire [21:0] _T_134 = tag_match_way0_expanded_p1_f[0] ? btb_bank0_rd_data_way0_p1_f : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5696 = _T_4160 ? btb_bank0_rd_data_way1_out_0 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5697 = _T_4162 ? btb_bank0_rd_data_way1_out_1 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5952 = _T_5696 | _T_5697; // @[Mux.scala 27:72]
  wire [21:0] _T_5698 = _T_4164 ? btb_bank0_rd_data_way1_out_2 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5953 = _T_5952 | _T_5698; // @[Mux.scala 27:72]
  wire [21:0] _T_5699 = _T_4166 ? btb_bank0_rd_data_way1_out_3 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5954 = _T_5953 | _T_5699; // @[Mux.scala 27:72]
  wire [21:0] _T_5700 = _T_4168 ? btb_bank0_rd_data_way1_out_4 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5955 = _T_5954 | _T_5700; // @[Mux.scala 27:72]
  wire [21:0] _T_5701 = _T_4170 ? btb_bank0_rd_data_way1_out_5 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5956 = _T_5955 | _T_5701; // @[Mux.scala 27:72]
  wire [21:0] _T_5702 = _T_4172 ? btb_bank0_rd_data_way1_out_6 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5957 = _T_5956 | _T_5702; // @[Mux.scala 27:72]
  wire [21:0] _T_5703 = _T_4174 ? btb_bank0_rd_data_way1_out_7 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5958 = _T_5957 | _T_5703; // @[Mux.scala 27:72]
  wire [21:0] _T_5704 = _T_4176 ? btb_bank0_rd_data_way1_out_8 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5959 = _T_5958 | _T_5704; // @[Mux.scala 27:72]
  wire [21:0] _T_5705 = _T_4178 ? btb_bank0_rd_data_way1_out_9 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5960 = _T_5959 | _T_5705; // @[Mux.scala 27:72]
  wire [21:0] _T_5706 = _T_4180 ? btb_bank0_rd_data_way1_out_10 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5961 = _T_5960 | _T_5706; // @[Mux.scala 27:72]
  wire [21:0] _T_5707 = _T_4182 ? btb_bank0_rd_data_way1_out_11 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5962 = _T_5961 | _T_5707; // @[Mux.scala 27:72]
  wire [21:0] _T_5708 = _T_4184 ? btb_bank0_rd_data_way1_out_12 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5963 = _T_5962 | _T_5708; // @[Mux.scala 27:72]
  wire [21:0] _T_5709 = _T_4186 ? btb_bank0_rd_data_way1_out_13 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5964 = _T_5963 | _T_5709; // @[Mux.scala 27:72]
  wire [21:0] _T_5710 = _T_4188 ? btb_bank0_rd_data_way1_out_14 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5965 = _T_5964 | _T_5710; // @[Mux.scala 27:72]
  wire [21:0] _T_5711 = _T_4190 ? btb_bank0_rd_data_way1_out_15 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5966 = _T_5965 | _T_5711; // @[Mux.scala 27:72]
  wire [21:0] _T_5712 = _T_4192 ? btb_bank0_rd_data_way1_out_16 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5967 = _T_5966 | _T_5712; // @[Mux.scala 27:72]
  wire [21:0] _T_5713 = _T_4194 ? btb_bank0_rd_data_way1_out_17 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5968 = _T_5967 | _T_5713; // @[Mux.scala 27:72]
  wire [21:0] _T_5714 = _T_4196 ? btb_bank0_rd_data_way1_out_18 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5969 = _T_5968 | _T_5714; // @[Mux.scala 27:72]
  wire [21:0] _T_5715 = _T_4198 ? btb_bank0_rd_data_way1_out_19 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5970 = _T_5969 | _T_5715; // @[Mux.scala 27:72]
  wire [21:0] _T_5716 = _T_4200 ? btb_bank0_rd_data_way1_out_20 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5971 = _T_5970 | _T_5716; // @[Mux.scala 27:72]
  wire [21:0] _T_5717 = _T_4202 ? btb_bank0_rd_data_way1_out_21 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5972 = _T_5971 | _T_5717; // @[Mux.scala 27:72]
  wire [21:0] _T_5718 = _T_4204 ? btb_bank0_rd_data_way1_out_22 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5973 = _T_5972 | _T_5718; // @[Mux.scala 27:72]
  wire [21:0] _T_5719 = _T_4206 ? btb_bank0_rd_data_way1_out_23 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5974 = _T_5973 | _T_5719; // @[Mux.scala 27:72]
  wire [21:0] _T_5720 = _T_4208 ? btb_bank0_rd_data_way1_out_24 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5975 = _T_5974 | _T_5720; // @[Mux.scala 27:72]
  wire [21:0] _T_5721 = _T_4210 ? btb_bank0_rd_data_way1_out_25 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5976 = _T_5975 | _T_5721; // @[Mux.scala 27:72]
  wire [21:0] _T_5722 = _T_4212 ? btb_bank0_rd_data_way1_out_26 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5977 = _T_5976 | _T_5722; // @[Mux.scala 27:72]
  wire [21:0] _T_5723 = _T_4214 ? btb_bank0_rd_data_way1_out_27 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5978 = _T_5977 | _T_5723; // @[Mux.scala 27:72]
  wire [21:0] _T_5724 = _T_4216 ? btb_bank0_rd_data_way1_out_28 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5979 = _T_5978 | _T_5724; // @[Mux.scala 27:72]
  wire [21:0] _T_5725 = _T_4218 ? btb_bank0_rd_data_way1_out_29 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5980 = _T_5979 | _T_5725; // @[Mux.scala 27:72]
  wire [21:0] _T_5726 = _T_4220 ? btb_bank0_rd_data_way1_out_30 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5981 = _T_5980 | _T_5726; // @[Mux.scala 27:72]
  wire [21:0] _T_5727 = _T_4222 ? btb_bank0_rd_data_way1_out_31 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5982 = _T_5981 | _T_5727; // @[Mux.scala 27:72]
  wire [21:0] _T_5728 = _T_4224 ? btb_bank0_rd_data_way1_out_32 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5983 = _T_5982 | _T_5728; // @[Mux.scala 27:72]
  wire [21:0] _T_5729 = _T_4226 ? btb_bank0_rd_data_way1_out_33 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5984 = _T_5983 | _T_5729; // @[Mux.scala 27:72]
  wire [21:0] _T_5730 = _T_4228 ? btb_bank0_rd_data_way1_out_34 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5985 = _T_5984 | _T_5730; // @[Mux.scala 27:72]
  wire [21:0] _T_5731 = _T_4230 ? btb_bank0_rd_data_way1_out_35 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5986 = _T_5985 | _T_5731; // @[Mux.scala 27:72]
  wire [21:0] _T_5732 = _T_4232 ? btb_bank0_rd_data_way1_out_36 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5987 = _T_5986 | _T_5732; // @[Mux.scala 27:72]
  wire [21:0] _T_5733 = _T_4234 ? btb_bank0_rd_data_way1_out_37 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5988 = _T_5987 | _T_5733; // @[Mux.scala 27:72]
  wire [21:0] _T_5734 = _T_4236 ? btb_bank0_rd_data_way1_out_38 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5989 = _T_5988 | _T_5734; // @[Mux.scala 27:72]
  wire [21:0] _T_5735 = _T_4238 ? btb_bank0_rd_data_way1_out_39 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5990 = _T_5989 | _T_5735; // @[Mux.scala 27:72]
  wire [21:0] _T_5736 = _T_4240 ? btb_bank0_rd_data_way1_out_40 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5991 = _T_5990 | _T_5736; // @[Mux.scala 27:72]
  wire [21:0] _T_5737 = _T_4242 ? btb_bank0_rd_data_way1_out_41 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5992 = _T_5991 | _T_5737; // @[Mux.scala 27:72]
  wire [21:0] _T_5738 = _T_4244 ? btb_bank0_rd_data_way1_out_42 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5993 = _T_5992 | _T_5738; // @[Mux.scala 27:72]
  wire [21:0] _T_5739 = _T_4246 ? btb_bank0_rd_data_way1_out_43 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5994 = _T_5993 | _T_5739; // @[Mux.scala 27:72]
  wire [21:0] _T_5740 = _T_4248 ? btb_bank0_rd_data_way1_out_44 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5995 = _T_5994 | _T_5740; // @[Mux.scala 27:72]
  wire [21:0] _T_5741 = _T_4250 ? btb_bank0_rd_data_way1_out_45 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5996 = _T_5995 | _T_5741; // @[Mux.scala 27:72]
  wire [21:0] _T_5742 = _T_4252 ? btb_bank0_rd_data_way1_out_46 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5997 = _T_5996 | _T_5742; // @[Mux.scala 27:72]
  wire [21:0] _T_5743 = _T_4254 ? btb_bank0_rd_data_way1_out_47 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5998 = _T_5997 | _T_5743; // @[Mux.scala 27:72]
  wire [21:0] _T_5744 = _T_4256 ? btb_bank0_rd_data_way1_out_48 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5999 = _T_5998 | _T_5744; // @[Mux.scala 27:72]
  wire [21:0] _T_5745 = _T_4258 ? btb_bank0_rd_data_way1_out_49 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6000 = _T_5999 | _T_5745; // @[Mux.scala 27:72]
  wire [21:0] _T_5746 = _T_4260 ? btb_bank0_rd_data_way1_out_50 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6001 = _T_6000 | _T_5746; // @[Mux.scala 27:72]
  wire [21:0] _T_5747 = _T_4262 ? btb_bank0_rd_data_way1_out_51 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6002 = _T_6001 | _T_5747; // @[Mux.scala 27:72]
  wire [21:0] _T_5748 = _T_4264 ? btb_bank0_rd_data_way1_out_52 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6003 = _T_6002 | _T_5748; // @[Mux.scala 27:72]
  wire [21:0] _T_5749 = _T_4266 ? btb_bank0_rd_data_way1_out_53 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6004 = _T_6003 | _T_5749; // @[Mux.scala 27:72]
  wire [21:0] _T_5750 = _T_4268 ? btb_bank0_rd_data_way1_out_54 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6005 = _T_6004 | _T_5750; // @[Mux.scala 27:72]
  wire [21:0] _T_5751 = _T_4270 ? btb_bank0_rd_data_way1_out_55 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6006 = _T_6005 | _T_5751; // @[Mux.scala 27:72]
  wire [21:0] _T_5752 = _T_4272 ? btb_bank0_rd_data_way1_out_56 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6007 = _T_6006 | _T_5752; // @[Mux.scala 27:72]
  wire [21:0] _T_5753 = _T_4274 ? btb_bank0_rd_data_way1_out_57 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6008 = _T_6007 | _T_5753; // @[Mux.scala 27:72]
  wire [21:0] _T_5754 = _T_4276 ? btb_bank0_rd_data_way1_out_58 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6009 = _T_6008 | _T_5754; // @[Mux.scala 27:72]
  wire [21:0] _T_5755 = _T_4278 ? btb_bank0_rd_data_way1_out_59 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6010 = _T_6009 | _T_5755; // @[Mux.scala 27:72]
  wire [21:0] _T_5756 = _T_4280 ? btb_bank0_rd_data_way1_out_60 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6011 = _T_6010 | _T_5756; // @[Mux.scala 27:72]
  wire [21:0] _T_5757 = _T_4282 ? btb_bank0_rd_data_way1_out_61 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6012 = _T_6011 | _T_5757; // @[Mux.scala 27:72]
  wire [21:0] _T_5758 = _T_4284 ? btb_bank0_rd_data_way1_out_62 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6013 = _T_6012 | _T_5758; // @[Mux.scala 27:72]
  wire [21:0] _T_5759 = _T_4286 ? btb_bank0_rd_data_way1_out_63 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6014 = _T_6013 | _T_5759; // @[Mux.scala 27:72]
  wire [21:0] _T_5760 = _T_4288 ? btb_bank0_rd_data_way1_out_64 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6015 = _T_6014 | _T_5760; // @[Mux.scala 27:72]
  wire [21:0] _T_5761 = _T_4290 ? btb_bank0_rd_data_way1_out_65 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6016 = _T_6015 | _T_5761; // @[Mux.scala 27:72]
  wire [21:0] _T_5762 = _T_4292 ? btb_bank0_rd_data_way1_out_66 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6017 = _T_6016 | _T_5762; // @[Mux.scala 27:72]
  wire [21:0] _T_5763 = _T_4294 ? btb_bank0_rd_data_way1_out_67 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6018 = _T_6017 | _T_5763; // @[Mux.scala 27:72]
  wire [21:0] _T_5764 = _T_4296 ? btb_bank0_rd_data_way1_out_68 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6019 = _T_6018 | _T_5764; // @[Mux.scala 27:72]
  wire [21:0] _T_5765 = _T_4298 ? btb_bank0_rd_data_way1_out_69 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6020 = _T_6019 | _T_5765; // @[Mux.scala 27:72]
  wire [21:0] _T_5766 = _T_4300 ? btb_bank0_rd_data_way1_out_70 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6021 = _T_6020 | _T_5766; // @[Mux.scala 27:72]
  wire [21:0] _T_5767 = _T_4302 ? btb_bank0_rd_data_way1_out_71 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6022 = _T_6021 | _T_5767; // @[Mux.scala 27:72]
  wire [21:0] _T_5768 = _T_4304 ? btb_bank0_rd_data_way1_out_72 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6023 = _T_6022 | _T_5768; // @[Mux.scala 27:72]
  wire [21:0] _T_5769 = _T_4306 ? btb_bank0_rd_data_way1_out_73 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6024 = _T_6023 | _T_5769; // @[Mux.scala 27:72]
  wire [21:0] _T_5770 = _T_4308 ? btb_bank0_rd_data_way1_out_74 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6025 = _T_6024 | _T_5770; // @[Mux.scala 27:72]
  wire [21:0] _T_5771 = _T_4310 ? btb_bank0_rd_data_way1_out_75 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6026 = _T_6025 | _T_5771; // @[Mux.scala 27:72]
  wire [21:0] _T_5772 = _T_4312 ? btb_bank0_rd_data_way1_out_76 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6027 = _T_6026 | _T_5772; // @[Mux.scala 27:72]
  wire [21:0] _T_5773 = _T_4314 ? btb_bank0_rd_data_way1_out_77 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6028 = _T_6027 | _T_5773; // @[Mux.scala 27:72]
  wire [21:0] _T_5774 = _T_4316 ? btb_bank0_rd_data_way1_out_78 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6029 = _T_6028 | _T_5774; // @[Mux.scala 27:72]
  wire [21:0] _T_5775 = _T_4318 ? btb_bank0_rd_data_way1_out_79 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6030 = _T_6029 | _T_5775; // @[Mux.scala 27:72]
  wire [21:0] _T_5776 = _T_4320 ? btb_bank0_rd_data_way1_out_80 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6031 = _T_6030 | _T_5776; // @[Mux.scala 27:72]
  wire [21:0] _T_5777 = _T_4322 ? btb_bank0_rd_data_way1_out_81 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6032 = _T_6031 | _T_5777; // @[Mux.scala 27:72]
  wire [21:0] _T_5778 = _T_4324 ? btb_bank0_rd_data_way1_out_82 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6033 = _T_6032 | _T_5778; // @[Mux.scala 27:72]
  wire [21:0] _T_5779 = _T_4326 ? btb_bank0_rd_data_way1_out_83 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6034 = _T_6033 | _T_5779; // @[Mux.scala 27:72]
  wire [21:0] _T_5780 = _T_4328 ? btb_bank0_rd_data_way1_out_84 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6035 = _T_6034 | _T_5780; // @[Mux.scala 27:72]
  wire [21:0] _T_5781 = _T_4330 ? btb_bank0_rd_data_way1_out_85 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6036 = _T_6035 | _T_5781; // @[Mux.scala 27:72]
  wire [21:0] _T_5782 = _T_4332 ? btb_bank0_rd_data_way1_out_86 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6037 = _T_6036 | _T_5782; // @[Mux.scala 27:72]
  wire [21:0] _T_5783 = _T_4334 ? btb_bank0_rd_data_way1_out_87 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6038 = _T_6037 | _T_5783; // @[Mux.scala 27:72]
  wire [21:0] _T_5784 = _T_4336 ? btb_bank0_rd_data_way1_out_88 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6039 = _T_6038 | _T_5784; // @[Mux.scala 27:72]
  wire [21:0] _T_5785 = _T_4338 ? btb_bank0_rd_data_way1_out_89 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6040 = _T_6039 | _T_5785; // @[Mux.scala 27:72]
  wire [21:0] _T_5786 = _T_4340 ? btb_bank0_rd_data_way1_out_90 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6041 = _T_6040 | _T_5786; // @[Mux.scala 27:72]
  wire [21:0] _T_5787 = _T_4342 ? btb_bank0_rd_data_way1_out_91 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6042 = _T_6041 | _T_5787; // @[Mux.scala 27:72]
  wire [21:0] _T_5788 = _T_4344 ? btb_bank0_rd_data_way1_out_92 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6043 = _T_6042 | _T_5788; // @[Mux.scala 27:72]
  wire [21:0] _T_5789 = _T_4346 ? btb_bank0_rd_data_way1_out_93 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6044 = _T_6043 | _T_5789; // @[Mux.scala 27:72]
  wire [21:0] _T_5790 = _T_4348 ? btb_bank0_rd_data_way1_out_94 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6045 = _T_6044 | _T_5790; // @[Mux.scala 27:72]
  wire [21:0] _T_5791 = _T_4350 ? btb_bank0_rd_data_way1_out_95 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6046 = _T_6045 | _T_5791; // @[Mux.scala 27:72]
  wire [21:0] _T_5792 = _T_4352 ? btb_bank0_rd_data_way1_out_96 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6047 = _T_6046 | _T_5792; // @[Mux.scala 27:72]
  wire [21:0] _T_5793 = _T_4354 ? btb_bank0_rd_data_way1_out_97 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6048 = _T_6047 | _T_5793; // @[Mux.scala 27:72]
  wire [21:0] _T_5794 = _T_4356 ? btb_bank0_rd_data_way1_out_98 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6049 = _T_6048 | _T_5794; // @[Mux.scala 27:72]
  wire [21:0] _T_5795 = _T_4358 ? btb_bank0_rd_data_way1_out_99 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6050 = _T_6049 | _T_5795; // @[Mux.scala 27:72]
  wire [21:0] _T_5796 = _T_4360 ? btb_bank0_rd_data_way1_out_100 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6051 = _T_6050 | _T_5796; // @[Mux.scala 27:72]
  wire [21:0] _T_5797 = _T_4362 ? btb_bank0_rd_data_way1_out_101 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6052 = _T_6051 | _T_5797; // @[Mux.scala 27:72]
  wire [21:0] _T_5798 = _T_4364 ? btb_bank0_rd_data_way1_out_102 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6053 = _T_6052 | _T_5798; // @[Mux.scala 27:72]
  wire [21:0] _T_5799 = _T_4366 ? btb_bank0_rd_data_way1_out_103 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6054 = _T_6053 | _T_5799; // @[Mux.scala 27:72]
  wire [21:0] _T_5800 = _T_4368 ? btb_bank0_rd_data_way1_out_104 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6055 = _T_6054 | _T_5800; // @[Mux.scala 27:72]
  wire [21:0] _T_5801 = _T_4370 ? btb_bank0_rd_data_way1_out_105 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6056 = _T_6055 | _T_5801; // @[Mux.scala 27:72]
  wire [21:0] _T_5802 = _T_4372 ? btb_bank0_rd_data_way1_out_106 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6057 = _T_6056 | _T_5802; // @[Mux.scala 27:72]
  wire [21:0] _T_5803 = _T_4374 ? btb_bank0_rd_data_way1_out_107 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6058 = _T_6057 | _T_5803; // @[Mux.scala 27:72]
  wire [21:0] _T_5804 = _T_4376 ? btb_bank0_rd_data_way1_out_108 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6059 = _T_6058 | _T_5804; // @[Mux.scala 27:72]
  wire [21:0] _T_5805 = _T_4378 ? btb_bank0_rd_data_way1_out_109 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6060 = _T_6059 | _T_5805; // @[Mux.scala 27:72]
  wire [21:0] _T_5806 = _T_4380 ? btb_bank0_rd_data_way1_out_110 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6061 = _T_6060 | _T_5806; // @[Mux.scala 27:72]
  wire [21:0] _T_5807 = _T_4382 ? btb_bank0_rd_data_way1_out_111 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6062 = _T_6061 | _T_5807; // @[Mux.scala 27:72]
  wire [21:0] _T_5808 = _T_4384 ? btb_bank0_rd_data_way1_out_112 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6063 = _T_6062 | _T_5808; // @[Mux.scala 27:72]
  wire [21:0] _T_5809 = _T_4386 ? btb_bank0_rd_data_way1_out_113 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6064 = _T_6063 | _T_5809; // @[Mux.scala 27:72]
  wire [21:0] _T_5810 = _T_4388 ? btb_bank0_rd_data_way1_out_114 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6065 = _T_6064 | _T_5810; // @[Mux.scala 27:72]
  wire [21:0] _T_5811 = _T_4390 ? btb_bank0_rd_data_way1_out_115 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6066 = _T_6065 | _T_5811; // @[Mux.scala 27:72]
  wire [21:0] _T_5812 = _T_4392 ? btb_bank0_rd_data_way1_out_116 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6067 = _T_6066 | _T_5812; // @[Mux.scala 27:72]
  wire [21:0] _T_5813 = _T_4394 ? btb_bank0_rd_data_way1_out_117 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6068 = _T_6067 | _T_5813; // @[Mux.scala 27:72]
  wire [21:0] _T_5814 = _T_4396 ? btb_bank0_rd_data_way1_out_118 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6069 = _T_6068 | _T_5814; // @[Mux.scala 27:72]
  wire [21:0] _T_5815 = _T_4398 ? btb_bank0_rd_data_way1_out_119 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6070 = _T_6069 | _T_5815; // @[Mux.scala 27:72]
  wire [21:0] _T_5816 = _T_4400 ? btb_bank0_rd_data_way1_out_120 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6071 = _T_6070 | _T_5816; // @[Mux.scala 27:72]
  wire [21:0] _T_5817 = _T_4402 ? btb_bank0_rd_data_way1_out_121 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6072 = _T_6071 | _T_5817; // @[Mux.scala 27:72]
  wire [21:0] _T_5818 = _T_4404 ? btb_bank0_rd_data_way1_out_122 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6073 = _T_6072 | _T_5818; // @[Mux.scala 27:72]
  wire [21:0] _T_5819 = _T_4406 ? btb_bank0_rd_data_way1_out_123 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6074 = _T_6073 | _T_5819; // @[Mux.scala 27:72]
  wire [21:0] _T_5820 = _T_4408 ? btb_bank0_rd_data_way1_out_124 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6075 = _T_6074 | _T_5820; // @[Mux.scala 27:72]
  wire [21:0] _T_5821 = _T_4410 ? btb_bank0_rd_data_way1_out_125 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6076 = _T_6075 | _T_5821; // @[Mux.scala 27:72]
  wire [21:0] _T_5822 = _T_4412 ? btb_bank0_rd_data_way1_out_126 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6077 = _T_6076 | _T_5822; // @[Mux.scala 27:72]
  wire [21:0] _T_5823 = _T_4414 ? btb_bank0_rd_data_way1_out_127 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6078 = _T_6077 | _T_5823; // @[Mux.scala 27:72]
  wire [21:0] _T_5824 = _T_4416 ? btb_bank0_rd_data_way1_out_128 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6079 = _T_6078 | _T_5824; // @[Mux.scala 27:72]
  wire [21:0] _T_5825 = _T_4418 ? btb_bank0_rd_data_way1_out_129 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6080 = _T_6079 | _T_5825; // @[Mux.scala 27:72]
  wire [21:0] _T_5826 = _T_4420 ? btb_bank0_rd_data_way1_out_130 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6081 = _T_6080 | _T_5826; // @[Mux.scala 27:72]
  wire [21:0] _T_5827 = _T_4422 ? btb_bank0_rd_data_way1_out_131 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6082 = _T_6081 | _T_5827; // @[Mux.scala 27:72]
  wire [21:0] _T_5828 = _T_4424 ? btb_bank0_rd_data_way1_out_132 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6083 = _T_6082 | _T_5828; // @[Mux.scala 27:72]
  wire [21:0] _T_5829 = _T_4426 ? btb_bank0_rd_data_way1_out_133 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6084 = _T_6083 | _T_5829; // @[Mux.scala 27:72]
  wire [21:0] _T_5830 = _T_4428 ? btb_bank0_rd_data_way1_out_134 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6085 = _T_6084 | _T_5830; // @[Mux.scala 27:72]
  wire [21:0] _T_5831 = _T_4430 ? btb_bank0_rd_data_way1_out_135 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6086 = _T_6085 | _T_5831; // @[Mux.scala 27:72]
  wire [21:0] _T_5832 = _T_4432 ? btb_bank0_rd_data_way1_out_136 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6087 = _T_6086 | _T_5832; // @[Mux.scala 27:72]
  wire [21:0] _T_5833 = _T_4434 ? btb_bank0_rd_data_way1_out_137 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6088 = _T_6087 | _T_5833; // @[Mux.scala 27:72]
  wire [21:0] _T_5834 = _T_4436 ? btb_bank0_rd_data_way1_out_138 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6089 = _T_6088 | _T_5834; // @[Mux.scala 27:72]
  wire [21:0] _T_5835 = _T_4438 ? btb_bank0_rd_data_way1_out_139 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6090 = _T_6089 | _T_5835; // @[Mux.scala 27:72]
  wire [21:0] _T_5836 = _T_4440 ? btb_bank0_rd_data_way1_out_140 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6091 = _T_6090 | _T_5836; // @[Mux.scala 27:72]
  wire [21:0] _T_5837 = _T_4442 ? btb_bank0_rd_data_way1_out_141 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6092 = _T_6091 | _T_5837; // @[Mux.scala 27:72]
  wire [21:0] _T_5838 = _T_4444 ? btb_bank0_rd_data_way1_out_142 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6093 = _T_6092 | _T_5838; // @[Mux.scala 27:72]
  wire [21:0] _T_5839 = _T_4446 ? btb_bank0_rd_data_way1_out_143 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6094 = _T_6093 | _T_5839; // @[Mux.scala 27:72]
  wire [21:0] _T_5840 = _T_4448 ? btb_bank0_rd_data_way1_out_144 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6095 = _T_6094 | _T_5840; // @[Mux.scala 27:72]
  wire [21:0] _T_5841 = _T_4450 ? btb_bank0_rd_data_way1_out_145 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6096 = _T_6095 | _T_5841; // @[Mux.scala 27:72]
  wire [21:0] _T_5842 = _T_4452 ? btb_bank0_rd_data_way1_out_146 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6097 = _T_6096 | _T_5842; // @[Mux.scala 27:72]
  wire [21:0] _T_5843 = _T_4454 ? btb_bank0_rd_data_way1_out_147 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6098 = _T_6097 | _T_5843; // @[Mux.scala 27:72]
  wire [21:0] _T_5844 = _T_4456 ? btb_bank0_rd_data_way1_out_148 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6099 = _T_6098 | _T_5844; // @[Mux.scala 27:72]
  wire [21:0] _T_5845 = _T_4458 ? btb_bank0_rd_data_way1_out_149 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6100 = _T_6099 | _T_5845; // @[Mux.scala 27:72]
  wire [21:0] _T_5846 = _T_4460 ? btb_bank0_rd_data_way1_out_150 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6101 = _T_6100 | _T_5846; // @[Mux.scala 27:72]
  wire [21:0] _T_5847 = _T_4462 ? btb_bank0_rd_data_way1_out_151 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6102 = _T_6101 | _T_5847; // @[Mux.scala 27:72]
  wire [21:0] _T_5848 = _T_4464 ? btb_bank0_rd_data_way1_out_152 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6103 = _T_6102 | _T_5848; // @[Mux.scala 27:72]
  wire [21:0] _T_5849 = _T_4466 ? btb_bank0_rd_data_way1_out_153 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6104 = _T_6103 | _T_5849; // @[Mux.scala 27:72]
  wire [21:0] _T_5850 = _T_4468 ? btb_bank0_rd_data_way1_out_154 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6105 = _T_6104 | _T_5850; // @[Mux.scala 27:72]
  wire [21:0] _T_5851 = _T_4470 ? btb_bank0_rd_data_way1_out_155 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6106 = _T_6105 | _T_5851; // @[Mux.scala 27:72]
  wire [21:0] _T_5852 = _T_4472 ? btb_bank0_rd_data_way1_out_156 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6107 = _T_6106 | _T_5852; // @[Mux.scala 27:72]
  wire [21:0] _T_5853 = _T_4474 ? btb_bank0_rd_data_way1_out_157 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6108 = _T_6107 | _T_5853; // @[Mux.scala 27:72]
  wire [21:0] _T_5854 = _T_4476 ? btb_bank0_rd_data_way1_out_158 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6109 = _T_6108 | _T_5854; // @[Mux.scala 27:72]
  wire [21:0] _T_5855 = _T_4478 ? btb_bank0_rd_data_way1_out_159 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6110 = _T_6109 | _T_5855; // @[Mux.scala 27:72]
  wire [21:0] _T_5856 = _T_4480 ? btb_bank0_rd_data_way1_out_160 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6111 = _T_6110 | _T_5856; // @[Mux.scala 27:72]
  wire [21:0] _T_5857 = _T_4482 ? btb_bank0_rd_data_way1_out_161 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6112 = _T_6111 | _T_5857; // @[Mux.scala 27:72]
  wire [21:0] _T_5858 = _T_4484 ? btb_bank0_rd_data_way1_out_162 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6113 = _T_6112 | _T_5858; // @[Mux.scala 27:72]
  wire [21:0] _T_5859 = _T_4486 ? btb_bank0_rd_data_way1_out_163 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6114 = _T_6113 | _T_5859; // @[Mux.scala 27:72]
  wire [21:0] _T_5860 = _T_4488 ? btb_bank0_rd_data_way1_out_164 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6115 = _T_6114 | _T_5860; // @[Mux.scala 27:72]
  wire [21:0] _T_5861 = _T_4490 ? btb_bank0_rd_data_way1_out_165 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6116 = _T_6115 | _T_5861; // @[Mux.scala 27:72]
  wire [21:0] _T_5862 = _T_4492 ? btb_bank0_rd_data_way1_out_166 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6117 = _T_6116 | _T_5862; // @[Mux.scala 27:72]
  wire [21:0] _T_5863 = _T_4494 ? btb_bank0_rd_data_way1_out_167 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6118 = _T_6117 | _T_5863; // @[Mux.scala 27:72]
  wire [21:0] _T_5864 = _T_4496 ? btb_bank0_rd_data_way1_out_168 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6119 = _T_6118 | _T_5864; // @[Mux.scala 27:72]
  wire [21:0] _T_5865 = _T_4498 ? btb_bank0_rd_data_way1_out_169 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6120 = _T_6119 | _T_5865; // @[Mux.scala 27:72]
  wire [21:0] _T_5866 = _T_4500 ? btb_bank0_rd_data_way1_out_170 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6121 = _T_6120 | _T_5866; // @[Mux.scala 27:72]
  wire [21:0] _T_5867 = _T_4502 ? btb_bank0_rd_data_way1_out_171 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6122 = _T_6121 | _T_5867; // @[Mux.scala 27:72]
  wire [21:0] _T_5868 = _T_4504 ? btb_bank0_rd_data_way1_out_172 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6123 = _T_6122 | _T_5868; // @[Mux.scala 27:72]
  wire [21:0] _T_5869 = _T_4506 ? btb_bank0_rd_data_way1_out_173 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6124 = _T_6123 | _T_5869; // @[Mux.scala 27:72]
  wire [21:0] _T_5870 = _T_4508 ? btb_bank0_rd_data_way1_out_174 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6125 = _T_6124 | _T_5870; // @[Mux.scala 27:72]
  wire [21:0] _T_5871 = _T_4510 ? btb_bank0_rd_data_way1_out_175 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6126 = _T_6125 | _T_5871; // @[Mux.scala 27:72]
  wire [21:0] _T_5872 = _T_4512 ? btb_bank0_rd_data_way1_out_176 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6127 = _T_6126 | _T_5872; // @[Mux.scala 27:72]
  wire [21:0] _T_5873 = _T_4514 ? btb_bank0_rd_data_way1_out_177 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6128 = _T_6127 | _T_5873; // @[Mux.scala 27:72]
  wire [21:0] _T_5874 = _T_4516 ? btb_bank0_rd_data_way1_out_178 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6129 = _T_6128 | _T_5874; // @[Mux.scala 27:72]
  wire [21:0] _T_5875 = _T_4518 ? btb_bank0_rd_data_way1_out_179 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6130 = _T_6129 | _T_5875; // @[Mux.scala 27:72]
  wire [21:0] _T_5876 = _T_4520 ? btb_bank0_rd_data_way1_out_180 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6131 = _T_6130 | _T_5876; // @[Mux.scala 27:72]
  wire [21:0] _T_5877 = _T_4522 ? btb_bank0_rd_data_way1_out_181 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6132 = _T_6131 | _T_5877; // @[Mux.scala 27:72]
  wire [21:0] _T_5878 = _T_4524 ? btb_bank0_rd_data_way1_out_182 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6133 = _T_6132 | _T_5878; // @[Mux.scala 27:72]
  wire [21:0] _T_5879 = _T_4526 ? btb_bank0_rd_data_way1_out_183 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6134 = _T_6133 | _T_5879; // @[Mux.scala 27:72]
  wire [21:0] _T_5880 = _T_4528 ? btb_bank0_rd_data_way1_out_184 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6135 = _T_6134 | _T_5880; // @[Mux.scala 27:72]
  wire [21:0] _T_5881 = _T_4530 ? btb_bank0_rd_data_way1_out_185 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6136 = _T_6135 | _T_5881; // @[Mux.scala 27:72]
  wire [21:0] _T_5882 = _T_4532 ? btb_bank0_rd_data_way1_out_186 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6137 = _T_6136 | _T_5882; // @[Mux.scala 27:72]
  wire [21:0] _T_5883 = _T_4534 ? btb_bank0_rd_data_way1_out_187 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6138 = _T_6137 | _T_5883; // @[Mux.scala 27:72]
  wire [21:0] _T_5884 = _T_4536 ? btb_bank0_rd_data_way1_out_188 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6139 = _T_6138 | _T_5884; // @[Mux.scala 27:72]
  wire [21:0] _T_5885 = _T_4538 ? btb_bank0_rd_data_way1_out_189 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6140 = _T_6139 | _T_5885; // @[Mux.scala 27:72]
  wire [21:0] _T_5886 = _T_4540 ? btb_bank0_rd_data_way1_out_190 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6141 = _T_6140 | _T_5886; // @[Mux.scala 27:72]
  wire [21:0] _T_5887 = _T_4542 ? btb_bank0_rd_data_way1_out_191 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6142 = _T_6141 | _T_5887; // @[Mux.scala 27:72]
  wire [21:0] _T_5888 = _T_4544 ? btb_bank0_rd_data_way1_out_192 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6143 = _T_6142 | _T_5888; // @[Mux.scala 27:72]
  wire [21:0] _T_5889 = _T_4546 ? btb_bank0_rd_data_way1_out_193 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6144 = _T_6143 | _T_5889; // @[Mux.scala 27:72]
  wire [21:0] _T_5890 = _T_4548 ? btb_bank0_rd_data_way1_out_194 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6145 = _T_6144 | _T_5890; // @[Mux.scala 27:72]
  wire [21:0] _T_5891 = _T_4550 ? btb_bank0_rd_data_way1_out_195 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6146 = _T_6145 | _T_5891; // @[Mux.scala 27:72]
  wire [21:0] _T_5892 = _T_4552 ? btb_bank0_rd_data_way1_out_196 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6147 = _T_6146 | _T_5892; // @[Mux.scala 27:72]
  wire [21:0] _T_5893 = _T_4554 ? btb_bank0_rd_data_way1_out_197 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6148 = _T_6147 | _T_5893; // @[Mux.scala 27:72]
  wire [21:0] _T_5894 = _T_4556 ? btb_bank0_rd_data_way1_out_198 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6149 = _T_6148 | _T_5894; // @[Mux.scala 27:72]
  wire [21:0] _T_5895 = _T_4558 ? btb_bank0_rd_data_way1_out_199 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6150 = _T_6149 | _T_5895; // @[Mux.scala 27:72]
  wire [21:0] _T_5896 = _T_4560 ? btb_bank0_rd_data_way1_out_200 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6151 = _T_6150 | _T_5896; // @[Mux.scala 27:72]
  wire [21:0] _T_5897 = _T_4562 ? btb_bank0_rd_data_way1_out_201 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6152 = _T_6151 | _T_5897; // @[Mux.scala 27:72]
  wire [21:0] _T_5898 = _T_4564 ? btb_bank0_rd_data_way1_out_202 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6153 = _T_6152 | _T_5898; // @[Mux.scala 27:72]
  wire [21:0] _T_5899 = _T_4566 ? btb_bank0_rd_data_way1_out_203 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6154 = _T_6153 | _T_5899; // @[Mux.scala 27:72]
  wire [21:0] _T_5900 = _T_4568 ? btb_bank0_rd_data_way1_out_204 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6155 = _T_6154 | _T_5900; // @[Mux.scala 27:72]
  wire [21:0] _T_5901 = _T_4570 ? btb_bank0_rd_data_way1_out_205 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6156 = _T_6155 | _T_5901; // @[Mux.scala 27:72]
  wire [21:0] _T_5902 = _T_4572 ? btb_bank0_rd_data_way1_out_206 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6157 = _T_6156 | _T_5902; // @[Mux.scala 27:72]
  wire [21:0] _T_5903 = _T_4574 ? btb_bank0_rd_data_way1_out_207 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6158 = _T_6157 | _T_5903; // @[Mux.scala 27:72]
  wire [21:0] _T_5904 = _T_4576 ? btb_bank0_rd_data_way1_out_208 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6159 = _T_6158 | _T_5904; // @[Mux.scala 27:72]
  wire [21:0] _T_5905 = _T_4578 ? btb_bank0_rd_data_way1_out_209 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6160 = _T_6159 | _T_5905; // @[Mux.scala 27:72]
  wire [21:0] _T_5906 = _T_4580 ? btb_bank0_rd_data_way1_out_210 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6161 = _T_6160 | _T_5906; // @[Mux.scala 27:72]
  wire [21:0] _T_5907 = _T_4582 ? btb_bank0_rd_data_way1_out_211 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6162 = _T_6161 | _T_5907; // @[Mux.scala 27:72]
  wire [21:0] _T_5908 = _T_4584 ? btb_bank0_rd_data_way1_out_212 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6163 = _T_6162 | _T_5908; // @[Mux.scala 27:72]
  wire [21:0] _T_5909 = _T_4586 ? btb_bank0_rd_data_way1_out_213 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6164 = _T_6163 | _T_5909; // @[Mux.scala 27:72]
  wire [21:0] _T_5910 = _T_4588 ? btb_bank0_rd_data_way1_out_214 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6165 = _T_6164 | _T_5910; // @[Mux.scala 27:72]
  wire [21:0] _T_5911 = _T_4590 ? btb_bank0_rd_data_way1_out_215 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6166 = _T_6165 | _T_5911; // @[Mux.scala 27:72]
  wire [21:0] _T_5912 = _T_4592 ? btb_bank0_rd_data_way1_out_216 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6167 = _T_6166 | _T_5912; // @[Mux.scala 27:72]
  wire [21:0] _T_5913 = _T_4594 ? btb_bank0_rd_data_way1_out_217 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6168 = _T_6167 | _T_5913; // @[Mux.scala 27:72]
  wire [21:0] _T_5914 = _T_4596 ? btb_bank0_rd_data_way1_out_218 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6169 = _T_6168 | _T_5914; // @[Mux.scala 27:72]
  wire [21:0] _T_5915 = _T_4598 ? btb_bank0_rd_data_way1_out_219 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6170 = _T_6169 | _T_5915; // @[Mux.scala 27:72]
  wire [21:0] _T_5916 = _T_4600 ? btb_bank0_rd_data_way1_out_220 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6171 = _T_6170 | _T_5916; // @[Mux.scala 27:72]
  wire [21:0] _T_5917 = _T_4602 ? btb_bank0_rd_data_way1_out_221 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6172 = _T_6171 | _T_5917; // @[Mux.scala 27:72]
  wire [21:0] _T_5918 = _T_4604 ? btb_bank0_rd_data_way1_out_222 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6173 = _T_6172 | _T_5918; // @[Mux.scala 27:72]
  wire [21:0] _T_5919 = _T_4606 ? btb_bank0_rd_data_way1_out_223 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6174 = _T_6173 | _T_5919; // @[Mux.scala 27:72]
  wire [21:0] _T_5920 = _T_4608 ? btb_bank0_rd_data_way1_out_224 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6175 = _T_6174 | _T_5920; // @[Mux.scala 27:72]
  wire [21:0] _T_5921 = _T_4610 ? btb_bank0_rd_data_way1_out_225 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6176 = _T_6175 | _T_5921; // @[Mux.scala 27:72]
  wire [21:0] _T_5922 = _T_4612 ? btb_bank0_rd_data_way1_out_226 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6177 = _T_6176 | _T_5922; // @[Mux.scala 27:72]
  wire [21:0] _T_5923 = _T_4614 ? btb_bank0_rd_data_way1_out_227 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6178 = _T_6177 | _T_5923; // @[Mux.scala 27:72]
  wire [21:0] _T_5924 = _T_4616 ? btb_bank0_rd_data_way1_out_228 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6179 = _T_6178 | _T_5924; // @[Mux.scala 27:72]
  wire [21:0] _T_5925 = _T_4618 ? btb_bank0_rd_data_way1_out_229 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6180 = _T_6179 | _T_5925; // @[Mux.scala 27:72]
  wire [21:0] _T_5926 = _T_4620 ? btb_bank0_rd_data_way1_out_230 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6181 = _T_6180 | _T_5926; // @[Mux.scala 27:72]
  wire [21:0] _T_5927 = _T_4622 ? btb_bank0_rd_data_way1_out_231 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6182 = _T_6181 | _T_5927; // @[Mux.scala 27:72]
  wire [21:0] _T_5928 = _T_4624 ? btb_bank0_rd_data_way1_out_232 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6183 = _T_6182 | _T_5928; // @[Mux.scala 27:72]
  wire [21:0] _T_5929 = _T_4626 ? btb_bank0_rd_data_way1_out_233 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6184 = _T_6183 | _T_5929; // @[Mux.scala 27:72]
  wire [21:0] _T_5930 = _T_4628 ? btb_bank0_rd_data_way1_out_234 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6185 = _T_6184 | _T_5930; // @[Mux.scala 27:72]
  wire [21:0] _T_5931 = _T_4630 ? btb_bank0_rd_data_way1_out_235 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6186 = _T_6185 | _T_5931; // @[Mux.scala 27:72]
  wire [21:0] _T_5932 = _T_4632 ? btb_bank0_rd_data_way1_out_236 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6187 = _T_6186 | _T_5932; // @[Mux.scala 27:72]
  wire [21:0] _T_5933 = _T_4634 ? btb_bank0_rd_data_way1_out_237 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6188 = _T_6187 | _T_5933; // @[Mux.scala 27:72]
  wire [21:0] _T_5934 = _T_4636 ? btb_bank0_rd_data_way1_out_238 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6189 = _T_6188 | _T_5934; // @[Mux.scala 27:72]
  wire [21:0] _T_5935 = _T_4638 ? btb_bank0_rd_data_way1_out_239 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6190 = _T_6189 | _T_5935; // @[Mux.scala 27:72]
  wire [21:0] _T_5936 = _T_4640 ? btb_bank0_rd_data_way1_out_240 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6191 = _T_6190 | _T_5936; // @[Mux.scala 27:72]
  wire [21:0] _T_5937 = _T_4642 ? btb_bank0_rd_data_way1_out_241 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6192 = _T_6191 | _T_5937; // @[Mux.scala 27:72]
  wire [21:0] _T_5938 = _T_4644 ? btb_bank0_rd_data_way1_out_242 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6193 = _T_6192 | _T_5938; // @[Mux.scala 27:72]
  wire [21:0] _T_5939 = _T_4646 ? btb_bank0_rd_data_way1_out_243 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6194 = _T_6193 | _T_5939; // @[Mux.scala 27:72]
  wire [21:0] _T_5940 = _T_4648 ? btb_bank0_rd_data_way1_out_244 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6195 = _T_6194 | _T_5940; // @[Mux.scala 27:72]
  wire [21:0] _T_5941 = _T_4650 ? btb_bank0_rd_data_way1_out_245 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6196 = _T_6195 | _T_5941; // @[Mux.scala 27:72]
  wire [21:0] _T_5942 = _T_4652 ? btb_bank0_rd_data_way1_out_246 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6197 = _T_6196 | _T_5942; // @[Mux.scala 27:72]
  wire [21:0] _T_5943 = _T_4654 ? btb_bank0_rd_data_way1_out_247 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6198 = _T_6197 | _T_5943; // @[Mux.scala 27:72]
  wire [21:0] _T_5944 = _T_4656 ? btb_bank0_rd_data_way1_out_248 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6199 = _T_6198 | _T_5944; // @[Mux.scala 27:72]
  wire [21:0] _T_5945 = _T_4658 ? btb_bank0_rd_data_way1_out_249 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6200 = _T_6199 | _T_5945; // @[Mux.scala 27:72]
  wire [21:0] _T_5946 = _T_4660 ? btb_bank0_rd_data_way1_out_250 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6201 = _T_6200 | _T_5946; // @[Mux.scala 27:72]
  wire [21:0] _T_5947 = _T_4662 ? btb_bank0_rd_data_way1_out_251 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6202 = _T_6201 | _T_5947; // @[Mux.scala 27:72]
  wire [21:0] _T_5948 = _T_4664 ? btb_bank0_rd_data_way1_out_252 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6203 = _T_6202 | _T_5948; // @[Mux.scala 27:72]
  wire [21:0] _T_5949 = _T_4666 ? btb_bank0_rd_data_way1_out_253 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6204 = _T_6203 | _T_5949; // @[Mux.scala 27:72]
  wire [21:0] _T_5950 = _T_4668 ? btb_bank0_rd_data_way1_out_254 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6205 = _T_6204 | _T_5950; // @[Mux.scala 27:72]
  wire [21:0] _T_5951 = _T_4670 ? btb_bank0_rd_data_way1_out_255 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] btb_bank0_rd_data_way1_p1_f = _T_6205 | _T_5951; // @[Mux.scala 27:72]
  wire  _T_73 = btb_bank0_rd_data_way1_p1_f[21:17] == fetch_rd_tag_p1_f; // @[ifu_bp_ctl.scala 138:106]
  wire  _T_74 = btb_bank0_rd_data_way1_p1_f[0] & _T_73; // @[ifu_bp_ctl.scala 138:61]
  wire  _T_77 = _T_74 & _T_67; // @[ifu_bp_ctl.scala 138:129]
  wire  _T_78 = _T_77 & io_ifc_fetch_req_f; // @[ifu_bp_ctl.scala 139:59]
  wire  tag_match_way1_p1_f = _T_78 & _T; // @[ifu_bp_ctl.scala 139:80]
  wire  _T_109 = btb_bank0_rd_data_way1_p1_f[3] ^ btb_bank0_rd_data_way1_p1_f[4]; // @[ifu_bp_ctl.scala 151:100]
  wire  _T_110 = tag_match_way1_p1_f & _T_109; // @[ifu_bp_ctl.scala 151:62]
  wire  _T_114 = ~_T_109; // @[ifu_bp_ctl.scala 152:64]
  wire  _T_115 = tag_match_way1_p1_f & _T_114; // @[ifu_bp_ctl.scala 152:62]
  wire [1:0] tag_match_way1_expanded_p1_f = {_T_110,_T_115}; // @[Cat.scala 29:58]
  wire [21:0] _T_135 = tag_match_way1_expanded_p1_f[0] ? btb_bank0_rd_data_way1_p1_f : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] btb_bank0e_rd_data_p1_f = _T_134 | _T_135; // @[Mux.scala 27:72]
  wire [21:0] _T_147 = io_ifc_fetch_addr_f[0] ? btb_bank0e_rd_data_p1_f : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] btb_vbank1_rd_data_f = _T_146 | _T_147; // @[Mux.scala 27:72]
  wire  _T_243 = btb_vbank1_rd_data_f[2] | btb_vbank1_rd_data_f[1]; // @[ifu_bp_ctl.scala 264:59]
  wire [21:0] _T_120 = tag_match_way0_expanded_f[0] ? btb_bank0_rd_data_way0_f : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_121 = tag_match_way1_expanded_f[0] ? btb_bank0_rd_data_way1_f : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] btb_bank0e_rd_data_f = _T_120 | _T_121; // @[Mux.scala 27:72]
  wire [21:0] _T_140 = _T_144 ? btb_bank0e_rd_data_f : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_141 = io_ifc_fetch_addr_f[0] ? btb_bank0o_rd_data_f : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] btb_vbank0_rd_data_f = _T_140 | _T_141; // @[Mux.scala 27:72]
  wire  _T_246 = btb_vbank0_rd_data_f[2] | btb_vbank0_rd_data_f[1]; // @[ifu_bp_ctl.scala 265:59]
  wire [1:0] bht_force_taken_f = {_T_243,_T_246}; // @[Cat.scala 29:58]
  wire [9:0] _T_570 = {btb_rd_addr_f,2'h0}; // @[Cat.scala 29:58]
  reg [7:0] fghr; // @[ifu_bp_ctl.scala 323:44]
  wire [7:0] bht_rd_addr_f = _T_570[9:2] ^ fghr; // @[lib.scala 56:35]
  wire  _T_21408 = bht_rd_addr_f == 8'h0; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_0; // @[Reg.scala 27:20]
  wire [1:0] _T_21920 = _T_21408 ? bht_bank_rd_data_out_1_0 : 2'h0; // @[Mux.scala 27:72]
  wire  _T_21410 = bht_rd_addr_f == 8'h1; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_1; // @[Reg.scala 27:20]
  wire [1:0] _T_21921 = _T_21410 ? bht_bank_rd_data_out_1_1 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22176 = _T_21920 | _T_21921; // @[Mux.scala 27:72]
  wire  _T_21412 = bht_rd_addr_f == 8'h2; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_2; // @[Reg.scala 27:20]
  wire [1:0] _T_21922 = _T_21412 ? bht_bank_rd_data_out_1_2 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22177 = _T_22176 | _T_21922; // @[Mux.scala 27:72]
  wire  _T_21414 = bht_rd_addr_f == 8'h3; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_3; // @[Reg.scala 27:20]
  wire [1:0] _T_21923 = _T_21414 ? bht_bank_rd_data_out_1_3 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22178 = _T_22177 | _T_21923; // @[Mux.scala 27:72]
  wire  _T_21416 = bht_rd_addr_f == 8'h4; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_4; // @[Reg.scala 27:20]
  wire [1:0] _T_21924 = _T_21416 ? bht_bank_rd_data_out_1_4 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22179 = _T_22178 | _T_21924; // @[Mux.scala 27:72]
  wire  _T_21418 = bht_rd_addr_f == 8'h5; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_5; // @[Reg.scala 27:20]
  wire [1:0] _T_21925 = _T_21418 ? bht_bank_rd_data_out_1_5 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22180 = _T_22179 | _T_21925; // @[Mux.scala 27:72]
  wire  _T_21420 = bht_rd_addr_f == 8'h6; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_6; // @[Reg.scala 27:20]
  wire [1:0] _T_21926 = _T_21420 ? bht_bank_rd_data_out_1_6 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22181 = _T_22180 | _T_21926; // @[Mux.scala 27:72]
  wire  _T_21422 = bht_rd_addr_f == 8'h7; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_7; // @[Reg.scala 27:20]
  wire [1:0] _T_21927 = _T_21422 ? bht_bank_rd_data_out_1_7 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22182 = _T_22181 | _T_21927; // @[Mux.scala 27:72]
  wire  _T_21424 = bht_rd_addr_f == 8'h8; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_8; // @[Reg.scala 27:20]
  wire [1:0] _T_21928 = _T_21424 ? bht_bank_rd_data_out_1_8 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22183 = _T_22182 | _T_21928; // @[Mux.scala 27:72]
  wire  _T_21426 = bht_rd_addr_f == 8'h9; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_9; // @[Reg.scala 27:20]
  wire [1:0] _T_21929 = _T_21426 ? bht_bank_rd_data_out_1_9 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22184 = _T_22183 | _T_21929; // @[Mux.scala 27:72]
  wire  _T_21428 = bht_rd_addr_f == 8'ha; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_10; // @[Reg.scala 27:20]
  wire [1:0] _T_21930 = _T_21428 ? bht_bank_rd_data_out_1_10 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22185 = _T_22184 | _T_21930; // @[Mux.scala 27:72]
  wire  _T_21430 = bht_rd_addr_f == 8'hb; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_11; // @[Reg.scala 27:20]
  wire [1:0] _T_21931 = _T_21430 ? bht_bank_rd_data_out_1_11 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22186 = _T_22185 | _T_21931; // @[Mux.scala 27:72]
  wire  _T_21432 = bht_rd_addr_f == 8'hc; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_12; // @[Reg.scala 27:20]
  wire [1:0] _T_21932 = _T_21432 ? bht_bank_rd_data_out_1_12 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22187 = _T_22186 | _T_21932; // @[Mux.scala 27:72]
  wire  _T_21434 = bht_rd_addr_f == 8'hd; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_13; // @[Reg.scala 27:20]
  wire [1:0] _T_21933 = _T_21434 ? bht_bank_rd_data_out_1_13 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22188 = _T_22187 | _T_21933; // @[Mux.scala 27:72]
  wire  _T_21436 = bht_rd_addr_f == 8'he; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_14; // @[Reg.scala 27:20]
  wire [1:0] _T_21934 = _T_21436 ? bht_bank_rd_data_out_1_14 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22189 = _T_22188 | _T_21934; // @[Mux.scala 27:72]
  wire  _T_21438 = bht_rd_addr_f == 8'hf; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_15; // @[Reg.scala 27:20]
  wire [1:0] _T_21935 = _T_21438 ? bht_bank_rd_data_out_1_15 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22190 = _T_22189 | _T_21935; // @[Mux.scala 27:72]
  wire  _T_21440 = bht_rd_addr_f == 8'h10; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_16; // @[Reg.scala 27:20]
  wire [1:0] _T_21936 = _T_21440 ? bht_bank_rd_data_out_1_16 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22191 = _T_22190 | _T_21936; // @[Mux.scala 27:72]
  wire  _T_21442 = bht_rd_addr_f == 8'h11; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_17; // @[Reg.scala 27:20]
  wire [1:0] _T_21937 = _T_21442 ? bht_bank_rd_data_out_1_17 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22192 = _T_22191 | _T_21937; // @[Mux.scala 27:72]
  wire  _T_21444 = bht_rd_addr_f == 8'h12; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_18; // @[Reg.scala 27:20]
  wire [1:0] _T_21938 = _T_21444 ? bht_bank_rd_data_out_1_18 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22193 = _T_22192 | _T_21938; // @[Mux.scala 27:72]
  wire  _T_21446 = bht_rd_addr_f == 8'h13; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_19; // @[Reg.scala 27:20]
  wire [1:0] _T_21939 = _T_21446 ? bht_bank_rd_data_out_1_19 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22194 = _T_22193 | _T_21939; // @[Mux.scala 27:72]
  wire  _T_21448 = bht_rd_addr_f == 8'h14; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_20; // @[Reg.scala 27:20]
  wire [1:0] _T_21940 = _T_21448 ? bht_bank_rd_data_out_1_20 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22195 = _T_22194 | _T_21940; // @[Mux.scala 27:72]
  wire  _T_21450 = bht_rd_addr_f == 8'h15; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_21; // @[Reg.scala 27:20]
  wire [1:0] _T_21941 = _T_21450 ? bht_bank_rd_data_out_1_21 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22196 = _T_22195 | _T_21941; // @[Mux.scala 27:72]
  wire  _T_21452 = bht_rd_addr_f == 8'h16; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_22; // @[Reg.scala 27:20]
  wire [1:0] _T_21942 = _T_21452 ? bht_bank_rd_data_out_1_22 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22197 = _T_22196 | _T_21942; // @[Mux.scala 27:72]
  wire  _T_21454 = bht_rd_addr_f == 8'h17; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_23; // @[Reg.scala 27:20]
  wire [1:0] _T_21943 = _T_21454 ? bht_bank_rd_data_out_1_23 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22198 = _T_22197 | _T_21943; // @[Mux.scala 27:72]
  wire  _T_21456 = bht_rd_addr_f == 8'h18; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_24; // @[Reg.scala 27:20]
  wire [1:0] _T_21944 = _T_21456 ? bht_bank_rd_data_out_1_24 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22199 = _T_22198 | _T_21944; // @[Mux.scala 27:72]
  wire  _T_21458 = bht_rd_addr_f == 8'h19; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_25; // @[Reg.scala 27:20]
  wire [1:0] _T_21945 = _T_21458 ? bht_bank_rd_data_out_1_25 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22200 = _T_22199 | _T_21945; // @[Mux.scala 27:72]
  wire  _T_21460 = bht_rd_addr_f == 8'h1a; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_26; // @[Reg.scala 27:20]
  wire [1:0] _T_21946 = _T_21460 ? bht_bank_rd_data_out_1_26 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22201 = _T_22200 | _T_21946; // @[Mux.scala 27:72]
  wire  _T_21462 = bht_rd_addr_f == 8'h1b; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_27; // @[Reg.scala 27:20]
  wire [1:0] _T_21947 = _T_21462 ? bht_bank_rd_data_out_1_27 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22202 = _T_22201 | _T_21947; // @[Mux.scala 27:72]
  wire  _T_21464 = bht_rd_addr_f == 8'h1c; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_28; // @[Reg.scala 27:20]
  wire [1:0] _T_21948 = _T_21464 ? bht_bank_rd_data_out_1_28 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22203 = _T_22202 | _T_21948; // @[Mux.scala 27:72]
  wire  _T_21466 = bht_rd_addr_f == 8'h1d; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_29; // @[Reg.scala 27:20]
  wire [1:0] _T_21949 = _T_21466 ? bht_bank_rd_data_out_1_29 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22204 = _T_22203 | _T_21949; // @[Mux.scala 27:72]
  wire  _T_21468 = bht_rd_addr_f == 8'h1e; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_30; // @[Reg.scala 27:20]
  wire [1:0] _T_21950 = _T_21468 ? bht_bank_rd_data_out_1_30 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22205 = _T_22204 | _T_21950; // @[Mux.scala 27:72]
  wire  _T_21470 = bht_rd_addr_f == 8'h1f; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_31; // @[Reg.scala 27:20]
  wire [1:0] _T_21951 = _T_21470 ? bht_bank_rd_data_out_1_31 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22206 = _T_22205 | _T_21951; // @[Mux.scala 27:72]
  wire  _T_21472 = bht_rd_addr_f == 8'h20; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_32; // @[Reg.scala 27:20]
  wire [1:0] _T_21952 = _T_21472 ? bht_bank_rd_data_out_1_32 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22207 = _T_22206 | _T_21952; // @[Mux.scala 27:72]
  wire  _T_21474 = bht_rd_addr_f == 8'h21; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_33; // @[Reg.scala 27:20]
  wire [1:0] _T_21953 = _T_21474 ? bht_bank_rd_data_out_1_33 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22208 = _T_22207 | _T_21953; // @[Mux.scala 27:72]
  wire  _T_21476 = bht_rd_addr_f == 8'h22; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_34; // @[Reg.scala 27:20]
  wire [1:0] _T_21954 = _T_21476 ? bht_bank_rd_data_out_1_34 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22209 = _T_22208 | _T_21954; // @[Mux.scala 27:72]
  wire  _T_21478 = bht_rd_addr_f == 8'h23; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_35; // @[Reg.scala 27:20]
  wire [1:0] _T_21955 = _T_21478 ? bht_bank_rd_data_out_1_35 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22210 = _T_22209 | _T_21955; // @[Mux.scala 27:72]
  wire  _T_21480 = bht_rd_addr_f == 8'h24; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_36; // @[Reg.scala 27:20]
  wire [1:0] _T_21956 = _T_21480 ? bht_bank_rd_data_out_1_36 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22211 = _T_22210 | _T_21956; // @[Mux.scala 27:72]
  wire  _T_21482 = bht_rd_addr_f == 8'h25; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_37; // @[Reg.scala 27:20]
  wire [1:0] _T_21957 = _T_21482 ? bht_bank_rd_data_out_1_37 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22212 = _T_22211 | _T_21957; // @[Mux.scala 27:72]
  wire  _T_21484 = bht_rd_addr_f == 8'h26; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_38; // @[Reg.scala 27:20]
  wire [1:0] _T_21958 = _T_21484 ? bht_bank_rd_data_out_1_38 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22213 = _T_22212 | _T_21958; // @[Mux.scala 27:72]
  wire  _T_21486 = bht_rd_addr_f == 8'h27; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_39; // @[Reg.scala 27:20]
  wire [1:0] _T_21959 = _T_21486 ? bht_bank_rd_data_out_1_39 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22214 = _T_22213 | _T_21959; // @[Mux.scala 27:72]
  wire  _T_21488 = bht_rd_addr_f == 8'h28; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_40; // @[Reg.scala 27:20]
  wire [1:0] _T_21960 = _T_21488 ? bht_bank_rd_data_out_1_40 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22215 = _T_22214 | _T_21960; // @[Mux.scala 27:72]
  wire  _T_21490 = bht_rd_addr_f == 8'h29; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_41; // @[Reg.scala 27:20]
  wire [1:0] _T_21961 = _T_21490 ? bht_bank_rd_data_out_1_41 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22216 = _T_22215 | _T_21961; // @[Mux.scala 27:72]
  wire  _T_21492 = bht_rd_addr_f == 8'h2a; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_42; // @[Reg.scala 27:20]
  wire [1:0] _T_21962 = _T_21492 ? bht_bank_rd_data_out_1_42 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22217 = _T_22216 | _T_21962; // @[Mux.scala 27:72]
  wire  _T_21494 = bht_rd_addr_f == 8'h2b; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_43; // @[Reg.scala 27:20]
  wire [1:0] _T_21963 = _T_21494 ? bht_bank_rd_data_out_1_43 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22218 = _T_22217 | _T_21963; // @[Mux.scala 27:72]
  wire  _T_21496 = bht_rd_addr_f == 8'h2c; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_44; // @[Reg.scala 27:20]
  wire [1:0] _T_21964 = _T_21496 ? bht_bank_rd_data_out_1_44 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22219 = _T_22218 | _T_21964; // @[Mux.scala 27:72]
  wire  _T_21498 = bht_rd_addr_f == 8'h2d; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_45; // @[Reg.scala 27:20]
  wire [1:0] _T_21965 = _T_21498 ? bht_bank_rd_data_out_1_45 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22220 = _T_22219 | _T_21965; // @[Mux.scala 27:72]
  wire  _T_21500 = bht_rd_addr_f == 8'h2e; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_46; // @[Reg.scala 27:20]
  wire [1:0] _T_21966 = _T_21500 ? bht_bank_rd_data_out_1_46 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22221 = _T_22220 | _T_21966; // @[Mux.scala 27:72]
  wire  _T_21502 = bht_rd_addr_f == 8'h2f; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_47; // @[Reg.scala 27:20]
  wire [1:0] _T_21967 = _T_21502 ? bht_bank_rd_data_out_1_47 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22222 = _T_22221 | _T_21967; // @[Mux.scala 27:72]
  wire  _T_21504 = bht_rd_addr_f == 8'h30; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_48; // @[Reg.scala 27:20]
  wire [1:0] _T_21968 = _T_21504 ? bht_bank_rd_data_out_1_48 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22223 = _T_22222 | _T_21968; // @[Mux.scala 27:72]
  wire  _T_21506 = bht_rd_addr_f == 8'h31; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_49; // @[Reg.scala 27:20]
  wire [1:0] _T_21969 = _T_21506 ? bht_bank_rd_data_out_1_49 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22224 = _T_22223 | _T_21969; // @[Mux.scala 27:72]
  wire  _T_21508 = bht_rd_addr_f == 8'h32; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_50; // @[Reg.scala 27:20]
  wire [1:0] _T_21970 = _T_21508 ? bht_bank_rd_data_out_1_50 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22225 = _T_22224 | _T_21970; // @[Mux.scala 27:72]
  wire  _T_21510 = bht_rd_addr_f == 8'h33; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_51; // @[Reg.scala 27:20]
  wire [1:0] _T_21971 = _T_21510 ? bht_bank_rd_data_out_1_51 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22226 = _T_22225 | _T_21971; // @[Mux.scala 27:72]
  wire  _T_21512 = bht_rd_addr_f == 8'h34; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_52; // @[Reg.scala 27:20]
  wire [1:0] _T_21972 = _T_21512 ? bht_bank_rd_data_out_1_52 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22227 = _T_22226 | _T_21972; // @[Mux.scala 27:72]
  wire  _T_21514 = bht_rd_addr_f == 8'h35; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_53; // @[Reg.scala 27:20]
  wire [1:0] _T_21973 = _T_21514 ? bht_bank_rd_data_out_1_53 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22228 = _T_22227 | _T_21973; // @[Mux.scala 27:72]
  wire  _T_21516 = bht_rd_addr_f == 8'h36; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_54; // @[Reg.scala 27:20]
  wire [1:0] _T_21974 = _T_21516 ? bht_bank_rd_data_out_1_54 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22229 = _T_22228 | _T_21974; // @[Mux.scala 27:72]
  wire  _T_21518 = bht_rd_addr_f == 8'h37; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_55; // @[Reg.scala 27:20]
  wire [1:0] _T_21975 = _T_21518 ? bht_bank_rd_data_out_1_55 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22230 = _T_22229 | _T_21975; // @[Mux.scala 27:72]
  wire  _T_21520 = bht_rd_addr_f == 8'h38; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_56; // @[Reg.scala 27:20]
  wire [1:0] _T_21976 = _T_21520 ? bht_bank_rd_data_out_1_56 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22231 = _T_22230 | _T_21976; // @[Mux.scala 27:72]
  wire  _T_21522 = bht_rd_addr_f == 8'h39; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_57; // @[Reg.scala 27:20]
  wire [1:0] _T_21977 = _T_21522 ? bht_bank_rd_data_out_1_57 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22232 = _T_22231 | _T_21977; // @[Mux.scala 27:72]
  wire  _T_21524 = bht_rd_addr_f == 8'h3a; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_58; // @[Reg.scala 27:20]
  wire [1:0] _T_21978 = _T_21524 ? bht_bank_rd_data_out_1_58 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22233 = _T_22232 | _T_21978; // @[Mux.scala 27:72]
  wire  _T_21526 = bht_rd_addr_f == 8'h3b; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_59; // @[Reg.scala 27:20]
  wire [1:0] _T_21979 = _T_21526 ? bht_bank_rd_data_out_1_59 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22234 = _T_22233 | _T_21979; // @[Mux.scala 27:72]
  wire  _T_21528 = bht_rd_addr_f == 8'h3c; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_60; // @[Reg.scala 27:20]
  wire [1:0] _T_21980 = _T_21528 ? bht_bank_rd_data_out_1_60 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22235 = _T_22234 | _T_21980; // @[Mux.scala 27:72]
  wire  _T_21530 = bht_rd_addr_f == 8'h3d; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_61; // @[Reg.scala 27:20]
  wire [1:0] _T_21981 = _T_21530 ? bht_bank_rd_data_out_1_61 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22236 = _T_22235 | _T_21981; // @[Mux.scala 27:72]
  wire  _T_21532 = bht_rd_addr_f == 8'h3e; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_62; // @[Reg.scala 27:20]
  wire [1:0] _T_21982 = _T_21532 ? bht_bank_rd_data_out_1_62 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22237 = _T_22236 | _T_21982; // @[Mux.scala 27:72]
  wire  _T_21534 = bht_rd_addr_f == 8'h3f; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_63; // @[Reg.scala 27:20]
  wire [1:0] _T_21983 = _T_21534 ? bht_bank_rd_data_out_1_63 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22238 = _T_22237 | _T_21983; // @[Mux.scala 27:72]
  wire  _T_21536 = bht_rd_addr_f == 8'h40; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_64; // @[Reg.scala 27:20]
  wire [1:0] _T_21984 = _T_21536 ? bht_bank_rd_data_out_1_64 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22239 = _T_22238 | _T_21984; // @[Mux.scala 27:72]
  wire  _T_21538 = bht_rd_addr_f == 8'h41; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_65; // @[Reg.scala 27:20]
  wire [1:0] _T_21985 = _T_21538 ? bht_bank_rd_data_out_1_65 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22240 = _T_22239 | _T_21985; // @[Mux.scala 27:72]
  wire  _T_21540 = bht_rd_addr_f == 8'h42; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_66; // @[Reg.scala 27:20]
  wire [1:0] _T_21986 = _T_21540 ? bht_bank_rd_data_out_1_66 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22241 = _T_22240 | _T_21986; // @[Mux.scala 27:72]
  wire  _T_21542 = bht_rd_addr_f == 8'h43; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_67; // @[Reg.scala 27:20]
  wire [1:0] _T_21987 = _T_21542 ? bht_bank_rd_data_out_1_67 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22242 = _T_22241 | _T_21987; // @[Mux.scala 27:72]
  wire  _T_21544 = bht_rd_addr_f == 8'h44; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_68; // @[Reg.scala 27:20]
  wire [1:0] _T_21988 = _T_21544 ? bht_bank_rd_data_out_1_68 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22243 = _T_22242 | _T_21988; // @[Mux.scala 27:72]
  wire  _T_21546 = bht_rd_addr_f == 8'h45; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_69; // @[Reg.scala 27:20]
  wire [1:0] _T_21989 = _T_21546 ? bht_bank_rd_data_out_1_69 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22244 = _T_22243 | _T_21989; // @[Mux.scala 27:72]
  wire  _T_21548 = bht_rd_addr_f == 8'h46; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_70; // @[Reg.scala 27:20]
  wire [1:0] _T_21990 = _T_21548 ? bht_bank_rd_data_out_1_70 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22245 = _T_22244 | _T_21990; // @[Mux.scala 27:72]
  wire  _T_21550 = bht_rd_addr_f == 8'h47; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_71; // @[Reg.scala 27:20]
  wire [1:0] _T_21991 = _T_21550 ? bht_bank_rd_data_out_1_71 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22246 = _T_22245 | _T_21991; // @[Mux.scala 27:72]
  wire  _T_21552 = bht_rd_addr_f == 8'h48; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_72; // @[Reg.scala 27:20]
  wire [1:0] _T_21992 = _T_21552 ? bht_bank_rd_data_out_1_72 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22247 = _T_22246 | _T_21992; // @[Mux.scala 27:72]
  wire  _T_21554 = bht_rd_addr_f == 8'h49; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_73; // @[Reg.scala 27:20]
  wire [1:0] _T_21993 = _T_21554 ? bht_bank_rd_data_out_1_73 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22248 = _T_22247 | _T_21993; // @[Mux.scala 27:72]
  wire  _T_21556 = bht_rd_addr_f == 8'h4a; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_74; // @[Reg.scala 27:20]
  wire [1:0] _T_21994 = _T_21556 ? bht_bank_rd_data_out_1_74 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22249 = _T_22248 | _T_21994; // @[Mux.scala 27:72]
  wire  _T_21558 = bht_rd_addr_f == 8'h4b; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_75; // @[Reg.scala 27:20]
  wire [1:0] _T_21995 = _T_21558 ? bht_bank_rd_data_out_1_75 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22250 = _T_22249 | _T_21995; // @[Mux.scala 27:72]
  wire  _T_21560 = bht_rd_addr_f == 8'h4c; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_76; // @[Reg.scala 27:20]
  wire [1:0] _T_21996 = _T_21560 ? bht_bank_rd_data_out_1_76 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22251 = _T_22250 | _T_21996; // @[Mux.scala 27:72]
  wire  _T_21562 = bht_rd_addr_f == 8'h4d; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_77; // @[Reg.scala 27:20]
  wire [1:0] _T_21997 = _T_21562 ? bht_bank_rd_data_out_1_77 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22252 = _T_22251 | _T_21997; // @[Mux.scala 27:72]
  wire  _T_21564 = bht_rd_addr_f == 8'h4e; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_78; // @[Reg.scala 27:20]
  wire [1:0] _T_21998 = _T_21564 ? bht_bank_rd_data_out_1_78 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22253 = _T_22252 | _T_21998; // @[Mux.scala 27:72]
  wire  _T_21566 = bht_rd_addr_f == 8'h4f; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_79; // @[Reg.scala 27:20]
  wire [1:0] _T_21999 = _T_21566 ? bht_bank_rd_data_out_1_79 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22254 = _T_22253 | _T_21999; // @[Mux.scala 27:72]
  wire  _T_21568 = bht_rd_addr_f == 8'h50; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_80; // @[Reg.scala 27:20]
  wire [1:0] _T_22000 = _T_21568 ? bht_bank_rd_data_out_1_80 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22255 = _T_22254 | _T_22000; // @[Mux.scala 27:72]
  wire  _T_21570 = bht_rd_addr_f == 8'h51; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_81; // @[Reg.scala 27:20]
  wire [1:0] _T_22001 = _T_21570 ? bht_bank_rd_data_out_1_81 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22256 = _T_22255 | _T_22001; // @[Mux.scala 27:72]
  wire  _T_21572 = bht_rd_addr_f == 8'h52; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_82; // @[Reg.scala 27:20]
  wire [1:0] _T_22002 = _T_21572 ? bht_bank_rd_data_out_1_82 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22257 = _T_22256 | _T_22002; // @[Mux.scala 27:72]
  wire  _T_21574 = bht_rd_addr_f == 8'h53; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_83; // @[Reg.scala 27:20]
  wire [1:0] _T_22003 = _T_21574 ? bht_bank_rd_data_out_1_83 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22258 = _T_22257 | _T_22003; // @[Mux.scala 27:72]
  wire  _T_21576 = bht_rd_addr_f == 8'h54; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_84; // @[Reg.scala 27:20]
  wire [1:0] _T_22004 = _T_21576 ? bht_bank_rd_data_out_1_84 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22259 = _T_22258 | _T_22004; // @[Mux.scala 27:72]
  wire  _T_21578 = bht_rd_addr_f == 8'h55; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_85; // @[Reg.scala 27:20]
  wire [1:0] _T_22005 = _T_21578 ? bht_bank_rd_data_out_1_85 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22260 = _T_22259 | _T_22005; // @[Mux.scala 27:72]
  wire  _T_21580 = bht_rd_addr_f == 8'h56; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_86; // @[Reg.scala 27:20]
  wire [1:0] _T_22006 = _T_21580 ? bht_bank_rd_data_out_1_86 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22261 = _T_22260 | _T_22006; // @[Mux.scala 27:72]
  wire  _T_21582 = bht_rd_addr_f == 8'h57; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_87; // @[Reg.scala 27:20]
  wire [1:0] _T_22007 = _T_21582 ? bht_bank_rd_data_out_1_87 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22262 = _T_22261 | _T_22007; // @[Mux.scala 27:72]
  wire  _T_21584 = bht_rd_addr_f == 8'h58; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_88; // @[Reg.scala 27:20]
  wire [1:0] _T_22008 = _T_21584 ? bht_bank_rd_data_out_1_88 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22263 = _T_22262 | _T_22008; // @[Mux.scala 27:72]
  wire  _T_21586 = bht_rd_addr_f == 8'h59; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_89; // @[Reg.scala 27:20]
  wire [1:0] _T_22009 = _T_21586 ? bht_bank_rd_data_out_1_89 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22264 = _T_22263 | _T_22009; // @[Mux.scala 27:72]
  wire  _T_21588 = bht_rd_addr_f == 8'h5a; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_90; // @[Reg.scala 27:20]
  wire [1:0] _T_22010 = _T_21588 ? bht_bank_rd_data_out_1_90 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22265 = _T_22264 | _T_22010; // @[Mux.scala 27:72]
  wire  _T_21590 = bht_rd_addr_f == 8'h5b; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_91; // @[Reg.scala 27:20]
  wire [1:0] _T_22011 = _T_21590 ? bht_bank_rd_data_out_1_91 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22266 = _T_22265 | _T_22011; // @[Mux.scala 27:72]
  wire  _T_21592 = bht_rd_addr_f == 8'h5c; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_92; // @[Reg.scala 27:20]
  wire [1:0] _T_22012 = _T_21592 ? bht_bank_rd_data_out_1_92 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22267 = _T_22266 | _T_22012; // @[Mux.scala 27:72]
  wire  _T_21594 = bht_rd_addr_f == 8'h5d; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_93; // @[Reg.scala 27:20]
  wire [1:0] _T_22013 = _T_21594 ? bht_bank_rd_data_out_1_93 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22268 = _T_22267 | _T_22013; // @[Mux.scala 27:72]
  wire  _T_21596 = bht_rd_addr_f == 8'h5e; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_94; // @[Reg.scala 27:20]
  wire [1:0] _T_22014 = _T_21596 ? bht_bank_rd_data_out_1_94 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22269 = _T_22268 | _T_22014; // @[Mux.scala 27:72]
  wire  _T_21598 = bht_rd_addr_f == 8'h5f; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_95; // @[Reg.scala 27:20]
  wire [1:0] _T_22015 = _T_21598 ? bht_bank_rd_data_out_1_95 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22270 = _T_22269 | _T_22015; // @[Mux.scala 27:72]
  wire  _T_21600 = bht_rd_addr_f == 8'h60; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_96; // @[Reg.scala 27:20]
  wire [1:0] _T_22016 = _T_21600 ? bht_bank_rd_data_out_1_96 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22271 = _T_22270 | _T_22016; // @[Mux.scala 27:72]
  wire  _T_21602 = bht_rd_addr_f == 8'h61; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_97; // @[Reg.scala 27:20]
  wire [1:0] _T_22017 = _T_21602 ? bht_bank_rd_data_out_1_97 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22272 = _T_22271 | _T_22017; // @[Mux.scala 27:72]
  wire  _T_21604 = bht_rd_addr_f == 8'h62; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_98; // @[Reg.scala 27:20]
  wire [1:0] _T_22018 = _T_21604 ? bht_bank_rd_data_out_1_98 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22273 = _T_22272 | _T_22018; // @[Mux.scala 27:72]
  wire  _T_21606 = bht_rd_addr_f == 8'h63; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_99; // @[Reg.scala 27:20]
  wire [1:0] _T_22019 = _T_21606 ? bht_bank_rd_data_out_1_99 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22274 = _T_22273 | _T_22019; // @[Mux.scala 27:72]
  wire  _T_21608 = bht_rd_addr_f == 8'h64; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_100; // @[Reg.scala 27:20]
  wire [1:0] _T_22020 = _T_21608 ? bht_bank_rd_data_out_1_100 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22275 = _T_22274 | _T_22020; // @[Mux.scala 27:72]
  wire  _T_21610 = bht_rd_addr_f == 8'h65; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_101; // @[Reg.scala 27:20]
  wire [1:0] _T_22021 = _T_21610 ? bht_bank_rd_data_out_1_101 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22276 = _T_22275 | _T_22021; // @[Mux.scala 27:72]
  wire  _T_21612 = bht_rd_addr_f == 8'h66; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_102; // @[Reg.scala 27:20]
  wire [1:0] _T_22022 = _T_21612 ? bht_bank_rd_data_out_1_102 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22277 = _T_22276 | _T_22022; // @[Mux.scala 27:72]
  wire  _T_21614 = bht_rd_addr_f == 8'h67; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_103; // @[Reg.scala 27:20]
  wire [1:0] _T_22023 = _T_21614 ? bht_bank_rd_data_out_1_103 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22278 = _T_22277 | _T_22023; // @[Mux.scala 27:72]
  wire  _T_21616 = bht_rd_addr_f == 8'h68; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_104; // @[Reg.scala 27:20]
  wire [1:0] _T_22024 = _T_21616 ? bht_bank_rd_data_out_1_104 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22279 = _T_22278 | _T_22024; // @[Mux.scala 27:72]
  wire  _T_21618 = bht_rd_addr_f == 8'h69; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_105; // @[Reg.scala 27:20]
  wire [1:0] _T_22025 = _T_21618 ? bht_bank_rd_data_out_1_105 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22280 = _T_22279 | _T_22025; // @[Mux.scala 27:72]
  wire  _T_21620 = bht_rd_addr_f == 8'h6a; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_106; // @[Reg.scala 27:20]
  wire [1:0] _T_22026 = _T_21620 ? bht_bank_rd_data_out_1_106 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22281 = _T_22280 | _T_22026; // @[Mux.scala 27:72]
  wire  _T_21622 = bht_rd_addr_f == 8'h6b; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_107; // @[Reg.scala 27:20]
  wire [1:0] _T_22027 = _T_21622 ? bht_bank_rd_data_out_1_107 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22282 = _T_22281 | _T_22027; // @[Mux.scala 27:72]
  wire  _T_21624 = bht_rd_addr_f == 8'h6c; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_108; // @[Reg.scala 27:20]
  wire [1:0] _T_22028 = _T_21624 ? bht_bank_rd_data_out_1_108 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22283 = _T_22282 | _T_22028; // @[Mux.scala 27:72]
  wire  _T_21626 = bht_rd_addr_f == 8'h6d; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_109; // @[Reg.scala 27:20]
  wire [1:0] _T_22029 = _T_21626 ? bht_bank_rd_data_out_1_109 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22284 = _T_22283 | _T_22029; // @[Mux.scala 27:72]
  wire  _T_21628 = bht_rd_addr_f == 8'h6e; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_110; // @[Reg.scala 27:20]
  wire [1:0] _T_22030 = _T_21628 ? bht_bank_rd_data_out_1_110 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22285 = _T_22284 | _T_22030; // @[Mux.scala 27:72]
  wire  _T_21630 = bht_rd_addr_f == 8'h6f; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_111; // @[Reg.scala 27:20]
  wire [1:0] _T_22031 = _T_21630 ? bht_bank_rd_data_out_1_111 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22286 = _T_22285 | _T_22031; // @[Mux.scala 27:72]
  wire  _T_21632 = bht_rd_addr_f == 8'h70; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_112; // @[Reg.scala 27:20]
  wire [1:0] _T_22032 = _T_21632 ? bht_bank_rd_data_out_1_112 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22287 = _T_22286 | _T_22032; // @[Mux.scala 27:72]
  wire  _T_21634 = bht_rd_addr_f == 8'h71; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_113; // @[Reg.scala 27:20]
  wire [1:0] _T_22033 = _T_21634 ? bht_bank_rd_data_out_1_113 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22288 = _T_22287 | _T_22033; // @[Mux.scala 27:72]
  wire  _T_21636 = bht_rd_addr_f == 8'h72; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_114; // @[Reg.scala 27:20]
  wire [1:0] _T_22034 = _T_21636 ? bht_bank_rd_data_out_1_114 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22289 = _T_22288 | _T_22034; // @[Mux.scala 27:72]
  wire  _T_21638 = bht_rd_addr_f == 8'h73; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_115; // @[Reg.scala 27:20]
  wire [1:0] _T_22035 = _T_21638 ? bht_bank_rd_data_out_1_115 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22290 = _T_22289 | _T_22035; // @[Mux.scala 27:72]
  wire  _T_21640 = bht_rd_addr_f == 8'h74; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_116; // @[Reg.scala 27:20]
  wire [1:0] _T_22036 = _T_21640 ? bht_bank_rd_data_out_1_116 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22291 = _T_22290 | _T_22036; // @[Mux.scala 27:72]
  wire  _T_21642 = bht_rd_addr_f == 8'h75; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_117; // @[Reg.scala 27:20]
  wire [1:0] _T_22037 = _T_21642 ? bht_bank_rd_data_out_1_117 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22292 = _T_22291 | _T_22037; // @[Mux.scala 27:72]
  wire  _T_21644 = bht_rd_addr_f == 8'h76; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_118; // @[Reg.scala 27:20]
  wire [1:0] _T_22038 = _T_21644 ? bht_bank_rd_data_out_1_118 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22293 = _T_22292 | _T_22038; // @[Mux.scala 27:72]
  wire  _T_21646 = bht_rd_addr_f == 8'h77; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_119; // @[Reg.scala 27:20]
  wire [1:0] _T_22039 = _T_21646 ? bht_bank_rd_data_out_1_119 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22294 = _T_22293 | _T_22039; // @[Mux.scala 27:72]
  wire  _T_21648 = bht_rd_addr_f == 8'h78; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_120; // @[Reg.scala 27:20]
  wire [1:0] _T_22040 = _T_21648 ? bht_bank_rd_data_out_1_120 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22295 = _T_22294 | _T_22040; // @[Mux.scala 27:72]
  wire  _T_21650 = bht_rd_addr_f == 8'h79; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_121; // @[Reg.scala 27:20]
  wire [1:0] _T_22041 = _T_21650 ? bht_bank_rd_data_out_1_121 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22296 = _T_22295 | _T_22041; // @[Mux.scala 27:72]
  wire  _T_21652 = bht_rd_addr_f == 8'h7a; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_122; // @[Reg.scala 27:20]
  wire [1:0] _T_22042 = _T_21652 ? bht_bank_rd_data_out_1_122 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22297 = _T_22296 | _T_22042; // @[Mux.scala 27:72]
  wire  _T_21654 = bht_rd_addr_f == 8'h7b; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_123; // @[Reg.scala 27:20]
  wire [1:0] _T_22043 = _T_21654 ? bht_bank_rd_data_out_1_123 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22298 = _T_22297 | _T_22043; // @[Mux.scala 27:72]
  wire  _T_21656 = bht_rd_addr_f == 8'h7c; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_124; // @[Reg.scala 27:20]
  wire [1:0] _T_22044 = _T_21656 ? bht_bank_rd_data_out_1_124 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22299 = _T_22298 | _T_22044; // @[Mux.scala 27:72]
  wire  _T_21658 = bht_rd_addr_f == 8'h7d; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_125; // @[Reg.scala 27:20]
  wire [1:0] _T_22045 = _T_21658 ? bht_bank_rd_data_out_1_125 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22300 = _T_22299 | _T_22045; // @[Mux.scala 27:72]
  wire  _T_21660 = bht_rd_addr_f == 8'h7e; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_126; // @[Reg.scala 27:20]
  wire [1:0] _T_22046 = _T_21660 ? bht_bank_rd_data_out_1_126 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22301 = _T_22300 | _T_22046; // @[Mux.scala 27:72]
  wire  _T_21662 = bht_rd_addr_f == 8'h7f; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_127; // @[Reg.scala 27:20]
  wire [1:0] _T_22047 = _T_21662 ? bht_bank_rd_data_out_1_127 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22302 = _T_22301 | _T_22047; // @[Mux.scala 27:72]
  wire  _T_21664 = bht_rd_addr_f == 8'h80; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_128; // @[Reg.scala 27:20]
  wire [1:0] _T_22048 = _T_21664 ? bht_bank_rd_data_out_1_128 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22303 = _T_22302 | _T_22048; // @[Mux.scala 27:72]
  wire  _T_21666 = bht_rd_addr_f == 8'h81; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_129; // @[Reg.scala 27:20]
  wire [1:0] _T_22049 = _T_21666 ? bht_bank_rd_data_out_1_129 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22304 = _T_22303 | _T_22049; // @[Mux.scala 27:72]
  wire  _T_21668 = bht_rd_addr_f == 8'h82; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_130; // @[Reg.scala 27:20]
  wire [1:0] _T_22050 = _T_21668 ? bht_bank_rd_data_out_1_130 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22305 = _T_22304 | _T_22050; // @[Mux.scala 27:72]
  wire  _T_21670 = bht_rd_addr_f == 8'h83; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_131; // @[Reg.scala 27:20]
  wire [1:0] _T_22051 = _T_21670 ? bht_bank_rd_data_out_1_131 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22306 = _T_22305 | _T_22051; // @[Mux.scala 27:72]
  wire  _T_21672 = bht_rd_addr_f == 8'h84; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_132; // @[Reg.scala 27:20]
  wire [1:0] _T_22052 = _T_21672 ? bht_bank_rd_data_out_1_132 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22307 = _T_22306 | _T_22052; // @[Mux.scala 27:72]
  wire  _T_21674 = bht_rd_addr_f == 8'h85; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_133; // @[Reg.scala 27:20]
  wire [1:0] _T_22053 = _T_21674 ? bht_bank_rd_data_out_1_133 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22308 = _T_22307 | _T_22053; // @[Mux.scala 27:72]
  wire  _T_21676 = bht_rd_addr_f == 8'h86; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_134; // @[Reg.scala 27:20]
  wire [1:0] _T_22054 = _T_21676 ? bht_bank_rd_data_out_1_134 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22309 = _T_22308 | _T_22054; // @[Mux.scala 27:72]
  wire  _T_21678 = bht_rd_addr_f == 8'h87; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_135; // @[Reg.scala 27:20]
  wire [1:0] _T_22055 = _T_21678 ? bht_bank_rd_data_out_1_135 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22310 = _T_22309 | _T_22055; // @[Mux.scala 27:72]
  wire  _T_21680 = bht_rd_addr_f == 8'h88; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_136; // @[Reg.scala 27:20]
  wire [1:0] _T_22056 = _T_21680 ? bht_bank_rd_data_out_1_136 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22311 = _T_22310 | _T_22056; // @[Mux.scala 27:72]
  wire  _T_21682 = bht_rd_addr_f == 8'h89; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_137; // @[Reg.scala 27:20]
  wire [1:0] _T_22057 = _T_21682 ? bht_bank_rd_data_out_1_137 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22312 = _T_22311 | _T_22057; // @[Mux.scala 27:72]
  wire  _T_21684 = bht_rd_addr_f == 8'h8a; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_138; // @[Reg.scala 27:20]
  wire [1:0] _T_22058 = _T_21684 ? bht_bank_rd_data_out_1_138 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22313 = _T_22312 | _T_22058; // @[Mux.scala 27:72]
  wire  _T_21686 = bht_rd_addr_f == 8'h8b; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_139; // @[Reg.scala 27:20]
  wire [1:0] _T_22059 = _T_21686 ? bht_bank_rd_data_out_1_139 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22314 = _T_22313 | _T_22059; // @[Mux.scala 27:72]
  wire  _T_21688 = bht_rd_addr_f == 8'h8c; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_140; // @[Reg.scala 27:20]
  wire [1:0] _T_22060 = _T_21688 ? bht_bank_rd_data_out_1_140 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22315 = _T_22314 | _T_22060; // @[Mux.scala 27:72]
  wire  _T_21690 = bht_rd_addr_f == 8'h8d; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_141; // @[Reg.scala 27:20]
  wire [1:0] _T_22061 = _T_21690 ? bht_bank_rd_data_out_1_141 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22316 = _T_22315 | _T_22061; // @[Mux.scala 27:72]
  wire  _T_21692 = bht_rd_addr_f == 8'h8e; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_142; // @[Reg.scala 27:20]
  wire [1:0] _T_22062 = _T_21692 ? bht_bank_rd_data_out_1_142 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22317 = _T_22316 | _T_22062; // @[Mux.scala 27:72]
  wire  _T_21694 = bht_rd_addr_f == 8'h8f; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_143; // @[Reg.scala 27:20]
  wire [1:0] _T_22063 = _T_21694 ? bht_bank_rd_data_out_1_143 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22318 = _T_22317 | _T_22063; // @[Mux.scala 27:72]
  wire  _T_21696 = bht_rd_addr_f == 8'h90; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_144; // @[Reg.scala 27:20]
  wire [1:0] _T_22064 = _T_21696 ? bht_bank_rd_data_out_1_144 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22319 = _T_22318 | _T_22064; // @[Mux.scala 27:72]
  wire  _T_21698 = bht_rd_addr_f == 8'h91; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_145; // @[Reg.scala 27:20]
  wire [1:0] _T_22065 = _T_21698 ? bht_bank_rd_data_out_1_145 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22320 = _T_22319 | _T_22065; // @[Mux.scala 27:72]
  wire  _T_21700 = bht_rd_addr_f == 8'h92; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_146; // @[Reg.scala 27:20]
  wire [1:0] _T_22066 = _T_21700 ? bht_bank_rd_data_out_1_146 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22321 = _T_22320 | _T_22066; // @[Mux.scala 27:72]
  wire  _T_21702 = bht_rd_addr_f == 8'h93; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_147; // @[Reg.scala 27:20]
  wire [1:0] _T_22067 = _T_21702 ? bht_bank_rd_data_out_1_147 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22322 = _T_22321 | _T_22067; // @[Mux.scala 27:72]
  wire  _T_21704 = bht_rd_addr_f == 8'h94; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_148; // @[Reg.scala 27:20]
  wire [1:0] _T_22068 = _T_21704 ? bht_bank_rd_data_out_1_148 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22323 = _T_22322 | _T_22068; // @[Mux.scala 27:72]
  wire  _T_21706 = bht_rd_addr_f == 8'h95; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_149; // @[Reg.scala 27:20]
  wire [1:0] _T_22069 = _T_21706 ? bht_bank_rd_data_out_1_149 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22324 = _T_22323 | _T_22069; // @[Mux.scala 27:72]
  wire  _T_21708 = bht_rd_addr_f == 8'h96; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_150; // @[Reg.scala 27:20]
  wire [1:0] _T_22070 = _T_21708 ? bht_bank_rd_data_out_1_150 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22325 = _T_22324 | _T_22070; // @[Mux.scala 27:72]
  wire  _T_21710 = bht_rd_addr_f == 8'h97; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_151; // @[Reg.scala 27:20]
  wire [1:0] _T_22071 = _T_21710 ? bht_bank_rd_data_out_1_151 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22326 = _T_22325 | _T_22071; // @[Mux.scala 27:72]
  wire  _T_21712 = bht_rd_addr_f == 8'h98; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_152; // @[Reg.scala 27:20]
  wire [1:0] _T_22072 = _T_21712 ? bht_bank_rd_data_out_1_152 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22327 = _T_22326 | _T_22072; // @[Mux.scala 27:72]
  wire  _T_21714 = bht_rd_addr_f == 8'h99; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_153; // @[Reg.scala 27:20]
  wire [1:0] _T_22073 = _T_21714 ? bht_bank_rd_data_out_1_153 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22328 = _T_22327 | _T_22073; // @[Mux.scala 27:72]
  wire  _T_21716 = bht_rd_addr_f == 8'h9a; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_154; // @[Reg.scala 27:20]
  wire [1:0] _T_22074 = _T_21716 ? bht_bank_rd_data_out_1_154 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22329 = _T_22328 | _T_22074; // @[Mux.scala 27:72]
  wire  _T_21718 = bht_rd_addr_f == 8'h9b; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_155; // @[Reg.scala 27:20]
  wire [1:0] _T_22075 = _T_21718 ? bht_bank_rd_data_out_1_155 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22330 = _T_22329 | _T_22075; // @[Mux.scala 27:72]
  wire  _T_21720 = bht_rd_addr_f == 8'h9c; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_156; // @[Reg.scala 27:20]
  wire [1:0] _T_22076 = _T_21720 ? bht_bank_rd_data_out_1_156 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22331 = _T_22330 | _T_22076; // @[Mux.scala 27:72]
  wire  _T_21722 = bht_rd_addr_f == 8'h9d; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_157; // @[Reg.scala 27:20]
  wire [1:0] _T_22077 = _T_21722 ? bht_bank_rd_data_out_1_157 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22332 = _T_22331 | _T_22077; // @[Mux.scala 27:72]
  wire  _T_21724 = bht_rd_addr_f == 8'h9e; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_158; // @[Reg.scala 27:20]
  wire [1:0] _T_22078 = _T_21724 ? bht_bank_rd_data_out_1_158 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22333 = _T_22332 | _T_22078; // @[Mux.scala 27:72]
  wire  _T_21726 = bht_rd_addr_f == 8'h9f; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_159; // @[Reg.scala 27:20]
  wire [1:0] _T_22079 = _T_21726 ? bht_bank_rd_data_out_1_159 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22334 = _T_22333 | _T_22079; // @[Mux.scala 27:72]
  wire  _T_21728 = bht_rd_addr_f == 8'ha0; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_160; // @[Reg.scala 27:20]
  wire [1:0] _T_22080 = _T_21728 ? bht_bank_rd_data_out_1_160 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22335 = _T_22334 | _T_22080; // @[Mux.scala 27:72]
  wire  _T_21730 = bht_rd_addr_f == 8'ha1; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_161; // @[Reg.scala 27:20]
  wire [1:0] _T_22081 = _T_21730 ? bht_bank_rd_data_out_1_161 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22336 = _T_22335 | _T_22081; // @[Mux.scala 27:72]
  wire  _T_21732 = bht_rd_addr_f == 8'ha2; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_162; // @[Reg.scala 27:20]
  wire [1:0] _T_22082 = _T_21732 ? bht_bank_rd_data_out_1_162 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22337 = _T_22336 | _T_22082; // @[Mux.scala 27:72]
  wire  _T_21734 = bht_rd_addr_f == 8'ha3; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_163; // @[Reg.scala 27:20]
  wire [1:0] _T_22083 = _T_21734 ? bht_bank_rd_data_out_1_163 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22338 = _T_22337 | _T_22083; // @[Mux.scala 27:72]
  wire  _T_21736 = bht_rd_addr_f == 8'ha4; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_164; // @[Reg.scala 27:20]
  wire [1:0] _T_22084 = _T_21736 ? bht_bank_rd_data_out_1_164 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22339 = _T_22338 | _T_22084; // @[Mux.scala 27:72]
  wire  _T_21738 = bht_rd_addr_f == 8'ha5; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_165; // @[Reg.scala 27:20]
  wire [1:0] _T_22085 = _T_21738 ? bht_bank_rd_data_out_1_165 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22340 = _T_22339 | _T_22085; // @[Mux.scala 27:72]
  wire  _T_21740 = bht_rd_addr_f == 8'ha6; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_166; // @[Reg.scala 27:20]
  wire [1:0] _T_22086 = _T_21740 ? bht_bank_rd_data_out_1_166 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22341 = _T_22340 | _T_22086; // @[Mux.scala 27:72]
  wire  _T_21742 = bht_rd_addr_f == 8'ha7; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_167; // @[Reg.scala 27:20]
  wire [1:0] _T_22087 = _T_21742 ? bht_bank_rd_data_out_1_167 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22342 = _T_22341 | _T_22087; // @[Mux.scala 27:72]
  wire  _T_21744 = bht_rd_addr_f == 8'ha8; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_168; // @[Reg.scala 27:20]
  wire [1:0] _T_22088 = _T_21744 ? bht_bank_rd_data_out_1_168 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22343 = _T_22342 | _T_22088; // @[Mux.scala 27:72]
  wire  _T_21746 = bht_rd_addr_f == 8'ha9; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_169; // @[Reg.scala 27:20]
  wire [1:0] _T_22089 = _T_21746 ? bht_bank_rd_data_out_1_169 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22344 = _T_22343 | _T_22089; // @[Mux.scala 27:72]
  wire  _T_21748 = bht_rd_addr_f == 8'haa; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_170; // @[Reg.scala 27:20]
  wire [1:0] _T_22090 = _T_21748 ? bht_bank_rd_data_out_1_170 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22345 = _T_22344 | _T_22090; // @[Mux.scala 27:72]
  wire  _T_21750 = bht_rd_addr_f == 8'hab; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_171; // @[Reg.scala 27:20]
  wire [1:0] _T_22091 = _T_21750 ? bht_bank_rd_data_out_1_171 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22346 = _T_22345 | _T_22091; // @[Mux.scala 27:72]
  wire  _T_21752 = bht_rd_addr_f == 8'hac; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_172; // @[Reg.scala 27:20]
  wire [1:0] _T_22092 = _T_21752 ? bht_bank_rd_data_out_1_172 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22347 = _T_22346 | _T_22092; // @[Mux.scala 27:72]
  wire  _T_21754 = bht_rd_addr_f == 8'had; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_173; // @[Reg.scala 27:20]
  wire [1:0] _T_22093 = _T_21754 ? bht_bank_rd_data_out_1_173 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22348 = _T_22347 | _T_22093; // @[Mux.scala 27:72]
  wire  _T_21756 = bht_rd_addr_f == 8'hae; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_174; // @[Reg.scala 27:20]
  wire [1:0] _T_22094 = _T_21756 ? bht_bank_rd_data_out_1_174 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22349 = _T_22348 | _T_22094; // @[Mux.scala 27:72]
  wire  _T_21758 = bht_rd_addr_f == 8'haf; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_175; // @[Reg.scala 27:20]
  wire [1:0] _T_22095 = _T_21758 ? bht_bank_rd_data_out_1_175 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22350 = _T_22349 | _T_22095; // @[Mux.scala 27:72]
  wire  _T_21760 = bht_rd_addr_f == 8'hb0; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_176; // @[Reg.scala 27:20]
  wire [1:0] _T_22096 = _T_21760 ? bht_bank_rd_data_out_1_176 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22351 = _T_22350 | _T_22096; // @[Mux.scala 27:72]
  wire  _T_21762 = bht_rd_addr_f == 8'hb1; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_177; // @[Reg.scala 27:20]
  wire [1:0] _T_22097 = _T_21762 ? bht_bank_rd_data_out_1_177 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22352 = _T_22351 | _T_22097; // @[Mux.scala 27:72]
  wire  _T_21764 = bht_rd_addr_f == 8'hb2; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_178; // @[Reg.scala 27:20]
  wire [1:0] _T_22098 = _T_21764 ? bht_bank_rd_data_out_1_178 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22353 = _T_22352 | _T_22098; // @[Mux.scala 27:72]
  wire  _T_21766 = bht_rd_addr_f == 8'hb3; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_179; // @[Reg.scala 27:20]
  wire [1:0] _T_22099 = _T_21766 ? bht_bank_rd_data_out_1_179 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22354 = _T_22353 | _T_22099; // @[Mux.scala 27:72]
  wire  _T_21768 = bht_rd_addr_f == 8'hb4; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_180; // @[Reg.scala 27:20]
  wire [1:0] _T_22100 = _T_21768 ? bht_bank_rd_data_out_1_180 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22355 = _T_22354 | _T_22100; // @[Mux.scala 27:72]
  wire  _T_21770 = bht_rd_addr_f == 8'hb5; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_181; // @[Reg.scala 27:20]
  wire [1:0] _T_22101 = _T_21770 ? bht_bank_rd_data_out_1_181 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22356 = _T_22355 | _T_22101; // @[Mux.scala 27:72]
  wire  _T_21772 = bht_rd_addr_f == 8'hb6; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_182; // @[Reg.scala 27:20]
  wire [1:0] _T_22102 = _T_21772 ? bht_bank_rd_data_out_1_182 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22357 = _T_22356 | _T_22102; // @[Mux.scala 27:72]
  wire  _T_21774 = bht_rd_addr_f == 8'hb7; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_183; // @[Reg.scala 27:20]
  wire [1:0] _T_22103 = _T_21774 ? bht_bank_rd_data_out_1_183 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22358 = _T_22357 | _T_22103; // @[Mux.scala 27:72]
  wire  _T_21776 = bht_rd_addr_f == 8'hb8; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_184; // @[Reg.scala 27:20]
  wire [1:0] _T_22104 = _T_21776 ? bht_bank_rd_data_out_1_184 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22359 = _T_22358 | _T_22104; // @[Mux.scala 27:72]
  wire  _T_21778 = bht_rd_addr_f == 8'hb9; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_185; // @[Reg.scala 27:20]
  wire [1:0] _T_22105 = _T_21778 ? bht_bank_rd_data_out_1_185 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22360 = _T_22359 | _T_22105; // @[Mux.scala 27:72]
  wire  _T_21780 = bht_rd_addr_f == 8'hba; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_186; // @[Reg.scala 27:20]
  wire [1:0] _T_22106 = _T_21780 ? bht_bank_rd_data_out_1_186 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22361 = _T_22360 | _T_22106; // @[Mux.scala 27:72]
  wire  _T_21782 = bht_rd_addr_f == 8'hbb; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_187; // @[Reg.scala 27:20]
  wire [1:0] _T_22107 = _T_21782 ? bht_bank_rd_data_out_1_187 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22362 = _T_22361 | _T_22107; // @[Mux.scala 27:72]
  wire  _T_21784 = bht_rd_addr_f == 8'hbc; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_188; // @[Reg.scala 27:20]
  wire [1:0] _T_22108 = _T_21784 ? bht_bank_rd_data_out_1_188 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22363 = _T_22362 | _T_22108; // @[Mux.scala 27:72]
  wire  _T_21786 = bht_rd_addr_f == 8'hbd; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_189; // @[Reg.scala 27:20]
  wire [1:0] _T_22109 = _T_21786 ? bht_bank_rd_data_out_1_189 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22364 = _T_22363 | _T_22109; // @[Mux.scala 27:72]
  wire  _T_21788 = bht_rd_addr_f == 8'hbe; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_190; // @[Reg.scala 27:20]
  wire [1:0] _T_22110 = _T_21788 ? bht_bank_rd_data_out_1_190 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22365 = _T_22364 | _T_22110; // @[Mux.scala 27:72]
  wire  _T_21790 = bht_rd_addr_f == 8'hbf; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_191; // @[Reg.scala 27:20]
  wire [1:0] _T_22111 = _T_21790 ? bht_bank_rd_data_out_1_191 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22366 = _T_22365 | _T_22111; // @[Mux.scala 27:72]
  wire  _T_21792 = bht_rd_addr_f == 8'hc0; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_192; // @[Reg.scala 27:20]
  wire [1:0] _T_22112 = _T_21792 ? bht_bank_rd_data_out_1_192 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22367 = _T_22366 | _T_22112; // @[Mux.scala 27:72]
  wire  _T_21794 = bht_rd_addr_f == 8'hc1; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_193; // @[Reg.scala 27:20]
  wire [1:0] _T_22113 = _T_21794 ? bht_bank_rd_data_out_1_193 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22368 = _T_22367 | _T_22113; // @[Mux.scala 27:72]
  wire  _T_21796 = bht_rd_addr_f == 8'hc2; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_194; // @[Reg.scala 27:20]
  wire [1:0] _T_22114 = _T_21796 ? bht_bank_rd_data_out_1_194 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22369 = _T_22368 | _T_22114; // @[Mux.scala 27:72]
  wire  _T_21798 = bht_rd_addr_f == 8'hc3; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_195; // @[Reg.scala 27:20]
  wire [1:0] _T_22115 = _T_21798 ? bht_bank_rd_data_out_1_195 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22370 = _T_22369 | _T_22115; // @[Mux.scala 27:72]
  wire  _T_21800 = bht_rd_addr_f == 8'hc4; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_196; // @[Reg.scala 27:20]
  wire [1:0] _T_22116 = _T_21800 ? bht_bank_rd_data_out_1_196 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22371 = _T_22370 | _T_22116; // @[Mux.scala 27:72]
  wire  _T_21802 = bht_rd_addr_f == 8'hc5; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_197; // @[Reg.scala 27:20]
  wire [1:0] _T_22117 = _T_21802 ? bht_bank_rd_data_out_1_197 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22372 = _T_22371 | _T_22117; // @[Mux.scala 27:72]
  wire  _T_21804 = bht_rd_addr_f == 8'hc6; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_198; // @[Reg.scala 27:20]
  wire [1:0] _T_22118 = _T_21804 ? bht_bank_rd_data_out_1_198 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22373 = _T_22372 | _T_22118; // @[Mux.scala 27:72]
  wire  _T_21806 = bht_rd_addr_f == 8'hc7; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_199; // @[Reg.scala 27:20]
  wire [1:0] _T_22119 = _T_21806 ? bht_bank_rd_data_out_1_199 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22374 = _T_22373 | _T_22119; // @[Mux.scala 27:72]
  wire  _T_21808 = bht_rd_addr_f == 8'hc8; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_200; // @[Reg.scala 27:20]
  wire [1:0] _T_22120 = _T_21808 ? bht_bank_rd_data_out_1_200 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22375 = _T_22374 | _T_22120; // @[Mux.scala 27:72]
  wire  _T_21810 = bht_rd_addr_f == 8'hc9; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_201; // @[Reg.scala 27:20]
  wire [1:0] _T_22121 = _T_21810 ? bht_bank_rd_data_out_1_201 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22376 = _T_22375 | _T_22121; // @[Mux.scala 27:72]
  wire  _T_21812 = bht_rd_addr_f == 8'hca; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_202; // @[Reg.scala 27:20]
  wire [1:0] _T_22122 = _T_21812 ? bht_bank_rd_data_out_1_202 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22377 = _T_22376 | _T_22122; // @[Mux.scala 27:72]
  wire  _T_21814 = bht_rd_addr_f == 8'hcb; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_203; // @[Reg.scala 27:20]
  wire [1:0] _T_22123 = _T_21814 ? bht_bank_rd_data_out_1_203 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22378 = _T_22377 | _T_22123; // @[Mux.scala 27:72]
  wire  _T_21816 = bht_rd_addr_f == 8'hcc; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_204; // @[Reg.scala 27:20]
  wire [1:0] _T_22124 = _T_21816 ? bht_bank_rd_data_out_1_204 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22379 = _T_22378 | _T_22124; // @[Mux.scala 27:72]
  wire  _T_21818 = bht_rd_addr_f == 8'hcd; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_205; // @[Reg.scala 27:20]
  wire [1:0] _T_22125 = _T_21818 ? bht_bank_rd_data_out_1_205 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22380 = _T_22379 | _T_22125; // @[Mux.scala 27:72]
  wire  _T_21820 = bht_rd_addr_f == 8'hce; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_206; // @[Reg.scala 27:20]
  wire [1:0] _T_22126 = _T_21820 ? bht_bank_rd_data_out_1_206 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22381 = _T_22380 | _T_22126; // @[Mux.scala 27:72]
  wire  _T_21822 = bht_rd_addr_f == 8'hcf; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_207; // @[Reg.scala 27:20]
  wire [1:0] _T_22127 = _T_21822 ? bht_bank_rd_data_out_1_207 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22382 = _T_22381 | _T_22127; // @[Mux.scala 27:72]
  wire  _T_21824 = bht_rd_addr_f == 8'hd0; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_208; // @[Reg.scala 27:20]
  wire [1:0] _T_22128 = _T_21824 ? bht_bank_rd_data_out_1_208 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22383 = _T_22382 | _T_22128; // @[Mux.scala 27:72]
  wire  _T_21826 = bht_rd_addr_f == 8'hd1; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_209; // @[Reg.scala 27:20]
  wire [1:0] _T_22129 = _T_21826 ? bht_bank_rd_data_out_1_209 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22384 = _T_22383 | _T_22129; // @[Mux.scala 27:72]
  wire  _T_21828 = bht_rd_addr_f == 8'hd2; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_210; // @[Reg.scala 27:20]
  wire [1:0] _T_22130 = _T_21828 ? bht_bank_rd_data_out_1_210 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22385 = _T_22384 | _T_22130; // @[Mux.scala 27:72]
  wire  _T_21830 = bht_rd_addr_f == 8'hd3; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_211; // @[Reg.scala 27:20]
  wire [1:0] _T_22131 = _T_21830 ? bht_bank_rd_data_out_1_211 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22386 = _T_22385 | _T_22131; // @[Mux.scala 27:72]
  wire  _T_21832 = bht_rd_addr_f == 8'hd4; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_212; // @[Reg.scala 27:20]
  wire [1:0] _T_22132 = _T_21832 ? bht_bank_rd_data_out_1_212 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22387 = _T_22386 | _T_22132; // @[Mux.scala 27:72]
  wire  _T_21834 = bht_rd_addr_f == 8'hd5; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_213; // @[Reg.scala 27:20]
  wire [1:0] _T_22133 = _T_21834 ? bht_bank_rd_data_out_1_213 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22388 = _T_22387 | _T_22133; // @[Mux.scala 27:72]
  wire  _T_21836 = bht_rd_addr_f == 8'hd6; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_214; // @[Reg.scala 27:20]
  wire [1:0] _T_22134 = _T_21836 ? bht_bank_rd_data_out_1_214 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22389 = _T_22388 | _T_22134; // @[Mux.scala 27:72]
  wire  _T_21838 = bht_rd_addr_f == 8'hd7; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_215; // @[Reg.scala 27:20]
  wire [1:0] _T_22135 = _T_21838 ? bht_bank_rd_data_out_1_215 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22390 = _T_22389 | _T_22135; // @[Mux.scala 27:72]
  wire  _T_21840 = bht_rd_addr_f == 8'hd8; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_216; // @[Reg.scala 27:20]
  wire [1:0] _T_22136 = _T_21840 ? bht_bank_rd_data_out_1_216 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22391 = _T_22390 | _T_22136; // @[Mux.scala 27:72]
  wire  _T_21842 = bht_rd_addr_f == 8'hd9; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_217; // @[Reg.scala 27:20]
  wire [1:0] _T_22137 = _T_21842 ? bht_bank_rd_data_out_1_217 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22392 = _T_22391 | _T_22137; // @[Mux.scala 27:72]
  wire  _T_21844 = bht_rd_addr_f == 8'hda; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_218; // @[Reg.scala 27:20]
  wire [1:0] _T_22138 = _T_21844 ? bht_bank_rd_data_out_1_218 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22393 = _T_22392 | _T_22138; // @[Mux.scala 27:72]
  wire  _T_21846 = bht_rd_addr_f == 8'hdb; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_219; // @[Reg.scala 27:20]
  wire [1:0] _T_22139 = _T_21846 ? bht_bank_rd_data_out_1_219 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22394 = _T_22393 | _T_22139; // @[Mux.scala 27:72]
  wire  _T_21848 = bht_rd_addr_f == 8'hdc; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_220; // @[Reg.scala 27:20]
  wire [1:0] _T_22140 = _T_21848 ? bht_bank_rd_data_out_1_220 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22395 = _T_22394 | _T_22140; // @[Mux.scala 27:72]
  wire  _T_21850 = bht_rd_addr_f == 8'hdd; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_221; // @[Reg.scala 27:20]
  wire [1:0] _T_22141 = _T_21850 ? bht_bank_rd_data_out_1_221 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22396 = _T_22395 | _T_22141; // @[Mux.scala 27:72]
  wire  _T_21852 = bht_rd_addr_f == 8'hde; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_222; // @[Reg.scala 27:20]
  wire [1:0] _T_22142 = _T_21852 ? bht_bank_rd_data_out_1_222 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22397 = _T_22396 | _T_22142; // @[Mux.scala 27:72]
  wire  _T_21854 = bht_rd_addr_f == 8'hdf; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_223; // @[Reg.scala 27:20]
  wire [1:0] _T_22143 = _T_21854 ? bht_bank_rd_data_out_1_223 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22398 = _T_22397 | _T_22143; // @[Mux.scala 27:72]
  wire  _T_21856 = bht_rd_addr_f == 8'he0; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_224; // @[Reg.scala 27:20]
  wire [1:0] _T_22144 = _T_21856 ? bht_bank_rd_data_out_1_224 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22399 = _T_22398 | _T_22144; // @[Mux.scala 27:72]
  wire  _T_21858 = bht_rd_addr_f == 8'he1; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_225; // @[Reg.scala 27:20]
  wire [1:0] _T_22145 = _T_21858 ? bht_bank_rd_data_out_1_225 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22400 = _T_22399 | _T_22145; // @[Mux.scala 27:72]
  wire  _T_21860 = bht_rd_addr_f == 8'he2; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_226; // @[Reg.scala 27:20]
  wire [1:0] _T_22146 = _T_21860 ? bht_bank_rd_data_out_1_226 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22401 = _T_22400 | _T_22146; // @[Mux.scala 27:72]
  wire  _T_21862 = bht_rd_addr_f == 8'he3; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_227; // @[Reg.scala 27:20]
  wire [1:0] _T_22147 = _T_21862 ? bht_bank_rd_data_out_1_227 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22402 = _T_22401 | _T_22147; // @[Mux.scala 27:72]
  wire  _T_21864 = bht_rd_addr_f == 8'he4; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_228; // @[Reg.scala 27:20]
  wire [1:0] _T_22148 = _T_21864 ? bht_bank_rd_data_out_1_228 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22403 = _T_22402 | _T_22148; // @[Mux.scala 27:72]
  wire  _T_21866 = bht_rd_addr_f == 8'he5; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_229; // @[Reg.scala 27:20]
  wire [1:0] _T_22149 = _T_21866 ? bht_bank_rd_data_out_1_229 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22404 = _T_22403 | _T_22149; // @[Mux.scala 27:72]
  wire  _T_21868 = bht_rd_addr_f == 8'he6; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_230; // @[Reg.scala 27:20]
  wire [1:0] _T_22150 = _T_21868 ? bht_bank_rd_data_out_1_230 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22405 = _T_22404 | _T_22150; // @[Mux.scala 27:72]
  wire  _T_21870 = bht_rd_addr_f == 8'he7; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_231; // @[Reg.scala 27:20]
  wire [1:0] _T_22151 = _T_21870 ? bht_bank_rd_data_out_1_231 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22406 = _T_22405 | _T_22151; // @[Mux.scala 27:72]
  wire  _T_21872 = bht_rd_addr_f == 8'he8; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_232; // @[Reg.scala 27:20]
  wire [1:0] _T_22152 = _T_21872 ? bht_bank_rd_data_out_1_232 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22407 = _T_22406 | _T_22152; // @[Mux.scala 27:72]
  wire  _T_21874 = bht_rd_addr_f == 8'he9; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_233; // @[Reg.scala 27:20]
  wire [1:0] _T_22153 = _T_21874 ? bht_bank_rd_data_out_1_233 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22408 = _T_22407 | _T_22153; // @[Mux.scala 27:72]
  wire  _T_21876 = bht_rd_addr_f == 8'hea; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_234; // @[Reg.scala 27:20]
  wire [1:0] _T_22154 = _T_21876 ? bht_bank_rd_data_out_1_234 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22409 = _T_22408 | _T_22154; // @[Mux.scala 27:72]
  wire  _T_21878 = bht_rd_addr_f == 8'heb; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_235; // @[Reg.scala 27:20]
  wire [1:0] _T_22155 = _T_21878 ? bht_bank_rd_data_out_1_235 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22410 = _T_22409 | _T_22155; // @[Mux.scala 27:72]
  wire  _T_21880 = bht_rd_addr_f == 8'hec; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_236; // @[Reg.scala 27:20]
  wire [1:0] _T_22156 = _T_21880 ? bht_bank_rd_data_out_1_236 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22411 = _T_22410 | _T_22156; // @[Mux.scala 27:72]
  wire  _T_21882 = bht_rd_addr_f == 8'hed; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_237; // @[Reg.scala 27:20]
  wire [1:0] _T_22157 = _T_21882 ? bht_bank_rd_data_out_1_237 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22412 = _T_22411 | _T_22157; // @[Mux.scala 27:72]
  wire  _T_21884 = bht_rd_addr_f == 8'hee; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_238; // @[Reg.scala 27:20]
  wire [1:0] _T_22158 = _T_21884 ? bht_bank_rd_data_out_1_238 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22413 = _T_22412 | _T_22158; // @[Mux.scala 27:72]
  wire  _T_21886 = bht_rd_addr_f == 8'hef; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_239; // @[Reg.scala 27:20]
  wire [1:0] _T_22159 = _T_21886 ? bht_bank_rd_data_out_1_239 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22414 = _T_22413 | _T_22159; // @[Mux.scala 27:72]
  wire  _T_21888 = bht_rd_addr_f == 8'hf0; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_240; // @[Reg.scala 27:20]
  wire [1:0] _T_22160 = _T_21888 ? bht_bank_rd_data_out_1_240 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22415 = _T_22414 | _T_22160; // @[Mux.scala 27:72]
  wire  _T_21890 = bht_rd_addr_f == 8'hf1; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_241; // @[Reg.scala 27:20]
  wire [1:0] _T_22161 = _T_21890 ? bht_bank_rd_data_out_1_241 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22416 = _T_22415 | _T_22161; // @[Mux.scala 27:72]
  wire  _T_21892 = bht_rd_addr_f == 8'hf2; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_242; // @[Reg.scala 27:20]
  wire [1:0] _T_22162 = _T_21892 ? bht_bank_rd_data_out_1_242 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22417 = _T_22416 | _T_22162; // @[Mux.scala 27:72]
  wire  _T_21894 = bht_rd_addr_f == 8'hf3; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_243; // @[Reg.scala 27:20]
  wire [1:0] _T_22163 = _T_21894 ? bht_bank_rd_data_out_1_243 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22418 = _T_22417 | _T_22163; // @[Mux.scala 27:72]
  wire  _T_21896 = bht_rd_addr_f == 8'hf4; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_244; // @[Reg.scala 27:20]
  wire [1:0] _T_22164 = _T_21896 ? bht_bank_rd_data_out_1_244 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22419 = _T_22418 | _T_22164; // @[Mux.scala 27:72]
  wire  _T_21898 = bht_rd_addr_f == 8'hf5; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_245; // @[Reg.scala 27:20]
  wire [1:0] _T_22165 = _T_21898 ? bht_bank_rd_data_out_1_245 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22420 = _T_22419 | _T_22165; // @[Mux.scala 27:72]
  wire  _T_21900 = bht_rd_addr_f == 8'hf6; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_246; // @[Reg.scala 27:20]
  wire [1:0] _T_22166 = _T_21900 ? bht_bank_rd_data_out_1_246 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22421 = _T_22420 | _T_22166; // @[Mux.scala 27:72]
  wire  _T_21902 = bht_rd_addr_f == 8'hf7; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_247; // @[Reg.scala 27:20]
  wire [1:0] _T_22167 = _T_21902 ? bht_bank_rd_data_out_1_247 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22422 = _T_22421 | _T_22167; // @[Mux.scala 27:72]
  wire  _T_21904 = bht_rd_addr_f == 8'hf8; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_248; // @[Reg.scala 27:20]
  wire [1:0] _T_22168 = _T_21904 ? bht_bank_rd_data_out_1_248 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22423 = _T_22422 | _T_22168; // @[Mux.scala 27:72]
  wire  _T_21906 = bht_rd_addr_f == 8'hf9; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_249; // @[Reg.scala 27:20]
  wire [1:0] _T_22169 = _T_21906 ? bht_bank_rd_data_out_1_249 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22424 = _T_22423 | _T_22169; // @[Mux.scala 27:72]
  wire  _T_21908 = bht_rd_addr_f == 8'hfa; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_250; // @[Reg.scala 27:20]
  wire [1:0] _T_22170 = _T_21908 ? bht_bank_rd_data_out_1_250 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22425 = _T_22424 | _T_22170; // @[Mux.scala 27:72]
  wire  _T_21910 = bht_rd_addr_f == 8'hfb; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_251; // @[Reg.scala 27:20]
  wire [1:0] _T_22171 = _T_21910 ? bht_bank_rd_data_out_1_251 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22426 = _T_22425 | _T_22171; // @[Mux.scala 27:72]
  wire  _T_21912 = bht_rd_addr_f == 8'hfc; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_252; // @[Reg.scala 27:20]
  wire [1:0] _T_22172 = _T_21912 ? bht_bank_rd_data_out_1_252 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22427 = _T_22426 | _T_22172; // @[Mux.scala 27:72]
  wire  _T_21914 = bht_rd_addr_f == 8'hfd; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_253; // @[Reg.scala 27:20]
  wire [1:0] _T_22173 = _T_21914 ? bht_bank_rd_data_out_1_253 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22428 = _T_22427 | _T_22173; // @[Mux.scala 27:72]
  wire  _T_21916 = bht_rd_addr_f == 8'hfe; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_254; // @[Reg.scala 27:20]
  wire [1:0] _T_22174 = _T_21916 ? bht_bank_rd_data_out_1_254 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22429 = _T_22428 | _T_22174; // @[Mux.scala 27:72]
  wire  _T_21918 = bht_rd_addr_f == 8'hff; // @[ifu_bp_ctl.scala 455:79]
  reg [1:0] bht_bank_rd_data_out_1_255; // @[Reg.scala 27:20]
  wire [1:0] _T_22175 = _T_21918 ? bht_bank_rd_data_out_1_255 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] bht_bank1_rd_data_f = _T_22429 | _T_22175; // @[Mux.scala 27:72]
  wire [1:0] _T_260 = _T_144 ? bht_bank1_rd_data_f : 2'h0; // @[Mux.scala 27:72]
  wire [9:0] _T_573 = {btb_rd_addr_p1_f,2'h0}; // @[Cat.scala 29:58]
  wire [7:0] bht_rd_addr_hashed_p1_f = _T_573[9:2] ^ fghr; // @[lib.scala 56:35]
  wire  _T_22432 = bht_rd_addr_hashed_p1_f == 8'h0; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_0; // @[Reg.scala 27:20]
  wire [1:0] _T_22944 = _T_22432 ? bht_bank_rd_data_out_0_0 : 2'h0; // @[Mux.scala 27:72]
  wire  _T_22434 = bht_rd_addr_hashed_p1_f == 8'h1; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_1; // @[Reg.scala 27:20]
  wire [1:0] _T_22945 = _T_22434 ? bht_bank_rd_data_out_0_1 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23200 = _T_22944 | _T_22945; // @[Mux.scala 27:72]
  wire  _T_22436 = bht_rd_addr_hashed_p1_f == 8'h2; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_2; // @[Reg.scala 27:20]
  wire [1:0] _T_22946 = _T_22436 ? bht_bank_rd_data_out_0_2 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23201 = _T_23200 | _T_22946; // @[Mux.scala 27:72]
  wire  _T_22438 = bht_rd_addr_hashed_p1_f == 8'h3; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_3; // @[Reg.scala 27:20]
  wire [1:0] _T_22947 = _T_22438 ? bht_bank_rd_data_out_0_3 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23202 = _T_23201 | _T_22947; // @[Mux.scala 27:72]
  wire  _T_22440 = bht_rd_addr_hashed_p1_f == 8'h4; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_4; // @[Reg.scala 27:20]
  wire [1:0] _T_22948 = _T_22440 ? bht_bank_rd_data_out_0_4 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23203 = _T_23202 | _T_22948; // @[Mux.scala 27:72]
  wire  _T_22442 = bht_rd_addr_hashed_p1_f == 8'h5; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_5; // @[Reg.scala 27:20]
  wire [1:0] _T_22949 = _T_22442 ? bht_bank_rd_data_out_0_5 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23204 = _T_23203 | _T_22949; // @[Mux.scala 27:72]
  wire  _T_22444 = bht_rd_addr_hashed_p1_f == 8'h6; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_6; // @[Reg.scala 27:20]
  wire [1:0] _T_22950 = _T_22444 ? bht_bank_rd_data_out_0_6 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23205 = _T_23204 | _T_22950; // @[Mux.scala 27:72]
  wire  _T_22446 = bht_rd_addr_hashed_p1_f == 8'h7; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_7; // @[Reg.scala 27:20]
  wire [1:0] _T_22951 = _T_22446 ? bht_bank_rd_data_out_0_7 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23206 = _T_23205 | _T_22951; // @[Mux.scala 27:72]
  wire  _T_22448 = bht_rd_addr_hashed_p1_f == 8'h8; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_8; // @[Reg.scala 27:20]
  wire [1:0] _T_22952 = _T_22448 ? bht_bank_rd_data_out_0_8 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23207 = _T_23206 | _T_22952; // @[Mux.scala 27:72]
  wire  _T_22450 = bht_rd_addr_hashed_p1_f == 8'h9; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_9; // @[Reg.scala 27:20]
  wire [1:0] _T_22953 = _T_22450 ? bht_bank_rd_data_out_0_9 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23208 = _T_23207 | _T_22953; // @[Mux.scala 27:72]
  wire  _T_22452 = bht_rd_addr_hashed_p1_f == 8'ha; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_10; // @[Reg.scala 27:20]
  wire [1:0] _T_22954 = _T_22452 ? bht_bank_rd_data_out_0_10 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23209 = _T_23208 | _T_22954; // @[Mux.scala 27:72]
  wire  _T_22454 = bht_rd_addr_hashed_p1_f == 8'hb; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_11; // @[Reg.scala 27:20]
  wire [1:0] _T_22955 = _T_22454 ? bht_bank_rd_data_out_0_11 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23210 = _T_23209 | _T_22955; // @[Mux.scala 27:72]
  wire  _T_22456 = bht_rd_addr_hashed_p1_f == 8'hc; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_12; // @[Reg.scala 27:20]
  wire [1:0] _T_22956 = _T_22456 ? bht_bank_rd_data_out_0_12 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23211 = _T_23210 | _T_22956; // @[Mux.scala 27:72]
  wire  _T_22458 = bht_rd_addr_hashed_p1_f == 8'hd; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_13; // @[Reg.scala 27:20]
  wire [1:0] _T_22957 = _T_22458 ? bht_bank_rd_data_out_0_13 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23212 = _T_23211 | _T_22957; // @[Mux.scala 27:72]
  wire  _T_22460 = bht_rd_addr_hashed_p1_f == 8'he; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_14; // @[Reg.scala 27:20]
  wire [1:0] _T_22958 = _T_22460 ? bht_bank_rd_data_out_0_14 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23213 = _T_23212 | _T_22958; // @[Mux.scala 27:72]
  wire  _T_22462 = bht_rd_addr_hashed_p1_f == 8'hf; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_15; // @[Reg.scala 27:20]
  wire [1:0] _T_22959 = _T_22462 ? bht_bank_rd_data_out_0_15 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23214 = _T_23213 | _T_22959; // @[Mux.scala 27:72]
  wire  _T_22464 = bht_rd_addr_hashed_p1_f == 8'h10; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_16; // @[Reg.scala 27:20]
  wire [1:0] _T_22960 = _T_22464 ? bht_bank_rd_data_out_0_16 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23215 = _T_23214 | _T_22960; // @[Mux.scala 27:72]
  wire  _T_22466 = bht_rd_addr_hashed_p1_f == 8'h11; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_17; // @[Reg.scala 27:20]
  wire [1:0] _T_22961 = _T_22466 ? bht_bank_rd_data_out_0_17 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23216 = _T_23215 | _T_22961; // @[Mux.scala 27:72]
  wire  _T_22468 = bht_rd_addr_hashed_p1_f == 8'h12; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_18; // @[Reg.scala 27:20]
  wire [1:0] _T_22962 = _T_22468 ? bht_bank_rd_data_out_0_18 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23217 = _T_23216 | _T_22962; // @[Mux.scala 27:72]
  wire  _T_22470 = bht_rd_addr_hashed_p1_f == 8'h13; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_19; // @[Reg.scala 27:20]
  wire [1:0] _T_22963 = _T_22470 ? bht_bank_rd_data_out_0_19 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23218 = _T_23217 | _T_22963; // @[Mux.scala 27:72]
  wire  _T_22472 = bht_rd_addr_hashed_p1_f == 8'h14; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_20; // @[Reg.scala 27:20]
  wire [1:0] _T_22964 = _T_22472 ? bht_bank_rd_data_out_0_20 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23219 = _T_23218 | _T_22964; // @[Mux.scala 27:72]
  wire  _T_22474 = bht_rd_addr_hashed_p1_f == 8'h15; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_21; // @[Reg.scala 27:20]
  wire [1:0] _T_22965 = _T_22474 ? bht_bank_rd_data_out_0_21 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23220 = _T_23219 | _T_22965; // @[Mux.scala 27:72]
  wire  _T_22476 = bht_rd_addr_hashed_p1_f == 8'h16; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_22; // @[Reg.scala 27:20]
  wire [1:0] _T_22966 = _T_22476 ? bht_bank_rd_data_out_0_22 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23221 = _T_23220 | _T_22966; // @[Mux.scala 27:72]
  wire  _T_22478 = bht_rd_addr_hashed_p1_f == 8'h17; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_23; // @[Reg.scala 27:20]
  wire [1:0] _T_22967 = _T_22478 ? bht_bank_rd_data_out_0_23 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23222 = _T_23221 | _T_22967; // @[Mux.scala 27:72]
  wire  _T_22480 = bht_rd_addr_hashed_p1_f == 8'h18; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_24; // @[Reg.scala 27:20]
  wire [1:0] _T_22968 = _T_22480 ? bht_bank_rd_data_out_0_24 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23223 = _T_23222 | _T_22968; // @[Mux.scala 27:72]
  wire  _T_22482 = bht_rd_addr_hashed_p1_f == 8'h19; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_25; // @[Reg.scala 27:20]
  wire [1:0] _T_22969 = _T_22482 ? bht_bank_rd_data_out_0_25 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23224 = _T_23223 | _T_22969; // @[Mux.scala 27:72]
  wire  _T_22484 = bht_rd_addr_hashed_p1_f == 8'h1a; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_26; // @[Reg.scala 27:20]
  wire [1:0] _T_22970 = _T_22484 ? bht_bank_rd_data_out_0_26 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23225 = _T_23224 | _T_22970; // @[Mux.scala 27:72]
  wire  _T_22486 = bht_rd_addr_hashed_p1_f == 8'h1b; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_27; // @[Reg.scala 27:20]
  wire [1:0] _T_22971 = _T_22486 ? bht_bank_rd_data_out_0_27 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23226 = _T_23225 | _T_22971; // @[Mux.scala 27:72]
  wire  _T_22488 = bht_rd_addr_hashed_p1_f == 8'h1c; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_28; // @[Reg.scala 27:20]
  wire [1:0] _T_22972 = _T_22488 ? bht_bank_rd_data_out_0_28 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23227 = _T_23226 | _T_22972; // @[Mux.scala 27:72]
  wire  _T_22490 = bht_rd_addr_hashed_p1_f == 8'h1d; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_29; // @[Reg.scala 27:20]
  wire [1:0] _T_22973 = _T_22490 ? bht_bank_rd_data_out_0_29 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23228 = _T_23227 | _T_22973; // @[Mux.scala 27:72]
  wire  _T_22492 = bht_rd_addr_hashed_p1_f == 8'h1e; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_30; // @[Reg.scala 27:20]
  wire [1:0] _T_22974 = _T_22492 ? bht_bank_rd_data_out_0_30 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23229 = _T_23228 | _T_22974; // @[Mux.scala 27:72]
  wire  _T_22494 = bht_rd_addr_hashed_p1_f == 8'h1f; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_31; // @[Reg.scala 27:20]
  wire [1:0] _T_22975 = _T_22494 ? bht_bank_rd_data_out_0_31 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23230 = _T_23229 | _T_22975; // @[Mux.scala 27:72]
  wire  _T_22496 = bht_rd_addr_hashed_p1_f == 8'h20; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_32; // @[Reg.scala 27:20]
  wire [1:0] _T_22976 = _T_22496 ? bht_bank_rd_data_out_0_32 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23231 = _T_23230 | _T_22976; // @[Mux.scala 27:72]
  wire  _T_22498 = bht_rd_addr_hashed_p1_f == 8'h21; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_33; // @[Reg.scala 27:20]
  wire [1:0] _T_22977 = _T_22498 ? bht_bank_rd_data_out_0_33 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23232 = _T_23231 | _T_22977; // @[Mux.scala 27:72]
  wire  _T_22500 = bht_rd_addr_hashed_p1_f == 8'h22; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_34; // @[Reg.scala 27:20]
  wire [1:0] _T_22978 = _T_22500 ? bht_bank_rd_data_out_0_34 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23233 = _T_23232 | _T_22978; // @[Mux.scala 27:72]
  wire  _T_22502 = bht_rd_addr_hashed_p1_f == 8'h23; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_35; // @[Reg.scala 27:20]
  wire [1:0] _T_22979 = _T_22502 ? bht_bank_rd_data_out_0_35 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23234 = _T_23233 | _T_22979; // @[Mux.scala 27:72]
  wire  _T_22504 = bht_rd_addr_hashed_p1_f == 8'h24; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_36; // @[Reg.scala 27:20]
  wire [1:0] _T_22980 = _T_22504 ? bht_bank_rd_data_out_0_36 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23235 = _T_23234 | _T_22980; // @[Mux.scala 27:72]
  wire  _T_22506 = bht_rd_addr_hashed_p1_f == 8'h25; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_37; // @[Reg.scala 27:20]
  wire [1:0] _T_22981 = _T_22506 ? bht_bank_rd_data_out_0_37 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23236 = _T_23235 | _T_22981; // @[Mux.scala 27:72]
  wire  _T_22508 = bht_rd_addr_hashed_p1_f == 8'h26; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_38; // @[Reg.scala 27:20]
  wire [1:0] _T_22982 = _T_22508 ? bht_bank_rd_data_out_0_38 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23237 = _T_23236 | _T_22982; // @[Mux.scala 27:72]
  wire  _T_22510 = bht_rd_addr_hashed_p1_f == 8'h27; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_39; // @[Reg.scala 27:20]
  wire [1:0] _T_22983 = _T_22510 ? bht_bank_rd_data_out_0_39 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23238 = _T_23237 | _T_22983; // @[Mux.scala 27:72]
  wire  _T_22512 = bht_rd_addr_hashed_p1_f == 8'h28; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_40; // @[Reg.scala 27:20]
  wire [1:0] _T_22984 = _T_22512 ? bht_bank_rd_data_out_0_40 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23239 = _T_23238 | _T_22984; // @[Mux.scala 27:72]
  wire  _T_22514 = bht_rd_addr_hashed_p1_f == 8'h29; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_41; // @[Reg.scala 27:20]
  wire [1:0] _T_22985 = _T_22514 ? bht_bank_rd_data_out_0_41 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23240 = _T_23239 | _T_22985; // @[Mux.scala 27:72]
  wire  _T_22516 = bht_rd_addr_hashed_p1_f == 8'h2a; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_42; // @[Reg.scala 27:20]
  wire [1:0] _T_22986 = _T_22516 ? bht_bank_rd_data_out_0_42 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23241 = _T_23240 | _T_22986; // @[Mux.scala 27:72]
  wire  _T_22518 = bht_rd_addr_hashed_p1_f == 8'h2b; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_43; // @[Reg.scala 27:20]
  wire [1:0] _T_22987 = _T_22518 ? bht_bank_rd_data_out_0_43 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23242 = _T_23241 | _T_22987; // @[Mux.scala 27:72]
  wire  _T_22520 = bht_rd_addr_hashed_p1_f == 8'h2c; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_44; // @[Reg.scala 27:20]
  wire [1:0] _T_22988 = _T_22520 ? bht_bank_rd_data_out_0_44 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23243 = _T_23242 | _T_22988; // @[Mux.scala 27:72]
  wire  _T_22522 = bht_rd_addr_hashed_p1_f == 8'h2d; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_45; // @[Reg.scala 27:20]
  wire [1:0] _T_22989 = _T_22522 ? bht_bank_rd_data_out_0_45 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23244 = _T_23243 | _T_22989; // @[Mux.scala 27:72]
  wire  _T_22524 = bht_rd_addr_hashed_p1_f == 8'h2e; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_46; // @[Reg.scala 27:20]
  wire [1:0] _T_22990 = _T_22524 ? bht_bank_rd_data_out_0_46 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23245 = _T_23244 | _T_22990; // @[Mux.scala 27:72]
  wire  _T_22526 = bht_rd_addr_hashed_p1_f == 8'h2f; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_47; // @[Reg.scala 27:20]
  wire [1:0] _T_22991 = _T_22526 ? bht_bank_rd_data_out_0_47 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23246 = _T_23245 | _T_22991; // @[Mux.scala 27:72]
  wire  _T_22528 = bht_rd_addr_hashed_p1_f == 8'h30; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_48; // @[Reg.scala 27:20]
  wire [1:0] _T_22992 = _T_22528 ? bht_bank_rd_data_out_0_48 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23247 = _T_23246 | _T_22992; // @[Mux.scala 27:72]
  wire  _T_22530 = bht_rd_addr_hashed_p1_f == 8'h31; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_49; // @[Reg.scala 27:20]
  wire [1:0] _T_22993 = _T_22530 ? bht_bank_rd_data_out_0_49 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23248 = _T_23247 | _T_22993; // @[Mux.scala 27:72]
  wire  _T_22532 = bht_rd_addr_hashed_p1_f == 8'h32; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_50; // @[Reg.scala 27:20]
  wire [1:0] _T_22994 = _T_22532 ? bht_bank_rd_data_out_0_50 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23249 = _T_23248 | _T_22994; // @[Mux.scala 27:72]
  wire  _T_22534 = bht_rd_addr_hashed_p1_f == 8'h33; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_51; // @[Reg.scala 27:20]
  wire [1:0] _T_22995 = _T_22534 ? bht_bank_rd_data_out_0_51 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23250 = _T_23249 | _T_22995; // @[Mux.scala 27:72]
  wire  _T_22536 = bht_rd_addr_hashed_p1_f == 8'h34; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_52; // @[Reg.scala 27:20]
  wire [1:0] _T_22996 = _T_22536 ? bht_bank_rd_data_out_0_52 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23251 = _T_23250 | _T_22996; // @[Mux.scala 27:72]
  wire  _T_22538 = bht_rd_addr_hashed_p1_f == 8'h35; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_53; // @[Reg.scala 27:20]
  wire [1:0] _T_22997 = _T_22538 ? bht_bank_rd_data_out_0_53 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23252 = _T_23251 | _T_22997; // @[Mux.scala 27:72]
  wire  _T_22540 = bht_rd_addr_hashed_p1_f == 8'h36; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_54; // @[Reg.scala 27:20]
  wire [1:0] _T_22998 = _T_22540 ? bht_bank_rd_data_out_0_54 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23253 = _T_23252 | _T_22998; // @[Mux.scala 27:72]
  wire  _T_22542 = bht_rd_addr_hashed_p1_f == 8'h37; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_55; // @[Reg.scala 27:20]
  wire [1:0] _T_22999 = _T_22542 ? bht_bank_rd_data_out_0_55 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23254 = _T_23253 | _T_22999; // @[Mux.scala 27:72]
  wire  _T_22544 = bht_rd_addr_hashed_p1_f == 8'h38; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_56; // @[Reg.scala 27:20]
  wire [1:0] _T_23000 = _T_22544 ? bht_bank_rd_data_out_0_56 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23255 = _T_23254 | _T_23000; // @[Mux.scala 27:72]
  wire  _T_22546 = bht_rd_addr_hashed_p1_f == 8'h39; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_57; // @[Reg.scala 27:20]
  wire [1:0] _T_23001 = _T_22546 ? bht_bank_rd_data_out_0_57 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23256 = _T_23255 | _T_23001; // @[Mux.scala 27:72]
  wire  _T_22548 = bht_rd_addr_hashed_p1_f == 8'h3a; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_58; // @[Reg.scala 27:20]
  wire [1:0] _T_23002 = _T_22548 ? bht_bank_rd_data_out_0_58 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23257 = _T_23256 | _T_23002; // @[Mux.scala 27:72]
  wire  _T_22550 = bht_rd_addr_hashed_p1_f == 8'h3b; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_59; // @[Reg.scala 27:20]
  wire [1:0] _T_23003 = _T_22550 ? bht_bank_rd_data_out_0_59 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23258 = _T_23257 | _T_23003; // @[Mux.scala 27:72]
  wire  _T_22552 = bht_rd_addr_hashed_p1_f == 8'h3c; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_60; // @[Reg.scala 27:20]
  wire [1:0] _T_23004 = _T_22552 ? bht_bank_rd_data_out_0_60 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23259 = _T_23258 | _T_23004; // @[Mux.scala 27:72]
  wire  _T_22554 = bht_rd_addr_hashed_p1_f == 8'h3d; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_61; // @[Reg.scala 27:20]
  wire [1:0] _T_23005 = _T_22554 ? bht_bank_rd_data_out_0_61 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23260 = _T_23259 | _T_23005; // @[Mux.scala 27:72]
  wire  _T_22556 = bht_rd_addr_hashed_p1_f == 8'h3e; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_62; // @[Reg.scala 27:20]
  wire [1:0] _T_23006 = _T_22556 ? bht_bank_rd_data_out_0_62 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23261 = _T_23260 | _T_23006; // @[Mux.scala 27:72]
  wire  _T_22558 = bht_rd_addr_hashed_p1_f == 8'h3f; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_63; // @[Reg.scala 27:20]
  wire [1:0] _T_23007 = _T_22558 ? bht_bank_rd_data_out_0_63 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23262 = _T_23261 | _T_23007; // @[Mux.scala 27:72]
  wire  _T_22560 = bht_rd_addr_hashed_p1_f == 8'h40; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_64; // @[Reg.scala 27:20]
  wire [1:0] _T_23008 = _T_22560 ? bht_bank_rd_data_out_0_64 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23263 = _T_23262 | _T_23008; // @[Mux.scala 27:72]
  wire  _T_22562 = bht_rd_addr_hashed_p1_f == 8'h41; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_65; // @[Reg.scala 27:20]
  wire [1:0] _T_23009 = _T_22562 ? bht_bank_rd_data_out_0_65 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23264 = _T_23263 | _T_23009; // @[Mux.scala 27:72]
  wire  _T_22564 = bht_rd_addr_hashed_p1_f == 8'h42; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_66; // @[Reg.scala 27:20]
  wire [1:0] _T_23010 = _T_22564 ? bht_bank_rd_data_out_0_66 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23265 = _T_23264 | _T_23010; // @[Mux.scala 27:72]
  wire  _T_22566 = bht_rd_addr_hashed_p1_f == 8'h43; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_67; // @[Reg.scala 27:20]
  wire [1:0] _T_23011 = _T_22566 ? bht_bank_rd_data_out_0_67 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23266 = _T_23265 | _T_23011; // @[Mux.scala 27:72]
  wire  _T_22568 = bht_rd_addr_hashed_p1_f == 8'h44; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_68; // @[Reg.scala 27:20]
  wire [1:0] _T_23012 = _T_22568 ? bht_bank_rd_data_out_0_68 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23267 = _T_23266 | _T_23012; // @[Mux.scala 27:72]
  wire  _T_22570 = bht_rd_addr_hashed_p1_f == 8'h45; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_69; // @[Reg.scala 27:20]
  wire [1:0] _T_23013 = _T_22570 ? bht_bank_rd_data_out_0_69 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23268 = _T_23267 | _T_23013; // @[Mux.scala 27:72]
  wire  _T_22572 = bht_rd_addr_hashed_p1_f == 8'h46; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_70; // @[Reg.scala 27:20]
  wire [1:0] _T_23014 = _T_22572 ? bht_bank_rd_data_out_0_70 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23269 = _T_23268 | _T_23014; // @[Mux.scala 27:72]
  wire  _T_22574 = bht_rd_addr_hashed_p1_f == 8'h47; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_71; // @[Reg.scala 27:20]
  wire [1:0] _T_23015 = _T_22574 ? bht_bank_rd_data_out_0_71 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23270 = _T_23269 | _T_23015; // @[Mux.scala 27:72]
  wire  _T_22576 = bht_rd_addr_hashed_p1_f == 8'h48; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_72; // @[Reg.scala 27:20]
  wire [1:0] _T_23016 = _T_22576 ? bht_bank_rd_data_out_0_72 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23271 = _T_23270 | _T_23016; // @[Mux.scala 27:72]
  wire  _T_22578 = bht_rd_addr_hashed_p1_f == 8'h49; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_73; // @[Reg.scala 27:20]
  wire [1:0] _T_23017 = _T_22578 ? bht_bank_rd_data_out_0_73 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23272 = _T_23271 | _T_23017; // @[Mux.scala 27:72]
  wire  _T_22580 = bht_rd_addr_hashed_p1_f == 8'h4a; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_74; // @[Reg.scala 27:20]
  wire [1:0] _T_23018 = _T_22580 ? bht_bank_rd_data_out_0_74 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23273 = _T_23272 | _T_23018; // @[Mux.scala 27:72]
  wire  _T_22582 = bht_rd_addr_hashed_p1_f == 8'h4b; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_75; // @[Reg.scala 27:20]
  wire [1:0] _T_23019 = _T_22582 ? bht_bank_rd_data_out_0_75 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23274 = _T_23273 | _T_23019; // @[Mux.scala 27:72]
  wire  _T_22584 = bht_rd_addr_hashed_p1_f == 8'h4c; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_76; // @[Reg.scala 27:20]
  wire [1:0] _T_23020 = _T_22584 ? bht_bank_rd_data_out_0_76 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23275 = _T_23274 | _T_23020; // @[Mux.scala 27:72]
  wire  _T_22586 = bht_rd_addr_hashed_p1_f == 8'h4d; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_77; // @[Reg.scala 27:20]
  wire [1:0] _T_23021 = _T_22586 ? bht_bank_rd_data_out_0_77 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23276 = _T_23275 | _T_23021; // @[Mux.scala 27:72]
  wire  _T_22588 = bht_rd_addr_hashed_p1_f == 8'h4e; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_78; // @[Reg.scala 27:20]
  wire [1:0] _T_23022 = _T_22588 ? bht_bank_rd_data_out_0_78 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23277 = _T_23276 | _T_23022; // @[Mux.scala 27:72]
  wire  _T_22590 = bht_rd_addr_hashed_p1_f == 8'h4f; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_79; // @[Reg.scala 27:20]
  wire [1:0] _T_23023 = _T_22590 ? bht_bank_rd_data_out_0_79 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23278 = _T_23277 | _T_23023; // @[Mux.scala 27:72]
  wire  _T_22592 = bht_rd_addr_hashed_p1_f == 8'h50; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_80; // @[Reg.scala 27:20]
  wire [1:0] _T_23024 = _T_22592 ? bht_bank_rd_data_out_0_80 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23279 = _T_23278 | _T_23024; // @[Mux.scala 27:72]
  wire  _T_22594 = bht_rd_addr_hashed_p1_f == 8'h51; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_81; // @[Reg.scala 27:20]
  wire [1:0] _T_23025 = _T_22594 ? bht_bank_rd_data_out_0_81 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23280 = _T_23279 | _T_23025; // @[Mux.scala 27:72]
  wire  _T_22596 = bht_rd_addr_hashed_p1_f == 8'h52; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_82; // @[Reg.scala 27:20]
  wire [1:0] _T_23026 = _T_22596 ? bht_bank_rd_data_out_0_82 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23281 = _T_23280 | _T_23026; // @[Mux.scala 27:72]
  wire  _T_22598 = bht_rd_addr_hashed_p1_f == 8'h53; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_83; // @[Reg.scala 27:20]
  wire [1:0] _T_23027 = _T_22598 ? bht_bank_rd_data_out_0_83 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23282 = _T_23281 | _T_23027; // @[Mux.scala 27:72]
  wire  _T_22600 = bht_rd_addr_hashed_p1_f == 8'h54; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_84; // @[Reg.scala 27:20]
  wire [1:0] _T_23028 = _T_22600 ? bht_bank_rd_data_out_0_84 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23283 = _T_23282 | _T_23028; // @[Mux.scala 27:72]
  wire  _T_22602 = bht_rd_addr_hashed_p1_f == 8'h55; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_85; // @[Reg.scala 27:20]
  wire [1:0] _T_23029 = _T_22602 ? bht_bank_rd_data_out_0_85 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23284 = _T_23283 | _T_23029; // @[Mux.scala 27:72]
  wire  _T_22604 = bht_rd_addr_hashed_p1_f == 8'h56; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_86; // @[Reg.scala 27:20]
  wire [1:0] _T_23030 = _T_22604 ? bht_bank_rd_data_out_0_86 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23285 = _T_23284 | _T_23030; // @[Mux.scala 27:72]
  wire  _T_22606 = bht_rd_addr_hashed_p1_f == 8'h57; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_87; // @[Reg.scala 27:20]
  wire [1:0] _T_23031 = _T_22606 ? bht_bank_rd_data_out_0_87 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23286 = _T_23285 | _T_23031; // @[Mux.scala 27:72]
  wire  _T_22608 = bht_rd_addr_hashed_p1_f == 8'h58; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_88; // @[Reg.scala 27:20]
  wire [1:0] _T_23032 = _T_22608 ? bht_bank_rd_data_out_0_88 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23287 = _T_23286 | _T_23032; // @[Mux.scala 27:72]
  wire  _T_22610 = bht_rd_addr_hashed_p1_f == 8'h59; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_89; // @[Reg.scala 27:20]
  wire [1:0] _T_23033 = _T_22610 ? bht_bank_rd_data_out_0_89 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23288 = _T_23287 | _T_23033; // @[Mux.scala 27:72]
  wire  _T_22612 = bht_rd_addr_hashed_p1_f == 8'h5a; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_90; // @[Reg.scala 27:20]
  wire [1:0] _T_23034 = _T_22612 ? bht_bank_rd_data_out_0_90 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23289 = _T_23288 | _T_23034; // @[Mux.scala 27:72]
  wire  _T_22614 = bht_rd_addr_hashed_p1_f == 8'h5b; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_91; // @[Reg.scala 27:20]
  wire [1:0] _T_23035 = _T_22614 ? bht_bank_rd_data_out_0_91 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23290 = _T_23289 | _T_23035; // @[Mux.scala 27:72]
  wire  _T_22616 = bht_rd_addr_hashed_p1_f == 8'h5c; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_92; // @[Reg.scala 27:20]
  wire [1:0] _T_23036 = _T_22616 ? bht_bank_rd_data_out_0_92 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23291 = _T_23290 | _T_23036; // @[Mux.scala 27:72]
  wire  _T_22618 = bht_rd_addr_hashed_p1_f == 8'h5d; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_93; // @[Reg.scala 27:20]
  wire [1:0] _T_23037 = _T_22618 ? bht_bank_rd_data_out_0_93 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23292 = _T_23291 | _T_23037; // @[Mux.scala 27:72]
  wire  _T_22620 = bht_rd_addr_hashed_p1_f == 8'h5e; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_94; // @[Reg.scala 27:20]
  wire [1:0] _T_23038 = _T_22620 ? bht_bank_rd_data_out_0_94 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23293 = _T_23292 | _T_23038; // @[Mux.scala 27:72]
  wire  _T_22622 = bht_rd_addr_hashed_p1_f == 8'h5f; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_95; // @[Reg.scala 27:20]
  wire [1:0] _T_23039 = _T_22622 ? bht_bank_rd_data_out_0_95 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23294 = _T_23293 | _T_23039; // @[Mux.scala 27:72]
  wire  _T_22624 = bht_rd_addr_hashed_p1_f == 8'h60; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_96; // @[Reg.scala 27:20]
  wire [1:0] _T_23040 = _T_22624 ? bht_bank_rd_data_out_0_96 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23295 = _T_23294 | _T_23040; // @[Mux.scala 27:72]
  wire  _T_22626 = bht_rd_addr_hashed_p1_f == 8'h61; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_97; // @[Reg.scala 27:20]
  wire [1:0] _T_23041 = _T_22626 ? bht_bank_rd_data_out_0_97 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23296 = _T_23295 | _T_23041; // @[Mux.scala 27:72]
  wire  _T_22628 = bht_rd_addr_hashed_p1_f == 8'h62; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_98; // @[Reg.scala 27:20]
  wire [1:0] _T_23042 = _T_22628 ? bht_bank_rd_data_out_0_98 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23297 = _T_23296 | _T_23042; // @[Mux.scala 27:72]
  wire  _T_22630 = bht_rd_addr_hashed_p1_f == 8'h63; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_99; // @[Reg.scala 27:20]
  wire [1:0] _T_23043 = _T_22630 ? bht_bank_rd_data_out_0_99 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23298 = _T_23297 | _T_23043; // @[Mux.scala 27:72]
  wire  _T_22632 = bht_rd_addr_hashed_p1_f == 8'h64; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_100; // @[Reg.scala 27:20]
  wire [1:0] _T_23044 = _T_22632 ? bht_bank_rd_data_out_0_100 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23299 = _T_23298 | _T_23044; // @[Mux.scala 27:72]
  wire  _T_22634 = bht_rd_addr_hashed_p1_f == 8'h65; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_101; // @[Reg.scala 27:20]
  wire [1:0] _T_23045 = _T_22634 ? bht_bank_rd_data_out_0_101 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23300 = _T_23299 | _T_23045; // @[Mux.scala 27:72]
  wire  _T_22636 = bht_rd_addr_hashed_p1_f == 8'h66; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_102; // @[Reg.scala 27:20]
  wire [1:0] _T_23046 = _T_22636 ? bht_bank_rd_data_out_0_102 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23301 = _T_23300 | _T_23046; // @[Mux.scala 27:72]
  wire  _T_22638 = bht_rd_addr_hashed_p1_f == 8'h67; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_103; // @[Reg.scala 27:20]
  wire [1:0] _T_23047 = _T_22638 ? bht_bank_rd_data_out_0_103 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23302 = _T_23301 | _T_23047; // @[Mux.scala 27:72]
  wire  _T_22640 = bht_rd_addr_hashed_p1_f == 8'h68; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_104; // @[Reg.scala 27:20]
  wire [1:0] _T_23048 = _T_22640 ? bht_bank_rd_data_out_0_104 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23303 = _T_23302 | _T_23048; // @[Mux.scala 27:72]
  wire  _T_22642 = bht_rd_addr_hashed_p1_f == 8'h69; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_105; // @[Reg.scala 27:20]
  wire [1:0] _T_23049 = _T_22642 ? bht_bank_rd_data_out_0_105 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23304 = _T_23303 | _T_23049; // @[Mux.scala 27:72]
  wire  _T_22644 = bht_rd_addr_hashed_p1_f == 8'h6a; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_106; // @[Reg.scala 27:20]
  wire [1:0] _T_23050 = _T_22644 ? bht_bank_rd_data_out_0_106 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23305 = _T_23304 | _T_23050; // @[Mux.scala 27:72]
  wire  _T_22646 = bht_rd_addr_hashed_p1_f == 8'h6b; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_107; // @[Reg.scala 27:20]
  wire [1:0] _T_23051 = _T_22646 ? bht_bank_rd_data_out_0_107 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23306 = _T_23305 | _T_23051; // @[Mux.scala 27:72]
  wire  _T_22648 = bht_rd_addr_hashed_p1_f == 8'h6c; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_108; // @[Reg.scala 27:20]
  wire [1:0] _T_23052 = _T_22648 ? bht_bank_rd_data_out_0_108 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23307 = _T_23306 | _T_23052; // @[Mux.scala 27:72]
  wire  _T_22650 = bht_rd_addr_hashed_p1_f == 8'h6d; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_109; // @[Reg.scala 27:20]
  wire [1:0] _T_23053 = _T_22650 ? bht_bank_rd_data_out_0_109 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23308 = _T_23307 | _T_23053; // @[Mux.scala 27:72]
  wire  _T_22652 = bht_rd_addr_hashed_p1_f == 8'h6e; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_110; // @[Reg.scala 27:20]
  wire [1:0] _T_23054 = _T_22652 ? bht_bank_rd_data_out_0_110 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23309 = _T_23308 | _T_23054; // @[Mux.scala 27:72]
  wire  _T_22654 = bht_rd_addr_hashed_p1_f == 8'h6f; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_111; // @[Reg.scala 27:20]
  wire [1:0] _T_23055 = _T_22654 ? bht_bank_rd_data_out_0_111 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23310 = _T_23309 | _T_23055; // @[Mux.scala 27:72]
  wire  _T_22656 = bht_rd_addr_hashed_p1_f == 8'h70; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_112; // @[Reg.scala 27:20]
  wire [1:0] _T_23056 = _T_22656 ? bht_bank_rd_data_out_0_112 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23311 = _T_23310 | _T_23056; // @[Mux.scala 27:72]
  wire  _T_22658 = bht_rd_addr_hashed_p1_f == 8'h71; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_113; // @[Reg.scala 27:20]
  wire [1:0] _T_23057 = _T_22658 ? bht_bank_rd_data_out_0_113 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23312 = _T_23311 | _T_23057; // @[Mux.scala 27:72]
  wire  _T_22660 = bht_rd_addr_hashed_p1_f == 8'h72; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_114; // @[Reg.scala 27:20]
  wire [1:0] _T_23058 = _T_22660 ? bht_bank_rd_data_out_0_114 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23313 = _T_23312 | _T_23058; // @[Mux.scala 27:72]
  wire  _T_22662 = bht_rd_addr_hashed_p1_f == 8'h73; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_115; // @[Reg.scala 27:20]
  wire [1:0] _T_23059 = _T_22662 ? bht_bank_rd_data_out_0_115 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23314 = _T_23313 | _T_23059; // @[Mux.scala 27:72]
  wire  _T_22664 = bht_rd_addr_hashed_p1_f == 8'h74; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_116; // @[Reg.scala 27:20]
  wire [1:0] _T_23060 = _T_22664 ? bht_bank_rd_data_out_0_116 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23315 = _T_23314 | _T_23060; // @[Mux.scala 27:72]
  wire  _T_22666 = bht_rd_addr_hashed_p1_f == 8'h75; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_117; // @[Reg.scala 27:20]
  wire [1:0] _T_23061 = _T_22666 ? bht_bank_rd_data_out_0_117 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23316 = _T_23315 | _T_23061; // @[Mux.scala 27:72]
  wire  _T_22668 = bht_rd_addr_hashed_p1_f == 8'h76; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_118; // @[Reg.scala 27:20]
  wire [1:0] _T_23062 = _T_22668 ? bht_bank_rd_data_out_0_118 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23317 = _T_23316 | _T_23062; // @[Mux.scala 27:72]
  wire  _T_22670 = bht_rd_addr_hashed_p1_f == 8'h77; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_119; // @[Reg.scala 27:20]
  wire [1:0] _T_23063 = _T_22670 ? bht_bank_rd_data_out_0_119 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23318 = _T_23317 | _T_23063; // @[Mux.scala 27:72]
  wire  _T_22672 = bht_rd_addr_hashed_p1_f == 8'h78; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_120; // @[Reg.scala 27:20]
  wire [1:0] _T_23064 = _T_22672 ? bht_bank_rd_data_out_0_120 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23319 = _T_23318 | _T_23064; // @[Mux.scala 27:72]
  wire  _T_22674 = bht_rd_addr_hashed_p1_f == 8'h79; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_121; // @[Reg.scala 27:20]
  wire [1:0] _T_23065 = _T_22674 ? bht_bank_rd_data_out_0_121 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23320 = _T_23319 | _T_23065; // @[Mux.scala 27:72]
  wire  _T_22676 = bht_rd_addr_hashed_p1_f == 8'h7a; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_122; // @[Reg.scala 27:20]
  wire [1:0] _T_23066 = _T_22676 ? bht_bank_rd_data_out_0_122 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23321 = _T_23320 | _T_23066; // @[Mux.scala 27:72]
  wire  _T_22678 = bht_rd_addr_hashed_p1_f == 8'h7b; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_123; // @[Reg.scala 27:20]
  wire [1:0] _T_23067 = _T_22678 ? bht_bank_rd_data_out_0_123 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23322 = _T_23321 | _T_23067; // @[Mux.scala 27:72]
  wire  _T_22680 = bht_rd_addr_hashed_p1_f == 8'h7c; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_124; // @[Reg.scala 27:20]
  wire [1:0] _T_23068 = _T_22680 ? bht_bank_rd_data_out_0_124 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23323 = _T_23322 | _T_23068; // @[Mux.scala 27:72]
  wire  _T_22682 = bht_rd_addr_hashed_p1_f == 8'h7d; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_125; // @[Reg.scala 27:20]
  wire [1:0] _T_23069 = _T_22682 ? bht_bank_rd_data_out_0_125 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23324 = _T_23323 | _T_23069; // @[Mux.scala 27:72]
  wire  _T_22684 = bht_rd_addr_hashed_p1_f == 8'h7e; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_126; // @[Reg.scala 27:20]
  wire [1:0] _T_23070 = _T_22684 ? bht_bank_rd_data_out_0_126 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23325 = _T_23324 | _T_23070; // @[Mux.scala 27:72]
  wire  _T_22686 = bht_rd_addr_hashed_p1_f == 8'h7f; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_127; // @[Reg.scala 27:20]
  wire [1:0] _T_23071 = _T_22686 ? bht_bank_rd_data_out_0_127 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23326 = _T_23325 | _T_23071; // @[Mux.scala 27:72]
  wire  _T_22688 = bht_rd_addr_hashed_p1_f == 8'h80; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_128; // @[Reg.scala 27:20]
  wire [1:0] _T_23072 = _T_22688 ? bht_bank_rd_data_out_0_128 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23327 = _T_23326 | _T_23072; // @[Mux.scala 27:72]
  wire  _T_22690 = bht_rd_addr_hashed_p1_f == 8'h81; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_129; // @[Reg.scala 27:20]
  wire [1:0] _T_23073 = _T_22690 ? bht_bank_rd_data_out_0_129 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23328 = _T_23327 | _T_23073; // @[Mux.scala 27:72]
  wire  _T_22692 = bht_rd_addr_hashed_p1_f == 8'h82; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_130; // @[Reg.scala 27:20]
  wire [1:0] _T_23074 = _T_22692 ? bht_bank_rd_data_out_0_130 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23329 = _T_23328 | _T_23074; // @[Mux.scala 27:72]
  wire  _T_22694 = bht_rd_addr_hashed_p1_f == 8'h83; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_131; // @[Reg.scala 27:20]
  wire [1:0] _T_23075 = _T_22694 ? bht_bank_rd_data_out_0_131 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23330 = _T_23329 | _T_23075; // @[Mux.scala 27:72]
  wire  _T_22696 = bht_rd_addr_hashed_p1_f == 8'h84; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_132; // @[Reg.scala 27:20]
  wire [1:0] _T_23076 = _T_22696 ? bht_bank_rd_data_out_0_132 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23331 = _T_23330 | _T_23076; // @[Mux.scala 27:72]
  wire  _T_22698 = bht_rd_addr_hashed_p1_f == 8'h85; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_133; // @[Reg.scala 27:20]
  wire [1:0] _T_23077 = _T_22698 ? bht_bank_rd_data_out_0_133 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23332 = _T_23331 | _T_23077; // @[Mux.scala 27:72]
  wire  _T_22700 = bht_rd_addr_hashed_p1_f == 8'h86; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_134; // @[Reg.scala 27:20]
  wire [1:0] _T_23078 = _T_22700 ? bht_bank_rd_data_out_0_134 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23333 = _T_23332 | _T_23078; // @[Mux.scala 27:72]
  wire  _T_22702 = bht_rd_addr_hashed_p1_f == 8'h87; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_135; // @[Reg.scala 27:20]
  wire [1:0] _T_23079 = _T_22702 ? bht_bank_rd_data_out_0_135 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23334 = _T_23333 | _T_23079; // @[Mux.scala 27:72]
  wire  _T_22704 = bht_rd_addr_hashed_p1_f == 8'h88; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_136; // @[Reg.scala 27:20]
  wire [1:0] _T_23080 = _T_22704 ? bht_bank_rd_data_out_0_136 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23335 = _T_23334 | _T_23080; // @[Mux.scala 27:72]
  wire  _T_22706 = bht_rd_addr_hashed_p1_f == 8'h89; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_137; // @[Reg.scala 27:20]
  wire [1:0] _T_23081 = _T_22706 ? bht_bank_rd_data_out_0_137 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23336 = _T_23335 | _T_23081; // @[Mux.scala 27:72]
  wire  _T_22708 = bht_rd_addr_hashed_p1_f == 8'h8a; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_138; // @[Reg.scala 27:20]
  wire [1:0] _T_23082 = _T_22708 ? bht_bank_rd_data_out_0_138 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23337 = _T_23336 | _T_23082; // @[Mux.scala 27:72]
  wire  _T_22710 = bht_rd_addr_hashed_p1_f == 8'h8b; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_139; // @[Reg.scala 27:20]
  wire [1:0] _T_23083 = _T_22710 ? bht_bank_rd_data_out_0_139 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23338 = _T_23337 | _T_23083; // @[Mux.scala 27:72]
  wire  _T_22712 = bht_rd_addr_hashed_p1_f == 8'h8c; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_140; // @[Reg.scala 27:20]
  wire [1:0] _T_23084 = _T_22712 ? bht_bank_rd_data_out_0_140 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23339 = _T_23338 | _T_23084; // @[Mux.scala 27:72]
  wire  _T_22714 = bht_rd_addr_hashed_p1_f == 8'h8d; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_141; // @[Reg.scala 27:20]
  wire [1:0] _T_23085 = _T_22714 ? bht_bank_rd_data_out_0_141 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23340 = _T_23339 | _T_23085; // @[Mux.scala 27:72]
  wire  _T_22716 = bht_rd_addr_hashed_p1_f == 8'h8e; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_142; // @[Reg.scala 27:20]
  wire [1:0] _T_23086 = _T_22716 ? bht_bank_rd_data_out_0_142 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23341 = _T_23340 | _T_23086; // @[Mux.scala 27:72]
  wire  _T_22718 = bht_rd_addr_hashed_p1_f == 8'h8f; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_143; // @[Reg.scala 27:20]
  wire [1:0] _T_23087 = _T_22718 ? bht_bank_rd_data_out_0_143 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23342 = _T_23341 | _T_23087; // @[Mux.scala 27:72]
  wire  _T_22720 = bht_rd_addr_hashed_p1_f == 8'h90; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_144; // @[Reg.scala 27:20]
  wire [1:0] _T_23088 = _T_22720 ? bht_bank_rd_data_out_0_144 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23343 = _T_23342 | _T_23088; // @[Mux.scala 27:72]
  wire  _T_22722 = bht_rd_addr_hashed_p1_f == 8'h91; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_145; // @[Reg.scala 27:20]
  wire [1:0] _T_23089 = _T_22722 ? bht_bank_rd_data_out_0_145 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23344 = _T_23343 | _T_23089; // @[Mux.scala 27:72]
  wire  _T_22724 = bht_rd_addr_hashed_p1_f == 8'h92; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_146; // @[Reg.scala 27:20]
  wire [1:0] _T_23090 = _T_22724 ? bht_bank_rd_data_out_0_146 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23345 = _T_23344 | _T_23090; // @[Mux.scala 27:72]
  wire  _T_22726 = bht_rd_addr_hashed_p1_f == 8'h93; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_147; // @[Reg.scala 27:20]
  wire [1:0] _T_23091 = _T_22726 ? bht_bank_rd_data_out_0_147 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23346 = _T_23345 | _T_23091; // @[Mux.scala 27:72]
  wire  _T_22728 = bht_rd_addr_hashed_p1_f == 8'h94; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_148; // @[Reg.scala 27:20]
  wire [1:0] _T_23092 = _T_22728 ? bht_bank_rd_data_out_0_148 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23347 = _T_23346 | _T_23092; // @[Mux.scala 27:72]
  wire  _T_22730 = bht_rd_addr_hashed_p1_f == 8'h95; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_149; // @[Reg.scala 27:20]
  wire [1:0] _T_23093 = _T_22730 ? bht_bank_rd_data_out_0_149 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23348 = _T_23347 | _T_23093; // @[Mux.scala 27:72]
  wire  _T_22732 = bht_rd_addr_hashed_p1_f == 8'h96; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_150; // @[Reg.scala 27:20]
  wire [1:0] _T_23094 = _T_22732 ? bht_bank_rd_data_out_0_150 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23349 = _T_23348 | _T_23094; // @[Mux.scala 27:72]
  wire  _T_22734 = bht_rd_addr_hashed_p1_f == 8'h97; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_151; // @[Reg.scala 27:20]
  wire [1:0] _T_23095 = _T_22734 ? bht_bank_rd_data_out_0_151 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23350 = _T_23349 | _T_23095; // @[Mux.scala 27:72]
  wire  _T_22736 = bht_rd_addr_hashed_p1_f == 8'h98; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_152; // @[Reg.scala 27:20]
  wire [1:0] _T_23096 = _T_22736 ? bht_bank_rd_data_out_0_152 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23351 = _T_23350 | _T_23096; // @[Mux.scala 27:72]
  wire  _T_22738 = bht_rd_addr_hashed_p1_f == 8'h99; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_153; // @[Reg.scala 27:20]
  wire [1:0] _T_23097 = _T_22738 ? bht_bank_rd_data_out_0_153 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23352 = _T_23351 | _T_23097; // @[Mux.scala 27:72]
  wire  _T_22740 = bht_rd_addr_hashed_p1_f == 8'h9a; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_154; // @[Reg.scala 27:20]
  wire [1:0] _T_23098 = _T_22740 ? bht_bank_rd_data_out_0_154 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23353 = _T_23352 | _T_23098; // @[Mux.scala 27:72]
  wire  _T_22742 = bht_rd_addr_hashed_p1_f == 8'h9b; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_155; // @[Reg.scala 27:20]
  wire [1:0] _T_23099 = _T_22742 ? bht_bank_rd_data_out_0_155 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23354 = _T_23353 | _T_23099; // @[Mux.scala 27:72]
  wire  _T_22744 = bht_rd_addr_hashed_p1_f == 8'h9c; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_156; // @[Reg.scala 27:20]
  wire [1:0] _T_23100 = _T_22744 ? bht_bank_rd_data_out_0_156 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23355 = _T_23354 | _T_23100; // @[Mux.scala 27:72]
  wire  _T_22746 = bht_rd_addr_hashed_p1_f == 8'h9d; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_157; // @[Reg.scala 27:20]
  wire [1:0] _T_23101 = _T_22746 ? bht_bank_rd_data_out_0_157 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23356 = _T_23355 | _T_23101; // @[Mux.scala 27:72]
  wire  _T_22748 = bht_rd_addr_hashed_p1_f == 8'h9e; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_158; // @[Reg.scala 27:20]
  wire [1:0] _T_23102 = _T_22748 ? bht_bank_rd_data_out_0_158 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23357 = _T_23356 | _T_23102; // @[Mux.scala 27:72]
  wire  _T_22750 = bht_rd_addr_hashed_p1_f == 8'h9f; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_159; // @[Reg.scala 27:20]
  wire [1:0] _T_23103 = _T_22750 ? bht_bank_rd_data_out_0_159 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23358 = _T_23357 | _T_23103; // @[Mux.scala 27:72]
  wire  _T_22752 = bht_rd_addr_hashed_p1_f == 8'ha0; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_160; // @[Reg.scala 27:20]
  wire [1:0] _T_23104 = _T_22752 ? bht_bank_rd_data_out_0_160 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23359 = _T_23358 | _T_23104; // @[Mux.scala 27:72]
  wire  _T_22754 = bht_rd_addr_hashed_p1_f == 8'ha1; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_161; // @[Reg.scala 27:20]
  wire [1:0] _T_23105 = _T_22754 ? bht_bank_rd_data_out_0_161 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23360 = _T_23359 | _T_23105; // @[Mux.scala 27:72]
  wire  _T_22756 = bht_rd_addr_hashed_p1_f == 8'ha2; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_162; // @[Reg.scala 27:20]
  wire [1:0] _T_23106 = _T_22756 ? bht_bank_rd_data_out_0_162 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23361 = _T_23360 | _T_23106; // @[Mux.scala 27:72]
  wire  _T_22758 = bht_rd_addr_hashed_p1_f == 8'ha3; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_163; // @[Reg.scala 27:20]
  wire [1:0] _T_23107 = _T_22758 ? bht_bank_rd_data_out_0_163 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23362 = _T_23361 | _T_23107; // @[Mux.scala 27:72]
  wire  _T_22760 = bht_rd_addr_hashed_p1_f == 8'ha4; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_164; // @[Reg.scala 27:20]
  wire [1:0] _T_23108 = _T_22760 ? bht_bank_rd_data_out_0_164 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23363 = _T_23362 | _T_23108; // @[Mux.scala 27:72]
  wire  _T_22762 = bht_rd_addr_hashed_p1_f == 8'ha5; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_165; // @[Reg.scala 27:20]
  wire [1:0] _T_23109 = _T_22762 ? bht_bank_rd_data_out_0_165 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23364 = _T_23363 | _T_23109; // @[Mux.scala 27:72]
  wire  _T_22764 = bht_rd_addr_hashed_p1_f == 8'ha6; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_166; // @[Reg.scala 27:20]
  wire [1:0] _T_23110 = _T_22764 ? bht_bank_rd_data_out_0_166 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23365 = _T_23364 | _T_23110; // @[Mux.scala 27:72]
  wire  _T_22766 = bht_rd_addr_hashed_p1_f == 8'ha7; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_167; // @[Reg.scala 27:20]
  wire [1:0] _T_23111 = _T_22766 ? bht_bank_rd_data_out_0_167 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23366 = _T_23365 | _T_23111; // @[Mux.scala 27:72]
  wire  _T_22768 = bht_rd_addr_hashed_p1_f == 8'ha8; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_168; // @[Reg.scala 27:20]
  wire [1:0] _T_23112 = _T_22768 ? bht_bank_rd_data_out_0_168 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23367 = _T_23366 | _T_23112; // @[Mux.scala 27:72]
  wire  _T_22770 = bht_rd_addr_hashed_p1_f == 8'ha9; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_169; // @[Reg.scala 27:20]
  wire [1:0] _T_23113 = _T_22770 ? bht_bank_rd_data_out_0_169 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23368 = _T_23367 | _T_23113; // @[Mux.scala 27:72]
  wire  _T_22772 = bht_rd_addr_hashed_p1_f == 8'haa; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_170; // @[Reg.scala 27:20]
  wire [1:0] _T_23114 = _T_22772 ? bht_bank_rd_data_out_0_170 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23369 = _T_23368 | _T_23114; // @[Mux.scala 27:72]
  wire  _T_22774 = bht_rd_addr_hashed_p1_f == 8'hab; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_171; // @[Reg.scala 27:20]
  wire [1:0] _T_23115 = _T_22774 ? bht_bank_rd_data_out_0_171 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23370 = _T_23369 | _T_23115; // @[Mux.scala 27:72]
  wire  _T_22776 = bht_rd_addr_hashed_p1_f == 8'hac; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_172; // @[Reg.scala 27:20]
  wire [1:0] _T_23116 = _T_22776 ? bht_bank_rd_data_out_0_172 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23371 = _T_23370 | _T_23116; // @[Mux.scala 27:72]
  wire  _T_22778 = bht_rd_addr_hashed_p1_f == 8'had; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_173; // @[Reg.scala 27:20]
  wire [1:0] _T_23117 = _T_22778 ? bht_bank_rd_data_out_0_173 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23372 = _T_23371 | _T_23117; // @[Mux.scala 27:72]
  wire  _T_22780 = bht_rd_addr_hashed_p1_f == 8'hae; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_174; // @[Reg.scala 27:20]
  wire [1:0] _T_23118 = _T_22780 ? bht_bank_rd_data_out_0_174 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23373 = _T_23372 | _T_23118; // @[Mux.scala 27:72]
  wire  _T_22782 = bht_rd_addr_hashed_p1_f == 8'haf; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_175; // @[Reg.scala 27:20]
  wire [1:0] _T_23119 = _T_22782 ? bht_bank_rd_data_out_0_175 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23374 = _T_23373 | _T_23119; // @[Mux.scala 27:72]
  wire  _T_22784 = bht_rd_addr_hashed_p1_f == 8'hb0; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_176; // @[Reg.scala 27:20]
  wire [1:0] _T_23120 = _T_22784 ? bht_bank_rd_data_out_0_176 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23375 = _T_23374 | _T_23120; // @[Mux.scala 27:72]
  wire  _T_22786 = bht_rd_addr_hashed_p1_f == 8'hb1; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_177; // @[Reg.scala 27:20]
  wire [1:0] _T_23121 = _T_22786 ? bht_bank_rd_data_out_0_177 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23376 = _T_23375 | _T_23121; // @[Mux.scala 27:72]
  wire  _T_22788 = bht_rd_addr_hashed_p1_f == 8'hb2; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_178; // @[Reg.scala 27:20]
  wire [1:0] _T_23122 = _T_22788 ? bht_bank_rd_data_out_0_178 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23377 = _T_23376 | _T_23122; // @[Mux.scala 27:72]
  wire  _T_22790 = bht_rd_addr_hashed_p1_f == 8'hb3; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_179; // @[Reg.scala 27:20]
  wire [1:0] _T_23123 = _T_22790 ? bht_bank_rd_data_out_0_179 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23378 = _T_23377 | _T_23123; // @[Mux.scala 27:72]
  wire  _T_22792 = bht_rd_addr_hashed_p1_f == 8'hb4; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_180; // @[Reg.scala 27:20]
  wire [1:0] _T_23124 = _T_22792 ? bht_bank_rd_data_out_0_180 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23379 = _T_23378 | _T_23124; // @[Mux.scala 27:72]
  wire  _T_22794 = bht_rd_addr_hashed_p1_f == 8'hb5; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_181; // @[Reg.scala 27:20]
  wire [1:0] _T_23125 = _T_22794 ? bht_bank_rd_data_out_0_181 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23380 = _T_23379 | _T_23125; // @[Mux.scala 27:72]
  wire  _T_22796 = bht_rd_addr_hashed_p1_f == 8'hb6; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_182; // @[Reg.scala 27:20]
  wire [1:0] _T_23126 = _T_22796 ? bht_bank_rd_data_out_0_182 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23381 = _T_23380 | _T_23126; // @[Mux.scala 27:72]
  wire  _T_22798 = bht_rd_addr_hashed_p1_f == 8'hb7; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_183; // @[Reg.scala 27:20]
  wire [1:0] _T_23127 = _T_22798 ? bht_bank_rd_data_out_0_183 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23382 = _T_23381 | _T_23127; // @[Mux.scala 27:72]
  wire  _T_22800 = bht_rd_addr_hashed_p1_f == 8'hb8; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_184; // @[Reg.scala 27:20]
  wire [1:0] _T_23128 = _T_22800 ? bht_bank_rd_data_out_0_184 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23383 = _T_23382 | _T_23128; // @[Mux.scala 27:72]
  wire  _T_22802 = bht_rd_addr_hashed_p1_f == 8'hb9; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_185; // @[Reg.scala 27:20]
  wire [1:0] _T_23129 = _T_22802 ? bht_bank_rd_data_out_0_185 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23384 = _T_23383 | _T_23129; // @[Mux.scala 27:72]
  wire  _T_22804 = bht_rd_addr_hashed_p1_f == 8'hba; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_186; // @[Reg.scala 27:20]
  wire [1:0] _T_23130 = _T_22804 ? bht_bank_rd_data_out_0_186 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23385 = _T_23384 | _T_23130; // @[Mux.scala 27:72]
  wire  _T_22806 = bht_rd_addr_hashed_p1_f == 8'hbb; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_187; // @[Reg.scala 27:20]
  wire [1:0] _T_23131 = _T_22806 ? bht_bank_rd_data_out_0_187 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23386 = _T_23385 | _T_23131; // @[Mux.scala 27:72]
  wire  _T_22808 = bht_rd_addr_hashed_p1_f == 8'hbc; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_188; // @[Reg.scala 27:20]
  wire [1:0] _T_23132 = _T_22808 ? bht_bank_rd_data_out_0_188 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23387 = _T_23386 | _T_23132; // @[Mux.scala 27:72]
  wire  _T_22810 = bht_rd_addr_hashed_p1_f == 8'hbd; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_189; // @[Reg.scala 27:20]
  wire [1:0] _T_23133 = _T_22810 ? bht_bank_rd_data_out_0_189 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23388 = _T_23387 | _T_23133; // @[Mux.scala 27:72]
  wire  _T_22812 = bht_rd_addr_hashed_p1_f == 8'hbe; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_190; // @[Reg.scala 27:20]
  wire [1:0] _T_23134 = _T_22812 ? bht_bank_rd_data_out_0_190 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23389 = _T_23388 | _T_23134; // @[Mux.scala 27:72]
  wire  _T_22814 = bht_rd_addr_hashed_p1_f == 8'hbf; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_191; // @[Reg.scala 27:20]
  wire [1:0] _T_23135 = _T_22814 ? bht_bank_rd_data_out_0_191 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23390 = _T_23389 | _T_23135; // @[Mux.scala 27:72]
  wire  _T_22816 = bht_rd_addr_hashed_p1_f == 8'hc0; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_192; // @[Reg.scala 27:20]
  wire [1:0] _T_23136 = _T_22816 ? bht_bank_rd_data_out_0_192 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23391 = _T_23390 | _T_23136; // @[Mux.scala 27:72]
  wire  _T_22818 = bht_rd_addr_hashed_p1_f == 8'hc1; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_193; // @[Reg.scala 27:20]
  wire [1:0] _T_23137 = _T_22818 ? bht_bank_rd_data_out_0_193 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23392 = _T_23391 | _T_23137; // @[Mux.scala 27:72]
  wire  _T_22820 = bht_rd_addr_hashed_p1_f == 8'hc2; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_194; // @[Reg.scala 27:20]
  wire [1:0] _T_23138 = _T_22820 ? bht_bank_rd_data_out_0_194 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23393 = _T_23392 | _T_23138; // @[Mux.scala 27:72]
  wire  _T_22822 = bht_rd_addr_hashed_p1_f == 8'hc3; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_195; // @[Reg.scala 27:20]
  wire [1:0] _T_23139 = _T_22822 ? bht_bank_rd_data_out_0_195 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23394 = _T_23393 | _T_23139; // @[Mux.scala 27:72]
  wire  _T_22824 = bht_rd_addr_hashed_p1_f == 8'hc4; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_196; // @[Reg.scala 27:20]
  wire [1:0] _T_23140 = _T_22824 ? bht_bank_rd_data_out_0_196 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23395 = _T_23394 | _T_23140; // @[Mux.scala 27:72]
  wire  _T_22826 = bht_rd_addr_hashed_p1_f == 8'hc5; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_197; // @[Reg.scala 27:20]
  wire [1:0] _T_23141 = _T_22826 ? bht_bank_rd_data_out_0_197 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23396 = _T_23395 | _T_23141; // @[Mux.scala 27:72]
  wire  _T_22828 = bht_rd_addr_hashed_p1_f == 8'hc6; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_198; // @[Reg.scala 27:20]
  wire [1:0] _T_23142 = _T_22828 ? bht_bank_rd_data_out_0_198 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23397 = _T_23396 | _T_23142; // @[Mux.scala 27:72]
  wire  _T_22830 = bht_rd_addr_hashed_p1_f == 8'hc7; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_199; // @[Reg.scala 27:20]
  wire [1:0] _T_23143 = _T_22830 ? bht_bank_rd_data_out_0_199 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23398 = _T_23397 | _T_23143; // @[Mux.scala 27:72]
  wire  _T_22832 = bht_rd_addr_hashed_p1_f == 8'hc8; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_200; // @[Reg.scala 27:20]
  wire [1:0] _T_23144 = _T_22832 ? bht_bank_rd_data_out_0_200 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23399 = _T_23398 | _T_23144; // @[Mux.scala 27:72]
  wire  _T_22834 = bht_rd_addr_hashed_p1_f == 8'hc9; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_201; // @[Reg.scala 27:20]
  wire [1:0] _T_23145 = _T_22834 ? bht_bank_rd_data_out_0_201 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23400 = _T_23399 | _T_23145; // @[Mux.scala 27:72]
  wire  _T_22836 = bht_rd_addr_hashed_p1_f == 8'hca; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_202; // @[Reg.scala 27:20]
  wire [1:0] _T_23146 = _T_22836 ? bht_bank_rd_data_out_0_202 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23401 = _T_23400 | _T_23146; // @[Mux.scala 27:72]
  wire  _T_22838 = bht_rd_addr_hashed_p1_f == 8'hcb; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_203; // @[Reg.scala 27:20]
  wire [1:0] _T_23147 = _T_22838 ? bht_bank_rd_data_out_0_203 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23402 = _T_23401 | _T_23147; // @[Mux.scala 27:72]
  wire  _T_22840 = bht_rd_addr_hashed_p1_f == 8'hcc; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_204; // @[Reg.scala 27:20]
  wire [1:0] _T_23148 = _T_22840 ? bht_bank_rd_data_out_0_204 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23403 = _T_23402 | _T_23148; // @[Mux.scala 27:72]
  wire  _T_22842 = bht_rd_addr_hashed_p1_f == 8'hcd; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_205; // @[Reg.scala 27:20]
  wire [1:0] _T_23149 = _T_22842 ? bht_bank_rd_data_out_0_205 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23404 = _T_23403 | _T_23149; // @[Mux.scala 27:72]
  wire  _T_22844 = bht_rd_addr_hashed_p1_f == 8'hce; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_206; // @[Reg.scala 27:20]
  wire [1:0] _T_23150 = _T_22844 ? bht_bank_rd_data_out_0_206 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23405 = _T_23404 | _T_23150; // @[Mux.scala 27:72]
  wire  _T_22846 = bht_rd_addr_hashed_p1_f == 8'hcf; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_207; // @[Reg.scala 27:20]
  wire [1:0] _T_23151 = _T_22846 ? bht_bank_rd_data_out_0_207 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23406 = _T_23405 | _T_23151; // @[Mux.scala 27:72]
  wire  _T_22848 = bht_rd_addr_hashed_p1_f == 8'hd0; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_208; // @[Reg.scala 27:20]
  wire [1:0] _T_23152 = _T_22848 ? bht_bank_rd_data_out_0_208 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23407 = _T_23406 | _T_23152; // @[Mux.scala 27:72]
  wire  _T_22850 = bht_rd_addr_hashed_p1_f == 8'hd1; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_209; // @[Reg.scala 27:20]
  wire [1:0] _T_23153 = _T_22850 ? bht_bank_rd_data_out_0_209 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23408 = _T_23407 | _T_23153; // @[Mux.scala 27:72]
  wire  _T_22852 = bht_rd_addr_hashed_p1_f == 8'hd2; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_210; // @[Reg.scala 27:20]
  wire [1:0] _T_23154 = _T_22852 ? bht_bank_rd_data_out_0_210 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23409 = _T_23408 | _T_23154; // @[Mux.scala 27:72]
  wire  _T_22854 = bht_rd_addr_hashed_p1_f == 8'hd3; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_211; // @[Reg.scala 27:20]
  wire [1:0] _T_23155 = _T_22854 ? bht_bank_rd_data_out_0_211 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23410 = _T_23409 | _T_23155; // @[Mux.scala 27:72]
  wire  _T_22856 = bht_rd_addr_hashed_p1_f == 8'hd4; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_212; // @[Reg.scala 27:20]
  wire [1:0] _T_23156 = _T_22856 ? bht_bank_rd_data_out_0_212 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23411 = _T_23410 | _T_23156; // @[Mux.scala 27:72]
  wire  _T_22858 = bht_rd_addr_hashed_p1_f == 8'hd5; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_213; // @[Reg.scala 27:20]
  wire [1:0] _T_23157 = _T_22858 ? bht_bank_rd_data_out_0_213 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23412 = _T_23411 | _T_23157; // @[Mux.scala 27:72]
  wire  _T_22860 = bht_rd_addr_hashed_p1_f == 8'hd6; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_214; // @[Reg.scala 27:20]
  wire [1:0] _T_23158 = _T_22860 ? bht_bank_rd_data_out_0_214 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23413 = _T_23412 | _T_23158; // @[Mux.scala 27:72]
  wire  _T_22862 = bht_rd_addr_hashed_p1_f == 8'hd7; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_215; // @[Reg.scala 27:20]
  wire [1:0] _T_23159 = _T_22862 ? bht_bank_rd_data_out_0_215 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23414 = _T_23413 | _T_23159; // @[Mux.scala 27:72]
  wire  _T_22864 = bht_rd_addr_hashed_p1_f == 8'hd8; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_216; // @[Reg.scala 27:20]
  wire [1:0] _T_23160 = _T_22864 ? bht_bank_rd_data_out_0_216 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23415 = _T_23414 | _T_23160; // @[Mux.scala 27:72]
  wire  _T_22866 = bht_rd_addr_hashed_p1_f == 8'hd9; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_217; // @[Reg.scala 27:20]
  wire [1:0] _T_23161 = _T_22866 ? bht_bank_rd_data_out_0_217 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23416 = _T_23415 | _T_23161; // @[Mux.scala 27:72]
  wire  _T_22868 = bht_rd_addr_hashed_p1_f == 8'hda; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_218; // @[Reg.scala 27:20]
  wire [1:0] _T_23162 = _T_22868 ? bht_bank_rd_data_out_0_218 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23417 = _T_23416 | _T_23162; // @[Mux.scala 27:72]
  wire  _T_22870 = bht_rd_addr_hashed_p1_f == 8'hdb; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_219; // @[Reg.scala 27:20]
  wire [1:0] _T_23163 = _T_22870 ? bht_bank_rd_data_out_0_219 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23418 = _T_23417 | _T_23163; // @[Mux.scala 27:72]
  wire  _T_22872 = bht_rd_addr_hashed_p1_f == 8'hdc; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_220; // @[Reg.scala 27:20]
  wire [1:0] _T_23164 = _T_22872 ? bht_bank_rd_data_out_0_220 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23419 = _T_23418 | _T_23164; // @[Mux.scala 27:72]
  wire  _T_22874 = bht_rd_addr_hashed_p1_f == 8'hdd; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_221; // @[Reg.scala 27:20]
  wire [1:0] _T_23165 = _T_22874 ? bht_bank_rd_data_out_0_221 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23420 = _T_23419 | _T_23165; // @[Mux.scala 27:72]
  wire  _T_22876 = bht_rd_addr_hashed_p1_f == 8'hde; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_222; // @[Reg.scala 27:20]
  wire [1:0] _T_23166 = _T_22876 ? bht_bank_rd_data_out_0_222 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23421 = _T_23420 | _T_23166; // @[Mux.scala 27:72]
  wire  _T_22878 = bht_rd_addr_hashed_p1_f == 8'hdf; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_223; // @[Reg.scala 27:20]
  wire [1:0] _T_23167 = _T_22878 ? bht_bank_rd_data_out_0_223 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23422 = _T_23421 | _T_23167; // @[Mux.scala 27:72]
  wire  _T_22880 = bht_rd_addr_hashed_p1_f == 8'he0; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_224; // @[Reg.scala 27:20]
  wire [1:0] _T_23168 = _T_22880 ? bht_bank_rd_data_out_0_224 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23423 = _T_23422 | _T_23168; // @[Mux.scala 27:72]
  wire  _T_22882 = bht_rd_addr_hashed_p1_f == 8'he1; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_225; // @[Reg.scala 27:20]
  wire [1:0] _T_23169 = _T_22882 ? bht_bank_rd_data_out_0_225 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23424 = _T_23423 | _T_23169; // @[Mux.scala 27:72]
  wire  _T_22884 = bht_rd_addr_hashed_p1_f == 8'he2; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_226; // @[Reg.scala 27:20]
  wire [1:0] _T_23170 = _T_22884 ? bht_bank_rd_data_out_0_226 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23425 = _T_23424 | _T_23170; // @[Mux.scala 27:72]
  wire  _T_22886 = bht_rd_addr_hashed_p1_f == 8'he3; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_227; // @[Reg.scala 27:20]
  wire [1:0] _T_23171 = _T_22886 ? bht_bank_rd_data_out_0_227 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23426 = _T_23425 | _T_23171; // @[Mux.scala 27:72]
  wire  _T_22888 = bht_rd_addr_hashed_p1_f == 8'he4; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_228; // @[Reg.scala 27:20]
  wire [1:0] _T_23172 = _T_22888 ? bht_bank_rd_data_out_0_228 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23427 = _T_23426 | _T_23172; // @[Mux.scala 27:72]
  wire  _T_22890 = bht_rd_addr_hashed_p1_f == 8'he5; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_229; // @[Reg.scala 27:20]
  wire [1:0] _T_23173 = _T_22890 ? bht_bank_rd_data_out_0_229 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23428 = _T_23427 | _T_23173; // @[Mux.scala 27:72]
  wire  _T_22892 = bht_rd_addr_hashed_p1_f == 8'he6; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_230; // @[Reg.scala 27:20]
  wire [1:0] _T_23174 = _T_22892 ? bht_bank_rd_data_out_0_230 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23429 = _T_23428 | _T_23174; // @[Mux.scala 27:72]
  wire  _T_22894 = bht_rd_addr_hashed_p1_f == 8'he7; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_231; // @[Reg.scala 27:20]
  wire [1:0] _T_23175 = _T_22894 ? bht_bank_rd_data_out_0_231 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23430 = _T_23429 | _T_23175; // @[Mux.scala 27:72]
  wire  _T_22896 = bht_rd_addr_hashed_p1_f == 8'he8; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_232; // @[Reg.scala 27:20]
  wire [1:0] _T_23176 = _T_22896 ? bht_bank_rd_data_out_0_232 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23431 = _T_23430 | _T_23176; // @[Mux.scala 27:72]
  wire  _T_22898 = bht_rd_addr_hashed_p1_f == 8'he9; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_233; // @[Reg.scala 27:20]
  wire [1:0] _T_23177 = _T_22898 ? bht_bank_rd_data_out_0_233 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23432 = _T_23431 | _T_23177; // @[Mux.scala 27:72]
  wire  _T_22900 = bht_rd_addr_hashed_p1_f == 8'hea; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_234; // @[Reg.scala 27:20]
  wire [1:0] _T_23178 = _T_22900 ? bht_bank_rd_data_out_0_234 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23433 = _T_23432 | _T_23178; // @[Mux.scala 27:72]
  wire  _T_22902 = bht_rd_addr_hashed_p1_f == 8'heb; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_235; // @[Reg.scala 27:20]
  wire [1:0] _T_23179 = _T_22902 ? bht_bank_rd_data_out_0_235 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23434 = _T_23433 | _T_23179; // @[Mux.scala 27:72]
  wire  _T_22904 = bht_rd_addr_hashed_p1_f == 8'hec; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_236; // @[Reg.scala 27:20]
  wire [1:0] _T_23180 = _T_22904 ? bht_bank_rd_data_out_0_236 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23435 = _T_23434 | _T_23180; // @[Mux.scala 27:72]
  wire  _T_22906 = bht_rd_addr_hashed_p1_f == 8'hed; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_237; // @[Reg.scala 27:20]
  wire [1:0] _T_23181 = _T_22906 ? bht_bank_rd_data_out_0_237 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23436 = _T_23435 | _T_23181; // @[Mux.scala 27:72]
  wire  _T_22908 = bht_rd_addr_hashed_p1_f == 8'hee; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_238; // @[Reg.scala 27:20]
  wire [1:0] _T_23182 = _T_22908 ? bht_bank_rd_data_out_0_238 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23437 = _T_23436 | _T_23182; // @[Mux.scala 27:72]
  wire  _T_22910 = bht_rd_addr_hashed_p1_f == 8'hef; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_239; // @[Reg.scala 27:20]
  wire [1:0] _T_23183 = _T_22910 ? bht_bank_rd_data_out_0_239 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23438 = _T_23437 | _T_23183; // @[Mux.scala 27:72]
  wire  _T_22912 = bht_rd_addr_hashed_p1_f == 8'hf0; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_240; // @[Reg.scala 27:20]
  wire [1:0] _T_23184 = _T_22912 ? bht_bank_rd_data_out_0_240 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23439 = _T_23438 | _T_23184; // @[Mux.scala 27:72]
  wire  _T_22914 = bht_rd_addr_hashed_p1_f == 8'hf1; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_241; // @[Reg.scala 27:20]
  wire [1:0] _T_23185 = _T_22914 ? bht_bank_rd_data_out_0_241 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23440 = _T_23439 | _T_23185; // @[Mux.scala 27:72]
  wire  _T_22916 = bht_rd_addr_hashed_p1_f == 8'hf2; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_242; // @[Reg.scala 27:20]
  wire [1:0] _T_23186 = _T_22916 ? bht_bank_rd_data_out_0_242 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23441 = _T_23440 | _T_23186; // @[Mux.scala 27:72]
  wire  _T_22918 = bht_rd_addr_hashed_p1_f == 8'hf3; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_243; // @[Reg.scala 27:20]
  wire [1:0] _T_23187 = _T_22918 ? bht_bank_rd_data_out_0_243 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23442 = _T_23441 | _T_23187; // @[Mux.scala 27:72]
  wire  _T_22920 = bht_rd_addr_hashed_p1_f == 8'hf4; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_244; // @[Reg.scala 27:20]
  wire [1:0] _T_23188 = _T_22920 ? bht_bank_rd_data_out_0_244 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23443 = _T_23442 | _T_23188; // @[Mux.scala 27:72]
  wire  _T_22922 = bht_rd_addr_hashed_p1_f == 8'hf5; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_245; // @[Reg.scala 27:20]
  wire [1:0] _T_23189 = _T_22922 ? bht_bank_rd_data_out_0_245 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23444 = _T_23443 | _T_23189; // @[Mux.scala 27:72]
  wire  _T_22924 = bht_rd_addr_hashed_p1_f == 8'hf6; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_246; // @[Reg.scala 27:20]
  wire [1:0] _T_23190 = _T_22924 ? bht_bank_rd_data_out_0_246 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23445 = _T_23444 | _T_23190; // @[Mux.scala 27:72]
  wire  _T_22926 = bht_rd_addr_hashed_p1_f == 8'hf7; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_247; // @[Reg.scala 27:20]
  wire [1:0] _T_23191 = _T_22926 ? bht_bank_rd_data_out_0_247 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23446 = _T_23445 | _T_23191; // @[Mux.scala 27:72]
  wire  _T_22928 = bht_rd_addr_hashed_p1_f == 8'hf8; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_248; // @[Reg.scala 27:20]
  wire [1:0] _T_23192 = _T_22928 ? bht_bank_rd_data_out_0_248 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23447 = _T_23446 | _T_23192; // @[Mux.scala 27:72]
  wire  _T_22930 = bht_rd_addr_hashed_p1_f == 8'hf9; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_249; // @[Reg.scala 27:20]
  wire [1:0] _T_23193 = _T_22930 ? bht_bank_rd_data_out_0_249 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23448 = _T_23447 | _T_23193; // @[Mux.scala 27:72]
  wire  _T_22932 = bht_rd_addr_hashed_p1_f == 8'hfa; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_250; // @[Reg.scala 27:20]
  wire [1:0] _T_23194 = _T_22932 ? bht_bank_rd_data_out_0_250 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23449 = _T_23448 | _T_23194; // @[Mux.scala 27:72]
  wire  _T_22934 = bht_rd_addr_hashed_p1_f == 8'hfb; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_251; // @[Reg.scala 27:20]
  wire [1:0] _T_23195 = _T_22934 ? bht_bank_rd_data_out_0_251 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23450 = _T_23449 | _T_23195; // @[Mux.scala 27:72]
  wire  _T_22936 = bht_rd_addr_hashed_p1_f == 8'hfc; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_252; // @[Reg.scala 27:20]
  wire [1:0] _T_23196 = _T_22936 ? bht_bank_rd_data_out_0_252 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23451 = _T_23450 | _T_23196; // @[Mux.scala 27:72]
  wire  _T_22938 = bht_rd_addr_hashed_p1_f == 8'hfd; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_253; // @[Reg.scala 27:20]
  wire [1:0] _T_23197 = _T_22938 ? bht_bank_rd_data_out_0_253 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23452 = _T_23451 | _T_23197; // @[Mux.scala 27:72]
  wire  _T_22940 = bht_rd_addr_hashed_p1_f == 8'hfe; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_254; // @[Reg.scala 27:20]
  wire [1:0] _T_23198 = _T_22940 ? bht_bank_rd_data_out_0_254 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23453 = _T_23452 | _T_23198; // @[Mux.scala 27:72]
  wire  _T_22942 = bht_rd_addr_hashed_p1_f == 8'hff; // @[ifu_bp_ctl.scala 456:85]
  reg [1:0] bht_bank_rd_data_out_0_255; // @[Reg.scala 27:20]
  wire [1:0] _T_23199 = _T_22942 ? bht_bank_rd_data_out_0_255 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] bht_bank0_rd_data_p1_f = _T_23453 | _T_23199; // @[Mux.scala 27:72]
  wire [1:0] _T_261 = io_ifc_fetch_addr_f[0] ? bht_bank0_rd_data_p1_f : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] bht_vbank1_rd_data_f = _T_260 | _T_261; // @[Mux.scala 27:72]
  wire  _T_265 = bht_force_taken_f[1] | bht_vbank1_rd_data_f[1]; // @[ifu_bp_ctl.scala 281:42]
  wire [1:0] wayhit_f = tag_match_way0_expanded_f | tag_match_way1_expanded_f; // @[ifu_bp_ctl.scala 155:44]
  wire [1:0] _T_159 = _T_144 ? wayhit_f : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] wayhit_p1_f = tag_match_way0_expanded_p1_f | tag_match_way1_expanded_p1_f; // @[ifu_bp_ctl.scala 157:50]
  wire [1:0] _T_158 = {wayhit_p1_f[0],wayhit_f[1]}; // @[Cat.scala 29:58]
  wire [1:0] _T_160 = io_ifc_fetch_addr_f[0] ? _T_158 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_161 = _T_159 | _T_160; // @[Mux.scala 27:72]
  wire  eoc_near = &io_ifc_fetch_addr_f[4:2]; // @[ifu_bp_ctl.scala 241:64]
  wire  _T_219 = ~eoc_near; // @[ifu_bp_ctl.scala 244:15]
  wire [1:0] _T_221 = ~io_ifc_fetch_addr_f[1:0]; // @[ifu_bp_ctl.scala 244:28]
  wire  _T_222 = |_T_221; // @[ifu_bp_ctl.scala 244:58]
  wire  eoc_mask = _T_219 | _T_222; // @[ifu_bp_ctl.scala 244:25]
  wire [1:0] _T_163 = {eoc_mask,1'h1}; // @[Cat.scala 29:58]
  wire [1:0] bht_valid_f = _T_161 & _T_163; // @[ifu_bp_ctl.scala 203:71]
  wire  _T_267 = _T_265 & bht_valid_f[1]; // @[ifu_bp_ctl.scala 281:69]
  wire [1:0] _T_20896 = _T_21408 ? bht_bank_rd_data_out_0_0 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20897 = _T_21410 ? bht_bank_rd_data_out_0_1 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21152 = _T_20896 | _T_20897; // @[Mux.scala 27:72]
  wire [1:0] _T_20898 = _T_21412 ? bht_bank_rd_data_out_0_2 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21153 = _T_21152 | _T_20898; // @[Mux.scala 27:72]
  wire [1:0] _T_20899 = _T_21414 ? bht_bank_rd_data_out_0_3 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21154 = _T_21153 | _T_20899; // @[Mux.scala 27:72]
  wire [1:0] _T_20900 = _T_21416 ? bht_bank_rd_data_out_0_4 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21155 = _T_21154 | _T_20900; // @[Mux.scala 27:72]
  wire [1:0] _T_20901 = _T_21418 ? bht_bank_rd_data_out_0_5 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21156 = _T_21155 | _T_20901; // @[Mux.scala 27:72]
  wire [1:0] _T_20902 = _T_21420 ? bht_bank_rd_data_out_0_6 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21157 = _T_21156 | _T_20902; // @[Mux.scala 27:72]
  wire [1:0] _T_20903 = _T_21422 ? bht_bank_rd_data_out_0_7 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21158 = _T_21157 | _T_20903; // @[Mux.scala 27:72]
  wire [1:0] _T_20904 = _T_21424 ? bht_bank_rd_data_out_0_8 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21159 = _T_21158 | _T_20904; // @[Mux.scala 27:72]
  wire [1:0] _T_20905 = _T_21426 ? bht_bank_rd_data_out_0_9 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21160 = _T_21159 | _T_20905; // @[Mux.scala 27:72]
  wire [1:0] _T_20906 = _T_21428 ? bht_bank_rd_data_out_0_10 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21161 = _T_21160 | _T_20906; // @[Mux.scala 27:72]
  wire [1:0] _T_20907 = _T_21430 ? bht_bank_rd_data_out_0_11 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21162 = _T_21161 | _T_20907; // @[Mux.scala 27:72]
  wire [1:0] _T_20908 = _T_21432 ? bht_bank_rd_data_out_0_12 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21163 = _T_21162 | _T_20908; // @[Mux.scala 27:72]
  wire [1:0] _T_20909 = _T_21434 ? bht_bank_rd_data_out_0_13 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21164 = _T_21163 | _T_20909; // @[Mux.scala 27:72]
  wire [1:0] _T_20910 = _T_21436 ? bht_bank_rd_data_out_0_14 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21165 = _T_21164 | _T_20910; // @[Mux.scala 27:72]
  wire [1:0] _T_20911 = _T_21438 ? bht_bank_rd_data_out_0_15 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21166 = _T_21165 | _T_20911; // @[Mux.scala 27:72]
  wire [1:0] _T_20912 = _T_21440 ? bht_bank_rd_data_out_0_16 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21167 = _T_21166 | _T_20912; // @[Mux.scala 27:72]
  wire [1:0] _T_20913 = _T_21442 ? bht_bank_rd_data_out_0_17 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21168 = _T_21167 | _T_20913; // @[Mux.scala 27:72]
  wire [1:0] _T_20914 = _T_21444 ? bht_bank_rd_data_out_0_18 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21169 = _T_21168 | _T_20914; // @[Mux.scala 27:72]
  wire [1:0] _T_20915 = _T_21446 ? bht_bank_rd_data_out_0_19 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21170 = _T_21169 | _T_20915; // @[Mux.scala 27:72]
  wire [1:0] _T_20916 = _T_21448 ? bht_bank_rd_data_out_0_20 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21171 = _T_21170 | _T_20916; // @[Mux.scala 27:72]
  wire [1:0] _T_20917 = _T_21450 ? bht_bank_rd_data_out_0_21 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21172 = _T_21171 | _T_20917; // @[Mux.scala 27:72]
  wire [1:0] _T_20918 = _T_21452 ? bht_bank_rd_data_out_0_22 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21173 = _T_21172 | _T_20918; // @[Mux.scala 27:72]
  wire [1:0] _T_20919 = _T_21454 ? bht_bank_rd_data_out_0_23 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21174 = _T_21173 | _T_20919; // @[Mux.scala 27:72]
  wire [1:0] _T_20920 = _T_21456 ? bht_bank_rd_data_out_0_24 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21175 = _T_21174 | _T_20920; // @[Mux.scala 27:72]
  wire [1:0] _T_20921 = _T_21458 ? bht_bank_rd_data_out_0_25 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21176 = _T_21175 | _T_20921; // @[Mux.scala 27:72]
  wire [1:0] _T_20922 = _T_21460 ? bht_bank_rd_data_out_0_26 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21177 = _T_21176 | _T_20922; // @[Mux.scala 27:72]
  wire [1:0] _T_20923 = _T_21462 ? bht_bank_rd_data_out_0_27 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21178 = _T_21177 | _T_20923; // @[Mux.scala 27:72]
  wire [1:0] _T_20924 = _T_21464 ? bht_bank_rd_data_out_0_28 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21179 = _T_21178 | _T_20924; // @[Mux.scala 27:72]
  wire [1:0] _T_20925 = _T_21466 ? bht_bank_rd_data_out_0_29 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21180 = _T_21179 | _T_20925; // @[Mux.scala 27:72]
  wire [1:0] _T_20926 = _T_21468 ? bht_bank_rd_data_out_0_30 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21181 = _T_21180 | _T_20926; // @[Mux.scala 27:72]
  wire [1:0] _T_20927 = _T_21470 ? bht_bank_rd_data_out_0_31 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21182 = _T_21181 | _T_20927; // @[Mux.scala 27:72]
  wire [1:0] _T_20928 = _T_21472 ? bht_bank_rd_data_out_0_32 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21183 = _T_21182 | _T_20928; // @[Mux.scala 27:72]
  wire [1:0] _T_20929 = _T_21474 ? bht_bank_rd_data_out_0_33 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21184 = _T_21183 | _T_20929; // @[Mux.scala 27:72]
  wire [1:0] _T_20930 = _T_21476 ? bht_bank_rd_data_out_0_34 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21185 = _T_21184 | _T_20930; // @[Mux.scala 27:72]
  wire [1:0] _T_20931 = _T_21478 ? bht_bank_rd_data_out_0_35 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21186 = _T_21185 | _T_20931; // @[Mux.scala 27:72]
  wire [1:0] _T_20932 = _T_21480 ? bht_bank_rd_data_out_0_36 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21187 = _T_21186 | _T_20932; // @[Mux.scala 27:72]
  wire [1:0] _T_20933 = _T_21482 ? bht_bank_rd_data_out_0_37 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21188 = _T_21187 | _T_20933; // @[Mux.scala 27:72]
  wire [1:0] _T_20934 = _T_21484 ? bht_bank_rd_data_out_0_38 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21189 = _T_21188 | _T_20934; // @[Mux.scala 27:72]
  wire [1:0] _T_20935 = _T_21486 ? bht_bank_rd_data_out_0_39 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21190 = _T_21189 | _T_20935; // @[Mux.scala 27:72]
  wire [1:0] _T_20936 = _T_21488 ? bht_bank_rd_data_out_0_40 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21191 = _T_21190 | _T_20936; // @[Mux.scala 27:72]
  wire [1:0] _T_20937 = _T_21490 ? bht_bank_rd_data_out_0_41 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21192 = _T_21191 | _T_20937; // @[Mux.scala 27:72]
  wire [1:0] _T_20938 = _T_21492 ? bht_bank_rd_data_out_0_42 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21193 = _T_21192 | _T_20938; // @[Mux.scala 27:72]
  wire [1:0] _T_20939 = _T_21494 ? bht_bank_rd_data_out_0_43 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21194 = _T_21193 | _T_20939; // @[Mux.scala 27:72]
  wire [1:0] _T_20940 = _T_21496 ? bht_bank_rd_data_out_0_44 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21195 = _T_21194 | _T_20940; // @[Mux.scala 27:72]
  wire [1:0] _T_20941 = _T_21498 ? bht_bank_rd_data_out_0_45 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21196 = _T_21195 | _T_20941; // @[Mux.scala 27:72]
  wire [1:0] _T_20942 = _T_21500 ? bht_bank_rd_data_out_0_46 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21197 = _T_21196 | _T_20942; // @[Mux.scala 27:72]
  wire [1:0] _T_20943 = _T_21502 ? bht_bank_rd_data_out_0_47 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21198 = _T_21197 | _T_20943; // @[Mux.scala 27:72]
  wire [1:0] _T_20944 = _T_21504 ? bht_bank_rd_data_out_0_48 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21199 = _T_21198 | _T_20944; // @[Mux.scala 27:72]
  wire [1:0] _T_20945 = _T_21506 ? bht_bank_rd_data_out_0_49 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21200 = _T_21199 | _T_20945; // @[Mux.scala 27:72]
  wire [1:0] _T_20946 = _T_21508 ? bht_bank_rd_data_out_0_50 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21201 = _T_21200 | _T_20946; // @[Mux.scala 27:72]
  wire [1:0] _T_20947 = _T_21510 ? bht_bank_rd_data_out_0_51 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21202 = _T_21201 | _T_20947; // @[Mux.scala 27:72]
  wire [1:0] _T_20948 = _T_21512 ? bht_bank_rd_data_out_0_52 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21203 = _T_21202 | _T_20948; // @[Mux.scala 27:72]
  wire [1:0] _T_20949 = _T_21514 ? bht_bank_rd_data_out_0_53 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21204 = _T_21203 | _T_20949; // @[Mux.scala 27:72]
  wire [1:0] _T_20950 = _T_21516 ? bht_bank_rd_data_out_0_54 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21205 = _T_21204 | _T_20950; // @[Mux.scala 27:72]
  wire [1:0] _T_20951 = _T_21518 ? bht_bank_rd_data_out_0_55 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21206 = _T_21205 | _T_20951; // @[Mux.scala 27:72]
  wire [1:0] _T_20952 = _T_21520 ? bht_bank_rd_data_out_0_56 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21207 = _T_21206 | _T_20952; // @[Mux.scala 27:72]
  wire [1:0] _T_20953 = _T_21522 ? bht_bank_rd_data_out_0_57 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21208 = _T_21207 | _T_20953; // @[Mux.scala 27:72]
  wire [1:0] _T_20954 = _T_21524 ? bht_bank_rd_data_out_0_58 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21209 = _T_21208 | _T_20954; // @[Mux.scala 27:72]
  wire [1:0] _T_20955 = _T_21526 ? bht_bank_rd_data_out_0_59 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21210 = _T_21209 | _T_20955; // @[Mux.scala 27:72]
  wire [1:0] _T_20956 = _T_21528 ? bht_bank_rd_data_out_0_60 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21211 = _T_21210 | _T_20956; // @[Mux.scala 27:72]
  wire [1:0] _T_20957 = _T_21530 ? bht_bank_rd_data_out_0_61 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21212 = _T_21211 | _T_20957; // @[Mux.scala 27:72]
  wire [1:0] _T_20958 = _T_21532 ? bht_bank_rd_data_out_0_62 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21213 = _T_21212 | _T_20958; // @[Mux.scala 27:72]
  wire [1:0] _T_20959 = _T_21534 ? bht_bank_rd_data_out_0_63 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21214 = _T_21213 | _T_20959; // @[Mux.scala 27:72]
  wire [1:0] _T_20960 = _T_21536 ? bht_bank_rd_data_out_0_64 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21215 = _T_21214 | _T_20960; // @[Mux.scala 27:72]
  wire [1:0] _T_20961 = _T_21538 ? bht_bank_rd_data_out_0_65 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21216 = _T_21215 | _T_20961; // @[Mux.scala 27:72]
  wire [1:0] _T_20962 = _T_21540 ? bht_bank_rd_data_out_0_66 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21217 = _T_21216 | _T_20962; // @[Mux.scala 27:72]
  wire [1:0] _T_20963 = _T_21542 ? bht_bank_rd_data_out_0_67 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21218 = _T_21217 | _T_20963; // @[Mux.scala 27:72]
  wire [1:0] _T_20964 = _T_21544 ? bht_bank_rd_data_out_0_68 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21219 = _T_21218 | _T_20964; // @[Mux.scala 27:72]
  wire [1:0] _T_20965 = _T_21546 ? bht_bank_rd_data_out_0_69 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21220 = _T_21219 | _T_20965; // @[Mux.scala 27:72]
  wire [1:0] _T_20966 = _T_21548 ? bht_bank_rd_data_out_0_70 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21221 = _T_21220 | _T_20966; // @[Mux.scala 27:72]
  wire [1:0] _T_20967 = _T_21550 ? bht_bank_rd_data_out_0_71 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21222 = _T_21221 | _T_20967; // @[Mux.scala 27:72]
  wire [1:0] _T_20968 = _T_21552 ? bht_bank_rd_data_out_0_72 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21223 = _T_21222 | _T_20968; // @[Mux.scala 27:72]
  wire [1:0] _T_20969 = _T_21554 ? bht_bank_rd_data_out_0_73 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21224 = _T_21223 | _T_20969; // @[Mux.scala 27:72]
  wire [1:0] _T_20970 = _T_21556 ? bht_bank_rd_data_out_0_74 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21225 = _T_21224 | _T_20970; // @[Mux.scala 27:72]
  wire [1:0] _T_20971 = _T_21558 ? bht_bank_rd_data_out_0_75 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21226 = _T_21225 | _T_20971; // @[Mux.scala 27:72]
  wire [1:0] _T_20972 = _T_21560 ? bht_bank_rd_data_out_0_76 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21227 = _T_21226 | _T_20972; // @[Mux.scala 27:72]
  wire [1:0] _T_20973 = _T_21562 ? bht_bank_rd_data_out_0_77 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21228 = _T_21227 | _T_20973; // @[Mux.scala 27:72]
  wire [1:0] _T_20974 = _T_21564 ? bht_bank_rd_data_out_0_78 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21229 = _T_21228 | _T_20974; // @[Mux.scala 27:72]
  wire [1:0] _T_20975 = _T_21566 ? bht_bank_rd_data_out_0_79 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21230 = _T_21229 | _T_20975; // @[Mux.scala 27:72]
  wire [1:0] _T_20976 = _T_21568 ? bht_bank_rd_data_out_0_80 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21231 = _T_21230 | _T_20976; // @[Mux.scala 27:72]
  wire [1:0] _T_20977 = _T_21570 ? bht_bank_rd_data_out_0_81 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21232 = _T_21231 | _T_20977; // @[Mux.scala 27:72]
  wire [1:0] _T_20978 = _T_21572 ? bht_bank_rd_data_out_0_82 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21233 = _T_21232 | _T_20978; // @[Mux.scala 27:72]
  wire [1:0] _T_20979 = _T_21574 ? bht_bank_rd_data_out_0_83 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21234 = _T_21233 | _T_20979; // @[Mux.scala 27:72]
  wire [1:0] _T_20980 = _T_21576 ? bht_bank_rd_data_out_0_84 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21235 = _T_21234 | _T_20980; // @[Mux.scala 27:72]
  wire [1:0] _T_20981 = _T_21578 ? bht_bank_rd_data_out_0_85 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21236 = _T_21235 | _T_20981; // @[Mux.scala 27:72]
  wire [1:0] _T_20982 = _T_21580 ? bht_bank_rd_data_out_0_86 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21237 = _T_21236 | _T_20982; // @[Mux.scala 27:72]
  wire [1:0] _T_20983 = _T_21582 ? bht_bank_rd_data_out_0_87 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21238 = _T_21237 | _T_20983; // @[Mux.scala 27:72]
  wire [1:0] _T_20984 = _T_21584 ? bht_bank_rd_data_out_0_88 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21239 = _T_21238 | _T_20984; // @[Mux.scala 27:72]
  wire [1:0] _T_20985 = _T_21586 ? bht_bank_rd_data_out_0_89 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21240 = _T_21239 | _T_20985; // @[Mux.scala 27:72]
  wire [1:0] _T_20986 = _T_21588 ? bht_bank_rd_data_out_0_90 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21241 = _T_21240 | _T_20986; // @[Mux.scala 27:72]
  wire [1:0] _T_20987 = _T_21590 ? bht_bank_rd_data_out_0_91 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21242 = _T_21241 | _T_20987; // @[Mux.scala 27:72]
  wire [1:0] _T_20988 = _T_21592 ? bht_bank_rd_data_out_0_92 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21243 = _T_21242 | _T_20988; // @[Mux.scala 27:72]
  wire [1:0] _T_20989 = _T_21594 ? bht_bank_rd_data_out_0_93 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21244 = _T_21243 | _T_20989; // @[Mux.scala 27:72]
  wire [1:0] _T_20990 = _T_21596 ? bht_bank_rd_data_out_0_94 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21245 = _T_21244 | _T_20990; // @[Mux.scala 27:72]
  wire [1:0] _T_20991 = _T_21598 ? bht_bank_rd_data_out_0_95 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21246 = _T_21245 | _T_20991; // @[Mux.scala 27:72]
  wire [1:0] _T_20992 = _T_21600 ? bht_bank_rd_data_out_0_96 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21247 = _T_21246 | _T_20992; // @[Mux.scala 27:72]
  wire [1:0] _T_20993 = _T_21602 ? bht_bank_rd_data_out_0_97 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21248 = _T_21247 | _T_20993; // @[Mux.scala 27:72]
  wire [1:0] _T_20994 = _T_21604 ? bht_bank_rd_data_out_0_98 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21249 = _T_21248 | _T_20994; // @[Mux.scala 27:72]
  wire [1:0] _T_20995 = _T_21606 ? bht_bank_rd_data_out_0_99 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21250 = _T_21249 | _T_20995; // @[Mux.scala 27:72]
  wire [1:0] _T_20996 = _T_21608 ? bht_bank_rd_data_out_0_100 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21251 = _T_21250 | _T_20996; // @[Mux.scala 27:72]
  wire [1:0] _T_20997 = _T_21610 ? bht_bank_rd_data_out_0_101 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21252 = _T_21251 | _T_20997; // @[Mux.scala 27:72]
  wire [1:0] _T_20998 = _T_21612 ? bht_bank_rd_data_out_0_102 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21253 = _T_21252 | _T_20998; // @[Mux.scala 27:72]
  wire [1:0] _T_20999 = _T_21614 ? bht_bank_rd_data_out_0_103 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21254 = _T_21253 | _T_20999; // @[Mux.scala 27:72]
  wire [1:0] _T_21000 = _T_21616 ? bht_bank_rd_data_out_0_104 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21255 = _T_21254 | _T_21000; // @[Mux.scala 27:72]
  wire [1:0] _T_21001 = _T_21618 ? bht_bank_rd_data_out_0_105 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21256 = _T_21255 | _T_21001; // @[Mux.scala 27:72]
  wire [1:0] _T_21002 = _T_21620 ? bht_bank_rd_data_out_0_106 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21257 = _T_21256 | _T_21002; // @[Mux.scala 27:72]
  wire [1:0] _T_21003 = _T_21622 ? bht_bank_rd_data_out_0_107 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21258 = _T_21257 | _T_21003; // @[Mux.scala 27:72]
  wire [1:0] _T_21004 = _T_21624 ? bht_bank_rd_data_out_0_108 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21259 = _T_21258 | _T_21004; // @[Mux.scala 27:72]
  wire [1:0] _T_21005 = _T_21626 ? bht_bank_rd_data_out_0_109 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21260 = _T_21259 | _T_21005; // @[Mux.scala 27:72]
  wire [1:0] _T_21006 = _T_21628 ? bht_bank_rd_data_out_0_110 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21261 = _T_21260 | _T_21006; // @[Mux.scala 27:72]
  wire [1:0] _T_21007 = _T_21630 ? bht_bank_rd_data_out_0_111 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21262 = _T_21261 | _T_21007; // @[Mux.scala 27:72]
  wire [1:0] _T_21008 = _T_21632 ? bht_bank_rd_data_out_0_112 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21263 = _T_21262 | _T_21008; // @[Mux.scala 27:72]
  wire [1:0] _T_21009 = _T_21634 ? bht_bank_rd_data_out_0_113 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21264 = _T_21263 | _T_21009; // @[Mux.scala 27:72]
  wire [1:0] _T_21010 = _T_21636 ? bht_bank_rd_data_out_0_114 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21265 = _T_21264 | _T_21010; // @[Mux.scala 27:72]
  wire [1:0] _T_21011 = _T_21638 ? bht_bank_rd_data_out_0_115 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21266 = _T_21265 | _T_21011; // @[Mux.scala 27:72]
  wire [1:0] _T_21012 = _T_21640 ? bht_bank_rd_data_out_0_116 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21267 = _T_21266 | _T_21012; // @[Mux.scala 27:72]
  wire [1:0] _T_21013 = _T_21642 ? bht_bank_rd_data_out_0_117 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21268 = _T_21267 | _T_21013; // @[Mux.scala 27:72]
  wire [1:0] _T_21014 = _T_21644 ? bht_bank_rd_data_out_0_118 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21269 = _T_21268 | _T_21014; // @[Mux.scala 27:72]
  wire [1:0] _T_21015 = _T_21646 ? bht_bank_rd_data_out_0_119 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21270 = _T_21269 | _T_21015; // @[Mux.scala 27:72]
  wire [1:0] _T_21016 = _T_21648 ? bht_bank_rd_data_out_0_120 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21271 = _T_21270 | _T_21016; // @[Mux.scala 27:72]
  wire [1:0] _T_21017 = _T_21650 ? bht_bank_rd_data_out_0_121 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21272 = _T_21271 | _T_21017; // @[Mux.scala 27:72]
  wire [1:0] _T_21018 = _T_21652 ? bht_bank_rd_data_out_0_122 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21273 = _T_21272 | _T_21018; // @[Mux.scala 27:72]
  wire [1:0] _T_21019 = _T_21654 ? bht_bank_rd_data_out_0_123 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21274 = _T_21273 | _T_21019; // @[Mux.scala 27:72]
  wire [1:0] _T_21020 = _T_21656 ? bht_bank_rd_data_out_0_124 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21275 = _T_21274 | _T_21020; // @[Mux.scala 27:72]
  wire [1:0] _T_21021 = _T_21658 ? bht_bank_rd_data_out_0_125 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21276 = _T_21275 | _T_21021; // @[Mux.scala 27:72]
  wire [1:0] _T_21022 = _T_21660 ? bht_bank_rd_data_out_0_126 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21277 = _T_21276 | _T_21022; // @[Mux.scala 27:72]
  wire [1:0] _T_21023 = _T_21662 ? bht_bank_rd_data_out_0_127 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21278 = _T_21277 | _T_21023; // @[Mux.scala 27:72]
  wire [1:0] _T_21024 = _T_21664 ? bht_bank_rd_data_out_0_128 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21279 = _T_21278 | _T_21024; // @[Mux.scala 27:72]
  wire [1:0] _T_21025 = _T_21666 ? bht_bank_rd_data_out_0_129 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21280 = _T_21279 | _T_21025; // @[Mux.scala 27:72]
  wire [1:0] _T_21026 = _T_21668 ? bht_bank_rd_data_out_0_130 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21281 = _T_21280 | _T_21026; // @[Mux.scala 27:72]
  wire [1:0] _T_21027 = _T_21670 ? bht_bank_rd_data_out_0_131 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21282 = _T_21281 | _T_21027; // @[Mux.scala 27:72]
  wire [1:0] _T_21028 = _T_21672 ? bht_bank_rd_data_out_0_132 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21283 = _T_21282 | _T_21028; // @[Mux.scala 27:72]
  wire [1:0] _T_21029 = _T_21674 ? bht_bank_rd_data_out_0_133 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21284 = _T_21283 | _T_21029; // @[Mux.scala 27:72]
  wire [1:0] _T_21030 = _T_21676 ? bht_bank_rd_data_out_0_134 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21285 = _T_21284 | _T_21030; // @[Mux.scala 27:72]
  wire [1:0] _T_21031 = _T_21678 ? bht_bank_rd_data_out_0_135 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21286 = _T_21285 | _T_21031; // @[Mux.scala 27:72]
  wire [1:0] _T_21032 = _T_21680 ? bht_bank_rd_data_out_0_136 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21287 = _T_21286 | _T_21032; // @[Mux.scala 27:72]
  wire [1:0] _T_21033 = _T_21682 ? bht_bank_rd_data_out_0_137 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21288 = _T_21287 | _T_21033; // @[Mux.scala 27:72]
  wire [1:0] _T_21034 = _T_21684 ? bht_bank_rd_data_out_0_138 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21289 = _T_21288 | _T_21034; // @[Mux.scala 27:72]
  wire [1:0] _T_21035 = _T_21686 ? bht_bank_rd_data_out_0_139 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21290 = _T_21289 | _T_21035; // @[Mux.scala 27:72]
  wire [1:0] _T_21036 = _T_21688 ? bht_bank_rd_data_out_0_140 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21291 = _T_21290 | _T_21036; // @[Mux.scala 27:72]
  wire [1:0] _T_21037 = _T_21690 ? bht_bank_rd_data_out_0_141 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21292 = _T_21291 | _T_21037; // @[Mux.scala 27:72]
  wire [1:0] _T_21038 = _T_21692 ? bht_bank_rd_data_out_0_142 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21293 = _T_21292 | _T_21038; // @[Mux.scala 27:72]
  wire [1:0] _T_21039 = _T_21694 ? bht_bank_rd_data_out_0_143 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21294 = _T_21293 | _T_21039; // @[Mux.scala 27:72]
  wire [1:0] _T_21040 = _T_21696 ? bht_bank_rd_data_out_0_144 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21295 = _T_21294 | _T_21040; // @[Mux.scala 27:72]
  wire [1:0] _T_21041 = _T_21698 ? bht_bank_rd_data_out_0_145 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21296 = _T_21295 | _T_21041; // @[Mux.scala 27:72]
  wire [1:0] _T_21042 = _T_21700 ? bht_bank_rd_data_out_0_146 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21297 = _T_21296 | _T_21042; // @[Mux.scala 27:72]
  wire [1:0] _T_21043 = _T_21702 ? bht_bank_rd_data_out_0_147 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21298 = _T_21297 | _T_21043; // @[Mux.scala 27:72]
  wire [1:0] _T_21044 = _T_21704 ? bht_bank_rd_data_out_0_148 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21299 = _T_21298 | _T_21044; // @[Mux.scala 27:72]
  wire [1:0] _T_21045 = _T_21706 ? bht_bank_rd_data_out_0_149 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21300 = _T_21299 | _T_21045; // @[Mux.scala 27:72]
  wire [1:0] _T_21046 = _T_21708 ? bht_bank_rd_data_out_0_150 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21301 = _T_21300 | _T_21046; // @[Mux.scala 27:72]
  wire [1:0] _T_21047 = _T_21710 ? bht_bank_rd_data_out_0_151 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21302 = _T_21301 | _T_21047; // @[Mux.scala 27:72]
  wire [1:0] _T_21048 = _T_21712 ? bht_bank_rd_data_out_0_152 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21303 = _T_21302 | _T_21048; // @[Mux.scala 27:72]
  wire [1:0] _T_21049 = _T_21714 ? bht_bank_rd_data_out_0_153 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21304 = _T_21303 | _T_21049; // @[Mux.scala 27:72]
  wire [1:0] _T_21050 = _T_21716 ? bht_bank_rd_data_out_0_154 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21305 = _T_21304 | _T_21050; // @[Mux.scala 27:72]
  wire [1:0] _T_21051 = _T_21718 ? bht_bank_rd_data_out_0_155 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21306 = _T_21305 | _T_21051; // @[Mux.scala 27:72]
  wire [1:0] _T_21052 = _T_21720 ? bht_bank_rd_data_out_0_156 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21307 = _T_21306 | _T_21052; // @[Mux.scala 27:72]
  wire [1:0] _T_21053 = _T_21722 ? bht_bank_rd_data_out_0_157 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21308 = _T_21307 | _T_21053; // @[Mux.scala 27:72]
  wire [1:0] _T_21054 = _T_21724 ? bht_bank_rd_data_out_0_158 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21309 = _T_21308 | _T_21054; // @[Mux.scala 27:72]
  wire [1:0] _T_21055 = _T_21726 ? bht_bank_rd_data_out_0_159 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21310 = _T_21309 | _T_21055; // @[Mux.scala 27:72]
  wire [1:0] _T_21056 = _T_21728 ? bht_bank_rd_data_out_0_160 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21311 = _T_21310 | _T_21056; // @[Mux.scala 27:72]
  wire [1:0] _T_21057 = _T_21730 ? bht_bank_rd_data_out_0_161 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21312 = _T_21311 | _T_21057; // @[Mux.scala 27:72]
  wire [1:0] _T_21058 = _T_21732 ? bht_bank_rd_data_out_0_162 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21313 = _T_21312 | _T_21058; // @[Mux.scala 27:72]
  wire [1:0] _T_21059 = _T_21734 ? bht_bank_rd_data_out_0_163 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21314 = _T_21313 | _T_21059; // @[Mux.scala 27:72]
  wire [1:0] _T_21060 = _T_21736 ? bht_bank_rd_data_out_0_164 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21315 = _T_21314 | _T_21060; // @[Mux.scala 27:72]
  wire [1:0] _T_21061 = _T_21738 ? bht_bank_rd_data_out_0_165 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21316 = _T_21315 | _T_21061; // @[Mux.scala 27:72]
  wire [1:0] _T_21062 = _T_21740 ? bht_bank_rd_data_out_0_166 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21317 = _T_21316 | _T_21062; // @[Mux.scala 27:72]
  wire [1:0] _T_21063 = _T_21742 ? bht_bank_rd_data_out_0_167 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21318 = _T_21317 | _T_21063; // @[Mux.scala 27:72]
  wire [1:0] _T_21064 = _T_21744 ? bht_bank_rd_data_out_0_168 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21319 = _T_21318 | _T_21064; // @[Mux.scala 27:72]
  wire [1:0] _T_21065 = _T_21746 ? bht_bank_rd_data_out_0_169 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21320 = _T_21319 | _T_21065; // @[Mux.scala 27:72]
  wire [1:0] _T_21066 = _T_21748 ? bht_bank_rd_data_out_0_170 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21321 = _T_21320 | _T_21066; // @[Mux.scala 27:72]
  wire [1:0] _T_21067 = _T_21750 ? bht_bank_rd_data_out_0_171 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21322 = _T_21321 | _T_21067; // @[Mux.scala 27:72]
  wire [1:0] _T_21068 = _T_21752 ? bht_bank_rd_data_out_0_172 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21323 = _T_21322 | _T_21068; // @[Mux.scala 27:72]
  wire [1:0] _T_21069 = _T_21754 ? bht_bank_rd_data_out_0_173 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21324 = _T_21323 | _T_21069; // @[Mux.scala 27:72]
  wire [1:0] _T_21070 = _T_21756 ? bht_bank_rd_data_out_0_174 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21325 = _T_21324 | _T_21070; // @[Mux.scala 27:72]
  wire [1:0] _T_21071 = _T_21758 ? bht_bank_rd_data_out_0_175 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21326 = _T_21325 | _T_21071; // @[Mux.scala 27:72]
  wire [1:0] _T_21072 = _T_21760 ? bht_bank_rd_data_out_0_176 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21327 = _T_21326 | _T_21072; // @[Mux.scala 27:72]
  wire [1:0] _T_21073 = _T_21762 ? bht_bank_rd_data_out_0_177 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21328 = _T_21327 | _T_21073; // @[Mux.scala 27:72]
  wire [1:0] _T_21074 = _T_21764 ? bht_bank_rd_data_out_0_178 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21329 = _T_21328 | _T_21074; // @[Mux.scala 27:72]
  wire [1:0] _T_21075 = _T_21766 ? bht_bank_rd_data_out_0_179 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21330 = _T_21329 | _T_21075; // @[Mux.scala 27:72]
  wire [1:0] _T_21076 = _T_21768 ? bht_bank_rd_data_out_0_180 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21331 = _T_21330 | _T_21076; // @[Mux.scala 27:72]
  wire [1:0] _T_21077 = _T_21770 ? bht_bank_rd_data_out_0_181 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21332 = _T_21331 | _T_21077; // @[Mux.scala 27:72]
  wire [1:0] _T_21078 = _T_21772 ? bht_bank_rd_data_out_0_182 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21333 = _T_21332 | _T_21078; // @[Mux.scala 27:72]
  wire [1:0] _T_21079 = _T_21774 ? bht_bank_rd_data_out_0_183 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21334 = _T_21333 | _T_21079; // @[Mux.scala 27:72]
  wire [1:0] _T_21080 = _T_21776 ? bht_bank_rd_data_out_0_184 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21335 = _T_21334 | _T_21080; // @[Mux.scala 27:72]
  wire [1:0] _T_21081 = _T_21778 ? bht_bank_rd_data_out_0_185 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21336 = _T_21335 | _T_21081; // @[Mux.scala 27:72]
  wire [1:0] _T_21082 = _T_21780 ? bht_bank_rd_data_out_0_186 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21337 = _T_21336 | _T_21082; // @[Mux.scala 27:72]
  wire [1:0] _T_21083 = _T_21782 ? bht_bank_rd_data_out_0_187 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21338 = _T_21337 | _T_21083; // @[Mux.scala 27:72]
  wire [1:0] _T_21084 = _T_21784 ? bht_bank_rd_data_out_0_188 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21339 = _T_21338 | _T_21084; // @[Mux.scala 27:72]
  wire [1:0] _T_21085 = _T_21786 ? bht_bank_rd_data_out_0_189 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21340 = _T_21339 | _T_21085; // @[Mux.scala 27:72]
  wire [1:0] _T_21086 = _T_21788 ? bht_bank_rd_data_out_0_190 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21341 = _T_21340 | _T_21086; // @[Mux.scala 27:72]
  wire [1:0] _T_21087 = _T_21790 ? bht_bank_rd_data_out_0_191 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21342 = _T_21341 | _T_21087; // @[Mux.scala 27:72]
  wire [1:0] _T_21088 = _T_21792 ? bht_bank_rd_data_out_0_192 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21343 = _T_21342 | _T_21088; // @[Mux.scala 27:72]
  wire [1:0] _T_21089 = _T_21794 ? bht_bank_rd_data_out_0_193 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21344 = _T_21343 | _T_21089; // @[Mux.scala 27:72]
  wire [1:0] _T_21090 = _T_21796 ? bht_bank_rd_data_out_0_194 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21345 = _T_21344 | _T_21090; // @[Mux.scala 27:72]
  wire [1:0] _T_21091 = _T_21798 ? bht_bank_rd_data_out_0_195 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21346 = _T_21345 | _T_21091; // @[Mux.scala 27:72]
  wire [1:0] _T_21092 = _T_21800 ? bht_bank_rd_data_out_0_196 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21347 = _T_21346 | _T_21092; // @[Mux.scala 27:72]
  wire [1:0] _T_21093 = _T_21802 ? bht_bank_rd_data_out_0_197 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21348 = _T_21347 | _T_21093; // @[Mux.scala 27:72]
  wire [1:0] _T_21094 = _T_21804 ? bht_bank_rd_data_out_0_198 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21349 = _T_21348 | _T_21094; // @[Mux.scala 27:72]
  wire [1:0] _T_21095 = _T_21806 ? bht_bank_rd_data_out_0_199 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21350 = _T_21349 | _T_21095; // @[Mux.scala 27:72]
  wire [1:0] _T_21096 = _T_21808 ? bht_bank_rd_data_out_0_200 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21351 = _T_21350 | _T_21096; // @[Mux.scala 27:72]
  wire [1:0] _T_21097 = _T_21810 ? bht_bank_rd_data_out_0_201 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21352 = _T_21351 | _T_21097; // @[Mux.scala 27:72]
  wire [1:0] _T_21098 = _T_21812 ? bht_bank_rd_data_out_0_202 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21353 = _T_21352 | _T_21098; // @[Mux.scala 27:72]
  wire [1:0] _T_21099 = _T_21814 ? bht_bank_rd_data_out_0_203 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21354 = _T_21353 | _T_21099; // @[Mux.scala 27:72]
  wire [1:0] _T_21100 = _T_21816 ? bht_bank_rd_data_out_0_204 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21355 = _T_21354 | _T_21100; // @[Mux.scala 27:72]
  wire [1:0] _T_21101 = _T_21818 ? bht_bank_rd_data_out_0_205 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21356 = _T_21355 | _T_21101; // @[Mux.scala 27:72]
  wire [1:0] _T_21102 = _T_21820 ? bht_bank_rd_data_out_0_206 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21357 = _T_21356 | _T_21102; // @[Mux.scala 27:72]
  wire [1:0] _T_21103 = _T_21822 ? bht_bank_rd_data_out_0_207 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21358 = _T_21357 | _T_21103; // @[Mux.scala 27:72]
  wire [1:0] _T_21104 = _T_21824 ? bht_bank_rd_data_out_0_208 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21359 = _T_21358 | _T_21104; // @[Mux.scala 27:72]
  wire [1:0] _T_21105 = _T_21826 ? bht_bank_rd_data_out_0_209 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21360 = _T_21359 | _T_21105; // @[Mux.scala 27:72]
  wire [1:0] _T_21106 = _T_21828 ? bht_bank_rd_data_out_0_210 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21361 = _T_21360 | _T_21106; // @[Mux.scala 27:72]
  wire [1:0] _T_21107 = _T_21830 ? bht_bank_rd_data_out_0_211 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21362 = _T_21361 | _T_21107; // @[Mux.scala 27:72]
  wire [1:0] _T_21108 = _T_21832 ? bht_bank_rd_data_out_0_212 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21363 = _T_21362 | _T_21108; // @[Mux.scala 27:72]
  wire [1:0] _T_21109 = _T_21834 ? bht_bank_rd_data_out_0_213 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21364 = _T_21363 | _T_21109; // @[Mux.scala 27:72]
  wire [1:0] _T_21110 = _T_21836 ? bht_bank_rd_data_out_0_214 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21365 = _T_21364 | _T_21110; // @[Mux.scala 27:72]
  wire [1:0] _T_21111 = _T_21838 ? bht_bank_rd_data_out_0_215 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21366 = _T_21365 | _T_21111; // @[Mux.scala 27:72]
  wire [1:0] _T_21112 = _T_21840 ? bht_bank_rd_data_out_0_216 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21367 = _T_21366 | _T_21112; // @[Mux.scala 27:72]
  wire [1:0] _T_21113 = _T_21842 ? bht_bank_rd_data_out_0_217 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21368 = _T_21367 | _T_21113; // @[Mux.scala 27:72]
  wire [1:0] _T_21114 = _T_21844 ? bht_bank_rd_data_out_0_218 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21369 = _T_21368 | _T_21114; // @[Mux.scala 27:72]
  wire [1:0] _T_21115 = _T_21846 ? bht_bank_rd_data_out_0_219 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21370 = _T_21369 | _T_21115; // @[Mux.scala 27:72]
  wire [1:0] _T_21116 = _T_21848 ? bht_bank_rd_data_out_0_220 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21371 = _T_21370 | _T_21116; // @[Mux.scala 27:72]
  wire [1:0] _T_21117 = _T_21850 ? bht_bank_rd_data_out_0_221 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21372 = _T_21371 | _T_21117; // @[Mux.scala 27:72]
  wire [1:0] _T_21118 = _T_21852 ? bht_bank_rd_data_out_0_222 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21373 = _T_21372 | _T_21118; // @[Mux.scala 27:72]
  wire [1:0] _T_21119 = _T_21854 ? bht_bank_rd_data_out_0_223 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21374 = _T_21373 | _T_21119; // @[Mux.scala 27:72]
  wire [1:0] _T_21120 = _T_21856 ? bht_bank_rd_data_out_0_224 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21375 = _T_21374 | _T_21120; // @[Mux.scala 27:72]
  wire [1:0] _T_21121 = _T_21858 ? bht_bank_rd_data_out_0_225 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21376 = _T_21375 | _T_21121; // @[Mux.scala 27:72]
  wire [1:0] _T_21122 = _T_21860 ? bht_bank_rd_data_out_0_226 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21377 = _T_21376 | _T_21122; // @[Mux.scala 27:72]
  wire [1:0] _T_21123 = _T_21862 ? bht_bank_rd_data_out_0_227 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21378 = _T_21377 | _T_21123; // @[Mux.scala 27:72]
  wire [1:0] _T_21124 = _T_21864 ? bht_bank_rd_data_out_0_228 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21379 = _T_21378 | _T_21124; // @[Mux.scala 27:72]
  wire [1:0] _T_21125 = _T_21866 ? bht_bank_rd_data_out_0_229 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21380 = _T_21379 | _T_21125; // @[Mux.scala 27:72]
  wire [1:0] _T_21126 = _T_21868 ? bht_bank_rd_data_out_0_230 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21381 = _T_21380 | _T_21126; // @[Mux.scala 27:72]
  wire [1:0] _T_21127 = _T_21870 ? bht_bank_rd_data_out_0_231 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21382 = _T_21381 | _T_21127; // @[Mux.scala 27:72]
  wire [1:0] _T_21128 = _T_21872 ? bht_bank_rd_data_out_0_232 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21383 = _T_21382 | _T_21128; // @[Mux.scala 27:72]
  wire [1:0] _T_21129 = _T_21874 ? bht_bank_rd_data_out_0_233 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21384 = _T_21383 | _T_21129; // @[Mux.scala 27:72]
  wire [1:0] _T_21130 = _T_21876 ? bht_bank_rd_data_out_0_234 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21385 = _T_21384 | _T_21130; // @[Mux.scala 27:72]
  wire [1:0] _T_21131 = _T_21878 ? bht_bank_rd_data_out_0_235 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21386 = _T_21385 | _T_21131; // @[Mux.scala 27:72]
  wire [1:0] _T_21132 = _T_21880 ? bht_bank_rd_data_out_0_236 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21387 = _T_21386 | _T_21132; // @[Mux.scala 27:72]
  wire [1:0] _T_21133 = _T_21882 ? bht_bank_rd_data_out_0_237 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21388 = _T_21387 | _T_21133; // @[Mux.scala 27:72]
  wire [1:0] _T_21134 = _T_21884 ? bht_bank_rd_data_out_0_238 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21389 = _T_21388 | _T_21134; // @[Mux.scala 27:72]
  wire [1:0] _T_21135 = _T_21886 ? bht_bank_rd_data_out_0_239 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21390 = _T_21389 | _T_21135; // @[Mux.scala 27:72]
  wire [1:0] _T_21136 = _T_21888 ? bht_bank_rd_data_out_0_240 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21391 = _T_21390 | _T_21136; // @[Mux.scala 27:72]
  wire [1:0] _T_21137 = _T_21890 ? bht_bank_rd_data_out_0_241 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21392 = _T_21391 | _T_21137; // @[Mux.scala 27:72]
  wire [1:0] _T_21138 = _T_21892 ? bht_bank_rd_data_out_0_242 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21393 = _T_21392 | _T_21138; // @[Mux.scala 27:72]
  wire [1:0] _T_21139 = _T_21894 ? bht_bank_rd_data_out_0_243 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21394 = _T_21393 | _T_21139; // @[Mux.scala 27:72]
  wire [1:0] _T_21140 = _T_21896 ? bht_bank_rd_data_out_0_244 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21395 = _T_21394 | _T_21140; // @[Mux.scala 27:72]
  wire [1:0] _T_21141 = _T_21898 ? bht_bank_rd_data_out_0_245 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21396 = _T_21395 | _T_21141; // @[Mux.scala 27:72]
  wire [1:0] _T_21142 = _T_21900 ? bht_bank_rd_data_out_0_246 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21397 = _T_21396 | _T_21142; // @[Mux.scala 27:72]
  wire [1:0] _T_21143 = _T_21902 ? bht_bank_rd_data_out_0_247 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21398 = _T_21397 | _T_21143; // @[Mux.scala 27:72]
  wire [1:0] _T_21144 = _T_21904 ? bht_bank_rd_data_out_0_248 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21399 = _T_21398 | _T_21144; // @[Mux.scala 27:72]
  wire [1:0] _T_21145 = _T_21906 ? bht_bank_rd_data_out_0_249 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21400 = _T_21399 | _T_21145; // @[Mux.scala 27:72]
  wire [1:0] _T_21146 = _T_21908 ? bht_bank_rd_data_out_0_250 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21401 = _T_21400 | _T_21146; // @[Mux.scala 27:72]
  wire [1:0] _T_21147 = _T_21910 ? bht_bank_rd_data_out_0_251 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21402 = _T_21401 | _T_21147; // @[Mux.scala 27:72]
  wire [1:0] _T_21148 = _T_21912 ? bht_bank_rd_data_out_0_252 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21403 = _T_21402 | _T_21148; // @[Mux.scala 27:72]
  wire [1:0] _T_21149 = _T_21914 ? bht_bank_rd_data_out_0_253 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21404 = _T_21403 | _T_21149; // @[Mux.scala 27:72]
  wire [1:0] _T_21150 = _T_21916 ? bht_bank_rd_data_out_0_254 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21405 = _T_21404 | _T_21150; // @[Mux.scala 27:72]
  wire [1:0] _T_21151 = _T_21918 ? bht_bank_rd_data_out_0_255 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] bht_bank0_rd_data_f = _T_21405 | _T_21151; // @[Mux.scala 27:72]
  wire [1:0] _T_252 = _T_144 ? bht_bank0_rd_data_f : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_253 = io_ifc_fetch_addr_f[0] ? bht_bank1_rd_data_f : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] bht_vbank0_rd_data_f = _T_252 | _T_253; // @[Mux.scala 27:72]
  wire  _T_270 = bht_force_taken_f[0] | bht_vbank0_rd_data_f[1]; // @[ifu_bp_ctl.scala 282:45]
  wire  _T_272 = _T_270 & bht_valid_f[0]; // @[ifu_bp_ctl.scala 282:72]
  wire [1:0] bht_dir_f = {_T_267,_T_272}; // @[Cat.scala 29:58]
  wire  _T_14 = ~bht_dir_f[0]; // @[ifu_bp_ctl.scala 96:23]
  wire [1:0] btb_sel_f = {_T_14,bht_dir_f[0]}; // @[Cat.scala 29:58]
  wire [1:0] fetch_start_f = {io_ifc_fetch_addr_f[0],_T_144}; // @[Cat.scala 29:58]
  wire  _T_32 = io_exu_bp_exu_mp_btag == fetch_rd_tag_f; // @[ifu_bp_ctl.scala 114:53]
  wire  _T_33 = _T_32 & exu_mp_valid; // @[ifu_bp_ctl.scala 114:73]
  wire  _T_34 = _T_33 & io_ifc_fetch_req_f; // @[ifu_bp_ctl.scala 114:88]
  wire  _T_35 = io_exu_bp_exu_mp_index == btb_rd_addr_f; // @[ifu_bp_ctl.scala 114:124]
  wire  fetch_mp_collision_f = _T_34 & _T_35; // @[ifu_bp_ctl.scala 114:109]
  wire  _T_36 = io_exu_bp_exu_mp_btag == fetch_rd_tag_p1_f; // @[ifu_bp_ctl.scala 115:56]
  wire  _T_37 = _T_36 & exu_mp_valid; // @[ifu_bp_ctl.scala 115:79]
  wire  _T_38 = _T_37 & io_ifc_fetch_req_f; // @[ifu_bp_ctl.scala 115:94]
  wire  _T_39 = io_exu_bp_exu_mp_index == btb_rd_addr_p1_f; // @[ifu_bp_ctl.scala 115:130]
  wire  fetch_mp_collision_p1_f = _T_38 & _T_39; // @[ifu_bp_ctl.scala 115:115]
  reg  exu_mp_way_f; // @[ifu_bp_ctl.scala 119:55]
  reg  exu_flush_final_d1; // @[ifu_bp_ctl.scala 120:61]
  wire [255:0] mp_wrindex_dec = 256'h1 << io_exu_bp_exu_mp_index; // @[ifu_bp_ctl.scala 191:28]
  wire [255:0] fetch_wrindex_dec = 256'h1 << btb_rd_addr_f; // @[ifu_bp_ctl.scala 194:31]
  wire [255:0] fetch_wrindex_p1_dec = 256'h1 << btb_rd_addr_p1_f; // @[ifu_bp_ctl.scala 197:34]
  wire [255:0] _T_150 = exu_mp_valid ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12]
  wire [255:0] mp_wrlru_b0 = mp_wrindex_dec & _T_150; // @[ifu_bp_ctl.scala 200:36]
  wire  _T_166 = bht_valid_f[0] | bht_valid_f[1]; // @[ifu_bp_ctl.scala 206:42]
  wire  _T_167 = _T_166 & io_ifc_fetch_req_f; // @[ifu_bp_ctl.scala 206:58]
  wire  lru_update_valid_f = _T_167 & _T; // @[ifu_bp_ctl.scala 206:79]
  wire [255:0] _T_170 = lru_update_valid_f ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12]
  wire [255:0] fetch_wrlru_b0 = fetch_wrindex_dec & _T_170; // @[ifu_bp_ctl.scala 208:42]
  wire [255:0] fetch_wrlru_p1_b0 = fetch_wrindex_p1_dec & _T_170; // @[ifu_bp_ctl.scala 209:48]
  wire [255:0] _T_173 = ~mp_wrlru_b0; // @[ifu_bp_ctl.scala 211:25]
  wire [255:0] _T_174 = ~fetch_wrlru_b0; // @[ifu_bp_ctl.scala 211:40]
  wire [255:0] btb_lru_b0_hold = _T_173 & _T_174; // @[ifu_bp_ctl.scala 211:38]
  wire  _T_176 = ~io_exu_bp_exu_mp_pkt_bits_way; // @[ifu_bp_ctl.scala 218:40]
  wire [255:0] _T_179 = _T_176 ? mp_wrlru_b0 : 256'h0; // @[Mux.scala 27:72]
  wire [255:0] _T_180 = tag_match_way0_f ? fetch_wrlru_b0 : 256'h0; // @[Mux.scala 27:72]
  wire [255:0] _T_181 = tag_match_way0_p1_f ? fetch_wrlru_p1_b0 : 256'h0; // @[Mux.scala 27:72]
  wire [255:0] _T_182 = _T_179 | _T_180; // @[Mux.scala 27:72]
  wire [255:0] _T_183 = _T_182 | _T_181; // @[Mux.scala 27:72]
  reg [255:0] btb_lru_b0_f; // @[lib.scala 374:16]
  wire [255:0] _T_185 = btb_lru_b0_hold & btb_lru_b0_f; // @[ifu_bp_ctl.scala 220:102]
  wire [255:0] _T_187 = fetch_wrindex_dec & btb_lru_b0_f; // @[ifu_bp_ctl.scala 223:78]
  wire  _T_188 = |_T_187; // @[ifu_bp_ctl.scala 223:94]
  wire  btb_lru_rd_f = fetch_mp_collision_f ? exu_mp_way_f : _T_188; // @[ifu_bp_ctl.scala 223:25]
  wire [255:0] _T_190 = fetch_wrindex_p1_dec & btb_lru_b0_f; // @[ifu_bp_ctl.scala 225:87]
  wire  _T_191 = |_T_190; // @[ifu_bp_ctl.scala 225:103]
  wire  btb_lru_rd_p1_f = fetch_mp_collision_p1_f ? exu_mp_way_f : _T_191; // @[ifu_bp_ctl.scala 225:28]
  wire [1:0] _T_194 = {btb_lru_rd_f,btb_lru_rd_f}; // @[Cat.scala 29:58]
  wire [1:0] _T_197 = {btb_lru_rd_p1_f,btb_lru_rd_f}; // @[Cat.scala 29:58]
  wire [1:0] _T_198 = _T_144 ? _T_194 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_199 = io_ifc_fetch_addr_f[0] ? _T_197 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] btb_vlru_rd_f = _T_198 | _T_199; // @[Mux.scala 27:72]
  wire [1:0] _T_208 = {tag_match_way1_expanded_p1_f[0],tag_match_way1_expanded_f[1]}; // @[Cat.scala 29:58]
  wire [1:0] _T_209 = _T_144 ? tag_match_way1_expanded_f : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_210 = io_ifc_fetch_addr_f[0] ? _T_208 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] tag_match_vway1_expanded_f = _T_209 | _T_210; // @[Mux.scala 27:72]
  wire [1:0] _T_212 = ~bht_valid_f; // @[ifu_bp_ctl.scala 235:52]
  wire [1:0] _T_213 = _T_212 & btb_vlru_rd_f; // @[ifu_bp_ctl.scala 235:63]
  wire [15:0] _T_230 = btb_sel_f[1] ? btb_vbank1_rd_data_f[16:1] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_231 = btb_sel_f[0] ? btb_vbank0_rd_data_f[16:1] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] btb_sel_data_f = _T_230 | _T_231; // @[Mux.scala 27:72]
  wire [11:0] btb_rd_tgt_f = btb_sel_data_f[15:4]; // @[ifu_bp_ctl.scala 251:36]
  wire  btb_rd_pc4_f = btb_sel_data_f[3]; // @[ifu_bp_ctl.scala 252:36]
  wire  btb_rd_call_f = btb_sel_data_f[1]; // @[ifu_bp_ctl.scala 253:37]
  wire  btb_rd_ret_f = btb_sel_data_f[0]; // @[ifu_bp_ctl.scala 254:36]
  wire [1:0] _T_280 = {bht_vbank1_rd_data_f[1],bht_vbank0_rd_data_f[1]}; // @[Cat.scala 29:58]
  wire [1:0] hist1_raw = bht_force_taken_f | _T_280; // @[ifu_bp_ctl.scala 288:34]
  wire [1:0] _T_234 = bht_valid_f & hist1_raw; // @[ifu_bp_ctl.scala 261:39]
  wire  _T_235 = |_T_234; // @[ifu_bp_ctl.scala 261:52]
  wire  _T_236 = _T_235 & io_ifc_fetch_req_f; // @[ifu_bp_ctl.scala 261:56]
  wire  _T_237 = ~leak_one_f_d1; // @[ifu_bp_ctl.scala 261:79]
  wire  _T_238 = _T_236 & _T_237; // @[ifu_bp_ctl.scala 261:77]
  wire  _T_239 = ~io_dec_bp_dec_tlu_bpred_disable; // @[ifu_bp_ctl.scala 261:96]
  wire  _T_275 = io_ifu_bp_hit_taken_f & btb_sel_f[1]; // @[ifu_bp_ctl.scala 285:51]
  wire  _T_276 = ~io_ifu_bp_hit_taken_f; // @[ifu_bp_ctl.scala 285:69]
  wire  _T_286 = bht_valid_f[1] & btb_vbank1_rd_data_f[4]; // @[ifu_bp_ctl.scala 294:34]
  wire  _T_289 = bht_valid_f[0] & btb_vbank0_rd_data_f[4]; // @[ifu_bp_ctl.scala 295:34]
  wire  _T_292 = ~btb_vbank1_rd_data_f[2]; // @[ifu_bp_ctl.scala 298:37]
  wire  _T_293 = bht_valid_f[1] & _T_292; // @[ifu_bp_ctl.scala 298:35]
  wire  _T_295 = _T_293 & btb_vbank1_rd_data_f[1]; // @[ifu_bp_ctl.scala 298:65]
  wire  _T_298 = ~btb_vbank0_rd_data_f[2]; // @[ifu_bp_ctl.scala 299:37]
  wire  _T_299 = bht_valid_f[0] & _T_298; // @[ifu_bp_ctl.scala 299:35]
  wire  _T_301 = _T_299 & btb_vbank0_rd_data_f[1]; // @[ifu_bp_ctl.scala 299:65]
  wire [1:0] num_valids = bht_valid_f[1] + bht_valid_f[0]; // @[ifu_bp_ctl.scala 302:35]
  wire [1:0] _T_304 = btb_sel_f & bht_dir_f; // @[ifu_bp_ctl.scala 305:28]
  wire  final_h = |_T_304; // @[ifu_bp_ctl.scala 305:41]
  wire  _T_305 = num_valids == 2'h2; // @[ifu_bp_ctl.scala 309:41]
  wire [7:0] _T_309 = {fghr[5:0],1'h0,final_h}; // @[Cat.scala 29:58]
  wire  _T_310 = num_valids == 2'h1; // @[ifu_bp_ctl.scala 310:41]
  wire [7:0] _T_313 = {fghr[6:0],final_h}; // @[Cat.scala 29:58]
  wire  _T_314 = num_valids == 2'h0; // @[ifu_bp_ctl.scala 311:41]
  wire [7:0] _T_317 = _T_305 ? _T_309 : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_318 = _T_310 ? _T_313 : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_319 = _T_314 ? fghr : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_320 = _T_317 | _T_318; // @[Mux.scala 27:72]
  wire [7:0] merged_ghr = _T_320 | _T_319; // @[Mux.scala 27:72]
  wire  _T_323 = ~exu_flush_final_d1; // @[ifu_bp_ctl.scala 320:27]
  wire  _T_324 = _T_323 & io_ifc_fetch_req_f; // @[ifu_bp_ctl.scala 320:47]
  wire  _T_325 = _T_324 & io_ic_hit_f; // @[ifu_bp_ctl.scala 320:70]
  wire  _T_327 = _T_325 & _T_237; // @[ifu_bp_ctl.scala 320:84]
  wire  _T_330 = io_ifc_fetch_req_f & io_ic_hit_f; // @[ifu_bp_ctl.scala 321:70]
  wire  _T_332 = _T_330 & _T_237; // @[ifu_bp_ctl.scala 321:84]
  wire  _T_333 = ~_T_332; // @[ifu_bp_ctl.scala 321:49]
  wire  _T_334 = _T_323 & _T_333; // @[ifu_bp_ctl.scala 321:47]
  wire [7:0] _T_336 = exu_flush_final_d1 ? io_exu_bp_exu_mp_fghr : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_337 = _T_327 ? merged_ghr : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_338 = _T_334 ? fghr : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_339 = _T_336 | _T_337; // @[Mux.scala 27:72]
  wire [1:0] _T_344 = io_dec_bp_dec_tlu_bpred_disable ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [1:0] _T_345 = ~_T_344; // @[ifu_bp_ctl.scala 330:36]
  wire  _T_349 = ~fetch_start_f[0]; // @[ifu_bp_ctl.scala 334:36]
  wire  _T_350 = bht_dir_f[0] & _T_349; // @[ifu_bp_ctl.scala 334:34]
  wire  _T_354 = _T_14 & fetch_start_f[0]; // @[ifu_bp_ctl.scala 334:72]
  wire  _T_355 = _T_350 | _T_354; // @[ifu_bp_ctl.scala 334:55]
  wire  _T_358 = bht_dir_f[0] & fetch_start_f[0]; // @[ifu_bp_ctl.scala 335:34]
  wire  _T_363 = _T_14 & _T_349; // @[ifu_bp_ctl.scala 335:71]
  wire  _T_364 = _T_358 | _T_363; // @[ifu_bp_ctl.scala 335:54]
  wire [1:0] bloc_f = {_T_355,_T_364}; // @[Cat.scala 29:58]
  wire  _T_368 = _T_14 & io_ifc_fetch_addr_f[0]; // @[ifu_bp_ctl.scala 337:35]
  wire  _T_369 = ~btb_rd_pc4_f; // @[ifu_bp_ctl.scala 337:62]
  wire  use_fa_plus = _T_368 & _T_369; // @[ifu_bp_ctl.scala 337:60]
  wire  _T_372 = fetch_start_f[0] & btb_sel_f[0]; // @[ifu_bp_ctl.scala 339:44]
  wire  btb_fg_crossing_f = _T_372 & btb_rd_pc4_f; // @[ifu_bp_ctl.scala 339:59]
  wire  bp_total_branch_offset_f = bloc_f[1] ^ btb_rd_pc4_f; // @[ifu_bp_ctl.scala 340:43]
  wire  _T_376 = io_ifc_fetch_req_f & _T_276; // @[ifu_bp_ctl.scala 342:85]
  reg [29:0] ifc_fetch_adder_prior; // @[lib.scala 374:16]
  wire  _T_381 = ~btb_fg_crossing_f; // @[ifu_bp_ctl.scala 348:32]
  wire  _T_382 = ~use_fa_plus; // @[ifu_bp_ctl.scala 348:53]
  wire  _T_383 = _T_381 & _T_382; // @[ifu_bp_ctl.scala 348:51]
  wire [29:0] _T_386 = use_fa_plus ? fetch_addr_p1_f : 30'h0; // @[Mux.scala 27:72]
  wire [29:0] _T_387 = btb_fg_crossing_f ? ifc_fetch_adder_prior : 30'h0; // @[Mux.scala 27:72]
  wire [29:0] _T_388 = _T_383 ? io_ifc_fetch_addr_f[30:1] : 30'h0; // @[Mux.scala 27:72]
  wire [29:0] _T_389 = _T_386 | _T_387; // @[Mux.scala 27:72]
  wire [29:0] adder_pc_in_f = _T_389 | _T_388; // @[Mux.scala 27:72]
  wire [31:0] _T_393 = {adder_pc_in_f,bp_total_branch_offset_f,1'h0}; // @[Cat.scala 29:58]
  wire [12:0] _T_394 = {btb_rd_tgt_f,1'h0}; // @[Cat.scala 29:58]
  wire [12:0] _T_397 = _T_393[12:1] + _T_394[12:1]; // @[lib.scala 68:31]
  wire [18:0] _T_400 = _T_393[31:13] + 19'h1; // @[lib.scala 69:27]
  wire [18:0] _T_403 = _T_393[31:13] - 19'h1; // @[lib.scala 70:27]
  wire  _T_406 = ~_T_397[12]; // @[lib.scala 72:28]
  wire  _T_407 = _T_394[12] ^ _T_406; // @[lib.scala 72:26]
  wire  _T_410 = ~_T_394[12]; // @[lib.scala 73:20]
  wire  _T_412 = _T_410 & _T_397[12]; // @[lib.scala 73:26]
  wire  _T_416 = _T_394[12] & _T_406; // @[lib.scala 74:26]
  wire [18:0] _T_418 = _T_407 ? _T_393[31:13] : 19'h0; // @[Mux.scala 27:72]
  wire [18:0] _T_419 = _T_412 ? _T_400 : 19'h0; // @[Mux.scala 27:72]
  wire [18:0] _T_420 = _T_416 ? _T_403 : 19'h0; // @[Mux.scala 27:72]
  wire [18:0] _T_421 = _T_418 | _T_419; // @[Mux.scala 27:72]
  wire [18:0] _T_422 = _T_421 | _T_420; // @[Mux.scala 27:72]
  wire [31:0] bp_btb_target_adder_f = {_T_422,_T_397[11:0],1'h0}; // @[Cat.scala 29:58]
  wire  _T_426 = ~btb_rd_call_f; // @[ifu_bp_ctl.scala 357:49]
  wire  _T_427 = btb_rd_ret_f & _T_426; // @[ifu_bp_ctl.scala 357:47]
  reg [31:0] rets_out_0; // @[lib.scala 374:16]
  wire  _T_429 = _T_427 & rets_out_0[0]; // @[ifu_bp_ctl.scala 357:64]
  wire [12:0] _T_440 = {11'h0,_T_369,1'h0}; // @[Cat.scala 29:58]
  wire [12:0] _T_443 = _T_393[12:1] + _T_440[12:1]; // @[lib.scala 68:31]
  wire  _T_452 = ~_T_443[12]; // @[lib.scala 72:28]
  wire  _T_453 = _T_440[12] ^ _T_452; // @[lib.scala 72:26]
  wire  _T_456 = ~_T_440[12]; // @[lib.scala 73:20]
  wire  _T_458 = _T_456 & _T_443[12]; // @[lib.scala 73:26]
  wire  _T_462 = _T_440[12] & _T_452; // @[lib.scala 74:26]
  wire [18:0] _T_464 = _T_453 ? _T_393[31:13] : 19'h0; // @[Mux.scala 27:72]
  wire [18:0] _T_465 = _T_458 ? _T_400 : 19'h0; // @[Mux.scala 27:72]
  wire [18:0] _T_466 = _T_462 ? _T_403 : 19'h0; // @[Mux.scala 27:72]
  wire [18:0] _T_467 = _T_464 | _T_465; // @[Mux.scala 27:72]
  wire [18:0] _T_468 = _T_467 | _T_466; // @[Mux.scala 27:72]
  wire [31:0] bp_rs_call_target_f = {_T_468,_T_443[11:0],1'h0}; // @[Cat.scala 29:58]
  wire  _T_472 = ~btb_rd_ret_f; // @[ifu_bp_ctl.scala 363:33]
  wire  _T_473 = btb_rd_call_f & _T_472; // @[ifu_bp_ctl.scala 363:31]
  wire  rs_push = _T_473 & io_ifu_bp_hit_taken_f; // @[ifu_bp_ctl.scala 363:47]
  wire  rs_pop = _T_427 & io_ifu_bp_hit_taken_f; // @[ifu_bp_ctl.scala 364:46]
  wire  _T_476 = ~rs_push; // @[ifu_bp_ctl.scala 365:17]
  wire  _T_477 = ~rs_pop; // @[ifu_bp_ctl.scala 365:28]
  wire  rs_hold = _T_476 & _T_477; // @[ifu_bp_ctl.scala 365:26]
  wire [31:0] _T_480 = {bp_rs_call_target_f[31:1],1'h1}; // @[Cat.scala 29:58]
  wire [31:0] _T_482 = rs_push ? _T_480 : 32'h0; // @[Mux.scala 27:72]
  reg [31:0] rets_out_1; // @[lib.scala 374:16]
  wire [31:0] _T_483 = rs_pop ? rets_out_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_487 = rs_push ? rets_out_0 : 32'h0; // @[Mux.scala 27:72]
  reg [31:0] rets_out_2; // @[lib.scala 374:16]
  wire [31:0] _T_488 = rs_pop ? rets_out_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_492 = rs_push ? rets_out_1 : 32'h0; // @[Mux.scala 27:72]
  reg [31:0] rets_out_3; // @[lib.scala 374:16]
  wire [31:0] _T_493 = rs_pop ? rets_out_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_497 = rs_push ? rets_out_2 : 32'h0; // @[Mux.scala 27:72]
  reg [31:0] rets_out_4; // @[lib.scala 374:16]
  wire [31:0] _T_498 = rs_pop ? rets_out_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_502 = rs_push ? rets_out_3 : 32'h0; // @[Mux.scala 27:72]
  reg [31:0] rets_out_5; // @[lib.scala 374:16]
  wire [31:0] _T_503 = rs_pop ? rets_out_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_507 = rs_push ? rets_out_4 : 32'h0; // @[Mux.scala 27:72]
  reg [31:0] rets_out_6; // @[lib.scala 374:16]
  wire [31:0] _T_508 = rs_pop ? rets_out_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_512 = rs_push ? rets_out_5 : 32'h0; // @[Mux.scala 27:72]
  reg [31:0] rets_out_7; // @[lib.scala 374:16]
  wire [31:0] _T_513 = rs_pop ? rets_out_7 : 32'h0; // @[Mux.scala 27:72]
  wire  _T_531 = ~dec_tlu_error_wb; // @[ifu_bp_ctl.scala 380:35]
  wire  btb_valid = exu_mp_valid & _T_531; // @[ifu_bp_ctl.scala 380:32]
  wire  _T_532 = io_exu_bp_exu_mp_pkt_bits_pcall | io_exu_bp_exu_mp_pkt_bits_pja; // @[ifu_bp_ctl.scala 384:89]
  wire  _T_533 = io_exu_bp_exu_mp_pkt_bits_pret | io_exu_bp_exu_mp_pkt_bits_pja; // @[ifu_bp_ctl.scala 384:113]
  wire [2:0] _T_535 = {_T_532,_T_533,btb_valid}; // @[Cat.scala 29:58]
  wire [18:0] _T_538 = {io_exu_bp_exu_mp_btag,io_exu_bp_exu_mp_pkt_bits_toffset,io_exu_bp_exu_mp_pkt_bits_pc4,io_exu_bp_exu_mp_pkt_bits_boffset}; // @[Cat.scala 29:58]
  wire  exu_mp_valid_write = exu_mp_valid & io_exu_bp_exu_mp_pkt_bits_ataken; // @[ifu_bp_ctl.scala 385:41]
  wire  _T_540 = _T_176 & exu_mp_valid_write; // @[ifu_bp_ctl.scala 388:39]
  wire  _T_542 = _T_540 & _T_531; // @[ifu_bp_ctl.scala 388:60]
  wire  _T_543 = ~io_dec_bp_dec_tlu_br0_r_pkt_bits_way; // @[ifu_bp_ctl.scala 388:87]
  wire  _T_544 = _T_543 & dec_tlu_error_wb; // @[ifu_bp_ctl.scala 388:104]
  wire  btb_wr_en_way0 = _T_542 | _T_544; // @[ifu_bp_ctl.scala 388:83]
  wire  _T_545 = io_exu_bp_exu_mp_pkt_bits_way & exu_mp_valid_write; // @[ifu_bp_ctl.scala 389:36]
  wire  _T_547 = _T_545 & _T_531; // @[ifu_bp_ctl.scala 389:57]
  wire  _T_548 = io_dec_bp_dec_tlu_br0_r_pkt_bits_way & dec_tlu_error_wb; // @[ifu_bp_ctl.scala 389:98]
  wire  btb_wr_en_way1 = _T_547 | _T_548; // @[ifu_bp_ctl.scala 389:80]
  wire [7:0] btb_wr_addr = dec_tlu_error_wb ? io_exu_bp_exu_i0_br_index_r : io_exu_bp_exu_mp_index; // @[ifu_bp_ctl.scala 392:24]
  wire  middle_of_bank = io_exu_bp_exu_mp_pkt_bits_pc4 ^ io_exu_bp_exu_mp_pkt_bits_boffset; // @[ifu_bp_ctl.scala 393:35]
  wire  _T_550 = ~io_exu_bp_exu_mp_pkt_bits_pcall; // @[ifu_bp_ctl.scala 396:43]
  wire  _T_551 = exu_mp_valid & _T_550; // @[ifu_bp_ctl.scala 396:41]
  wire  _T_552 = ~io_exu_bp_exu_mp_pkt_bits_pret; // @[ifu_bp_ctl.scala 396:58]
  wire  _T_553 = _T_551 & _T_552; // @[ifu_bp_ctl.scala 396:56]
  wire  _T_554 = ~io_exu_bp_exu_mp_pkt_bits_pja; // @[ifu_bp_ctl.scala 396:72]
  wire  _T_555 = _T_553 & _T_554; // @[ifu_bp_ctl.scala 396:70]
  wire [1:0] _T_557 = _T_555 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire  _T_558 = ~middle_of_bank; // @[ifu_bp_ctl.scala 396:106]
  wire [1:0] _T_559 = {middle_of_bank,_T_558}; // @[Cat.scala 29:58]
  wire [1:0] bht_wr_en0 = _T_557 & _T_559; // @[ifu_bp_ctl.scala 396:84]
  wire [1:0] _T_561 = io_dec_bp_dec_tlu_br0_r_pkt_valid ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire  _T_562 = ~io_dec_bp_dec_tlu_br0_r_pkt_bits_middle; // @[ifu_bp_ctl.scala 397:75]
  wire [1:0] _T_563 = {io_dec_bp_dec_tlu_br0_r_pkt_bits_middle,_T_562}; // @[Cat.scala 29:58]
  wire [1:0] bht_wr_en2 = _T_561 & _T_563; // @[ifu_bp_ctl.scala 397:46]
  wire [9:0] _T_564 = {io_exu_bp_exu_mp_index,2'h0}; // @[Cat.scala 29:58]
  wire [7:0] bht_wr_addr0 = _T_564[9:2] ^ io_exu_bp_exu_mp_eghr; // @[lib.scala 56:35]
  wire [9:0] _T_567 = {io_exu_bp_exu_i0_br_index_r,2'h0}; // @[Cat.scala 29:58]
  wire [7:0] bht_wr_addr2 = _T_567[9:2] ^ io_exu_bp_exu_i0_br_fghr_r; // @[lib.scala 56:35]
  wire  _T_576 = btb_wr_addr == 8'h0; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_579 = btb_wr_addr == 8'h1; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_582 = btb_wr_addr == 8'h2; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_585 = btb_wr_addr == 8'h3; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_588 = btb_wr_addr == 8'h4; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_591 = btb_wr_addr == 8'h5; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_594 = btb_wr_addr == 8'h6; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_597 = btb_wr_addr == 8'h7; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_600 = btb_wr_addr == 8'h8; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_603 = btb_wr_addr == 8'h9; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_606 = btb_wr_addr == 8'ha; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_609 = btb_wr_addr == 8'hb; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_612 = btb_wr_addr == 8'hc; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_615 = btb_wr_addr == 8'hd; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_618 = btb_wr_addr == 8'he; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_621 = btb_wr_addr == 8'hf; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_624 = btb_wr_addr == 8'h10; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_627 = btb_wr_addr == 8'h11; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_630 = btb_wr_addr == 8'h12; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_633 = btb_wr_addr == 8'h13; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_636 = btb_wr_addr == 8'h14; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_639 = btb_wr_addr == 8'h15; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_642 = btb_wr_addr == 8'h16; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_645 = btb_wr_addr == 8'h17; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_648 = btb_wr_addr == 8'h18; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_651 = btb_wr_addr == 8'h19; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_654 = btb_wr_addr == 8'h1a; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_657 = btb_wr_addr == 8'h1b; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_660 = btb_wr_addr == 8'h1c; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_663 = btb_wr_addr == 8'h1d; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_666 = btb_wr_addr == 8'h1e; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_669 = btb_wr_addr == 8'h1f; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_672 = btb_wr_addr == 8'h20; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_675 = btb_wr_addr == 8'h21; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_678 = btb_wr_addr == 8'h22; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_681 = btb_wr_addr == 8'h23; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_684 = btb_wr_addr == 8'h24; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_687 = btb_wr_addr == 8'h25; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_690 = btb_wr_addr == 8'h26; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_693 = btb_wr_addr == 8'h27; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_696 = btb_wr_addr == 8'h28; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_699 = btb_wr_addr == 8'h29; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_702 = btb_wr_addr == 8'h2a; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_705 = btb_wr_addr == 8'h2b; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_708 = btb_wr_addr == 8'h2c; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_711 = btb_wr_addr == 8'h2d; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_714 = btb_wr_addr == 8'h2e; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_717 = btb_wr_addr == 8'h2f; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_720 = btb_wr_addr == 8'h30; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_723 = btb_wr_addr == 8'h31; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_726 = btb_wr_addr == 8'h32; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_729 = btb_wr_addr == 8'h33; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_732 = btb_wr_addr == 8'h34; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_735 = btb_wr_addr == 8'h35; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_738 = btb_wr_addr == 8'h36; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_741 = btb_wr_addr == 8'h37; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_744 = btb_wr_addr == 8'h38; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_747 = btb_wr_addr == 8'h39; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_750 = btb_wr_addr == 8'h3a; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_753 = btb_wr_addr == 8'h3b; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_756 = btb_wr_addr == 8'h3c; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_759 = btb_wr_addr == 8'h3d; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_762 = btb_wr_addr == 8'h3e; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_765 = btb_wr_addr == 8'h3f; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_768 = btb_wr_addr == 8'h40; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_771 = btb_wr_addr == 8'h41; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_774 = btb_wr_addr == 8'h42; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_777 = btb_wr_addr == 8'h43; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_780 = btb_wr_addr == 8'h44; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_783 = btb_wr_addr == 8'h45; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_786 = btb_wr_addr == 8'h46; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_789 = btb_wr_addr == 8'h47; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_792 = btb_wr_addr == 8'h48; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_795 = btb_wr_addr == 8'h49; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_798 = btb_wr_addr == 8'h4a; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_801 = btb_wr_addr == 8'h4b; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_804 = btb_wr_addr == 8'h4c; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_807 = btb_wr_addr == 8'h4d; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_810 = btb_wr_addr == 8'h4e; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_813 = btb_wr_addr == 8'h4f; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_816 = btb_wr_addr == 8'h50; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_819 = btb_wr_addr == 8'h51; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_822 = btb_wr_addr == 8'h52; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_825 = btb_wr_addr == 8'h53; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_828 = btb_wr_addr == 8'h54; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_831 = btb_wr_addr == 8'h55; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_834 = btb_wr_addr == 8'h56; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_837 = btb_wr_addr == 8'h57; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_840 = btb_wr_addr == 8'h58; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_843 = btb_wr_addr == 8'h59; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_846 = btb_wr_addr == 8'h5a; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_849 = btb_wr_addr == 8'h5b; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_852 = btb_wr_addr == 8'h5c; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_855 = btb_wr_addr == 8'h5d; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_858 = btb_wr_addr == 8'h5e; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_861 = btb_wr_addr == 8'h5f; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_864 = btb_wr_addr == 8'h60; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_867 = btb_wr_addr == 8'h61; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_870 = btb_wr_addr == 8'h62; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_873 = btb_wr_addr == 8'h63; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_876 = btb_wr_addr == 8'h64; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_879 = btb_wr_addr == 8'h65; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_882 = btb_wr_addr == 8'h66; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_885 = btb_wr_addr == 8'h67; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_888 = btb_wr_addr == 8'h68; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_891 = btb_wr_addr == 8'h69; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_894 = btb_wr_addr == 8'h6a; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_897 = btb_wr_addr == 8'h6b; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_900 = btb_wr_addr == 8'h6c; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_903 = btb_wr_addr == 8'h6d; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_906 = btb_wr_addr == 8'h6e; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_909 = btb_wr_addr == 8'h6f; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_912 = btb_wr_addr == 8'h70; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_915 = btb_wr_addr == 8'h71; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_918 = btb_wr_addr == 8'h72; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_921 = btb_wr_addr == 8'h73; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_924 = btb_wr_addr == 8'h74; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_927 = btb_wr_addr == 8'h75; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_930 = btb_wr_addr == 8'h76; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_933 = btb_wr_addr == 8'h77; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_936 = btb_wr_addr == 8'h78; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_939 = btb_wr_addr == 8'h79; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_942 = btb_wr_addr == 8'h7a; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_945 = btb_wr_addr == 8'h7b; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_948 = btb_wr_addr == 8'h7c; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_951 = btb_wr_addr == 8'h7d; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_954 = btb_wr_addr == 8'h7e; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_957 = btb_wr_addr == 8'h7f; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_960 = btb_wr_addr == 8'h80; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_963 = btb_wr_addr == 8'h81; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_966 = btb_wr_addr == 8'h82; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_969 = btb_wr_addr == 8'h83; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_972 = btb_wr_addr == 8'h84; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_975 = btb_wr_addr == 8'h85; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_978 = btb_wr_addr == 8'h86; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_981 = btb_wr_addr == 8'h87; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_984 = btb_wr_addr == 8'h88; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_987 = btb_wr_addr == 8'h89; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_990 = btb_wr_addr == 8'h8a; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_993 = btb_wr_addr == 8'h8b; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_996 = btb_wr_addr == 8'h8c; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_999 = btb_wr_addr == 8'h8d; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1002 = btb_wr_addr == 8'h8e; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1005 = btb_wr_addr == 8'h8f; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1008 = btb_wr_addr == 8'h90; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1011 = btb_wr_addr == 8'h91; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1014 = btb_wr_addr == 8'h92; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1017 = btb_wr_addr == 8'h93; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1020 = btb_wr_addr == 8'h94; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1023 = btb_wr_addr == 8'h95; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1026 = btb_wr_addr == 8'h96; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1029 = btb_wr_addr == 8'h97; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1032 = btb_wr_addr == 8'h98; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1035 = btb_wr_addr == 8'h99; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1038 = btb_wr_addr == 8'h9a; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1041 = btb_wr_addr == 8'h9b; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1044 = btb_wr_addr == 8'h9c; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1047 = btb_wr_addr == 8'h9d; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1050 = btb_wr_addr == 8'h9e; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1053 = btb_wr_addr == 8'h9f; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1056 = btb_wr_addr == 8'ha0; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1059 = btb_wr_addr == 8'ha1; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1062 = btb_wr_addr == 8'ha2; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1065 = btb_wr_addr == 8'ha3; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1068 = btb_wr_addr == 8'ha4; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1071 = btb_wr_addr == 8'ha5; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1074 = btb_wr_addr == 8'ha6; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1077 = btb_wr_addr == 8'ha7; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1080 = btb_wr_addr == 8'ha8; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1083 = btb_wr_addr == 8'ha9; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1086 = btb_wr_addr == 8'haa; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1089 = btb_wr_addr == 8'hab; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1092 = btb_wr_addr == 8'hac; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1095 = btb_wr_addr == 8'had; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1098 = btb_wr_addr == 8'hae; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1101 = btb_wr_addr == 8'haf; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1104 = btb_wr_addr == 8'hb0; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1107 = btb_wr_addr == 8'hb1; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1110 = btb_wr_addr == 8'hb2; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1113 = btb_wr_addr == 8'hb3; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1116 = btb_wr_addr == 8'hb4; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1119 = btb_wr_addr == 8'hb5; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1122 = btb_wr_addr == 8'hb6; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1125 = btb_wr_addr == 8'hb7; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1128 = btb_wr_addr == 8'hb8; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1131 = btb_wr_addr == 8'hb9; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1134 = btb_wr_addr == 8'hba; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1137 = btb_wr_addr == 8'hbb; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1140 = btb_wr_addr == 8'hbc; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1143 = btb_wr_addr == 8'hbd; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1146 = btb_wr_addr == 8'hbe; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1149 = btb_wr_addr == 8'hbf; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1152 = btb_wr_addr == 8'hc0; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1155 = btb_wr_addr == 8'hc1; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1158 = btb_wr_addr == 8'hc2; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1161 = btb_wr_addr == 8'hc3; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1164 = btb_wr_addr == 8'hc4; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1167 = btb_wr_addr == 8'hc5; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1170 = btb_wr_addr == 8'hc6; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1173 = btb_wr_addr == 8'hc7; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1176 = btb_wr_addr == 8'hc8; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1179 = btb_wr_addr == 8'hc9; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1182 = btb_wr_addr == 8'hca; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1185 = btb_wr_addr == 8'hcb; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1188 = btb_wr_addr == 8'hcc; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1191 = btb_wr_addr == 8'hcd; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1194 = btb_wr_addr == 8'hce; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1197 = btb_wr_addr == 8'hcf; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1200 = btb_wr_addr == 8'hd0; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1203 = btb_wr_addr == 8'hd1; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1206 = btb_wr_addr == 8'hd2; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1209 = btb_wr_addr == 8'hd3; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1212 = btb_wr_addr == 8'hd4; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1215 = btb_wr_addr == 8'hd5; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1218 = btb_wr_addr == 8'hd6; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1221 = btb_wr_addr == 8'hd7; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1224 = btb_wr_addr == 8'hd8; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1227 = btb_wr_addr == 8'hd9; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1230 = btb_wr_addr == 8'hda; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1233 = btb_wr_addr == 8'hdb; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1236 = btb_wr_addr == 8'hdc; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1239 = btb_wr_addr == 8'hdd; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1242 = btb_wr_addr == 8'hde; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1245 = btb_wr_addr == 8'hdf; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1248 = btb_wr_addr == 8'he0; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1251 = btb_wr_addr == 8'he1; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1254 = btb_wr_addr == 8'he2; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1257 = btb_wr_addr == 8'he3; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1260 = btb_wr_addr == 8'he4; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1263 = btb_wr_addr == 8'he5; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1266 = btb_wr_addr == 8'he6; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1269 = btb_wr_addr == 8'he7; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1272 = btb_wr_addr == 8'he8; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1275 = btb_wr_addr == 8'he9; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1278 = btb_wr_addr == 8'hea; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1281 = btb_wr_addr == 8'heb; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1284 = btb_wr_addr == 8'hec; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1287 = btb_wr_addr == 8'hed; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1290 = btb_wr_addr == 8'hee; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1293 = btb_wr_addr == 8'hef; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1296 = btb_wr_addr == 8'hf0; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1299 = btb_wr_addr == 8'hf1; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1302 = btb_wr_addr == 8'hf2; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1305 = btb_wr_addr == 8'hf3; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1308 = btb_wr_addr == 8'hf4; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1311 = btb_wr_addr == 8'hf5; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1314 = btb_wr_addr == 8'hf6; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1317 = btb_wr_addr == 8'hf7; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1320 = btb_wr_addr == 8'hf8; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1323 = btb_wr_addr == 8'hf9; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1326 = btb_wr_addr == 8'hfa; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1329 = btb_wr_addr == 8'hfb; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1332 = btb_wr_addr == 8'hfc; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1335 = btb_wr_addr == 8'hfd; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1338 = btb_wr_addr == 8'hfe; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_1341 = btb_wr_addr == 8'hff; // @[ifu_bp_ctl.scala 415:95]
  wire  _T_6210 = bht_wr_addr0[7:4] == 4'h0; // @[ifu_bp_ctl.scala 429:109]
  wire  _T_6212 = bht_wr_en0[0] & _T_6210; // @[ifu_bp_ctl.scala 429:44]
  wire  _T_6215 = bht_wr_addr2[7:4] == 4'h0; // @[ifu_bp_ctl.scala 430:109]
  wire  _T_6217 = bht_wr_en2[0] & _T_6215; // @[ifu_bp_ctl.scala 430:44]
  wire  _T_6221 = bht_wr_addr0[7:4] == 4'h1; // @[ifu_bp_ctl.scala 429:109]
  wire  _T_6223 = bht_wr_en0[0] & _T_6221; // @[ifu_bp_ctl.scala 429:44]
  wire  _T_6226 = bht_wr_addr2[7:4] == 4'h1; // @[ifu_bp_ctl.scala 430:109]
  wire  _T_6228 = bht_wr_en2[0] & _T_6226; // @[ifu_bp_ctl.scala 430:44]
  wire  _T_6232 = bht_wr_addr0[7:4] == 4'h2; // @[ifu_bp_ctl.scala 429:109]
  wire  _T_6234 = bht_wr_en0[0] & _T_6232; // @[ifu_bp_ctl.scala 429:44]
  wire  _T_6237 = bht_wr_addr2[7:4] == 4'h2; // @[ifu_bp_ctl.scala 430:109]
  wire  _T_6239 = bht_wr_en2[0] & _T_6237; // @[ifu_bp_ctl.scala 430:44]
  wire  _T_6243 = bht_wr_addr0[7:4] == 4'h3; // @[ifu_bp_ctl.scala 429:109]
  wire  _T_6245 = bht_wr_en0[0] & _T_6243; // @[ifu_bp_ctl.scala 429:44]
  wire  _T_6248 = bht_wr_addr2[7:4] == 4'h3; // @[ifu_bp_ctl.scala 430:109]
  wire  _T_6250 = bht_wr_en2[0] & _T_6248; // @[ifu_bp_ctl.scala 430:44]
  wire  _T_6254 = bht_wr_addr0[7:4] == 4'h4; // @[ifu_bp_ctl.scala 429:109]
  wire  _T_6256 = bht_wr_en0[0] & _T_6254; // @[ifu_bp_ctl.scala 429:44]
  wire  _T_6259 = bht_wr_addr2[7:4] == 4'h4; // @[ifu_bp_ctl.scala 430:109]
  wire  _T_6261 = bht_wr_en2[0] & _T_6259; // @[ifu_bp_ctl.scala 430:44]
  wire  _T_6265 = bht_wr_addr0[7:4] == 4'h5; // @[ifu_bp_ctl.scala 429:109]
  wire  _T_6267 = bht_wr_en0[0] & _T_6265; // @[ifu_bp_ctl.scala 429:44]
  wire  _T_6270 = bht_wr_addr2[7:4] == 4'h5; // @[ifu_bp_ctl.scala 430:109]
  wire  _T_6272 = bht_wr_en2[0] & _T_6270; // @[ifu_bp_ctl.scala 430:44]
  wire  _T_6276 = bht_wr_addr0[7:4] == 4'h6; // @[ifu_bp_ctl.scala 429:109]
  wire  _T_6278 = bht_wr_en0[0] & _T_6276; // @[ifu_bp_ctl.scala 429:44]
  wire  _T_6281 = bht_wr_addr2[7:4] == 4'h6; // @[ifu_bp_ctl.scala 430:109]
  wire  _T_6283 = bht_wr_en2[0] & _T_6281; // @[ifu_bp_ctl.scala 430:44]
  wire  _T_6287 = bht_wr_addr0[7:4] == 4'h7; // @[ifu_bp_ctl.scala 429:109]
  wire  _T_6289 = bht_wr_en0[0] & _T_6287; // @[ifu_bp_ctl.scala 429:44]
  wire  _T_6292 = bht_wr_addr2[7:4] == 4'h7; // @[ifu_bp_ctl.scala 430:109]
  wire  _T_6294 = bht_wr_en2[0] & _T_6292; // @[ifu_bp_ctl.scala 430:44]
  wire  _T_6298 = bht_wr_addr0[7:4] == 4'h8; // @[ifu_bp_ctl.scala 429:109]
  wire  _T_6300 = bht_wr_en0[0] & _T_6298; // @[ifu_bp_ctl.scala 429:44]
  wire  _T_6303 = bht_wr_addr2[7:4] == 4'h8; // @[ifu_bp_ctl.scala 430:109]
  wire  _T_6305 = bht_wr_en2[0] & _T_6303; // @[ifu_bp_ctl.scala 430:44]
  wire  _T_6309 = bht_wr_addr0[7:4] == 4'h9; // @[ifu_bp_ctl.scala 429:109]
  wire  _T_6311 = bht_wr_en0[0] & _T_6309; // @[ifu_bp_ctl.scala 429:44]
  wire  _T_6314 = bht_wr_addr2[7:4] == 4'h9; // @[ifu_bp_ctl.scala 430:109]
  wire  _T_6316 = bht_wr_en2[0] & _T_6314; // @[ifu_bp_ctl.scala 430:44]
  wire  _T_6320 = bht_wr_addr0[7:4] == 4'ha; // @[ifu_bp_ctl.scala 429:109]
  wire  _T_6322 = bht_wr_en0[0] & _T_6320; // @[ifu_bp_ctl.scala 429:44]
  wire  _T_6325 = bht_wr_addr2[7:4] == 4'ha; // @[ifu_bp_ctl.scala 430:109]
  wire  _T_6327 = bht_wr_en2[0] & _T_6325; // @[ifu_bp_ctl.scala 430:44]
  wire  _T_6331 = bht_wr_addr0[7:4] == 4'hb; // @[ifu_bp_ctl.scala 429:109]
  wire  _T_6333 = bht_wr_en0[0] & _T_6331; // @[ifu_bp_ctl.scala 429:44]
  wire  _T_6336 = bht_wr_addr2[7:4] == 4'hb; // @[ifu_bp_ctl.scala 430:109]
  wire  _T_6338 = bht_wr_en2[0] & _T_6336; // @[ifu_bp_ctl.scala 430:44]
  wire  _T_6342 = bht_wr_addr0[7:4] == 4'hc; // @[ifu_bp_ctl.scala 429:109]
  wire  _T_6344 = bht_wr_en0[0] & _T_6342; // @[ifu_bp_ctl.scala 429:44]
  wire  _T_6347 = bht_wr_addr2[7:4] == 4'hc; // @[ifu_bp_ctl.scala 430:109]
  wire  _T_6349 = bht_wr_en2[0] & _T_6347; // @[ifu_bp_ctl.scala 430:44]
  wire  _T_6353 = bht_wr_addr0[7:4] == 4'hd; // @[ifu_bp_ctl.scala 429:109]
  wire  _T_6355 = bht_wr_en0[0] & _T_6353; // @[ifu_bp_ctl.scala 429:44]
  wire  _T_6358 = bht_wr_addr2[7:4] == 4'hd; // @[ifu_bp_ctl.scala 430:109]
  wire  _T_6360 = bht_wr_en2[0] & _T_6358; // @[ifu_bp_ctl.scala 430:44]
  wire  _T_6364 = bht_wr_addr0[7:4] == 4'he; // @[ifu_bp_ctl.scala 429:109]
  wire  _T_6366 = bht_wr_en0[0] & _T_6364; // @[ifu_bp_ctl.scala 429:44]
  wire  _T_6369 = bht_wr_addr2[7:4] == 4'he; // @[ifu_bp_ctl.scala 430:109]
  wire  _T_6371 = bht_wr_en2[0] & _T_6369; // @[ifu_bp_ctl.scala 430:44]
  wire  _T_6375 = bht_wr_addr0[7:4] == 4'hf; // @[ifu_bp_ctl.scala 429:109]
  wire  _T_6377 = bht_wr_en0[0] & _T_6375; // @[ifu_bp_ctl.scala 429:44]
  wire  _T_6380 = bht_wr_addr2[7:4] == 4'hf; // @[ifu_bp_ctl.scala 430:109]
  wire  _T_6382 = bht_wr_en2[0] & _T_6380; // @[ifu_bp_ctl.scala 430:44]
  wire  _T_6388 = bht_wr_en0[1] & _T_6210; // @[ifu_bp_ctl.scala 429:44]
  wire  _T_6393 = bht_wr_en2[1] & _T_6215; // @[ifu_bp_ctl.scala 430:44]
  wire  _T_6399 = bht_wr_en0[1] & _T_6221; // @[ifu_bp_ctl.scala 429:44]
  wire  _T_6404 = bht_wr_en2[1] & _T_6226; // @[ifu_bp_ctl.scala 430:44]
  wire  _T_6410 = bht_wr_en0[1] & _T_6232; // @[ifu_bp_ctl.scala 429:44]
  wire  _T_6415 = bht_wr_en2[1] & _T_6237; // @[ifu_bp_ctl.scala 430:44]
  wire  _T_6421 = bht_wr_en0[1] & _T_6243; // @[ifu_bp_ctl.scala 429:44]
  wire  _T_6426 = bht_wr_en2[1] & _T_6248; // @[ifu_bp_ctl.scala 430:44]
  wire  _T_6432 = bht_wr_en0[1] & _T_6254; // @[ifu_bp_ctl.scala 429:44]
  wire  _T_6437 = bht_wr_en2[1] & _T_6259; // @[ifu_bp_ctl.scala 430:44]
  wire  _T_6443 = bht_wr_en0[1] & _T_6265; // @[ifu_bp_ctl.scala 429:44]
  wire  _T_6448 = bht_wr_en2[1] & _T_6270; // @[ifu_bp_ctl.scala 430:44]
  wire  _T_6454 = bht_wr_en0[1] & _T_6276; // @[ifu_bp_ctl.scala 429:44]
  wire  _T_6459 = bht_wr_en2[1] & _T_6281; // @[ifu_bp_ctl.scala 430:44]
  wire  _T_6465 = bht_wr_en0[1] & _T_6287; // @[ifu_bp_ctl.scala 429:44]
  wire  _T_6470 = bht_wr_en2[1] & _T_6292; // @[ifu_bp_ctl.scala 430:44]
  wire  _T_6476 = bht_wr_en0[1] & _T_6298; // @[ifu_bp_ctl.scala 429:44]
  wire  _T_6481 = bht_wr_en2[1] & _T_6303; // @[ifu_bp_ctl.scala 430:44]
  wire  _T_6487 = bht_wr_en0[1] & _T_6309; // @[ifu_bp_ctl.scala 429:44]
  wire  _T_6492 = bht_wr_en2[1] & _T_6314; // @[ifu_bp_ctl.scala 430:44]
  wire  _T_6498 = bht_wr_en0[1] & _T_6320; // @[ifu_bp_ctl.scala 429:44]
  wire  _T_6503 = bht_wr_en2[1] & _T_6325; // @[ifu_bp_ctl.scala 430:44]
  wire  _T_6509 = bht_wr_en0[1] & _T_6331; // @[ifu_bp_ctl.scala 429:44]
  wire  _T_6514 = bht_wr_en2[1] & _T_6336; // @[ifu_bp_ctl.scala 430:44]
  wire  _T_6520 = bht_wr_en0[1] & _T_6342; // @[ifu_bp_ctl.scala 429:44]
  wire  _T_6525 = bht_wr_en2[1] & _T_6347; // @[ifu_bp_ctl.scala 430:44]
  wire  _T_6531 = bht_wr_en0[1] & _T_6353; // @[ifu_bp_ctl.scala 429:44]
  wire  _T_6536 = bht_wr_en2[1] & _T_6358; // @[ifu_bp_ctl.scala 430:44]
  wire  _T_6542 = bht_wr_en0[1] & _T_6364; // @[ifu_bp_ctl.scala 429:44]
  wire  _T_6547 = bht_wr_en2[1] & _T_6369; // @[ifu_bp_ctl.scala 430:44]
  wire  _T_6553 = bht_wr_en0[1] & _T_6375; // @[ifu_bp_ctl.scala 429:44]
  wire  _T_6558 = bht_wr_en2[1] & _T_6380; // @[ifu_bp_ctl.scala 430:44]
  wire  _T_6562 = bht_wr_addr2[3:0] == 4'h0; // @[ifu_bp_ctl.scala 435:74]
  wire  _T_6563 = bht_wr_en2[0] & _T_6562; // @[ifu_bp_ctl.scala 435:23]
  wire  _T_6566 = _T_6563 & _T_6215; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_6571 = bht_wr_addr2[3:0] == 4'h1; // @[ifu_bp_ctl.scala 435:74]
  wire  _T_6572 = bht_wr_en2[0] & _T_6571; // @[ifu_bp_ctl.scala 435:23]
  wire  _T_6575 = _T_6572 & _T_6215; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_6580 = bht_wr_addr2[3:0] == 4'h2; // @[ifu_bp_ctl.scala 435:74]
  wire  _T_6581 = bht_wr_en2[0] & _T_6580; // @[ifu_bp_ctl.scala 435:23]
  wire  _T_6584 = _T_6581 & _T_6215; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_6589 = bht_wr_addr2[3:0] == 4'h3; // @[ifu_bp_ctl.scala 435:74]
  wire  _T_6590 = bht_wr_en2[0] & _T_6589; // @[ifu_bp_ctl.scala 435:23]
  wire  _T_6593 = _T_6590 & _T_6215; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_6598 = bht_wr_addr2[3:0] == 4'h4; // @[ifu_bp_ctl.scala 435:74]
  wire  _T_6599 = bht_wr_en2[0] & _T_6598; // @[ifu_bp_ctl.scala 435:23]
  wire  _T_6602 = _T_6599 & _T_6215; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_6607 = bht_wr_addr2[3:0] == 4'h5; // @[ifu_bp_ctl.scala 435:74]
  wire  _T_6608 = bht_wr_en2[0] & _T_6607; // @[ifu_bp_ctl.scala 435:23]
  wire  _T_6611 = _T_6608 & _T_6215; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_6616 = bht_wr_addr2[3:0] == 4'h6; // @[ifu_bp_ctl.scala 435:74]
  wire  _T_6617 = bht_wr_en2[0] & _T_6616; // @[ifu_bp_ctl.scala 435:23]
  wire  _T_6620 = _T_6617 & _T_6215; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_6625 = bht_wr_addr2[3:0] == 4'h7; // @[ifu_bp_ctl.scala 435:74]
  wire  _T_6626 = bht_wr_en2[0] & _T_6625; // @[ifu_bp_ctl.scala 435:23]
  wire  _T_6629 = _T_6626 & _T_6215; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_6634 = bht_wr_addr2[3:0] == 4'h8; // @[ifu_bp_ctl.scala 435:74]
  wire  _T_6635 = bht_wr_en2[0] & _T_6634; // @[ifu_bp_ctl.scala 435:23]
  wire  _T_6638 = _T_6635 & _T_6215; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_6643 = bht_wr_addr2[3:0] == 4'h9; // @[ifu_bp_ctl.scala 435:74]
  wire  _T_6644 = bht_wr_en2[0] & _T_6643; // @[ifu_bp_ctl.scala 435:23]
  wire  _T_6647 = _T_6644 & _T_6215; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_6652 = bht_wr_addr2[3:0] == 4'ha; // @[ifu_bp_ctl.scala 435:74]
  wire  _T_6653 = bht_wr_en2[0] & _T_6652; // @[ifu_bp_ctl.scala 435:23]
  wire  _T_6656 = _T_6653 & _T_6215; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_6661 = bht_wr_addr2[3:0] == 4'hb; // @[ifu_bp_ctl.scala 435:74]
  wire  _T_6662 = bht_wr_en2[0] & _T_6661; // @[ifu_bp_ctl.scala 435:23]
  wire  _T_6665 = _T_6662 & _T_6215; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_6670 = bht_wr_addr2[3:0] == 4'hc; // @[ifu_bp_ctl.scala 435:74]
  wire  _T_6671 = bht_wr_en2[0] & _T_6670; // @[ifu_bp_ctl.scala 435:23]
  wire  _T_6674 = _T_6671 & _T_6215; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_6679 = bht_wr_addr2[3:0] == 4'hd; // @[ifu_bp_ctl.scala 435:74]
  wire  _T_6680 = bht_wr_en2[0] & _T_6679; // @[ifu_bp_ctl.scala 435:23]
  wire  _T_6683 = _T_6680 & _T_6215; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_6688 = bht_wr_addr2[3:0] == 4'he; // @[ifu_bp_ctl.scala 435:74]
  wire  _T_6689 = bht_wr_en2[0] & _T_6688; // @[ifu_bp_ctl.scala 435:23]
  wire  _T_6692 = _T_6689 & _T_6215; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_6697 = bht_wr_addr2[3:0] == 4'hf; // @[ifu_bp_ctl.scala 435:74]
  wire  _T_6698 = bht_wr_en2[0] & _T_6697; // @[ifu_bp_ctl.scala 435:23]
  wire  _T_6701 = _T_6698 & _T_6215; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_6710 = _T_6563 & _T_6226; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_6719 = _T_6572 & _T_6226; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_6728 = _T_6581 & _T_6226; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_6737 = _T_6590 & _T_6226; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_6746 = _T_6599 & _T_6226; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_6755 = _T_6608 & _T_6226; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_6764 = _T_6617 & _T_6226; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_6773 = _T_6626 & _T_6226; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_6782 = _T_6635 & _T_6226; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_6791 = _T_6644 & _T_6226; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_6800 = _T_6653 & _T_6226; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_6809 = _T_6662 & _T_6226; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_6818 = _T_6671 & _T_6226; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_6827 = _T_6680 & _T_6226; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_6836 = _T_6689 & _T_6226; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_6845 = _T_6698 & _T_6226; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_6854 = _T_6563 & _T_6237; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_6863 = _T_6572 & _T_6237; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_6872 = _T_6581 & _T_6237; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_6881 = _T_6590 & _T_6237; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_6890 = _T_6599 & _T_6237; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_6899 = _T_6608 & _T_6237; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_6908 = _T_6617 & _T_6237; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_6917 = _T_6626 & _T_6237; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_6926 = _T_6635 & _T_6237; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_6935 = _T_6644 & _T_6237; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_6944 = _T_6653 & _T_6237; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_6953 = _T_6662 & _T_6237; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_6962 = _T_6671 & _T_6237; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_6971 = _T_6680 & _T_6237; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_6980 = _T_6689 & _T_6237; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_6989 = _T_6698 & _T_6237; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_6998 = _T_6563 & _T_6248; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7007 = _T_6572 & _T_6248; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7016 = _T_6581 & _T_6248; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7025 = _T_6590 & _T_6248; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7034 = _T_6599 & _T_6248; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7043 = _T_6608 & _T_6248; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7052 = _T_6617 & _T_6248; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7061 = _T_6626 & _T_6248; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7070 = _T_6635 & _T_6248; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7079 = _T_6644 & _T_6248; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7088 = _T_6653 & _T_6248; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7097 = _T_6662 & _T_6248; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7106 = _T_6671 & _T_6248; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7115 = _T_6680 & _T_6248; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7124 = _T_6689 & _T_6248; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7133 = _T_6698 & _T_6248; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7142 = _T_6563 & _T_6259; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7151 = _T_6572 & _T_6259; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7160 = _T_6581 & _T_6259; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7169 = _T_6590 & _T_6259; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7178 = _T_6599 & _T_6259; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7187 = _T_6608 & _T_6259; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7196 = _T_6617 & _T_6259; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7205 = _T_6626 & _T_6259; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7214 = _T_6635 & _T_6259; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7223 = _T_6644 & _T_6259; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7232 = _T_6653 & _T_6259; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7241 = _T_6662 & _T_6259; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7250 = _T_6671 & _T_6259; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7259 = _T_6680 & _T_6259; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7268 = _T_6689 & _T_6259; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7277 = _T_6698 & _T_6259; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7286 = _T_6563 & _T_6270; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7295 = _T_6572 & _T_6270; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7304 = _T_6581 & _T_6270; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7313 = _T_6590 & _T_6270; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7322 = _T_6599 & _T_6270; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7331 = _T_6608 & _T_6270; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7340 = _T_6617 & _T_6270; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7349 = _T_6626 & _T_6270; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7358 = _T_6635 & _T_6270; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7367 = _T_6644 & _T_6270; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7376 = _T_6653 & _T_6270; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7385 = _T_6662 & _T_6270; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7394 = _T_6671 & _T_6270; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7403 = _T_6680 & _T_6270; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7412 = _T_6689 & _T_6270; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7421 = _T_6698 & _T_6270; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7430 = _T_6563 & _T_6281; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7439 = _T_6572 & _T_6281; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7448 = _T_6581 & _T_6281; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7457 = _T_6590 & _T_6281; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7466 = _T_6599 & _T_6281; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7475 = _T_6608 & _T_6281; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7484 = _T_6617 & _T_6281; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7493 = _T_6626 & _T_6281; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7502 = _T_6635 & _T_6281; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7511 = _T_6644 & _T_6281; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7520 = _T_6653 & _T_6281; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7529 = _T_6662 & _T_6281; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7538 = _T_6671 & _T_6281; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7547 = _T_6680 & _T_6281; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7556 = _T_6689 & _T_6281; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7565 = _T_6698 & _T_6281; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7574 = _T_6563 & _T_6292; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7583 = _T_6572 & _T_6292; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7592 = _T_6581 & _T_6292; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7601 = _T_6590 & _T_6292; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7610 = _T_6599 & _T_6292; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7619 = _T_6608 & _T_6292; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7628 = _T_6617 & _T_6292; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7637 = _T_6626 & _T_6292; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7646 = _T_6635 & _T_6292; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7655 = _T_6644 & _T_6292; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7664 = _T_6653 & _T_6292; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7673 = _T_6662 & _T_6292; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7682 = _T_6671 & _T_6292; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7691 = _T_6680 & _T_6292; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7700 = _T_6689 & _T_6292; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7709 = _T_6698 & _T_6292; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7718 = _T_6563 & _T_6303; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7727 = _T_6572 & _T_6303; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7736 = _T_6581 & _T_6303; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7745 = _T_6590 & _T_6303; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7754 = _T_6599 & _T_6303; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7763 = _T_6608 & _T_6303; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7772 = _T_6617 & _T_6303; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7781 = _T_6626 & _T_6303; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7790 = _T_6635 & _T_6303; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7799 = _T_6644 & _T_6303; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7808 = _T_6653 & _T_6303; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7817 = _T_6662 & _T_6303; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7826 = _T_6671 & _T_6303; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7835 = _T_6680 & _T_6303; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7844 = _T_6689 & _T_6303; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7853 = _T_6698 & _T_6303; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7862 = _T_6563 & _T_6314; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7871 = _T_6572 & _T_6314; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7880 = _T_6581 & _T_6314; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7889 = _T_6590 & _T_6314; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7898 = _T_6599 & _T_6314; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7907 = _T_6608 & _T_6314; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7916 = _T_6617 & _T_6314; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7925 = _T_6626 & _T_6314; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7934 = _T_6635 & _T_6314; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7943 = _T_6644 & _T_6314; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7952 = _T_6653 & _T_6314; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7961 = _T_6662 & _T_6314; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7970 = _T_6671 & _T_6314; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7979 = _T_6680 & _T_6314; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7988 = _T_6689 & _T_6314; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_7997 = _T_6698 & _T_6314; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8006 = _T_6563 & _T_6325; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8015 = _T_6572 & _T_6325; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8024 = _T_6581 & _T_6325; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8033 = _T_6590 & _T_6325; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8042 = _T_6599 & _T_6325; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8051 = _T_6608 & _T_6325; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8060 = _T_6617 & _T_6325; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8069 = _T_6626 & _T_6325; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8078 = _T_6635 & _T_6325; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8087 = _T_6644 & _T_6325; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8096 = _T_6653 & _T_6325; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8105 = _T_6662 & _T_6325; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8114 = _T_6671 & _T_6325; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8123 = _T_6680 & _T_6325; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8132 = _T_6689 & _T_6325; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8141 = _T_6698 & _T_6325; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8150 = _T_6563 & _T_6336; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8159 = _T_6572 & _T_6336; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8168 = _T_6581 & _T_6336; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8177 = _T_6590 & _T_6336; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8186 = _T_6599 & _T_6336; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8195 = _T_6608 & _T_6336; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8204 = _T_6617 & _T_6336; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8213 = _T_6626 & _T_6336; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8222 = _T_6635 & _T_6336; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8231 = _T_6644 & _T_6336; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8240 = _T_6653 & _T_6336; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8249 = _T_6662 & _T_6336; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8258 = _T_6671 & _T_6336; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8267 = _T_6680 & _T_6336; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8276 = _T_6689 & _T_6336; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8285 = _T_6698 & _T_6336; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8294 = _T_6563 & _T_6347; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8303 = _T_6572 & _T_6347; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8312 = _T_6581 & _T_6347; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8321 = _T_6590 & _T_6347; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8330 = _T_6599 & _T_6347; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8339 = _T_6608 & _T_6347; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8348 = _T_6617 & _T_6347; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8357 = _T_6626 & _T_6347; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8366 = _T_6635 & _T_6347; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8375 = _T_6644 & _T_6347; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8384 = _T_6653 & _T_6347; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8393 = _T_6662 & _T_6347; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8402 = _T_6671 & _T_6347; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8411 = _T_6680 & _T_6347; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8420 = _T_6689 & _T_6347; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8429 = _T_6698 & _T_6347; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8438 = _T_6563 & _T_6358; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8447 = _T_6572 & _T_6358; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8456 = _T_6581 & _T_6358; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8465 = _T_6590 & _T_6358; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8474 = _T_6599 & _T_6358; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8483 = _T_6608 & _T_6358; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8492 = _T_6617 & _T_6358; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8501 = _T_6626 & _T_6358; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8510 = _T_6635 & _T_6358; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8519 = _T_6644 & _T_6358; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8528 = _T_6653 & _T_6358; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8537 = _T_6662 & _T_6358; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8546 = _T_6671 & _T_6358; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8555 = _T_6680 & _T_6358; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8564 = _T_6689 & _T_6358; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8573 = _T_6698 & _T_6358; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8582 = _T_6563 & _T_6369; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8591 = _T_6572 & _T_6369; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8600 = _T_6581 & _T_6369; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8609 = _T_6590 & _T_6369; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8618 = _T_6599 & _T_6369; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8627 = _T_6608 & _T_6369; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8636 = _T_6617 & _T_6369; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8645 = _T_6626 & _T_6369; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8654 = _T_6635 & _T_6369; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8663 = _T_6644 & _T_6369; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8672 = _T_6653 & _T_6369; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8681 = _T_6662 & _T_6369; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8690 = _T_6671 & _T_6369; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8699 = _T_6680 & _T_6369; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8708 = _T_6689 & _T_6369; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8717 = _T_6698 & _T_6369; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8726 = _T_6563 & _T_6380; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8735 = _T_6572 & _T_6380; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8744 = _T_6581 & _T_6380; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8753 = _T_6590 & _T_6380; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8762 = _T_6599 & _T_6380; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8771 = _T_6608 & _T_6380; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8780 = _T_6617 & _T_6380; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8789 = _T_6626 & _T_6380; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8798 = _T_6635 & _T_6380; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8807 = _T_6644 & _T_6380; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8816 = _T_6653 & _T_6380; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8825 = _T_6662 & _T_6380; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8834 = _T_6671 & _T_6380; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8843 = _T_6680 & _T_6380; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8852 = _T_6689 & _T_6380; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8861 = _T_6698 & _T_6380; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8867 = bht_wr_en2[1] & _T_6562; // @[ifu_bp_ctl.scala 435:23]
  wire  _T_8870 = _T_8867 & _T_6215; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8876 = bht_wr_en2[1] & _T_6571; // @[ifu_bp_ctl.scala 435:23]
  wire  _T_8879 = _T_8876 & _T_6215; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8885 = bht_wr_en2[1] & _T_6580; // @[ifu_bp_ctl.scala 435:23]
  wire  _T_8888 = _T_8885 & _T_6215; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8894 = bht_wr_en2[1] & _T_6589; // @[ifu_bp_ctl.scala 435:23]
  wire  _T_8897 = _T_8894 & _T_6215; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8903 = bht_wr_en2[1] & _T_6598; // @[ifu_bp_ctl.scala 435:23]
  wire  _T_8906 = _T_8903 & _T_6215; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8912 = bht_wr_en2[1] & _T_6607; // @[ifu_bp_ctl.scala 435:23]
  wire  _T_8915 = _T_8912 & _T_6215; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8921 = bht_wr_en2[1] & _T_6616; // @[ifu_bp_ctl.scala 435:23]
  wire  _T_8924 = _T_8921 & _T_6215; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8930 = bht_wr_en2[1] & _T_6625; // @[ifu_bp_ctl.scala 435:23]
  wire  _T_8933 = _T_8930 & _T_6215; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8939 = bht_wr_en2[1] & _T_6634; // @[ifu_bp_ctl.scala 435:23]
  wire  _T_8942 = _T_8939 & _T_6215; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8948 = bht_wr_en2[1] & _T_6643; // @[ifu_bp_ctl.scala 435:23]
  wire  _T_8951 = _T_8948 & _T_6215; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8957 = bht_wr_en2[1] & _T_6652; // @[ifu_bp_ctl.scala 435:23]
  wire  _T_8960 = _T_8957 & _T_6215; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8966 = bht_wr_en2[1] & _T_6661; // @[ifu_bp_ctl.scala 435:23]
  wire  _T_8969 = _T_8966 & _T_6215; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8975 = bht_wr_en2[1] & _T_6670; // @[ifu_bp_ctl.scala 435:23]
  wire  _T_8978 = _T_8975 & _T_6215; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8984 = bht_wr_en2[1] & _T_6679; // @[ifu_bp_ctl.scala 435:23]
  wire  _T_8987 = _T_8984 & _T_6215; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_8993 = bht_wr_en2[1] & _T_6688; // @[ifu_bp_ctl.scala 435:23]
  wire  _T_8996 = _T_8993 & _T_6215; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9002 = bht_wr_en2[1] & _T_6697; // @[ifu_bp_ctl.scala 435:23]
  wire  _T_9005 = _T_9002 & _T_6215; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9014 = _T_8867 & _T_6226; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9023 = _T_8876 & _T_6226; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9032 = _T_8885 & _T_6226; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9041 = _T_8894 & _T_6226; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9050 = _T_8903 & _T_6226; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9059 = _T_8912 & _T_6226; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9068 = _T_8921 & _T_6226; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9077 = _T_8930 & _T_6226; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9086 = _T_8939 & _T_6226; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9095 = _T_8948 & _T_6226; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9104 = _T_8957 & _T_6226; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9113 = _T_8966 & _T_6226; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9122 = _T_8975 & _T_6226; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9131 = _T_8984 & _T_6226; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9140 = _T_8993 & _T_6226; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9149 = _T_9002 & _T_6226; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9158 = _T_8867 & _T_6237; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9167 = _T_8876 & _T_6237; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9176 = _T_8885 & _T_6237; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9185 = _T_8894 & _T_6237; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9194 = _T_8903 & _T_6237; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9203 = _T_8912 & _T_6237; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9212 = _T_8921 & _T_6237; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9221 = _T_8930 & _T_6237; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9230 = _T_8939 & _T_6237; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9239 = _T_8948 & _T_6237; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9248 = _T_8957 & _T_6237; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9257 = _T_8966 & _T_6237; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9266 = _T_8975 & _T_6237; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9275 = _T_8984 & _T_6237; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9284 = _T_8993 & _T_6237; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9293 = _T_9002 & _T_6237; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9302 = _T_8867 & _T_6248; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9311 = _T_8876 & _T_6248; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9320 = _T_8885 & _T_6248; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9329 = _T_8894 & _T_6248; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9338 = _T_8903 & _T_6248; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9347 = _T_8912 & _T_6248; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9356 = _T_8921 & _T_6248; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9365 = _T_8930 & _T_6248; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9374 = _T_8939 & _T_6248; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9383 = _T_8948 & _T_6248; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9392 = _T_8957 & _T_6248; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9401 = _T_8966 & _T_6248; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9410 = _T_8975 & _T_6248; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9419 = _T_8984 & _T_6248; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9428 = _T_8993 & _T_6248; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9437 = _T_9002 & _T_6248; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9446 = _T_8867 & _T_6259; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9455 = _T_8876 & _T_6259; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9464 = _T_8885 & _T_6259; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9473 = _T_8894 & _T_6259; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9482 = _T_8903 & _T_6259; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9491 = _T_8912 & _T_6259; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9500 = _T_8921 & _T_6259; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9509 = _T_8930 & _T_6259; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9518 = _T_8939 & _T_6259; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9527 = _T_8948 & _T_6259; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9536 = _T_8957 & _T_6259; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9545 = _T_8966 & _T_6259; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9554 = _T_8975 & _T_6259; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9563 = _T_8984 & _T_6259; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9572 = _T_8993 & _T_6259; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9581 = _T_9002 & _T_6259; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9590 = _T_8867 & _T_6270; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9599 = _T_8876 & _T_6270; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9608 = _T_8885 & _T_6270; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9617 = _T_8894 & _T_6270; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9626 = _T_8903 & _T_6270; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9635 = _T_8912 & _T_6270; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9644 = _T_8921 & _T_6270; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9653 = _T_8930 & _T_6270; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9662 = _T_8939 & _T_6270; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9671 = _T_8948 & _T_6270; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9680 = _T_8957 & _T_6270; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9689 = _T_8966 & _T_6270; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9698 = _T_8975 & _T_6270; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9707 = _T_8984 & _T_6270; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9716 = _T_8993 & _T_6270; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9725 = _T_9002 & _T_6270; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9734 = _T_8867 & _T_6281; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9743 = _T_8876 & _T_6281; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9752 = _T_8885 & _T_6281; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9761 = _T_8894 & _T_6281; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9770 = _T_8903 & _T_6281; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9779 = _T_8912 & _T_6281; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9788 = _T_8921 & _T_6281; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9797 = _T_8930 & _T_6281; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9806 = _T_8939 & _T_6281; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9815 = _T_8948 & _T_6281; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9824 = _T_8957 & _T_6281; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9833 = _T_8966 & _T_6281; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9842 = _T_8975 & _T_6281; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9851 = _T_8984 & _T_6281; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9860 = _T_8993 & _T_6281; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9869 = _T_9002 & _T_6281; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9878 = _T_8867 & _T_6292; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9887 = _T_8876 & _T_6292; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9896 = _T_8885 & _T_6292; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9905 = _T_8894 & _T_6292; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9914 = _T_8903 & _T_6292; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9923 = _T_8912 & _T_6292; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9932 = _T_8921 & _T_6292; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9941 = _T_8930 & _T_6292; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9950 = _T_8939 & _T_6292; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9959 = _T_8948 & _T_6292; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9968 = _T_8957 & _T_6292; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9977 = _T_8966 & _T_6292; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9986 = _T_8975 & _T_6292; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_9995 = _T_8984 & _T_6292; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10004 = _T_8993 & _T_6292; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10013 = _T_9002 & _T_6292; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10022 = _T_8867 & _T_6303; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10031 = _T_8876 & _T_6303; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10040 = _T_8885 & _T_6303; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10049 = _T_8894 & _T_6303; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10058 = _T_8903 & _T_6303; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10067 = _T_8912 & _T_6303; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10076 = _T_8921 & _T_6303; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10085 = _T_8930 & _T_6303; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10094 = _T_8939 & _T_6303; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10103 = _T_8948 & _T_6303; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10112 = _T_8957 & _T_6303; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10121 = _T_8966 & _T_6303; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10130 = _T_8975 & _T_6303; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10139 = _T_8984 & _T_6303; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10148 = _T_8993 & _T_6303; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10157 = _T_9002 & _T_6303; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10166 = _T_8867 & _T_6314; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10175 = _T_8876 & _T_6314; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10184 = _T_8885 & _T_6314; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10193 = _T_8894 & _T_6314; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10202 = _T_8903 & _T_6314; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10211 = _T_8912 & _T_6314; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10220 = _T_8921 & _T_6314; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10229 = _T_8930 & _T_6314; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10238 = _T_8939 & _T_6314; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10247 = _T_8948 & _T_6314; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10256 = _T_8957 & _T_6314; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10265 = _T_8966 & _T_6314; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10274 = _T_8975 & _T_6314; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10283 = _T_8984 & _T_6314; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10292 = _T_8993 & _T_6314; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10301 = _T_9002 & _T_6314; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10310 = _T_8867 & _T_6325; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10319 = _T_8876 & _T_6325; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10328 = _T_8885 & _T_6325; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10337 = _T_8894 & _T_6325; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10346 = _T_8903 & _T_6325; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10355 = _T_8912 & _T_6325; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10364 = _T_8921 & _T_6325; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10373 = _T_8930 & _T_6325; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10382 = _T_8939 & _T_6325; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10391 = _T_8948 & _T_6325; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10400 = _T_8957 & _T_6325; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10409 = _T_8966 & _T_6325; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10418 = _T_8975 & _T_6325; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10427 = _T_8984 & _T_6325; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10436 = _T_8993 & _T_6325; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10445 = _T_9002 & _T_6325; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10454 = _T_8867 & _T_6336; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10463 = _T_8876 & _T_6336; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10472 = _T_8885 & _T_6336; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10481 = _T_8894 & _T_6336; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10490 = _T_8903 & _T_6336; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10499 = _T_8912 & _T_6336; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10508 = _T_8921 & _T_6336; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10517 = _T_8930 & _T_6336; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10526 = _T_8939 & _T_6336; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10535 = _T_8948 & _T_6336; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10544 = _T_8957 & _T_6336; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10553 = _T_8966 & _T_6336; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10562 = _T_8975 & _T_6336; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10571 = _T_8984 & _T_6336; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10580 = _T_8993 & _T_6336; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10589 = _T_9002 & _T_6336; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10598 = _T_8867 & _T_6347; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10607 = _T_8876 & _T_6347; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10616 = _T_8885 & _T_6347; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10625 = _T_8894 & _T_6347; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10634 = _T_8903 & _T_6347; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10643 = _T_8912 & _T_6347; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10652 = _T_8921 & _T_6347; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10661 = _T_8930 & _T_6347; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10670 = _T_8939 & _T_6347; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10679 = _T_8948 & _T_6347; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10688 = _T_8957 & _T_6347; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10697 = _T_8966 & _T_6347; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10706 = _T_8975 & _T_6347; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10715 = _T_8984 & _T_6347; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10724 = _T_8993 & _T_6347; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10733 = _T_9002 & _T_6347; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10742 = _T_8867 & _T_6358; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10751 = _T_8876 & _T_6358; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10760 = _T_8885 & _T_6358; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10769 = _T_8894 & _T_6358; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10778 = _T_8903 & _T_6358; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10787 = _T_8912 & _T_6358; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10796 = _T_8921 & _T_6358; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10805 = _T_8930 & _T_6358; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10814 = _T_8939 & _T_6358; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10823 = _T_8948 & _T_6358; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10832 = _T_8957 & _T_6358; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10841 = _T_8966 & _T_6358; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10850 = _T_8975 & _T_6358; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10859 = _T_8984 & _T_6358; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10868 = _T_8993 & _T_6358; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10877 = _T_9002 & _T_6358; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10886 = _T_8867 & _T_6369; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10895 = _T_8876 & _T_6369; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10904 = _T_8885 & _T_6369; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10913 = _T_8894 & _T_6369; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10922 = _T_8903 & _T_6369; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10931 = _T_8912 & _T_6369; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10940 = _T_8921 & _T_6369; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10949 = _T_8930 & _T_6369; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10958 = _T_8939 & _T_6369; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10967 = _T_8948 & _T_6369; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10976 = _T_8957 & _T_6369; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10985 = _T_8966 & _T_6369; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_10994 = _T_8975 & _T_6369; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_11003 = _T_8984 & _T_6369; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_11012 = _T_8993 & _T_6369; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_11021 = _T_9002 & _T_6369; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_11030 = _T_8867 & _T_6380; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_11039 = _T_8876 & _T_6380; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_11048 = _T_8885 & _T_6380; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_11057 = _T_8894 & _T_6380; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_11066 = _T_8903 & _T_6380; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_11075 = _T_8912 & _T_6380; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_11084 = _T_8921 & _T_6380; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_11093 = _T_8930 & _T_6380; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_11102 = _T_8939 & _T_6380; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_11111 = _T_8948 & _T_6380; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_11120 = _T_8957 & _T_6380; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_11129 = _T_8966 & _T_6380; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_11138 = _T_8975 & _T_6380; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_11147 = _T_8984 & _T_6380; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_11156 = _T_8993 & _T_6380; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_11165 = _T_9002 & _T_6380; // @[ifu_bp_ctl.scala 435:81]
  wire  _T_11170 = bht_wr_addr0[3:0] == 4'h0; // @[ifu_bp_ctl.scala 443:97]
  wire  _T_11171 = bht_wr_en0[0] & _T_11170; // @[ifu_bp_ctl.scala 443:45]
  wire  _T_11175 = _T_11171 & _T_6210; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_0_0 = _T_11175 | _T_6566; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_11187 = bht_wr_addr0[3:0] == 4'h1; // @[ifu_bp_ctl.scala 443:97]
  wire  _T_11188 = bht_wr_en0[0] & _T_11187; // @[ifu_bp_ctl.scala 443:45]
  wire  _T_11192 = _T_11188 & _T_6210; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_0_1 = _T_11192 | _T_6575; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_11204 = bht_wr_addr0[3:0] == 4'h2; // @[ifu_bp_ctl.scala 443:97]
  wire  _T_11205 = bht_wr_en0[0] & _T_11204; // @[ifu_bp_ctl.scala 443:45]
  wire  _T_11209 = _T_11205 & _T_6210; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_0_2 = _T_11209 | _T_6584; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_11221 = bht_wr_addr0[3:0] == 4'h3; // @[ifu_bp_ctl.scala 443:97]
  wire  _T_11222 = bht_wr_en0[0] & _T_11221; // @[ifu_bp_ctl.scala 443:45]
  wire  _T_11226 = _T_11222 & _T_6210; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_0_3 = _T_11226 | _T_6593; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_11238 = bht_wr_addr0[3:0] == 4'h4; // @[ifu_bp_ctl.scala 443:97]
  wire  _T_11239 = bht_wr_en0[0] & _T_11238; // @[ifu_bp_ctl.scala 443:45]
  wire  _T_11243 = _T_11239 & _T_6210; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_0_4 = _T_11243 | _T_6602; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_11255 = bht_wr_addr0[3:0] == 4'h5; // @[ifu_bp_ctl.scala 443:97]
  wire  _T_11256 = bht_wr_en0[0] & _T_11255; // @[ifu_bp_ctl.scala 443:45]
  wire  _T_11260 = _T_11256 & _T_6210; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_0_5 = _T_11260 | _T_6611; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_11272 = bht_wr_addr0[3:0] == 4'h6; // @[ifu_bp_ctl.scala 443:97]
  wire  _T_11273 = bht_wr_en0[0] & _T_11272; // @[ifu_bp_ctl.scala 443:45]
  wire  _T_11277 = _T_11273 & _T_6210; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_0_6 = _T_11277 | _T_6620; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_11289 = bht_wr_addr0[3:0] == 4'h7; // @[ifu_bp_ctl.scala 443:97]
  wire  _T_11290 = bht_wr_en0[0] & _T_11289; // @[ifu_bp_ctl.scala 443:45]
  wire  _T_11294 = _T_11290 & _T_6210; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_0_7 = _T_11294 | _T_6629; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_11306 = bht_wr_addr0[3:0] == 4'h8; // @[ifu_bp_ctl.scala 443:97]
  wire  _T_11307 = bht_wr_en0[0] & _T_11306; // @[ifu_bp_ctl.scala 443:45]
  wire  _T_11311 = _T_11307 & _T_6210; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_0_8 = _T_11311 | _T_6638; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_11323 = bht_wr_addr0[3:0] == 4'h9; // @[ifu_bp_ctl.scala 443:97]
  wire  _T_11324 = bht_wr_en0[0] & _T_11323; // @[ifu_bp_ctl.scala 443:45]
  wire  _T_11328 = _T_11324 & _T_6210; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_0_9 = _T_11328 | _T_6647; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_11340 = bht_wr_addr0[3:0] == 4'ha; // @[ifu_bp_ctl.scala 443:97]
  wire  _T_11341 = bht_wr_en0[0] & _T_11340; // @[ifu_bp_ctl.scala 443:45]
  wire  _T_11345 = _T_11341 & _T_6210; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_0_10 = _T_11345 | _T_6656; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_11357 = bht_wr_addr0[3:0] == 4'hb; // @[ifu_bp_ctl.scala 443:97]
  wire  _T_11358 = bht_wr_en0[0] & _T_11357; // @[ifu_bp_ctl.scala 443:45]
  wire  _T_11362 = _T_11358 & _T_6210; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_0_11 = _T_11362 | _T_6665; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_11374 = bht_wr_addr0[3:0] == 4'hc; // @[ifu_bp_ctl.scala 443:97]
  wire  _T_11375 = bht_wr_en0[0] & _T_11374; // @[ifu_bp_ctl.scala 443:45]
  wire  _T_11379 = _T_11375 & _T_6210; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_0_12 = _T_11379 | _T_6674; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_11391 = bht_wr_addr0[3:0] == 4'hd; // @[ifu_bp_ctl.scala 443:97]
  wire  _T_11392 = bht_wr_en0[0] & _T_11391; // @[ifu_bp_ctl.scala 443:45]
  wire  _T_11396 = _T_11392 & _T_6210; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_0_13 = _T_11396 | _T_6683; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_11408 = bht_wr_addr0[3:0] == 4'he; // @[ifu_bp_ctl.scala 443:97]
  wire  _T_11409 = bht_wr_en0[0] & _T_11408; // @[ifu_bp_ctl.scala 443:45]
  wire  _T_11413 = _T_11409 & _T_6210; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_0_14 = _T_11413 | _T_6692; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_11425 = bht_wr_addr0[3:0] == 4'hf; // @[ifu_bp_ctl.scala 443:97]
  wire  _T_11426 = bht_wr_en0[0] & _T_11425; // @[ifu_bp_ctl.scala 443:45]
  wire  _T_11430 = _T_11426 & _T_6210; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_0_15 = _T_11430 | _T_6701; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_11447 = _T_11171 & _T_6221; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_1_0 = _T_11447 | _T_6710; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_11464 = _T_11188 & _T_6221; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_1_1 = _T_11464 | _T_6719; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_11481 = _T_11205 & _T_6221; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_1_2 = _T_11481 | _T_6728; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_11498 = _T_11222 & _T_6221; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_1_3 = _T_11498 | _T_6737; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_11515 = _T_11239 & _T_6221; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_1_4 = _T_11515 | _T_6746; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_11532 = _T_11256 & _T_6221; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_1_5 = _T_11532 | _T_6755; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_11549 = _T_11273 & _T_6221; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_1_6 = _T_11549 | _T_6764; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_11566 = _T_11290 & _T_6221; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_1_7 = _T_11566 | _T_6773; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_11583 = _T_11307 & _T_6221; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_1_8 = _T_11583 | _T_6782; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_11600 = _T_11324 & _T_6221; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_1_9 = _T_11600 | _T_6791; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_11617 = _T_11341 & _T_6221; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_1_10 = _T_11617 | _T_6800; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_11634 = _T_11358 & _T_6221; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_1_11 = _T_11634 | _T_6809; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_11651 = _T_11375 & _T_6221; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_1_12 = _T_11651 | _T_6818; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_11668 = _T_11392 & _T_6221; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_1_13 = _T_11668 | _T_6827; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_11685 = _T_11409 & _T_6221; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_1_14 = _T_11685 | _T_6836; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_11702 = _T_11426 & _T_6221; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_1_15 = _T_11702 | _T_6845; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_11719 = _T_11171 & _T_6232; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_2_0 = _T_11719 | _T_6854; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_11736 = _T_11188 & _T_6232; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_2_1 = _T_11736 | _T_6863; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_11753 = _T_11205 & _T_6232; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_2_2 = _T_11753 | _T_6872; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_11770 = _T_11222 & _T_6232; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_2_3 = _T_11770 | _T_6881; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_11787 = _T_11239 & _T_6232; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_2_4 = _T_11787 | _T_6890; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_11804 = _T_11256 & _T_6232; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_2_5 = _T_11804 | _T_6899; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_11821 = _T_11273 & _T_6232; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_2_6 = _T_11821 | _T_6908; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_11838 = _T_11290 & _T_6232; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_2_7 = _T_11838 | _T_6917; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_11855 = _T_11307 & _T_6232; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_2_8 = _T_11855 | _T_6926; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_11872 = _T_11324 & _T_6232; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_2_9 = _T_11872 | _T_6935; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_11889 = _T_11341 & _T_6232; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_2_10 = _T_11889 | _T_6944; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_11906 = _T_11358 & _T_6232; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_2_11 = _T_11906 | _T_6953; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_11923 = _T_11375 & _T_6232; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_2_12 = _T_11923 | _T_6962; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_11940 = _T_11392 & _T_6232; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_2_13 = _T_11940 | _T_6971; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_11957 = _T_11409 & _T_6232; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_2_14 = _T_11957 | _T_6980; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_11974 = _T_11426 & _T_6232; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_2_15 = _T_11974 | _T_6989; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_11991 = _T_11171 & _T_6243; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_3_0 = _T_11991 | _T_6998; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12008 = _T_11188 & _T_6243; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_3_1 = _T_12008 | _T_7007; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12025 = _T_11205 & _T_6243; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_3_2 = _T_12025 | _T_7016; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12042 = _T_11222 & _T_6243; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_3_3 = _T_12042 | _T_7025; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12059 = _T_11239 & _T_6243; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_3_4 = _T_12059 | _T_7034; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12076 = _T_11256 & _T_6243; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_3_5 = _T_12076 | _T_7043; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12093 = _T_11273 & _T_6243; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_3_6 = _T_12093 | _T_7052; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12110 = _T_11290 & _T_6243; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_3_7 = _T_12110 | _T_7061; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12127 = _T_11307 & _T_6243; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_3_8 = _T_12127 | _T_7070; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12144 = _T_11324 & _T_6243; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_3_9 = _T_12144 | _T_7079; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12161 = _T_11341 & _T_6243; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_3_10 = _T_12161 | _T_7088; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12178 = _T_11358 & _T_6243; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_3_11 = _T_12178 | _T_7097; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12195 = _T_11375 & _T_6243; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_3_12 = _T_12195 | _T_7106; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12212 = _T_11392 & _T_6243; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_3_13 = _T_12212 | _T_7115; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12229 = _T_11409 & _T_6243; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_3_14 = _T_12229 | _T_7124; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12246 = _T_11426 & _T_6243; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_3_15 = _T_12246 | _T_7133; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12263 = _T_11171 & _T_6254; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_4_0 = _T_12263 | _T_7142; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12280 = _T_11188 & _T_6254; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_4_1 = _T_12280 | _T_7151; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12297 = _T_11205 & _T_6254; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_4_2 = _T_12297 | _T_7160; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12314 = _T_11222 & _T_6254; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_4_3 = _T_12314 | _T_7169; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12331 = _T_11239 & _T_6254; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_4_4 = _T_12331 | _T_7178; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12348 = _T_11256 & _T_6254; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_4_5 = _T_12348 | _T_7187; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12365 = _T_11273 & _T_6254; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_4_6 = _T_12365 | _T_7196; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12382 = _T_11290 & _T_6254; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_4_7 = _T_12382 | _T_7205; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12399 = _T_11307 & _T_6254; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_4_8 = _T_12399 | _T_7214; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12416 = _T_11324 & _T_6254; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_4_9 = _T_12416 | _T_7223; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12433 = _T_11341 & _T_6254; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_4_10 = _T_12433 | _T_7232; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12450 = _T_11358 & _T_6254; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_4_11 = _T_12450 | _T_7241; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12467 = _T_11375 & _T_6254; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_4_12 = _T_12467 | _T_7250; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12484 = _T_11392 & _T_6254; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_4_13 = _T_12484 | _T_7259; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12501 = _T_11409 & _T_6254; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_4_14 = _T_12501 | _T_7268; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12518 = _T_11426 & _T_6254; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_4_15 = _T_12518 | _T_7277; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12535 = _T_11171 & _T_6265; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_5_0 = _T_12535 | _T_7286; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12552 = _T_11188 & _T_6265; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_5_1 = _T_12552 | _T_7295; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12569 = _T_11205 & _T_6265; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_5_2 = _T_12569 | _T_7304; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12586 = _T_11222 & _T_6265; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_5_3 = _T_12586 | _T_7313; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12603 = _T_11239 & _T_6265; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_5_4 = _T_12603 | _T_7322; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12620 = _T_11256 & _T_6265; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_5_5 = _T_12620 | _T_7331; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12637 = _T_11273 & _T_6265; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_5_6 = _T_12637 | _T_7340; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12654 = _T_11290 & _T_6265; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_5_7 = _T_12654 | _T_7349; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12671 = _T_11307 & _T_6265; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_5_8 = _T_12671 | _T_7358; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12688 = _T_11324 & _T_6265; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_5_9 = _T_12688 | _T_7367; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12705 = _T_11341 & _T_6265; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_5_10 = _T_12705 | _T_7376; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12722 = _T_11358 & _T_6265; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_5_11 = _T_12722 | _T_7385; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12739 = _T_11375 & _T_6265; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_5_12 = _T_12739 | _T_7394; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12756 = _T_11392 & _T_6265; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_5_13 = _T_12756 | _T_7403; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12773 = _T_11409 & _T_6265; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_5_14 = _T_12773 | _T_7412; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12790 = _T_11426 & _T_6265; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_5_15 = _T_12790 | _T_7421; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12807 = _T_11171 & _T_6276; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_6_0 = _T_12807 | _T_7430; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12824 = _T_11188 & _T_6276; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_6_1 = _T_12824 | _T_7439; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12841 = _T_11205 & _T_6276; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_6_2 = _T_12841 | _T_7448; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12858 = _T_11222 & _T_6276; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_6_3 = _T_12858 | _T_7457; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12875 = _T_11239 & _T_6276; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_6_4 = _T_12875 | _T_7466; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12892 = _T_11256 & _T_6276; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_6_5 = _T_12892 | _T_7475; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12909 = _T_11273 & _T_6276; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_6_6 = _T_12909 | _T_7484; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12926 = _T_11290 & _T_6276; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_6_7 = _T_12926 | _T_7493; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12943 = _T_11307 & _T_6276; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_6_8 = _T_12943 | _T_7502; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12960 = _T_11324 & _T_6276; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_6_9 = _T_12960 | _T_7511; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12977 = _T_11341 & _T_6276; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_6_10 = _T_12977 | _T_7520; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_12994 = _T_11358 & _T_6276; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_6_11 = _T_12994 | _T_7529; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13011 = _T_11375 & _T_6276; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_6_12 = _T_13011 | _T_7538; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13028 = _T_11392 & _T_6276; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_6_13 = _T_13028 | _T_7547; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13045 = _T_11409 & _T_6276; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_6_14 = _T_13045 | _T_7556; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13062 = _T_11426 & _T_6276; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_6_15 = _T_13062 | _T_7565; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13079 = _T_11171 & _T_6287; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_7_0 = _T_13079 | _T_7574; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13096 = _T_11188 & _T_6287; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_7_1 = _T_13096 | _T_7583; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13113 = _T_11205 & _T_6287; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_7_2 = _T_13113 | _T_7592; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13130 = _T_11222 & _T_6287; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_7_3 = _T_13130 | _T_7601; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13147 = _T_11239 & _T_6287; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_7_4 = _T_13147 | _T_7610; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13164 = _T_11256 & _T_6287; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_7_5 = _T_13164 | _T_7619; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13181 = _T_11273 & _T_6287; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_7_6 = _T_13181 | _T_7628; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13198 = _T_11290 & _T_6287; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_7_7 = _T_13198 | _T_7637; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13215 = _T_11307 & _T_6287; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_7_8 = _T_13215 | _T_7646; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13232 = _T_11324 & _T_6287; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_7_9 = _T_13232 | _T_7655; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13249 = _T_11341 & _T_6287; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_7_10 = _T_13249 | _T_7664; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13266 = _T_11358 & _T_6287; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_7_11 = _T_13266 | _T_7673; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13283 = _T_11375 & _T_6287; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_7_12 = _T_13283 | _T_7682; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13300 = _T_11392 & _T_6287; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_7_13 = _T_13300 | _T_7691; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13317 = _T_11409 & _T_6287; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_7_14 = _T_13317 | _T_7700; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13334 = _T_11426 & _T_6287; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_7_15 = _T_13334 | _T_7709; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13351 = _T_11171 & _T_6298; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_8_0 = _T_13351 | _T_7718; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13368 = _T_11188 & _T_6298; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_8_1 = _T_13368 | _T_7727; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13385 = _T_11205 & _T_6298; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_8_2 = _T_13385 | _T_7736; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13402 = _T_11222 & _T_6298; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_8_3 = _T_13402 | _T_7745; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13419 = _T_11239 & _T_6298; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_8_4 = _T_13419 | _T_7754; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13436 = _T_11256 & _T_6298; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_8_5 = _T_13436 | _T_7763; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13453 = _T_11273 & _T_6298; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_8_6 = _T_13453 | _T_7772; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13470 = _T_11290 & _T_6298; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_8_7 = _T_13470 | _T_7781; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13487 = _T_11307 & _T_6298; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_8_8 = _T_13487 | _T_7790; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13504 = _T_11324 & _T_6298; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_8_9 = _T_13504 | _T_7799; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13521 = _T_11341 & _T_6298; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_8_10 = _T_13521 | _T_7808; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13538 = _T_11358 & _T_6298; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_8_11 = _T_13538 | _T_7817; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13555 = _T_11375 & _T_6298; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_8_12 = _T_13555 | _T_7826; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13572 = _T_11392 & _T_6298; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_8_13 = _T_13572 | _T_7835; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13589 = _T_11409 & _T_6298; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_8_14 = _T_13589 | _T_7844; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13606 = _T_11426 & _T_6298; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_8_15 = _T_13606 | _T_7853; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13623 = _T_11171 & _T_6309; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_9_0 = _T_13623 | _T_7862; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13640 = _T_11188 & _T_6309; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_9_1 = _T_13640 | _T_7871; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13657 = _T_11205 & _T_6309; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_9_2 = _T_13657 | _T_7880; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13674 = _T_11222 & _T_6309; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_9_3 = _T_13674 | _T_7889; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13691 = _T_11239 & _T_6309; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_9_4 = _T_13691 | _T_7898; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13708 = _T_11256 & _T_6309; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_9_5 = _T_13708 | _T_7907; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13725 = _T_11273 & _T_6309; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_9_6 = _T_13725 | _T_7916; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13742 = _T_11290 & _T_6309; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_9_7 = _T_13742 | _T_7925; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13759 = _T_11307 & _T_6309; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_9_8 = _T_13759 | _T_7934; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13776 = _T_11324 & _T_6309; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_9_9 = _T_13776 | _T_7943; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13793 = _T_11341 & _T_6309; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_9_10 = _T_13793 | _T_7952; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13810 = _T_11358 & _T_6309; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_9_11 = _T_13810 | _T_7961; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13827 = _T_11375 & _T_6309; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_9_12 = _T_13827 | _T_7970; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13844 = _T_11392 & _T_6309; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_9_13 = _T_13844 | _T_7979; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13861 = _T_11409 & _T_6309; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_9_14 = _T_13861 | _T_7988; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13878 = _T_11426 & _T_6309; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_9_15 = _T_13878 | _T_7997; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13895 = _T_11171 & _T_6320; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_10_0 = _T_13895 | _T_8006; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13912 = _T_11188 & _T_6320; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_10_1 = _T_13912 | _T_8015; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13929 = _T_11205 & _T_6320; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_10_2 = _T_13929 | _T_8024; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13946 = _T_11222 & _T_6320; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_10_3 = _T_13946 | _T_8033; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13963 = _T_11239 & _T_6320; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_10_4 = _T_13963 | _T_8042; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13980 = _T_11256 & _T_6320; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_10_5 = _T_13980 | _T_8051; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_13997 = _T_11273 & _T_6320; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_10_6 = _T_13997 | _T_8060; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14014 = _T_11290 & _T_6320; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_10_7 = _T_14014 | _T_8069; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14031 = _T_11307 & _T_6320; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_10_8 = _T_14031 | _T_8078; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14048 = _T_11324 & _T_6320; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_10_9 = _T_14048 | _T_8087; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14065 = _T_11341 & _T_6320; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_10_10 = _T_14065 | _T_8096; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14082 = _T_11358 & _T_6320; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_10_11 = _T_14082 | _T_8105; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14099 = _T_11375 & _T_6320; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_10_12 = _T_14099 | _T_8114; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14116 = _T_11392 & _T_6320; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_10_13 = _T_14116 | _T_8123; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14133 = _T_11409 & _T_6320; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_10_14 = _T_14133 | _T_8132; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14150 = _T_11426 & _T_6320; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_10_15 = _T_14150 | _T_8141; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14167 = _T_11171 & _T_6331; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_11_0 = _T_14167 | _T_8150; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14184 = _T_11188 & _T_6331; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_11_1 = _T_14184 | _T_8159; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14201 = _T_11205 & _T_6331; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_11_2 = _T_14201 | _T_8168; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14218 = _T_11222 & _T_6331; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_11_3 = _T_14218 | _T_8177; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14235 = _T_11239 & _T_6331; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_11_4 = _T_14235 | _T_8186; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14252 = _T_11256 & _T_6331; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_11_5 = _T_14252 | _T_8195; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14269 = _T_11273 & _T_6331; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_11_6 = _T_14269 | _T_8204; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14286 = _T_11290 & _T_6331; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_11_7 = _T_14286 | _T_8213; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14303 = _T_11307 & _T_6331; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_11_8 = _T_14303 | _T_8222; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14320 = _T_11324 & _T_6331; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_11_9 = _T_14320 | _T_8231; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14337 = _T_11341 & _T_6331; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_11_10 = _T_14337 | _T_8240; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14354 = _T_11358 & _T_6331; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_11_11 = _T_14354 | _T_8249; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14371 = _T_11375 & _T_6331; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_11_12 = _T_14371 | _T_8258; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14388 = _T_11392 & _T_6331; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_11_13 = _T_14388 | _T_8267; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14405 = _T_11409 & _T_6331; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_11_14 = _T_14405 | _T_8276; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14422 = _T_11426 & _T_6331; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_11_15 = _T_14422 | _T_8285; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14439 = _T_11171 & _T_6342; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_12_0 = _T_14439 | _T_8294; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14456 = _T_11188 & _T_6342; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_12_1 = _T_14456 | _T_8303; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14473 = _T_11205 & _T_6342; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_12_2 = _T_14473 | _T_8312; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14490 = _T_11222 & _T_6342; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_12_3 = _T_14490 | _T_8321; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14507 = _T_11239 & _T_6342; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_12_4 = _T_14507 | _T_8330; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14524 = _T_11256 & _T_6342; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_12_5 = _T_14524 | _T_8339; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14541 = _T_11273 & _T_6342; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_12_6 = _T_14541 | _T_8348; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14558 = _T_11290 & _T_6342; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_12_7 = _T_14558 | _T_8357; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14575 = _T_11307 & _T_6342; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_12_8 = _T_14575 | _T_8366; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14592 = _T_11324 & _T_6342; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_12_9 = _T_14592 | _T_8375; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14609 = _T_11341 & _T_6342; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_12_10 = _T_14609 | _T_8384; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14626 = _T_11358 & _T_6342; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_12_11 = _T_14626 | _T_8393; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14643 = _T_11375 & _T_6342; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_12_12 = _T_14643 | _T_8402; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14660 = _T_11392 & _T_6342; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_12_13 = _T_14660 | _T_8411; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14677 = _T_11409 & _T_6342; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_12_14 = _T_14677 | _T_8420; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14694 = _T_11426 & _T_6342; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_12_15 = _T_14694 | _T_8429; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14711 = _T_11171 & _T_6353; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_13_0 = _T_14711 | _T_8438; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14728 = _T_11188 & _T_6353; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_13_1 = _T_14728 | _T_8447; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14745 = _T_11205 & _T_6353; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_13_2 = _T_14745 | _T_8456; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14762 = _T_11222 & _T_6353; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_13_3 = _T_14762 | _T_8465; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14779 = _T_11239 & _T_6353; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_13_4 = _T_14779 | _T_8474; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14796 = _T_11256 & _T_6353; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_13_5 = _T_14796 | _T_8483; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14813 = _T_11273 & _T_6353; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_13_6 = _T_14813 | _T_8492; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14830 = _T_11290 & _T_6353; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_13_7 = _T_14830 | _T_8501; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14847 = _T_11307 & _T_6353; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_13_8 = _T_14847 | _T_8510; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14864 = _T_11324 & _T_6353; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_13_9 = _T_14864 | _T_8519; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14881 = _T_11341 & _T_6353; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_13_10 = _T_14881 | _T_8528; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14898 = _T_11358 & _T_6353; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_13_11 = _T_14898 | _T_8537; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14915 = _T_11375 & _T_6353; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_13_12 = _T_14915 | _T_8546; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14932 = _T_11392 & _T_6353; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_13_13 = _T_14932 | _T_8555; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14949 = _T_11409 & _T_6353; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_13_14 = _T_14949 | _T_8564; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14966 = _T_11426 & _T_6353; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_13_15 = _T_14966 | _T_8573; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_14983 = _T_11171 & _T_6364; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_14_0 = _T_14983 | _T_8582; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15000 = _T_11188 & _T_6364; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_14_1 = _T_15000 | _T_8591; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15017 = _T_11205 & _T_6364; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_14_2 = _T_15017 | _T_8600; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15034 = _T_11222 & _T_6364; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_14_3 = _T_15034 | _T_8609; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15051 = _T_11239 & _T_6364; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_14_4 = _T_15051 | _T_8618; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15068 = _T_11256 & _T_6364; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_14_5 = _T_15068 | _T_8627; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15085 = _T_11273 & _T_6364; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_14_6 = _T_15085 | _T_8636; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15102 = _T_11290 & _T_6364; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_14_7 = _T_15102 | _T_8645; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15119 = _T_11307 & _T_6364; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_14_8 = _T_15119 | _T_8654; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15136 = _T_11324 & _T_6364; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_14_9 = _T_15136 | _T_8663; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15153 = _T_11341 & _T_6364; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_14_10 = _T_15153 | _T_8672; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15170 = _T_11358 & _T_6364; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_14_11 = _T_15170 | _T_8681; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15187 = _T_11375 & _T_6364; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_14_12 = _T_15187 | _T_8690; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15204 = _T_11392 & _T_6364; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_14_13 = _T_15204 | _T_8699; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15221 = _T_11409 & _T_6364; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_14_14 = _T_15221 | _T_8708; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15238 = _T_11426 & _T_6364; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_14_15 = _T_15238 | _T_8717; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15255 = _T_11171 & _T_6375; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_15_0 = _T_15255 | _T_8726; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15272 = _T_11188 & _T_6375; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_15_1 = _T_15272 | _T_8735; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15289 = _T_11205 & _T_6375; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_15_2 = _T_15289 | _T_8744; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15306 = _T_11222 & _T_6375; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_15_3 = _T_15306 | _T_8753; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15323 = _T_11239 & _T_6375; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_15_4 = _T_15323 | _T_8762; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15340 = _T_11256 & _T_6375; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_15_5 = _T_15340 | _T_8771; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15357 = _T_11273 & _T_6375; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_15_6 = _T_15357 | _T_8780; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15374 = _T_11290 & _T_6375; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_15_7 = _T_15374 | _T_8789; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15391 = _T_11307 & _T_6375; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_15_8 = _T_15391 | _T_8798; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15408 = _T_11324 & _T_6375; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_15_9 = _T_15408 | _T_8807; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15425 = _T_11341 & _T_6375; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_15_10 = _T_15425 | _T_8816; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15442 = _T_11358 & _T_6375; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_15_11 = _T_15442 | _T_8825; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15459 = _T_11375 & _T_6375; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_15_12 = _T_15459 | _T_8834; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15476 = _T_11392 & _T_6375; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_15_13 = _T_15476 | _T_8843; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15493 = _T_11409 & _T_6375; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_15_14 = _T_15493 | _T_8852; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15510 = _T_11426 & _T_6375; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_0_15_15 = _T_15510 | _T_8861; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15523 = bht_wr_en0[1] & _T_11170; // @[ifu_bp_ctl.scala 443:45]
  wire  _T_15527 = _T_15523 & _T_6210; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_0_0 = _T_15527 | _T_8870; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15540 = bht_wr_en0[1] & _T_11187; // @[ifu_bp_ctl.scala 443:45]
  wire  _T_15544 = _T_15540 & _T_6210; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_0_1 = _T_15544 | _T_8879; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15557 = bht_wr_en0[1] & _T_11204; // @[ifu_bp_ctl.scala 443:45]
  wire  _T_15561 = _T_15557 & _T_6210; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_0_2 = _T_15561 | _T_8888; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15574 = bht_wr_en0[1] & _T_11221; // @[ifu_bp_ctl.scala 443:45]
  wire  _T_15578 = _T_15574 & _T_6210; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_0_3 = _T_15578 | _T_8897; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15591 = bht_wr_en0[1] & _T_11238; // @[ifu_bp_ctl.scala 443:45]
  wire  _T_15595 = _T_15591 & _T_6210; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_0_4 = _T_15595 | _T_8906; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15608 = bht_wr_en0[1] & _T_11255; // @[ifu_bp_ctl.scala 443:45]
  wire  _T_15612 = _T_15608 & _T_6210; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_0_5 = _T_15612 | _T_8915; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15625 = bht_wr_en0[1] & _T_11272; // @[ifu_bp_ctl.scala 443:45]
  wire  _T_15629 = _T_15625 & _T_6210; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_0_6 = _T_15629 | _T_8924; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15642 = bht_wr_en0[1] & _T_11289; // @[ifu_bp_ctl.scala 443:45]
  wire  _T_15646 = _T_15642 & _T_6210; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_0_7 = _T_15646 | _T_8933; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15659 = bht_wr_en0[1] & _T_11306; // @[ifu_bp_ctl.scala 443:45]
  wire  _T_15663 = _T_15659 & _T_6210; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_0_8 = _T_15663 | _T_8942; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15676 = bht_wr_en0[1] & _T_11323; // @[ifu_bp_ctl.scala 443:45]
  wire  _T_15680 = _T_15676 & _T_6210; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_0_9 = _T_15680 | _T_8951; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15693 = bht_wr_en0[1] & _T_11340; // @[ifu_bp_ctl.scala 443:45]
  wire  _T_15697 = _T_15693 & _T_6210; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_0_10 = _T_15697 | _T_8960; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15710 = bht_wr_en0[1] & _T_11357; // @[ifu_bp_ctl.scala 443:45]
  wire  _T_15714 = _T_15710 & _T_6210; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_0_11 = _T_15714 | _T_8969; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15727 = bht_wr_en0[1] & _T_11374; // @[ifu_bp_ctl.scala 443:45]
  wire  _T_15731 = _T_15727 & _T_6210; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_0_12 = _T_15731 | _T_8978; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15744 = bht_wr_en0[1] & _T_11391; // @[ifu_bp_ctl.scala 443:45]
  wire  _T_15748 = _T_15744 & _T_6210; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_0_13 = _T_15748 | _T_8987; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15761 = bht_wr_en0[1] & _T_11408; // @[ifu_bp_ctl.scala 443:45]
  wire  _T_15765 = _T_15761 & _T_6210; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_0_14 = _T_15765 | _T_8996; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15778 = bht_wr_en0[1] & _T_11425; // @[ifu_bp_ctl.scala 443:45]
  wire  _T_15782 = _T_15778 & _T_6210; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_0_15 = _T_15782 | _T_9005; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15799 = _T_15523 & _T_6221; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_1_0 = _T_15799 | _T_9014; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15816 = _T_15540 & _T_6221; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_1_1 = _T_15816 | _T_9023; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15833 = _T_15557 & _T_6221; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_1_2 = _T_15833 | _T_9032; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15850 = _T_15574 & _T_6221; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_1_3 = _T_15850 | _T_9041; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15867 = _T_15591 & _T_6221; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_1_4 = _T_15867 | _T_9050; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15884 = _T_15608 & _T_6221; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_1_5 = _T_15884 | _T_9059; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15901 = _T_15625 & _T_6221; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_1_6 = _T_15901 | _T_9068; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15918 = _T_15642 & _T_6221; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_1_7 = _T_15918 | _T_9077; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15935 = _T_15659 & _T_6221; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_1_8 = _T_15935 | _T_9086; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15952 = _T_15676 & _T_6221; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_1_9 = _T_15952 | _T_9095; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15969 = _T_15693 & _T_6221; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_1_10 = _T_15969 | _T_9104; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_15986 = _T_15710 & _T_6221; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_1_11 = _T_15986 | _T_9113; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16003 = _T_15727 & _T_6221; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_1_12 = _T_16003 | _T_9122; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16020 = _T_15744 & _T_6221; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_1_13 = _T_16020 | _T_9131; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16037 = _T_15761 & _T_6221; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_1_14 = _T_16037 | _T_9140; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16054 = _T_15778 & _T_6221; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_1_15 = _T_16054 | _T_9149; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16071 = _T_15523 & _T_6232; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_2_0 = _T_16071 | _T_9158; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16088 = _T_15540 & _T_6232; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_2_1 = _T_16088 | _T_9167; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16105 = _T_15557 & _T_6232; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_2_2 = _T_16105 | _T_9176; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16122 = _T_15574 & _T_6232; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_2_3 = _T_16122 | _T_9185; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16139 = _T_15591 & _T_6232; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_2_4 = _T_16139 | _T_9194; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16156 = _T_15608 & _T_6232; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_2_5 = _T_16156 | _T_9203; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16173 = _T_15625 & _T_6232; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_2_6 = _T_16173 | _T_9212; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16190 = _T_15642 & _T_6232; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_2_7 = _T_16190 | _T_9221; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16207 = _T_15659 & _T_6232; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_2_8 = _T_16207 | _T_9230; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16224 = _T_15676 & _T_6232; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_2_9 = _T_16224 | _T_9239; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16241 = _T_15693 & _T_6232; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_2_10 = _T_16241 | _T_9248; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16258 = _T_15710 & _T_6232; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_2_11 = _T_16258 | _T_9257; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16275 = _T_15727 & _T_6232; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_2_12 = _T_16275 | _T_9266; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16292 = _T_15744 & _T_6232; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_2_13 = _T_16292 | _T_9275; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16309 = _T_15761 & _T_6232; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_2_14 = _T_16309 | _T_9284; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16326 = _T_15778 & _T_6232; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_2_15 = _T_16326 | _T_9293; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16343 = _T_15523 & _T_6243; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_3_0 = _T_16343 | _T_9302; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16360 = _T_15540 & _T_6243; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_3_1 = _T_16360 | _T_9311; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16377 = _T_15557 & _T_6243; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_3_2 = _T_16377 | _T_9320; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16394 = _T_15574 & _T_6243; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_3_3 = _T_16394 | _T_9329; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16411 = _T_15591 & _T_6243; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_3_4 = _T_16411 | _T_9338; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16428 = _T_15608 & _T_6243; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_3_5 = _T_16428 | _T_9347; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16445 = _T_15625 & _T_6243; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_3_6 = _T_16445 | _T_9356; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16462 = _T_15642 & _T_6243; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_3_7 = _T_16462 | _T_9365; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16479 = _T_15659 & _T_6243; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_3_8 = _T_16479 | _T_9374; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16496 = _T_15676 & _T_6243; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_3_9 = _T_16496 | _T_9383; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16513 = _T_15693 & _T_6243; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_3_10 = _T_16513 | _T_9392; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16530 = _T_15710 & _T_6243; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_3_11 = _T_16530 | _T_9401; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16547 = _T_15727 & _T_6243; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_3_12 = _T_16547 | _T_9410; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16564 = _T_15744 & _T_6243; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_3_13 = _T_16564 | _T_9419; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16581 = _T_15761 & _T_6243; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_3_14 = _T_16581 | _T_9428; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16598 = _T_15778 & _T_6243; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_3_15 = _T_16598 | _T_9437; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16615 = _T_15523 & _T_6254; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_4_0 = _T_16615 | _T_9446; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16632 = _T_15540 & _T_6254; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_4_1 = _T_16632 | _T_9455; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16649 = _T_15557 & _T_6254; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_4_2 = _T_16649 | _T_9464; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16666 = _T_15574 & _T_6254; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_4_3 = _T_16666 | _T_9473; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16683 = _T_15591 & _T_6254; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_4_4 = _T_16683 | _T_9482; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16700 = _T_15608 & _T_6254; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_4_5 = _T_16700 | _T_9491; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16717 = _T_15625 & _T_6254; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_4_6 = _T_16717 | _T_9500; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16734 = _T_15642 & _T_6254; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_4_7 = _T_16734 | _T_9509; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16751 = _T_15659 & _T_6254; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_4_8 = _T_16751 | _T_9518; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16768 = _T_15676 & _T_6254; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_4_9 = _T_16768 | _T_9527; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16785 = _T_15693 & _T_6254; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_4_10 = _T_16785 | _T_9536; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16802 = _T_15710 & _T_6254; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_4_11 = _T_16802 | _T_9545; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16819 = _T_15727 & _T_6254; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_4_12 = _T_16819 | _T_9554; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16836 = _T_15744 & _T_6254; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_4_13 = _T_16836 | _T_9563; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16853 = _T_15761 & _T_6254; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_4_14 = _T_16853 | _T_9572; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16870 = _T_15778 & _T_6254; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_4_15 = _T_16870 | _T_9581; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16887 = _T_15523 & _T_6265; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_5_0 = _T_16887 | _T_9590; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16904 = _T_15540 & _T_6265; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_5_1 = _T_16904 | _T_9599; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16921 = _T_15557 & _T_6265; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_5_2 = _T_16921 | _T_9608; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16938 = _T_15574 & _T_6265; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_5_3 = _T_16938 | _T_9617; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16955 = _T_15591 & _T_6265; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_5_4 = _T_16955 | _T_9626; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16972 = _T_15608 & _T_6265; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_5_5 = _T_16972 | _T_9635; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_16989 = _T_15625 & _T_6265; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_5_6 = _T_16989 | _T_9644; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17006 = _T_15642 & _T_6265; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_5_7 = _T_17006 | _T_9653; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17023 = _T_15659 & _T_6265; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_5_8 = _T_17023 | _T_9662; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17040 = _T_15676 & _T_6265; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_5_9 = _T_17040 | _T_9671; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17057 = _T_15693 & _T_6265; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_5_10 = _T_17057 | _T_9680; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17074 = _T_15710 & _T_6265; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_5_11 = _T_17074 | _T_9689; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17091 = _T_15727 & _T_6265; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_5_12 = _T_17091 | _T_9698; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17108 = _T_15744 & _T_6265; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_5_13 = _T_17108 | _T_9707; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17125 = _T_15761 & _T_6265; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_5_14 = _T_17125 | _T_9716; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17142 = _T_15778 & _T_6265; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_5_15 = _T_17142 | _T_9725; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17159 = _T_15523 & _T_6276; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_6_0 = _T_17159 | _T_9734; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17176 = _T_15540 & _T_6276; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_6_1 = _T_17176 | _T_9743; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17193 = _T_15557 & _T_6276; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_6_2 = _T_17193 | _T_9752; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17210 = _T_15574 & _T_6276; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_6_3 = _T_17210 | _T_9761; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17227 = _T_15591 & _T_6276; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_6_4 = _T_17227 | _T_9770; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17244 = _T_15608 & _T_6276; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_6_5 = _T_17244 | _T_9779; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17261 = _T_15625 & _T_6276; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_6_6 = _T_17261 | _T_9788; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17278 = _T_15642 & _T_6276; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_6_7 = _T_17278 | _T_9797; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17295 = _T_15659 & _T_6276; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_6_8 = _T_17295 | _T_9806; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17312 = _T_15676 & _T_6276; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_6_9 = _T_17312 | _T_9815; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17329 = _T_15693 & _T_6276; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_6_10 = _T_17329 | _T_9824; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17346 = _T_15710 & _T_6276; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_6_11 = _T_17346 | _T_9833; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17363 = _T_15727 & _T_6276; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_6_12 = _T_17363 | _T_9842; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17380 = _T_15744 & _T_6276; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_6_13 = _T_17380 | _T_9851; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17397 = _T_15761 & _T_6276; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_6_14 = _T_17397 | _T_9860; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17414 = _T_15778 & _T_6276; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_6_15 = _T_17414 | _T_9869; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17431 = _T_15523 & _T_6287; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_7_0 = _T_17431 | _T_9878; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17448 = _T_15540 & _T_6287; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_7_1 = _T_17448 | _T_9887; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17465 = _T_15557 & _T_6287; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_7_2 = _T_17465 | _T_9896; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17482 = _T_15574 & _T_6287; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_7_3 = _T_17482 | _T_9905; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17499 = _T_15591 & _T_6287; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_7_4 = _T_17499 | _T_9914; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17516 = _T_15608 & _T_6287; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_7_5 = _T_17516 | _T_9923; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17533 = _T_15625 & _T_6287; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_7_6 = _T_17533 | _T_9932; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17550 = _T_15642 & _T_6287; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_7_7 = _T_17550 | _T_9941; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17567 = _T_15659 & _T_6287; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_7_8 = _T_17567 | _T_9950; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17584 = _T_15676 & _T_6287; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_7_9 = _T_17584 | _T_9959; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17601 = _T_15693 & _T_6287; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_7_10 = _T_17601 | _T_9968; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17618 = _T_15710 & _T_6287; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_7_11 = _T_17618 | _T_9977; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17635 = _T_15727 & _T_6287; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_7_12 = _T_17635 | _T_9986; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17652 = _T_15744 & _T_6287; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_7_13 = _T_17652 | _T_9995; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17669 = _T_15761 & _T_6287; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_7_14 = _T_17669 | _T_10004; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17686 = _T_15778 & _T_6287; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_7_15 = _T_17686 | _T_10013; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17703 = _T_15523 & _T_6298; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_8_0 = _T_17703 | _T_10022; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17720 = _T_15540 & _T_6298; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_8_1 = _T_17720 | _T_10031; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17737 = _T_15557 & _T_6298; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_8_2 = _T_17737 | _T_10040; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17754 = _T_15574 & _T_6298; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_8_3 = _T_17754 | _T_10049; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17771 = _T_15591 & _T_6298; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_8_4 = _T_17771 | _T_10058; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17788 = _T_15608 & _T_6298; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_8_5 = _T_17788 | _T_10067; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17805 = _T_15625 & _T_6298; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_8_6 = _T_17805 | _T_10076; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17822 = _T_15642 & _T_6298; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_8_7 = _T_17822 | _T_10085; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17839 = _T_15659 & _T_6298; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_8_8 = _T_17839 | _T_10094; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17856 = _T_15676 & _T_6298; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_8_9 = _T_17856 | _T_10103; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17873 = _T_15693 & _T_6298; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_8_10 = _T_17873 | _T_10112; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17890 = _T_15710 & _T_6298; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_8_11 = _T_17890 | _T_10121; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17907 = _T_15727 & _T_6298; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_8_12 = _T_17907 | _T_10130; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17924 = _T_15744 & _T_6298; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_8_13 = _T_17924 | _T_10139; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17941 = _T_15761 & _T_6298; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_8_14 = _T_17941 | _T_10148; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17958 = _T_15778 & _T_6298; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_8_15 = _T_17958 | _T_10157; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17975 = _T_15523 & _T_6309; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_9_0 = _T_17975 | _T_10166; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_17992 = _T_15540 & _T_6309; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_9_1 = _T_17992 | _T_10175; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18009 = _T_15557 & _T_6309; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_9_2 = _T_18009 | _T_10184; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18026 = _T_15574 & _T_6309; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_9_3 = _T_18026 | _T_10193; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18043 = _T_15591 & _T_6309; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_9_4 = _T_18043 | _T_10202; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18060 = _T_15608 & _T_6309; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_9_5 = _T_18060 | _T_10211; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18077 = _T_15625 & _T_6309; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_9_6 = _T_18077 | _T_10220; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18094 = _T_15642 & _T_6309; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_9_7 = _T_18094 | _T_10229; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18111 = _T_15659 & _T_6309; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_9_8 = _T_18111 | _T_10238; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18128 = _T_15676 & _T_6309; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_9_9 = _T_18128 | _T_10247; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18145 = _T_15693 & _T_6309; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_9_10 = _T_18145 | _T_10256; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18162 = _T_15710 & _T_6309; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_9_11 = _T_18162 | _T_10265; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18179 = _T_15727 & _T_6309; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_9_12 = _T_18179 | _T_10274; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18196 = _T_15744 & _T_6309; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_9_13 = _T_18196 | _T_10283; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18213 = _T_15761 & _T_6309; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_9_14 = _T_18213 | _T_10292; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18230 = _T_15778 & _T_6309; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_9_15 = _T_18230 | _T_10301; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18247 = _T_15523 & _T_6320; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_10_0 = _T_18247 | _T_10310; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18264 = _T_15540 & _T_6320; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_10_1 = _T_18264 | _T_10319; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18281 = _T_15557 & _T_6320; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_10_2 = _T_18281 | _T_10328; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18298 = _T_15574 & _T_6320; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_10_3 = _T_18298 | _T_10337; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18315 = _T_15591 & _T_6320; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_10_4 = _T_18315 | _T_10346; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18332 = _T_15608 & _T_6320; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_10_5 = _T_18332 | _T_10355; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18349 = _T_15625 & _T_6320; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_10_6 = _T_18349 | _T_10364; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18366 = _T_15642 & _T_6320; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_10_7 = _T_18366 | _T_10373; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18383 = _T_15659 & _T_6320; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_10_8 = _T_18383 | _T_10382; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18400 = _T_15676 & _T_6320; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_10_9 = _T_18400 | _T_10391; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18417 = _T_15693 & _T_6320; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_10_10 = _T_18417 | _T_10400; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18434 = _T_15710 & _T_6320; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_10_11 = _T_18434 | _T_10409; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18451 = _T_15727 & _T_6320; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_10_12 = _T_18451 | _T_10418; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18468 = _T_15744 & _T_6320; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_10_13 = _T_18468 | _T_10427; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18485 = _T_15761 & _T_6320; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_10_14 = _T_18485 | _T_10436; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18502 = _T_15778 & _T_6320; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_10_15 = _T_18502 | _T_10445; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18519 = _T_15523 & _T_6331; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_11_0 = _T_18519 | _T_10454; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18536 = _T_15540 & _T_6331; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_11_1 = _T_18536 | _T_10463; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18553 = _T_15557 & _T_6331; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_11_2 = _T_18553 | _T_10472; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18570 = _T_15574 & _T_6331; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_11_3 = _T_18570 | _T_10481; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18587 = _T_15591 & _T_6331; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_11_4 = _T_18587 | _T_10490; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18604 = _T_15608 & _T_6331; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_11_5 = _T_18604 | _T_10499; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18621 = _T_15625 & _T_6331; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_11_6 = _T_18621 | _T_10508; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18638 = _T_15642 & _T_6331; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_11_7 = _T_18638 | _T_10517; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18655 = _T_15659 & _T_6331; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_11_8 = _T_18655 | _T_10526; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18672 = _T_15676 & _T_6331; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_11_9 = _T_18672 | _T_10535; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18689 = _T_15693 & _T_6331; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_11_10 = _T_18689 | _T_10544; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18706 = _T_15710 & _T_6331; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_11_11 = _T_18706 | _T_10553; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18723 = _T_15727 & _T_6331; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_11_12 = _T_18723 | _T_10562; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18740 = _T_15744 & _T_6331; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_11_13 = _T_18740 | _T_10571; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18757 = _T_15761 & _T_6331; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_11_14 = _T_18757 | _T_10580; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18774 = _T_15778 & _T_6331; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_11_15 = _T_18774 | _T_10589; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18791 = _T_15523 & _T_6342; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_12_0 = _T_18791 | _T_10598; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18808 = _T_15540 & _T_6342; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_12_1 = _T_18808 | _T_10607; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18825 = _T_15557 & _T_6342; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_12_2 = _T_18825 | _T_10616; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18842 = _T_15574 & _T_6342; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_12_3 = _T_18842 | _T_10625; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18859 = _T_15591 & _T_6342; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_12_4 = _T_18859 | _T_10634; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18876 = _T_15608 & _T_6342; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_12_5 = _T_18876 | _T_10643; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18893 = _T_15625 & _T_6342; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_12_6 = _T_18893 | _T_10652; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18910 = _T_15642 & _T_6342; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_12_7 = _T_18910 | _T_10661; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18927 = _T_15659 & _T_6342; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_12_8 = _T_18927 | _T_10670; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18944 = _T_15676 & _T_6342; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_12_9 = _T_18944 | _T_10679; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18961 = _T_15693 & _T_6342; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_12_10 = _T_18961 | _T_10688; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18978 = _T_15710 & _T_6342; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_12_11 = _T_18978 | _T_10697; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_18995 = _T_15727 & _T_6342; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_12_12 = _T_18995 | _T_10706; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_19012 = _T_15744 & _T_6342; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_12_13 = _T_19012 | _T_10715; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_19029 = _T_15761 & _T_6342; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_12_14 = _T_19029 | _T_10724; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_19046 = _T_15778 & _T_6342; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_12_15 = _T_19046 | _T_10733; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_19063 = _T_15523 & _T_6353; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_13_0 = _T_19063 | _T_10742; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_19080 = _T_15540 & _T_6353; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_13_1 = _T_19080 | _T_10751; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_19097 = _T_15557 & _T_6353; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_13_2 = _T_19097 | _T_10760; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_19114 = _T_15574 & _T_6353; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_13_3 = _T_19114 | _T_10769; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_19131 = _T_15591 & _T_6353; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_13_4 = _T_19131 | _T_10778; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_19148 = _T_15608 & _T_6353; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_13_5 = _T_19148 | _T_10787; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_19165 = _T_15625 & _T_6353; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_13_6 = _T_19165 | _T_10796; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_19182 = _T_15642 & _T_6353; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_13_7 = _T_19182 | _T_10805; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_19199 = _T_15659 & _T_6353; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_13_8 = _T_19199 | _T_10814; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_19216 = _T_15676 & _T_6353; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_13_9 = _T_19216 | _T_10823; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_19233 = _T_15693 & _T_6353; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_13_10 = _T_19233 | _T_10832; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_19250 = _T_15710 & _T_6353; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_13_11 = _T_19250 | _T_10841; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_19267 = _T_15727 & _T_6353; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_13_12 = _T_19267 | _T_10850; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_19284 = _T_15744 & _T_6353; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_13_13 = _T_19284 | _T_10859; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_19301 = _T_15761 & _T_6353; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_13_14 = _T_19301 | _T_10868; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_19318 = _T_15778 & _T_6353; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_13_15 = _T_19318 | _T_10877; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_19335 = _T_15523 & _T_6364; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_14_0 = _T_19335 | _T_10886; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_19352 = _T_15540 & _T_6364; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_14_1 = _T_19352 | _T_10895; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_19369 = _T_15557 & _T_6364; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_14_2 = _T_19369 | _T_10904; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_19386 = _T_15574 & _T_6364; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_14_3 = _T_19386 | _T_10913; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_19403 = _T_15591 & _T_6364; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_14_4 = _T_19403 | _T_10922; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_19420 = _T_15608 & _T_6364; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_14_5 = _T_19420 | _T_10931; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_19437 = _T_15625 & _T_6364; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_14_6 = _T_19437 | _T_10940; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_19454 = _T_15642 & _T_6364; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_14_7 = _T_19454 | _T_10949; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_19471 = _T_15659 & _T_6364; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_14_8 = _T_19471 | _T_10958; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_19488 = _T_15676 & _T_6364; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_14_9 = _T_19488 | _T_10967; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_19505 = _T_15693 & _T_6364; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_14_10 = _T_19505 | _T_10976; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_19522 = _T_15710 & _T_6364; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_14_11 = _T_19522 | _T_10985; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_19539 = _T_15727 & _T_6364; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_14_12 = _T_19539 | _T_10994; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_19556 = _T_15744 & _T_6364; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_14_13 = _T_19556 | _T_11003; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_19573 = _T_15761 & _T_6364; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_14_14 = _T_19573 | _T_11012; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_19590 = _T_15778 & _T_6364; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_14_15 = _T_19590 | _T_11021; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_19607 = _T_15523 & _T_6375; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_15_0 = _T_19607 | _T_11030; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_19624 = _T_15540 & _T_6375; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_15_1 = _T_19624 | _T_11039; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_19641 = _T_15557 & _T_6375; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_15_2 = _T_19641 | _T_11048; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_19658 = _T_15574 & _T_6375; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_15_3 = _T_19658 | _T_11057; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_19675 = _T_15591 & _T_6375; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_15_4 = _T_19675 | _T_11066; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_19692 = _T_15608 & _T_6375; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_15_5 = _T_19692 | _T_11075; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_19709 = _T_15625 & _T_6375; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_15_6 = _T_19709 | _T_11084; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_19726 = _T_15642 & _T_6375; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_15_7 = _T_19726 | _T_11093; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_19743 = _T_15659 & _T_6375; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_15_8 = _T_19743 | _T_11102; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_19760 = _T_15676 & _T_6375; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_15_9 = _T_19760 | _T_11111; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_19777 = _T_15693 & _T_6375; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_15_10 = _T_19777 | _T_11120; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_19794 = _T_15710 & _T_6375; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_15_11 = _T_19794 | _T_11129; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_19811 = _T_15727 & _T_6375; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_15_12 = _T_19811 | _T_11138; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_19828 = _T_15744 & _T_6375; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_15_13 = _T_19828 | _T_11147; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_19845 = _T_15761 & _T_6375; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_15_14 = _T_19845 | _T_11156; // @[ifu_bp_ctl.scala 443:223]
  wire  _T_19862 = _T_15778 & _T_6375; // @[ifu_bp_ctl.scala 443:110]
  wire  bht_bank_sel_1_15_15 = _T_19862 | _T_11165; // @[ifu_bp_ctl.scala 443:223]
  rvclkhdr rvclkhdr ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_io_l1clk),
    .io_clk(rvclkhdr_io_clk),
    .io_en(rvclkhdr_io_en),
    .io_scan_mode(rvclkhdr_io_scan_mode)
  );
  rvclkhdr rvclkhdr_1 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_1_io_l1clk),
    .io_clk(rvclkhdr_1_io_clk),
    .io_en(rvclkhdr_1_io_en),
    .io_scan_mode(rvclkhdr_1_io_scan_mode)
  );
  rvclkhdr rvclkhdr_2 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_2_io_l1clk),
    .io_clk(rvclkhdr_2_io_clk),
    .io_en(rvclkhdr_2_io_en),
    .io_scan_mode(rvclkhdr_2_io_scan_mode)
  );
  rvclkhdr rvclkhdr_3 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_3_io_l1clk),
    .io_clk(rvclkhdr_3_io_clk),
    .io_en(rvclkhdr_3_io_en),
    .io_scan_mode(rvclkhdr_3_io_scan_mode)
  );
  rvclkhdr rvclkhdr_4 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_4_io_l1clk),
    .io_clk(rvclkhdr_4_io_clk),
    .io_en(rvclkhdr_4_io_en),
    .io_scan_mode(rvclkhdr_4_io_scan_mode)
  );
  rvclkhdr rvclkhdr_5 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_5_io_l1clk),
    .io_clk(rvclkhdr_5_io_clk),
    .io_en(rvclkhdr_5_io_en),
    .io_scan_mode(rvclkhdr_5_io_scan_mode)
  );
  rvclkhdr rvclkhdr_6 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_6_io_l1clk),
    .io_clk(rvclkhdr_6_io_clk),
    .io_en(rvclkhdr_6_io_en),
    .io_scan_mode(rvclkhdr_6_io_scan_mode)
  );
  rvclkhdr rvclkhdr_7 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_7_io_l1clk),
    .io_clk(rvclkhdr_7_io_clk),
    .io_en(rvclkhdr_7_io_en),
    .io_scan_mode(rvclkhdr_7_io_scan_mode)
  );
  rvclkhdr rvclkhdr_8 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_8_io_l1clk),
    .io_clk(rvclkhdr_8_io_clk),
    .io_en(rvclkhdr_8_io_en),
    .io_scan_mode(rvclkhdr_8_io_scan_mode)
  );
  rvclkhdr rvclkhdr_9 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_9_io_l1clk),
    .io_clk(rvclkhdr_9_io_clk),
    .io_en(rvclkhdr_9_io_en),
    .io_scan_mode(rvclkhdr_9_io_scan_mode)
  );
  rvclkhdr rvclkhdr_10 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_10_io_l1clk),
    .io_clk(rvclkhdr_10_io_clk),
    .io_en(rvclkhdr_10_io_en),
    .io_scan_mode(rvclkhdr_10_io_scan_mode)
  );
  rvclkhdr rvclkhdr_11 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_11_io_l1clk),
    .io_clk(rvclkhdr_11_io_clk),
    .io_en(rvclkhdr_11_io_en),
    .io_scan_mode(rvclkhdr_11_io_scan_mode)
  );
  rvclkhdr rvclkhdr_12 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_12_io_l1clk),
    .io_clk(rvclkhdr_12_io_clk),
    .io_en(rvclkhdr_12_io_en),
    .io_scan_mode(rvclkhdr_12_io_scan_mode)
  );
  rvclkhdr rvclkhdr_13 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_13_io_l1clk),
    .io_clk(rvclkhdr_13_io_clk),
    .io_en(rvclkhdr_13_io_en),
    .io_scan_mode(rvclkhdr_13_io_scan_mode)
  );
  rvclkhdr rvclkhdr_14 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_14_io_l1clk),
    .io_clk(rvclkhdr_14_io_clk),
    .io_en(rvclkhdr_14_io_en),
    .io_scan_mode(rvclkhdr_14_io_scan_mode)
  );
  rvclkhdr rvclkhdr_15 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_15_io_l1clk),
    .io_clk(rvclkhdr_15_io_clk),
    .io_en(rvclkhdr_15_io_en),
    .io_scan_mode(rvclkhdr_15_io_scan_mode)
  );
  rvclkhdr rvclkhdr_16 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_16_io_l1clk),
    .io_clk(rvclkhdr_16_io_clk),
    .io_en(rvclkhdr_16_io_en),
    .io_scan_mode(rvclkhdr_16_io_scan_mode)
  );
  rvclkhdr rvclkhdr_17 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_17_io_l1clk),
    .io_clk(rvclkhdr_17_io_clk),
    .io_en(rvclkhdr_17_io_en),
    .io_scan_mode(rvclkhdr_17_io_scan_mode)
  );
  rvclkhdr rvclkhdr_18 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_18_io_l1clk),
    .io_clk(rvclkhdr_18_io_clk),
    .io_en(rvclkhdr_18_io_en),
    .io_scan_mode(rvclkhdr_18_io_scan_mode)
  );
  rvclkhdr rvclkhdr_19 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_19_io_l1clk),
    .io_clk(rvclkhdr_19_io_clk),
    .io_en(rvclkhdr_19_io_en),
    .io_scan_mode(rvclkhdr_19_io_scan_mode)
  );
  rvclkhdr rvclkhdr_20 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_20_io_l1clk),
    .io_clk(rvclkhdr_20_io_clk),
    .io_en(rvclkhdr_20_io_en),
    .io_scan_mode(rvclkhdr_20_io_scan_mode)
  );
  rvclkhdr rvclkhdr_21 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_21_io_l1clk),
    .io_clk(rvclkhdr_21_io_clk),
    .io_en(rvclkhdr_21_io_en),
    .io_scan_mode(rvclkhdr_21_io_scan_mode)
  );
  rvclkhdr rvclkhdr_22 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_22_io_l1clk),
    .io_clk(rvclkhdr_22_io_clk),
    .io_en(rvclkhdr_22_io_en),
    .io_scan_mode(rvclkhdr_22_io_scan_mode)
  );
  rvclkhdr rvclkhdr_23 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_23_io_l1clk),
    .io_clk(rvclkhdr_23_io_clk),
    .io_en(rvclkhdr_23_io_en),
    .io_scan_mode(rvclkhdr_23_io_scan_mode)
  );
  rvclkhdr rvclkhdr_24 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_24_io_l1clk),
    .io_clk(rvclkhdr_24_io_clk),
    .io_en(rvclkhdr_24_io_en),
    .io_scan_mode(rvclkhdr_24_io_scan_mode)
  );
  rvclkhdr rvclkhdr_25 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_25_io_l1clk),
    .io_clk(rvclkhdr_25_io_clk),
    .io_en(rvclkhdr_25_io_en),
    .io_scan_mode(rvclkhdr_25_io_scan_mode)
  );
  rvclkhdr rvclkhdr_26 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_26_io_l1clk),
    .io_clk(rvclkhdr_26_io_clk),
    .io_en(rvclkhdr_26_io_en),
    .io_scan_mode(rvclkhdr_26_io_scan_mode)
  );
  rvclkhdr rvclkhdr_27 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_27_io_l1clk),
    .io_clk(rvclkhdr_27_io_clk),
    .io_en(rvclkhdr_27_io_en),
    .io_scan_mode(rvclkhdr_27_io_scan_mode)
  );
  rvclkhdr rvclkhdr_28 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_28_io_l1clk),
    .io_clk(rvclkhdr_28_io_clk),
    .io_en(rvclkhdr_28_io_en),
    .io_scan_mode(rvclkhdr_28_io_scan_mode)
  );
  rvclkhdr rvclkhdr_29 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_29_io_l1clk),
    .io_clk(rvclkhdr_29_io_clk),
    .io_en(rvclkhdr_29_io_en),
    .io_scan_mode(rvclkhdr_29_io_scan_mode)
  );
  rvclkhdr rvclkhdr_30 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_30_io_l1clk),
    .io_clk(rvclkhdr_30_io_clk),
    .io_en(rvclkhdr_30_io_en),
    .io_scan_mode(rvclkhdr_30_io_scan_mode)
  );
  rvclkhdr rvclkhdr_31 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_31_io_l1clk),
    .io_clk(rvclkhdr_31_io_clk),
    .io_en(rvclkhdr_31_io_en),
    .io_scan_mode(rvclkhdr_31_io_scan_mode)
  );
  rvclkhdr rvclkhdr_32 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_32_io_l1clk),
    .io_clk(rvclkhdr_32_io_clk),
    .io_en(rvclkhdr_32_io_en),
    .io_scan_mode(rvclkhdr_32_io_scan_mode)
  );
  rvclkhdr rvclkhdr_33 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_33_io_l1clk),
    .io_clk(rvclkhdr_33_io_clk),
    .io_en(rvclkhdr_33_io_en),
    .io_scan_mode(rvclkhdr_33_io_scan_mode)
  );
  rvclkhdr rvclkhdr_34 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_34_io_l1clk),
    .io_clk(rvclkhdr_34_io_clk),
    .io_en(rvclkhdr_34_io_en),
    .io_scan_mode(rvclkhdr_34_io_scan_mode)
  );
  rvclkhdr rvclkhdr_35 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_35_io_l1clk),
    .io_clk(rvclkhdr_35_io_clk),
    .io_en(rvclkhdr_35_io_en),
    .io_scan_mode(rvclkhdr_35_io_scan_mode)
  );
  rvclkhdr rvclkhdr_36 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_36_io_l1clk),
    .io_clk(rvclkhdr_36_io_clk),
    .io_en(rvclkhdr_36_io_en),
    .io_scan_mode(rvclkhdr_36_io_scan_mode)
  );
  rvclkhdr rvclkhdr_37 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_37_io_l1clk),
    .io_clk(rvclkhdr_37_io_clk),
    .io_en(rvclkhdr_37_io_en),
    .io_scan_mode(rvclkhdr_37_io_scan_mode)
  );
  rvclkhdr rvclkhdr_38 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_38_io_l1clk),
    .io_clk(rvclkhdr_38_io_clk),
    .io_en(rvclkhdr_38_io_en),
    .io_scan_mode(rvclkhdr_38_io_scan_mode)
  );
  rvclkhdr rvclkhdr_39 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_39_io_l1clk),
    .io_clk(rvclkhdr_39_io_clk),
    .io_en(rvclkhdr_39_io_en),
    .io_scan_mode(rvclkhdr_39_io_scan_mode)
  );
  rvclkhdr rvclkhdr_40 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_40_io_l1clk),
    .io_clk(rvclkhdr_40_io_clk),
    .io_en(rvclkhdr_40_io_en),
    .io_scan_mode(rvclkhdr_40_io_scan_mode)
  );
  rvclkhdr rvclkhdr_41 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_41_io_l1clk),
    .io_clk(rvclkhdr_41_io_clk),
    .io_en(rvclkhdr_41_io_en),
    .io_scan_mode(rvclkhdr_41_io_scan_mode)
  );
  rvclkhdr rvclkhdr_42 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_42_io_l1clk),
    .io_clk(rvclkhdr_42_io_clk),
    .io_en(rvclkhdr_42_io_en),
    .io_scan_mode(rvclkhdr_42_io_scan_mode)
  );
  rvclkhdr rvclkhdr_43 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_43_io_l1clk),
    .io_clk(rvclkhdr_43_io_clk),
    .io_en(rvclkhdr_43_io_en),
    .io_scan_mode(rvclkhdr_43_io_scan_mode)
  );
  rvclkhdr rvclkhdr_44 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_44_io_l1clk),
    .io_clk(rvclkhdr_44_io_clk),
    .io_en(rvclkhdr_44_io_en),
    .io_scan_mode(rvclkhdr_44_io_scan_mode)
  );
  rvclkhdr rvclkhdr_45 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_45_io_l1clk),
    .io_clk(rvclkhdr_45_io_clk),
    .io_en(rvclkhdr_45_io_en),
    .io_scan_mode(rvclkhdr_45_io_scan_mode)
  );
  rvclkhdr rvclkhdr_46 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_46_io_l1clk),
    .io_clk(rvclkhdr_46_io_clk),
    .io_en(rvclkhdr_46_io_en),
    .io_scan_mode(rvclkhdr_46_io_scan_mode)
  );
  rvclkhdr rvclkhdr_47 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_47_io_l1clk),
    .io_clk(rvclkhdr_47_io_clk),
    .io_en(rvclkhdr_47_io_en),
    .io_scan_mode(rvclkhdr_47_io_scan_mode)
  );
  rvclkhdr rvclkhdr_48 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_48_io_l1clk),
    .io_clk(rvclkhdr_48_io_clk),
    .io_en(rvclkhdr_48_io_en),
    .io_scan_mode(rvclkhdr_48_io_scan_mode)
  );
  rvclkhdr rvclkhdr_49 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_49_io_l1clk),
    .io_clk(rvclkhdr_49_io_clk),
    .io_en(rvclkhdr_49_io_en),
    .io_scan_mode(rvclkhdr_49_io_scan_mode)
  );
  rvclkhdr rvclkhdr_50 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_50_io_l1clk),
    .io_clk(rvclkhdr_50_io_clk),
    .io_en(rvclkhdr_50_io_en),
    .io_scan_mode(rvclkhdr_50_io_scan_mode)
  );
  rvclkhdr rvclkhdr_51 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_51_io_l1clk),
    .io_clk(rvclkhdr_51_io_clk),
    .io_en(rvclkhdr_51_io_en),
    .io_scan_mode(rvclkhdr_51_io_scan_mode)
  );
  rvclkhdr rvclkhdr_52 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_52_io_l1clk),
    .io_clk(rvclkhdr_52_io_clk),
    .io_en(rvclkhdr_52_io_en),
    .io_scan_mode(rvclkhdr_52_io_scan_mode)
  );
  rvclkhdr rvclkhdr_53 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_53_io_l1clk),
    .io_clk(rvclkhdr_53_io_clk),
    .io_en(rvclkhdr_53_io_en),
    .io_scan_mode(rvclkhdr_53_io_scan_mode)
  );
  rvclkhdr rvclkhdr_54 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_54_io_l1clk),
    .io_clk(rvclkhdr_54_io_clk),
    .io_en(rvclkhdr_54_io_en),
    .io_scan_mode(rvclkhdr_54_io_scan_mode)
  );
  rvclkhdr rvclkhdr_55 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_55_io_l1clk),
    .io_clk(rvclkhdr_55_io_clk),
    .io_en(rvclkhdr_55_io_en),
    .io_scan_mode(rvclkhdr_55_io_scan_mode)
  );
  rvclkhdr rvclkhdr_56 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_56_io_l1clk),
    .io_clk(rvclkhdr_56_io_clk),
    .io_en(rvclkhdr_56_io_en),
    .io_scan_mode(rvclkhdr_56_io_scan_mode)
  );
  rvclkhdr rvclkhdr_57 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_57_io_l1clk),
    .io_clk(rvclkhdr_57_io_clk),
    .io_en(rvclkhdr_57_io_en),
    .io_scan_mode(rvclkhdr_57_io_scan_mode)
  );
  rvclkhdr rvclkhdr_58 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_58_io_l1clk),
    .io_clk(rvclkhdr_58_io_clk),
    .io_en(rvclkhdr_58_io_en),
    .io_scan_mode(rvclkhdr_58_io_scan_mode)
  );
  rvclkhdr rvclkhdr_59 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_59_io_l1clk),
    .io_clk(rvclkhdr_59_io_clk),
    .io_en(rvclkhdr_59_io_en),
    .io_scan_mode(rvclkhdr_59_io_scan_mode)
  );
  rvclkhdr rvclkhdr_60 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_60_io_l1clk),
    .io_clk(rvclkhdr_60_io_clk),
    .io_en(rvclkhdr_60_io_en),
    .io_scan_mode(rvclkhdr_60_io_scan_mode)
  );
  rvclkhdr rvclkhdr_61 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_61_io_l1clk),
    .io_clk(rvclkhdr_61_io_clk),
    .io_en(rvclkhdr_61_io_en),
    .io_scan_mode(rvclkhdr_61_io_scan_mode)
  );
  rvclkhdr rvclkhdr_62 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_62_io_l1clk),
    .io_clk(rvclkhdr_62_io_clk),
    .io_en(rvclkhdr_62_io_en),
    .io_scan_mode(rvclkhdr_62_io_scan_mode)
  );
  rvclkhdr rvclkhdr_63 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_63_io_l1clk),
    .io_clk(rvclkhdr_63_io_clk),
    .io_en(rvclkhdr_63_io_en),
    .io_scan_mode(rvclkhdr_63_io_scan_mode)
  );
  rvclkhdr rvclkhdr_64 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_64_io_l1clk),
    .io_clk(rvclkhdr_64_io_clk),
    .io_en(rvclkhdr_64_io_en),
    .io_scan_mode(rvclkhdr_64_io_scan_mode)
  );
  rvclkhdr rvclkhdr_65 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_65_io_l1clk),
    .io_clk(rvclkhdr_65_io_clk),
    .io_en(rvclkhdr_65_io_en),
    .io_scan_mode(rvclkhdr_65_io_scan_mode)
  );
  rvclkhdr rvclkhdr_66 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_66_io_l1clk),
    .io_clk(rvclkhdr_66_io_clk),
    .io_en(rvclkhdr_66_io_en),
    .io_scan_mode(rvclkhdr_66_io_scan_mode)
  );
  rvclkhdr rvclkhdr_67 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_67_io_l1clk),
    .io_clk(rvclkhdr_67_io_clk),
    .io_en(rvclkhdr_67_io_en),
    .io_scan_mode(rvclkhdr_67_io_scan_mode)
  );
  rvclkhdr rvclkhdr_68 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_68_io_l1clk),
    .io_clk(rvclkhdr_68_io_clk),
    .io_en(rvclkhdr_68_io_en),
    .io_scan_mode(rvclkhdr_68_io_scan_mode)
  );
  rvclkhdr rvclkhdr_69 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_69_io_l1clk),
    .io_clk(rvclkhdr_69_io_clk),
    .io_en(rvclkhdr_69_io_en),
    .io_scan_mode(rvclkhdr_69_io_scan_mode)
  );
  rvclkhdr rvclkhdr_70 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_70_io_l1clk),
    .io_clk(rvclkhdr_70_io_clk),
    .io_en(rvclkhdr_70_io_en),
    .io_scan_mode(rvclkhdr_70_io_scan_mode)
  );
  rvclkhdr rvclkhdr_71 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_71_io_l1clk),
    .io_clk(rvclkhdr_71_io_clk),
    .io_en(rvclkhdr_71_io_en),
    .io_scan_mode(rvclkhdr_71_io_scan_mode)
  );
  rvclkhdr rvclkhdr_72 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_72_io_l1clk),
    .io_clk(rvclkhdr_72_io_clk),
    .io_en(rvclkhdr_72_io_en),
    .io_scan_mode(rvclkhdr_72_io_scan_mode)
  );
  rvclkhdr rvclkhdr_73 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_73_io_l1clk),
    .io_clk(rvclkhdr_73_io_clk),
    .io_en(rvclkhdr_73_io_en),
    .io_scan_mode(rvclkhdr_73_io_scan_mode)
  );
  rvclkhdr rvclkhdr_74 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_74_io_l1clk),
    .io_clk(rvclkhdr_74_io_clk),
    .io_en(rvclkhdr_74_io_en),
    .io_scan_mode(rvclkhdr_74_io_scan_mode)
  );
  rvclkhdr rvclkhdr_75 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_75_io_l1clk),
    .io_clk(rvclkhdr_75_io_clk),
    .io_en(rvclkhdr_75_io_en),
    .io_scan_mode(rvclkhdr_75_io_scan_mode)
  );
  rvclkhdr rvclkhdr_76 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_76_io_l1clk),
    .io_clk(rvclkhdr_76_io_clk),
    .io_en(rvclkhdr_76_io_en),
    .io_scan_mode(rvclkhdr_76_io_scan_mode)
  );
  rvclkhdr rvclkhdr_77 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_77_io_l1clk),
    .io_clk(rvclkhdr_77_io_clk),
    .io_en(rvclkhdr_77_io_en),
    .io_scan_mode(rvclkhdr_77_io_scan_mode)
  );
  rvclkhdr rvclkhdr_78 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_78_io_l1clk),
    .io_clk(rvclkhdr_78_io_clk),
    .io_en(rvclkhdr_78_io_en),
    .io_scan_mode(rvclkhdr_78_io_scan_mode)
  );
  rvclkhdr rvclkhdr_79 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_79_io_l1clk),
    .io_clk(rvclkhdr_79_io_clk),
    .io_en(rvclkhdr_79_io_en),
    .io_scan_mode(rvclkhdr_79_io_scan_mode)
  );
  rvclkhdr rvclkhdr_80 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_80_io_l1clk),
    .io_clk(rvclkhdr_80_io_clk),
    .io_en(rvclkhdr_80_io_en),
    .io_scan_mode(rvclkhdr_80_io_scan_mode)
  );
  rvclkhdr rvclkhdr_81 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_81_io_l1clk),
    .io_clk(rvclkhdr_81_io_clk),
    .io_en(rvclkhdr_81_io_en),
    .io_scan_mode(rvclkhdr_81_io_scan_mode)
  );
  rvclkhdr rvclkhdr_82 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_82_io_l1clk),
    .io_clk(rvclkhdr_82_io_clk),
    .io_en(rvclkhdr_82_io_en),
    .io_scan_mode(rvclkhdr_82_io_scan_mode)
  );
  rvclkhdr rvclkhdr_83 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_83_io_l1clk),
    .io_clk(rvclkhdr_83_io_clk),
    .io_en(rvclkhdr_83_io_en),
    .io_scan_mode(rvclkhdr_83_io_scan_mode)
  );
  rvclkhdr rvclkhdr_84 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_84_io_l1clk),
    .io_clk(rvclkhdr_84_io_clk),
    .io_en(rvclkhdr_84_io_en),
    .io_scan_mode(rvclkhdr_84_io_scan_mode)
  );
  rvclkhdr rvclkhdr_85 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_85_io_l1clk),
    .io_clk(rvclkhdr_85_io_clk),
    .io_en(rvclkhdr_85_io_en),
    .io_scan_mode(rvclkhdr_85_io_scan_mode)
  );
  rvclkhdr rvclkhdr_86 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_86_io_l1clk),
    .io_clk(rvclkhdr_86_io_clk),
    .io_en(rvclkhdr_86_io_en),
    .io_scan_mode(rvclkhdr_86_io_scan_mode)
  );
  rvclkhdr rvclkhdr_87 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_87_io_l1clk),
    .io_clk(rvclkhdr_87_io_clk),
    .io_en(rvclkhdr_87_io_en),
    .io_scan_mode(rvclkhdr_87_io_scan_mode)
  );
  rvclkhdr rvclkhdr_88 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_88_io_l1clk),
    .io_clk(rvclkhdr_88_io_clk),
    .io_en(rvclkhdr_88_io_en),
    .io_scan_mode(rvclkhdr_88_io_scan_mode)
  );
  rvclkhdr rvclkhdr_89 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_89_io_l1clk),
    .io_clk(rvclkhdr_89_io_clk),
    .io_en(rvclkhdr_89_io_en),
    .io_scan_mode(rvclkhdr_89_io_scan_mode)
  );
  rvclkhdr rvclkhdr_90 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_90_io_l1clk),
    .io_clk(rvclkhdr_90_io_clk),
    .io_en(rvclkhdr_90_io_en),
    .io_scan_mode(rvclkhdr_90_io_scan_mode)
  );
  rvclkhdr rvclkhdr_91 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_91_io_l1clk),
    .io_clk(rvclkhdr_91_io_clk),
    .io_en(rvclkhdr_91_io_en),
    .io_scan_mode(rvclkhdr_91_io_scan_mode)
  );
  rvclkhdr rvclkhdr_92 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_92_io_l1clk),
    .io_clk(rvclkhdr_92_io_clk),
    .io_en(rvclkhdr_92_io_en),
    .io_scan_mode(rvclkhdr_92_io_scan_mode)
  );
  rvclkhdr rvclkhdr_93 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_93_io_l1clk),
    .io_clk(rvclkhdr_93_io_clk),
    .io_en(rvclkhdr_93_io_en),
    .io_scan_mode(rvclkhdr_93_io_scan_mode)
  );
  rvclkhdr rvclkhdr_94 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_94_io_l1clk),
    .io_clk(rvclkhdr_94_io_clk),
    .io_en(rvclkhdr_94_io_en),
    .io_scan_mode(rvclkhdr_94_io_scan_mode)
  );
  rvclkhdr rvclkhdr_95 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_95_io_l1clk),
    .io_clk(rvclkhdr_95_io_clk),
    .io_en(rvclkhdr_95_io_en),
    .io_scan_mode(rvclkhdr_95_io_scan_mode)
  );
  rvclkhdr rvclkhdr_96 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_96_io_l1clk),
    .io_clk(rvclkhdr_96_io_clk),
    .io_en(rvclkhdr_96_io_en),
    .io_scan_mode(rvclkhdr_96_io_scan_mode)
  );
  rvclkhdr rvclkhdr_97 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_97_io_l1clk),
    .io_clk(rvclkhdr_97_io_clk),
    .io_en(rvclkhdr_97_io_en),
    .io_scan_mode(rvclkhdr_97_io_scan_mode)
  );
  rvclkhdr rvclkhdr_98 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_98_io_l1clk),
    .io_clk(rvclkhdr_98_io_clk),
    .io_en(rvclkhdr_98_io_en),
    .io_scan_mode(rvclkhdr_98_io_scan_mode)
  );
  rvclkhdr rvclkhdr_99 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_99_io_l1clk),
    .io_clk(rvclkhdr_99_io_clk),
    .io_en(rvclkhdr_99_io_en),
    .io_scan_mode(rvclkhdr_99_io_scan_mode)
  );
  rvclkhdr rvclkhdr_100 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_100_io_l1clk),
    .io_clk(rvclkhdr_100_io_clk),
    .io_en(rvclkhdr_100_io_en),
    .io_scan_mode(rvclkhdr_100_io_scan_mode)
  );
  rvclkhdr rvclkhdr_101 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_101_io_l1clk),
    .io_clk(rvclkhdr_101_io_clk),
    .io_en(rvclkhdr_101_io_en),
    .io_scan_mode(rvclkhdr_101_io_scan_mode)
  );
  rvclkhdr rvclkhdr_102 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_102_io_l1clk),
    .io_clk(rvclkhdr_102_io_clk),
    .io_en(rvclkhdr_102_io_en),
    .io_scan_mode(rvclkhdr_102_io_scan_mode)
  );
  rvclkhdr rvclkhdr_103 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_103_io_l1clk),
    .io_clk(rvclkhdr_103_io_clk),
    .io_en(rvclkhdr_103_io_en),
    .io_scan_mode(rvclkhdr_103_io_scan_mode)
  );
  rvclkhdr rvclkhdr_104 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_104_io_l1clk),
    .io_clk(rvclkhdr_104_io_clk),
    .io_en(rvclkhdr_104_io_en),
    .io_scan_mode(rvclkhdr_104_io_scan_mode)
  );
  rvclkhdr rvclkhdr_105 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_105_io_l1clk),
    .io_clk(rvclkhdr_105_io_clk),
    .io_en(rvclkhdr_105_io_en),
    .io_scan_mode(rvclkhdr_105_io_scan_mode)
  );
  rvclkhdr rvclkhdr_106 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_106_io_l1clk),
    .io_clk(rvclkhdr_106_io_clk),
    .io_en(rvclkhdr_106_io_en),
    .io_scan_mode(rvclkhdr_106_io_scan_mode)
  );
  rvclkhdr rvclkhdr_107 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_107_io_l1clk),
    .io_clk(rvclkhdr_107_io_clk),
    .io_en(rvclkhdr_107_io_en),
    .io_scan_mode(rvclkhdr_107_io_scan_mode)
  );
  rvclkhdr rvclkhdr_108 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_108_io_l1clk),
    .io_clk(rvclkhdr_108_io_clk),
    .io_en(rvclkhdr_108_io_en),
    .io_scan_mode(rvclkhdr_108_io_scan_mode)
  );
  rvclkhdr rvclkhdr_109 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_109_io_l1clk),
    .io_clk(rvclkhdr_109_io_clk),
    .io_en(rvclkhdr_109_io_en),
    .io_scan_mode(rvclkhdr_109_io_scan_mode)
  );
  rvclkhdr rvclkhdr_110 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_110_io_l1clk),
    .io_clk(rvclkhdr_110_io_clk),
    .io_en(rvclkhdr_110_io_en),
    .io_scan_mode(rvclkhdr_110_io_scan_mode)
  );
  rvclkhdr rvclkhdr_111 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_111_io_l1clk),
    .io_clk(rvclkhdr_111_io_clk),
    .io_en(rvclkhdr_111_io_en),
    .io_scan_mode(rvclkhdr_111_io_scan_mode)
  );
  rvclkhdr rvclkhdr_112 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_112_io_l1clk),
    .io_clk(rvclkhdr_112_io_clk),
    .io_en(rvclkhdr_112_io_en),
    .io_scan_mode(rvclkhdr_112_io_scan_mode)
  );
  rvclkhdr rvclkhdr_113 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_113_io_l1clk),
    .io_clk(rvclkhdr_113_io_clk),
    .io_en(rvclkhdr_113_io_en),
    .io_scan_mode(rvclkhdr_113_io_scan_mode)
  );
  rvclkhdr rvclkhdr_114 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_114_io_l1clk),
    .io_clk(rvclkhdr_114_io_clk),
    .io_en(rvclkhdr_114_io_en),
    .io_scan_mode(rvclkhdr_114_io_scan_mode)
  );
  rvclkhdr rvclkhdr_115 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_115_io_l1clk),
    .io_clk(rvclkhdr_115_io_clk),
    .io_en(rvclkhdr_115_io_en),
    .io_scan_mode(rvclkhdr_115_io_scan_mode)
  );
  rvclkhdr rvclkhdr_116 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_116_io_l1clk),
    .io_clk(rvclkhdr_116_io_clk),
    .io_en(rvclkhdr_116_io_en),
    .io_scan_mode(rvclkhdr_116_io_scan_mode)
  );
  rvclkhdr rvclkhdr_117 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_117_io_l1clk),
    .io_clk(rvclkhdr_117_io_clk),
    .io_en(rvclkhdr_117_io_en),
    .io_scan_mode(rvclkhdr_117_io_scan_mode)
  );
  rvclkhdr rvclkhdr_118 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_118_io_l1clk),
    .io_clk(rvclkhdr_118_io_clk),
    .io_en(rvclkhdr_118_io_en),
    .io_scan_mode(rvclkhdr_118_io_scan_mode)
  );
  rvclkhdr rvclkhdr_119 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_119_io_l1clk),
    .io_clk(rvclkhdr_119_io_clk),
    .io_en(rvclkhdr_119_io_en),
    .io_scan_mode(rvclkhdr_119_io_scan_mode)
  );
  rvclkhdr rvclkhdr_120 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_120_io_l1clk),
    .io_clk(rvclkhdr_120_io_clk),
    .io_en(rvclkhdr_120_io_en),
    .io_scan_mode(rvclkhdr_120_io_scan_mode)
  );
  rvclkhdr rvclkhdr_121 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_121_io_l1clk),
    .io_clk(rvclkhdr_121_io_clk),
    .io_en(rvclkhdr_121_io_en),
    .io_scan_mode(rvclkhdr_121_io_scan_mode)
  );
  rvclkhdr rvclkhdr_122 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_122_io_l1clk),
    .io_clk(rvclkhdr_122_io_clk),
    .io_en(rvclkhdr_122_io_en),
    .io_scan_mode(rvclkhdr_122_io_scan_mode)
  );
  rvclkhdr rvclkhdr_123 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_123_io_l1clk),
    .io_clk(rvclkhdr_123_io_clk),
    .io_en(rvclkhdr_123_io_en),
    .io_scan_mode(rvclkhdr_123_io_scan_mode)
  );
  rvclkhdr rvclkhdr_124 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_124_io_l1clk),
    .io_clk(rvclkhdr_124_io_clk),
    .io_en(rvclkhdr_124_io_en),
    .io_scan_mode(rvclkhdr_124_io_scan_mode)
  );
  rvclkhdr rvclkhdr_125 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_125_io_l1clk),
    .io_clk(rvclkhdr_125_io_clk),
    .io_en(rvclkhdr_125_io_en),
    .io_scan_mode(rvclkhdr_125_io_scan_mode)
  );
  rvclkhdr rvclkhdr_126 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_126_io_l1clk),
    .io_clk(rvclkhdr_126_io_clk),
    .io_en(rvclkhdr_126_io_en),
    .io_scan_mode(rvclkhdr_126_io_scan_mode)
  );
  rvclkhdr rvclkhdr_127 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_127_io_l1clk),
    .io_clk(rvclkhdr_127_io_clk),
    .io_en(rvclkhdr_127_io_en),
    .io_scan_mode(rvclkhdr_127_io_scan_mode)
  );
  rvclkhdr rvclkhdr_128 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_128_io_l1clk),
    .io_clk(rvclkhdr_128_io_clk),
    .io_en(rvclkhdr_128_io_en),
    .io_scan_mode(rvclkhdr_128_io_scan_mode)
  );
  rvclkhdr rvclkhdr_129 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_129_io_l1clk),
    .io_clk(rvclkhdr_129_io_clk),
    .io_en(rvclkhdr_129_io_en),
    .io_scan_mode(rvclkhdr_129_io_scan_mode)
  );
  rvclkhdr rvclkhdr_130 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_130_io_l1clk),
    .io_clk(rvclkhdr_130_io_clk),
    .io_en(rvclkhdr_130_io_en),
    .io_scan_mode(rvclkhdr_130_io_scan_mode)
  );
  rvclkhdr rvclkhdr_131 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_131_io_l1clk),
    .io_clk(rvclkhdr_131_io_clk),
    .io_en(rvclkhdr_131_io_en),
    .io_scan_mode(rvclkhdr_131_io_scan_mode)
  );
  rvclkhdr rvclkhdr_132 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_132_io_l1clk),
    .io_clk(rvclkhdr_132_io_clk),
    .io_en(rvclkhdr_132_io_en),
    .io_scan_mode(rvclkhdr_132_io_scan_mode)
  );
  rvclkhdr rvclkhdr_133 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_133_io_l1clk),
    .io_clk(rvclkhdr_133_io_clk),
    .io_en(rvclkhdr_133_io_en),
    .io_scan_mode(rvclkhdr_133_io_scan_mode)
  );
  rvclkhdr rvclkhdr_134 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_134_io_l1clk),
    .io_clk(rvclkhdr_134_io_clk),
    .io_en(rvclkhdr_134_io_en),
    .io_scan_mode(rvclkhdr_134_io_scan_mode)
  );
  rvclkhdr rvclkhdr_135 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_135_io_l1clk),
    .io_clk(rvclkhdr_135_io_clk),
    .io_en(rvclkhdr_135_io_en),
    .io_scan_mode(rvclkhdr_135_io_scan_mode)
  );
  rvclkhdr rvclkhdr_136 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_136_io_l1clk),
    .io_clk(rvclkhdr_136_io_clk),
    .io_en(rvclkhdr_136_io_en),
    .io_scan_mode(rvclkhdr_136_io_scan_mode)
  );
  rvclkhdr rvclkhdr_137 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_137_io_l1clk),
    .io_clk(rvclkhdr_137_io_clk),
    .io_en(rvclkhdr_137_io_en),
    .io_scan_mode(rvclkhdr_137_io_scan_mode)
  );
  rvclkhdr rvclkhdr_138 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_138_io_l1clk),
    .io_clk(rvclkhdr_138_io_clk),
    .io_en(rvclkhdr_138_io_en),
    .io_scan_mode(rvclkhdr_138_io_scan_mode)
  );
  rvclkhdr rvclkhdr_139 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_139_io_l1clk),
    .io_clk(rvclkhdr_139_io_clk),
    .io_en(rvclkhdr_139_io_en),
    .io_scan_mode(rvclkhdr_139_io_scan_mode)
  );
  rvclkhdr rvclkhdr_140 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_140_io_l1clk),
    .io_clk(rvclkhdr_140_io_clk),
    .io_en(rvclkhdr_140_io_en),
    .io_scan_mode(rvclkhdr_140_io_scan_mode)
  );
  rvclkhdr rvclkhdr_141 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_141_io_l1clk),
    .io_clk(rvclkhdr_141_io_clk),
    .io_en(rvclkhdr_141_io_en),
    .io_scan_mode(rvclkhdr_141_io_scan_mode)
  );
  rvclkhdr rvclkhdr_142 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_142_io_l1clk),
    .io_clk(rvclkhdr_142_io_clk),
    .io_en(rvclkhdr_142_io_en),
    .io_scan_mode(rvclkhdr_142_io_scan_mode)
  );
  rvclkhdr rvclkhdr_143 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_143_io_l1clk),
    .io_clk(rvclkhdr_143_io_clk),
    .io_en(rvclkhdr_143_io_en),
    .io_scan_mode(rvclkhdr_143_io_scan_mode)
  );
  rvclkhdr rvclkhdr_144 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_144_io_l1clk),
    .io_clk(rvclkhdr_144_io_clk),
    .io_en(rvclkhdr_144_io_en),
    .io_scan_mode(rvclkhdr_144_io_scan_mode)
  );
  rvclkhdr rvclkhdr_145 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_145_io_l1clk),
    .io_clk(rvclkhdr_145_io_clk),
    .io_en(rvclkhdr_145_io_en),
    .io_scan_mode(rvclkhdr_145_io_scan_mode)
  );
  rvclkhdr rvclkhdr_146 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_146_io_l1clk),
    .io_clk(rvclkhdr_146_io_clk),
    .io_en(rvclkhdr_146_io_en),
    .io_scan_mode(rvclkhdr_146_io_scan_mode)
  );
  rvclkhdr rvclkhdr_147 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_147_io_l1clk),
    .io_clk(rvclkhdr_147_io_clk),
    .io_en(rvclkhdr_147_io_en),
    .io_scan_mode(rvclkhdr_147_io_scan_mode)
  );
  rvclkhdr rvclkhdr_148 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_148_io_l1clk),
    .io_clk(rvclkhdr_148_io_clk),
    .io_en(rvclkhdr_148_io_en),
    .io_scan_mode(rvclkhdr_148_io_scan_mode)
  );
  rvclkhdr rvclkhdr_149 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_149_io_l1clk),
    .io_clk(rvclkhdr_149_io_clk),
    .io_en(rvclkhdr_149_io_en),
    .io_scan_mode(rvclkhdr_149_io_scan_mode)
  );
  rvclkhdr rvclkhdr_150 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_150_io_l1clk),
    .io_clk(rvclkhdr_150_io_clk),
    .io_en(rvclkhdr_150_io_en),
    .io_scan_mode(rvclkhdr_150_io_scan_mode)
  );
  rvclkhdr rvclkhdr_151 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_151_io_l1clk),
    .io_clk(rvclkhdr_151_io_clk),
    .io_en(rvclkhdr_151_io_en),
    .io_scan_mode(rvclkhdr_151_io_scan_mode)
  );
  rvclkhdr rvclkhdr_152 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_152_io_l1clk),
    .io_clk(rvclkhdr_152_io_clk),
    .io_en(rvclkhdr_152_io_en),
    .io_scan_mode(rvclkhdr_152_io_scan_mode)
  );
  rvclkhdr rvclkhdr_153 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_153_io_l1clk),
    .io_clk(rvclkhdr_153_io_clk),
    .io_en(rvclkhdr_153_io_en),
    .io_scan_mode(rvclkhdr_153_io_scan_mode)
  );
  rvclkhdr rvclkhdr_154 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_154_io_l1clk),
    .io_clk(rvclkhdr_154_io_clk),
    .io_en(rvclkhdr_154_io_en),
    .io_scan_mode(rvclkhdr_154_io_scan_mode)
  );
  rvclkhdr rvclkhdr_155 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_155_io_l1clk),
    .io_clk(rvclkhdr_155_io_clk),
    .io_en(rvclkhdr_155_io_en),
    .io_scan_mode(rvclkhdr_155_io_scan_mode)
  );
  rvclkhdr rvclkhdr_156 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_156_io_l1clk),
    .io_clk(rvclkhdr_156_io_clk),
    .io_en(rvclkhdr_156_io_en),
    .io_scan_mode(rvclkhdr_156_io_scan_mode)
  );
  rvclkhdr rvclkhdr_157 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_157_io_l1clk),
    .io_clk(rvclkhdr_157_io_clk),
    .io_en(rvclkhdr_157_io_en),
    .io_scan_mode(rvclkhdr_157_io_scan_mode)
  );
  rvclkhdr rvclkhdr_158 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_158_io_l1clk),
    .io_clk(rvclkhdr_158_io_clk),
    .io_en(rvclkhdr_158_io_en),
    .io_scan_mode(rvclkhdr_158_io_scan_mode)
  );
  rvclkhdr rvclkhdr_159 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_159_io_l1clk),
    .io_clk(rvclkhdr_159_io_clk),
    .io_en(rvclkhdr_159_io_en),
    .io_scan_mode(rvclkhdr_159_io_scan_mode)
  );
  rvclkhdr rvclkhdr_160 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_160_io_l1clk),
    .io_clk(rvclkhdr_160_io_clk),
    .io_en(rvclkhdr_160_io_en),
    .io_scan_mode(rvclkhdr_160_io_scan_mode)
  );
  rvclkhdr rvclkhdr_161 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_161_io_l1clk),
    .io_clk(rvclkhdr_161_io_clk),
    .io_en(rvclkhdr_161_io_en),
    .io_scan_mode(rvclkhdr_161_io_scan_mode)
  );
  rvclkhdr rvclkhdr_162 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_162_io_l1clk),
    .io_clk(rvclkhdr_162_io_clk),
    .io_en(rvclkhdr_162_io_en),
    .io_scan_mode(rvclkhdr_162_io_scan_mode)
  );
  rvclkhdr rvclkhdr_163 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_163_io_l1clk),
    .io_clk(rvclkhdr_163_io_clk),
    .io_en(rvclkhdr_163_io_en),
    .io_scan_mode(rvclkhdr_163_io_scan_mode)
  );
  rvclkhdr rvclkhdr_164 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_164_io_l1clk),
    .io_clk(rvclkhdr_164_io_clk),
    .io_en(rvclkhdr_164_io_en),
    .io_scan_mode(rvclkhdr_164_io_scan_mode)
  );
  rvclkhdr rvclkhdr_165 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_165_io_l1clk),
    .io_clk(rvclkhdr_165_io_clk),
    .io_en(rvclkhdr_165_io_en),
    .io_scan_mode(rvclkhdr_165_io_scan_mode)
  );
  rvclkhdr rvclkhdr_166 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_166_io_l1clk),
    .io_clk(rvclkhdr_166_io_clk),
    .io_en(rvclkhdr_166_io_en),
    .io_scan_mode(rvclkhdr_166_io_scan_mode)
  );
  rvclkhdr rvclkhdr_167 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_167_io_l1clk),
    .io_clk(rvclkhdr_167_io_clk),
    .io_en(rvclkhdr_167_io_en),
    .io_scan_mode(rvclkhdr_167_io_scan_mode)
  );
  rvclkhdr rvclkhdr_168 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_168_io_l1clk),
    .io_clk(rvclkhdr_168_io_clk),
    .io_en(rvclkhdr_168_io_en),
    .io_scan_mode(rvclkhdr_168_io_scan_mode)
  );
  rvclkhdr rvclkhdr_169 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_169_io_l1clk),
    .io_clk(rvclkhdr_169_io_clk),
    .io_en(rvclkhdr_169_io_en),
    .io_scan_mode(rvclkhdr_169_io_scan_mode)
  );
  rvclkhdr rvclkhdr_170 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_170_io_l1clk),
    .io_clk(rvclkhdr_170_io_clk),
    .io_en(rvclkhdr_170_io_en),
    .io_scan_mode(rvclkhdr_170_io_scan_mode)
  );
  rvclkhdr rvclkhdr_171 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_171_io_l1clk),
    .io_clk(rvclkhdr_171_io_clk),
    .io_en(rvclkhdr_171_io_en),
    .io_scan_mode(rvclkhdr_171_io_scan_mode)
  );
  rvclkhdr rvclkhdr_172 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_172_io_l1clk),
    .io_clk(rvclkhdr_172_io_clk),
    .io_en(rvclkhdr_172_io_en),
    .io_scan_mode(rvclkhdr_172_io_scan_mode)
  );
  rvclkhdr rvclkhdr_173 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_173_io_l1clk),
    .io_clk(rvclkhdr_173_io_clk),
    .io_en(rvclkhdr_173_io_en),
    .io_scan_mode(rvclkhdr_173_io_scan_mode)
  );
  rvclkhdr rvclkhdr_174 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_174_io_l1clk),
    .io_clk(rvclkhdr_174_io_clk),
    .io_en(rvclkhdr_174_io_en),
    .io_scan_mode(rvclkhdr_174_io_scan_mode)
  );
  rvclkhdr rvclkhdr_175 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_175_io_l1clk),
    .io_clk(rvclkhdr_175_io_clk),
    .io_en(rvclkhdr_175_io_en),
    .io_scan_mode(rvclkhdr_175_io_scan_mode)
  );
  rvclkhdr rvclkhdr_176 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_176_io_l1clk),
    .io_clk(rvclkhdr_176_io_clk),
    .io_en(rvclkhdr_176_io_en),
    .io_scan_mode(rvclkhdr_176_io_scan_mode)
  );
  rvclkhdr rvclkhdr_177 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_177_io_l1clk),
    .io_clk(rvclkhdr_177_io_clk),
    .io_en(rvclkhdr_177_io_en),
    .io_scan_mode(rvclkhdr_177_io_scan_mode)
  );
  rvclkhdr rvclkhdr_178 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_178_io_l1clk),
    .io_clk(rvclkhdr_178_io_clk),
    .io_en(rvclkhdr_178_io_en),
    .io_scan_mode(rvclkhdr_178_io_scan_mode)
  );
  rvclkhdr rvclkhdr_179 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_179_io_l1clk),
    .io_clk(rvclkhdr_179_io_clk),
    .io_en(rvclkhdr_179_io_en),
    .io_scan_mode(rvclkhdr_179_io_scan_mode)
  );
  rvclkhdr rvclkhdr_180 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_180_io_l1clk),
    .io_clk(rvclkhdr_180_io_clk),
    .io_en(rvclkhdr_180_io_en),
    .io_scan_mode(rvclkhdr_180_io_scan_mode)
  );
  rvclkhdr rvclkhdr_181 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_181_io_l1clk),
    .io_clk(rvclkhdr_181_io_clk),
    .io_en(rvclkhdr_181_io_en),
    .io_scan_mode(rvclkhdr_181_io_scan_mode)
  );
  rvclkhdr rvclkhdr_182 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_182_io_l1clk),
    .io_clk(rvclkhdr_182_io_clk),
    .io_en(rvclkhdr_182_io_en),
    .io_scan_mode(rvclkhdr_182_io_scan_mode)
  );
  rvclkhdr rvclkhdr_183 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_183_io_l1clk),
    .io_clk(rvclkhdr_183_io_clk),
    .io_en(rvclkhdr_183_io_en),
    .io_scan_mode(rvclkhdr_183_io_scan_mode)
  );
  rvclkhdr rvclkhdr_184 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_184_io_l1clk),
    .io_clk(rvclkhdr_184_io_clk),
    .io_en(rvclkhdr_184_io_en),
    .io_scan_mode(rvclkhdr_184_io_scan_mode)
  );
  rvclkhdr rvclkhdr_185 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_185_io_l1clk),
    .io_clk(rvclkhdr_185_io_clk),
    .io_en(rvclkhdr_185_io_en),
    .io_scan_mode(rvclkhdr_185_io_scan_mode)
  );
  rvclkhdr rvclkhdr_186 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_186_io_l1clk),
    .io_clk(rvclkhdr_186_io_clk),
    .io_en(rvclkhdr_186_io_en),
    .io_scan_mode(rvclkhdr_186_io_scan_mode)
  );
  rvclkhdr rvclkhdr_187 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_187_io_l1clk),
    .io_clk(rvclkhdr_187_io_clk),
    .io_en(rvclkhdr_187_io_en),
    .io_scan_mode(rvclkhdr_187_io_scan_mode)
  );
  rvclkhdr rvclkhdr_188 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_188_io_l1clk),
    .io_clk(rvclkhdr_188_io_clk),
    .io_en(rvclkhdr_188_io_en),
    .io_scan_mode(rvclkhdr_188_io_scan_mode)
  );
  rvclkhdr rvclkhdr_189 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_189_io_l1clk),
    .io_clk(rvclkhdr_189_io_clk),
    .io_en(rvclkhdr_189_io_en),
    .io_scan_mode(rvclkhdr_189_io_scan_mode)
  );
  rvclkhdr rvclkhdr_190 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_190_io_l1clk),
    .io_clk(rvclkhdr_190_io_clk),
    .io_en(rvclkhdr_190_io_en),
    .io_scan_mode(rvclkhdr_190_io_scan_mode)
  );
  rvclkhdr rvclkhdr_191 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_191_io_l1clk),
    .io_clk(rvclkhdr_191_io_clk),
    .io_en(rvclkhdr_191_io_en),
    .io_scan_mode(rvclkhdr_191_io_scan_mode)
  );
  rvclkhdr rvclkhdr_192 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_192_io_l1clk),
    .io_clk(rvclkhdr_192_io_clk),
    .io_en(rvclkhdr_192_io_en),
    .io_scan_mode(rvclkhdr_192_io_scan_mode)
  );
  rvclkhdr rvclkhdr_193 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_193_io_l1clk),
    .io_clk(rvclkhdr_193_io_clk),
    .io_en(rvclkhdr_193_io_en),
    .io_scan_mode(rvclkhdr_193_io_scan_mode)
  );
  rvclkhdr rvclkhdr_194 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_194_io_l1clk),
    .io_clk(rvclkhdr_194_io_clk),
    .io_en(rvclkhdr_194_io_en),
    .io_scan_mode(rvclkhdr_194_io_scan_mode)
  );
  rvclkhdr rvclkhdr_195 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_195_io_l1clk),
    .io_clk(rvclkhdr_195_io_clk),
    .io_en(rvclkhdr_195_io_en),
    .io_scan_mode(rvclkhdr_195_io_scan_mode)
  );
  rvclkhdr rvclkhdr_196 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_196_io_l1clk),
    .io_clk(rvclkhdr_196_io_clk),
    .io_en(rvclkhdr_196_io_en),
    .io_scan_mode(rvclkhdr_196_io_scan_mode)
  );
  rvclkhdr rvclkhdr_197 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_197_io_l1clk),
    .io_clk(rvclkhdr_197_io_clk),
    .io_en(rvclkhdr_197_io_en),
    .io_scan_mode(rvclkhdr_197_io_scan_mode)
  );
  rvclkhdr rvclkhdr_198 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_198_io_l1clk),
    .io_clk(rvclkhdr_198_io_clk),
    .io_en(rvclkhdr_198_io_en),
    .io_scan_mode(rvclkhdr_198_io_scan_mode)
  );
  rvclkhdr rvclkhdr_199 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_199_io_l1clk),
    .io_clk(rvclkhdr_199_io_clk),
    .io_en(rvclkhdr_199_io_en),
    .io_scan_mode(rvclkhdr_199_io_scan_mode)
  );
  rvclkhdr rvclkhdr_200 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_200_io_l1clk),
    .io_clk(rvclkhdr_200_io_clk),
    .io_en(rvclkhdr_200_io_en),
    .io_scan_mode(rvclkhdr_200_io_scan_mode)
  );
  rvclkhdr rvclkhdr_201 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_201_io_l1clk),
    .io_clk(rvclkhdr_201_io_clk),
    .io_en(rvclkhdr_201_io_en),
    .io_scan_mode(rvclkhdr_201_io_scan_mode)
  );
  rvclkhdr rvclkhdr_202 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_202_io_l1clk),
    .io_clk(rvclkhdr_202_io_clk),
    .io_en(rvclkhdr_202_io_en),
    .io_scan_mode(rvclkhdr_202_io_scan_mode)
  );
  rvclkhdr rvclkhdr_203 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_203_io_l1clk),
    .io_clk(rvclkhdr_203_io_clk),
    .io_en(rvclkhdr_203_io_en),
    .io_scan_mode(rvclkhdr_203_io_scan_mode)
  );
  rvclkhdr rvclkhdr_204 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_204_io_l1clk),
    .io_clk(rvclkhdr_204_io_clk),
    .io_en(rvclkhdr_204_io_en),
    .io_scan_mode(rvclkhdr_204_io_scan_mode)
  );
  rvclkhdr rvclkhdr_205 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_205_io_l1clk),
    .io_clk(rvclkhdr_205_io_clk),
    .io_en(rvclkhdr_205_io_en),
    .io_scan_mode(rvclkhdr_205_io_scan_mode)
  );
  rvclkhdr rvclkhdr_206 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_206_io_l1clk),
    .io_clk(rvclkhdr_206_io_clk),
    .io_en(rvclkhdr_206_io_en),
    .io_scan_mode(rvclkhdr_206_io_scan_mode)
  );
  rvclkhdr rvclkhdr_207 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_207_io_l1clk),
    .io_clk(rvclkhdr_207_io_clk),
    .io_en(rvclkhdr_207_io_en),
    .io_scan_mode(rvclkhdr_207_io_scan_mode)
  );
  rvclkhdr rvclkhdr_208 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_208_io_l1clk),
    .io_clk(rvclkhdr_208_io_clk),
    .io_en(rvclkhdr_208_io_en),
    .io_scan_mode(rvclkhdr_208_io_scan_mode)
  );
  rvclkhdr rvclkhdr_209 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_209_io_l1clk),
    .io_clk(rvclkhdr_209_io_clk),
    .io_en(rvclkhdr_209_io_en),
    .io_scan_mode(rvclkhdr_209_io_scan_mode)
  );
  rvclkhdr rvclkhdr_210 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_210_io_l1clk),
    .io_clk(rvclkhdr_210_io_clk),
    .io_en(rvclkhdr_210_io_en),
    .io_scan_mode(rvclkhdr_210_io_scan_mode)
  );
  rvclkhdr rvclkhdr_211 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_211_io_l1clk),
    .io_clk(rvclkhdr_211_io_clk),
    .io_en(rvclkhdr_211_io_en),
    .io_scan_mode(rvclkhdr_211_io_scan_mode)
  );
  rvclkhdr rvclkhdr_212 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_212_io_l1clk),
    .io_clk(rvclkhdr_212_io_clk),
    .io_en(rvclkhdr_212_io_en),
    .io_scan_mode(rvclkhdr_212_io_scan_mode)
  );
  rvclkhdr rvclkhdr_213 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_213_io_l1clk),
    .io_clk(rvclkhdr_213_io_clk),
    .io_en(rvclkhdr_213_io_en),
    .io_scan_mode(rvclkhdr_213_io_scan_mode)
  );
  rvclkhdr rvclkhdr_214 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_214_io_l1clk),
    .io_clk(rvclkhdr_214_io_clk),
    .io_en(rvclkhdr_214_io_en),
    .io_scan_mode(rvclkhdr_214_io_scan_mode)
  );
  rvclkhdr rvclkhdr_215 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_215_io_l1clk),
    .io_clk(rvclkhdr_215_io_clk),
    .io_en(rvclkhdr_215_io_en),
    .io_scan_mode(rvclkhdr_215_io_scan_mode)
  );
  rvclkhdr rvclkhdr_216 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_216_io_l1clk),
    .io_clk(rvclkhdr_216_io_clk),
    .io_en(rvclkhdr_216_io_en),
    .io_scan_mode(rvclkhdr_216_io_scan_mode)
  );
  rvclkhdr rvclkhdr_217 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_217_io_l1clk),
    .io_clk(rvclkhdr_217_io_clk),
    .io_en(rvclkhdr_217_io_en),
    .io_scan_mode(rvclkhdr_217_io_scan_mode)
  );
  rvclkhdr rvclkhdr_218 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_218_io_l1clk),
    .io_clk(rvclkhdr_218_io_clk),
    .io_en(rvclkhdr_218_io_en),
    .io_scan_mode(rvclkhdr_218_io_scan_mode)
  );
  rvclkhdr rvclkhdr_219 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_219_io_l1clk),
    .io_clk(rvclkhdr_219_io_clk),
    .io_en(rvclkhdr_219_io_en),
    .io_scan_mode(rvclkhdr_219_io_scan_mode)
  );
  rvclkhdr rvclkhdr_220 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_220_io_l1clk),
    .io_clk(rvclkhdr_220_io_clk),
    .io_en(rvclkhdr_220_io_en),
    .io_scan_mode(rvclkhdr_220_io_scan_mode)
  );
  rvclkhdr rvclkhdr_221 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_221_io_l1clk),
    .io_clk(rvclkhdr_221_io_clk),
    .io_en(rvclkhdr_221_io_en),
    .io_scan_mode(rvclkhdr_221_io_scan_mode)
  );
  rvclkhdr rvclkhdr_222 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_222_io_l1clk),
    .io_clk(rvclkhdr_222_io_clk),
    .io_en(rvclkhdr_222_io_en),
    .io_scan_mode(rvclkhdr_222_io_scan_mode)
  );
  rvclkhdr rvclkhdr_223 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_223_io_l1clk),
    .io_clk(rvclkhdr_223_io_clk),
    .io_en(rvclkhdr_223_io_en),
    .io_scan_mode(rvclkhdr_223_io_scan_mode)
  );
  rvclkhdr rvclkhdr_224 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_224_io_l1clk),
    .io_clk(rvclkhdr_224_io_clk),
    .io_en(rvclkhdr_224_io_en),
    .io_scan_mode(rvclkhdr_224_io_scan_mode)
  );
  rvclkhdr rvclkhdr_225 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_225_io_l1clk),
    .io_clk(rvclkhdr_225_io_clk),
    .io_en(rvclkhdr_225_io_en),
    .io_scan_mode(rvclkhdr_225_io_scan_mode)
  );
  rvclkhdr rvclkhdr_226 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_226_io_l1clk),
    .io_clk(rvclkhdr_226_io_clk),
    .io_en(rvclkhdr_226_io_en),
    .io_scan_mode(rvclkhdr_226_io_scan_mode)
  );
  rvclkhdr rvclkhdr_227 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_227_io_l1clk),
    .io_clk(rvclkhdr_227_io_clk),
    .io_en(rvclkhdr_227_io_en),
    .io_scan_mode(rvclkhdr_227_io_scan_mode)
  );
  rvclkhdr rvclkhdr_228 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_228_io_l1clk),
    .io_clk(rvclkhdr_228_io_clk),
    .io_en(rvclkhdr_228_io_en),
    .io_scan_mode(rvclkhdr_228_io_scan_mode)
  );
  rvclkhdr rvclkhdr_229 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_229_io_l1clk),
    .io_clk(rvclkhdr_229_io_clk),
    .io_en(rvclkhdr_229_io_en),
    .io_scan_mode(rvclkhdr_229_io_scan_mode)
  );
  rvclkhdr rvclkhdr_230 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_230_io_l1clk),
    .io_clk(rvclkhdr_230_io_clk),
    .io_en(rvclkhdr_230_io_en),
    .io_scan_mode(rvclkhdr_230_io_scan_mode)
  );
  rvclkhdr rvclkhdr_231 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_231_io_l1clk),
    .io_clk(rvclkhdr_231_io_clk),
    .io_en(rvclkhdr_231_io_en),
    .io_scan_mode(rvclkhdr_231_io_scan_mode)
  );
  rvclkhdr rvclkhdr_232 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_232_io_l1clk),
    .io_clk(rvclkhdr_232_io_clk),
    .io_en(rvclkhdr_232_io_en),
    .io_scan_mode(rvclkhdr_232_io_scan_mode)
  );
  rvclkhdr rvclkhdr_233 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_233_io_l1clk),
    .io_clk(rvclkhdr_233_io_clk),
    .io_en(rvclkhdr_233_io_en),
    .io_scan_mode(rvclkhdr_233_io_scan_mode)
  );
  rvclkhdr rvclkhdr_234 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_234_io_l1clk),
    .io_clk(rvclkhdr_234_io_clk),
    .io_en(rvclkhdr_234_io_en),
    .io_scan_mode(rvclkhdr_234_io_scan_mode)
  );
  rvclkhdr rvclkhdr_235 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_235_io_l1clk),
    .io_clk(rvclkhdr_235_io_clk),
    .io_en(rvclkhdr_235_io_en),
    .io_scan_mode(rvclkhdr_235_io_scan_mode)
  );
  rvclkhdr rvclkhdr_236 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_236_io_l1clk),
    .io_clk(rvclkhdr_236_io_clk),
    .io_en(rvclkhdr_236_io_en),
    .io_scan_mode(rvclkhdr_236_io_scan_mode)
  );
  rvclkhdr rvclkhdr_237 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_237_io_l1clk),
    .io_clk(rvclkhdr_237_io_clk),
    .io_en(rvclkhdr_237_io_en),
    .io_scan_mode(rvclkhdr_237_io_scan_mode)
  );
  rvclkhdr rvclkhdr_238 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_238_io_l1clk),
    .io_clk(rvclkhdr_238_io_clk),
    .io_en(rvclkhdr_238_io_en),
    .io_scan_mode(rvclkhdr_238_io_scan_mode)
  );
  rvclkhdr rvclkhdr_239 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_239_io_l1clk),
    .io_clk(rvclkhdr_239_io_clk),
    .io_en(rvclkhdr_239_io_en),
    .io_scan_mode(rvclkhdr_239_io_scan_mode)
  );
  rvclkhdr rvclkhdr_240 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_240_io_l1clk),
    .io_clk(rvclkhdr_240_io_clk),
    .io_en(rvclkhdr_240_io_en),
    .io_scan_mode(rvclkhdr_240_io_scan_mode)
  );
  rvclkhdr rvclkhdr_241 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_241_io_l1clk),
    .io_clk(rvclkhdr_241_io_clk),
    .io_en(rvclkhdr_241_io_en),
    .io_scan_mode(rvclkhdr_241_io_scan_mode)
  );
  rvclkhdr rvclkhdr_242 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_242_io_l1clk),
    .io_clk(rvclkhdr_242_io_clk),
    .io_en(rvclkhdr_242_io_en),
    .io_scan_mode(rvclkhdr_242_io_scan_mode)
  );
  rvclkhdr rvclkhdr_243 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_243_io_l1clk),
    .io_clk(rvclkhdr_243_io_clk),
    .io_en(rvclkhdr_243_io_en),
    .io_scan_mode(rvclkhdr_243_io_scan_mode)
  );
  rvclkhdr rvclkhdr_244 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_244_io_l1clk),
    .io_clk(rvclkhdr_244_io_clk),
    .io_en(rvclkhdr_244_io_en),
    .io_scan_mode(rvclkhdr_244_io_scan_mode)
  );
  rvclkhdr rvclkhdr_245 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_245_io_l1clk),
    .io_clk(rvclkhdr_245_io_clk),
    .io_en(rvclkhdr_245_io_en),
    .io_scan_mode(rvclkhdr_245_io_scan_mode)
  );
  rvclkhdr rvclkhdr_246 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_246_io_l1clk),
    .io_clk(rvclkhdr_246_io_clk),
    .io_en(rvclkhdr_246_io_en),
    .io_scan_mode(rvclkhdr_246_io_scan_mode)
  );
  rvclkhdr rvclkhdr_247 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_247_io_l1clk),
    .io_clk(rvclkhdr_247_io_clk),
    .io_en(rvclkhdr_247_io_en),
    .io_scan_mode(rvclkhdr_247_io_scan_mode)
  );
  rvclkhdr rvclkhdr_248 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_248_io_l1clk),
    .io_clk(rvclkhdr_248_io_clk),
    .io_en(rvclkhdr_248_io_en),
    .io_scan_mode(rvclkhdr_248_io_scan_mode)
  );
  rvclkhdr rvclkhdr_249 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_249_io_l1clk),
    .io_clk(rvclkhdr_249_io_clk),
    .io_en(rvclkhdr_249_io_en),
    .io_scan_mode(rvclkhdr_249_io_scan_mode)
  );
  rvclkhdr rvclkhdr_250 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_250_io_l1clk),
    .io_clk(rvclkhdr_250_io_clk),
    .io_en(rvclkhdr_250_io_en),
    .io_scan_mode(rvclkhdr_250_io_scan_mode)
  );
  rvclkhdr rvclkhdr_251 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_251_io_l1clk),
    .io_clk(rvclkhdr_251_io_clk),
    .io_en(rvclkhdr_251_io_en),
    .io_scan_mode(rvclkhdr_251_io_scan_mode)
  );
  rvclkhdr rvclkhdr_252 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_252_io_l1clk),
    .io_clk(rvclkhdr_252_io_clk),
    .io_en(rvclkhdr_252_io_en),
    .io_scan_mode(rvclkhdr_252_io_scan_mode)
  );
  rvclkhdr rvclkhdr_253 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_253_io_l1clk),
    .io_clk(rvclkhdr_253_io_clk),
    .io_en(rvclkhdr_253_io_en),
    .io_scan_mode(rvclkhdr_253_io_scan_mode)
  );
  rvclkhdr rvclkhdr_254 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_254_io_l1clk),
    .io_clk(rvclkhdr_254_io_clk),
    .io_en(rvclkhdr_254_io_en),
    .io_scan_mode(rvclkhdr_254_io_scan_mode)
  );
  rvclkhdr rvclkhdr_255 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_255_io_l1clk),
    .io_clk(rvclkhdr_255_io_clk),
    .io_en(rvclkhdr_255_io_en),
    .io_scan_mode(rvclkhdr_255_io_scan_mode)
  );
  rvclkhdr rvclkhdr_256 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_256_io_l1clk),
    .io_clk(rvclkhdr_256_io_clk),
    .io_en(rvclkhdr_256_io_en),
    .io_scan_mode(rvclkhdr_256_io_scan_mode)
  );
  rvclkhdr rvclkhdr_257 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_257_io_l1clk),
    .io_clk(rvclkhdr_257_io_clk),
    .io_en(rvclkhdr_257_io_en),
    .io_scan_mode(rvclkhdr_257_io_scan_mode)
  );
  rvclkhdr rvclkhdr_258 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_258_io_l1clk),
    .io_clk(rvclkhdr_258_io_clk),
    .io_en(rvclkhdr_258_io_en),
    .io_scan_mode(rvclkhdr_258_io_scan_mode)
  );
  rvclkhdr rvclkhdr_259 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_259_io_l1clk),
    .io_clk(rvclkhdr_259_io_clk),
    .io_en(rvclkhdr_259_io_en),
    .io_scan_mode(rvclkhdr_259_io_scan_mode)
  );
  rvclkhdr rvclkhdr_260 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_260_io_l1clk),
    .io_clk(rvclkhdr_260_io_clk),
    .io_en(rvclkhdr_260_io_en),
    .io_scan_mode(rvclkhdr_260_io_scan_mode)
  );
  rvclkhdr rvclkhdr_261 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_261_io_l1clk),
    .io_clk(rvclkhdr_261_io_clk),
    .io_en(rvclkhdr_261_io_en),
    .io_scan_mode(rvclkhdr_261_io_scan_mode)
  );
  rvclkhdr rvclkhdr_262 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_262_io_l1clk),
    .io_clk(rvclkhdr_262_io_clk),
    .io_en(rvclkhdr_262_io_en),
    .io_scan_mode(rvclkhdr_262_io_scan_mode)
  );
  rvclkhdr rvclkhdr_263 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_263_io_l1clk),
    .io_clk(rvclkhdr_263_io_clk),
    .io_en(rvclkhdr_263_io_en),
    .io_scan_mode(rvclkhdr_263_io_scan_mode)
  );
  rvclkhdr rvclkhdr_264 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_264_io_l1clk),
    .io_clk(rvclkhdr_264_io_clk),
    .io_en(rvclkhdr_264_io_en),
    .io_scan_mode(rvclkhdr_264_io_scan_mode)
  );
  rvclkhdr rvclkhdr_265 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_265_io_l1clk),
    .io_clk(rvclkhdr_265_io_clk),
    .io_en(rvclkhdr_265_io_en),
    .io_scan_mode(rvclkhdr_265_io_scan_mode)
  );
  rvclkhdr rvclkhdr_266 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_266_io_l1clk),
    .io_clk(rvclkhdr_266_io_clk),
    .io_en(rvclkhdr_266_io_en),
    .io_scan_mode(rvclkhdr_266_io_scan_mode)
  );
  rvclkhdr rvclkhdr_267 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_267_io_l1clk),
    .io_clk(rvclkhdr_267_io_clk),
    .io_en(rvclkhdr_267_io_en),
    .io_scan_mode(rvclkhdr_267_io_scan_mode)
  );
  rvclkhdr rvclkhdr_268 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_268_io_l1clk),
    .io_clk(rvclkhdr_268_io_clk),
    .io_en(rvclkhdr_268_io_en),
    .io_scan_mode(rvclkhdr_268_io_scan_mode)
  );
  rvclkhdr rvclkhdr_269 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_269_io_l1clk),
    .io_clk(rvclkhdr_269_io_clk),
    .io_en(rvclkhdr_269_io_en),
    .io_scan_mode(rvclkhdr_269_io_scan_mode)
  );
  rvclkhdr rvclkhdr_270 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_270_io_l1clk),
    .io_clk(rvclkhdr_270_io_clk),
    .io_en(rvclkhdr_270_io_en),
    .io_scan_mode(rvclkhdr_270_io_scan_mode)
  );
  rvclkhdr rvclkhdr_271 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_271_io_l1clk),
    .io_clk(rvclkhdr_271_io_clk),
    .io_en(rvclkhdr_271_io_en),
    .io_scan_mode(rvclkhdr_271_io_scan_mode)
  );
  rvclkhdr rvclkhdr_272 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_272_io_l1clk),
    .io_clk(rvclkhdr_272_io_clk),
    .io_en(rvclkhdr_272_io_en),
    .io_scan_mode(rvclkhdr_272_io_scan_mode)
  );
  rvclkhdr rvclkhdr_273 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_273_io_l1clk),
    .io_clk(rvclkhdr_273_io_clk),
    .io_en(rvclkhdr_273_io_en),
    .io_scan_mode(rvclkhdr_273_io_scan_mode)
  );
  rvclkhdr rvclkhdr_274 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_274_io_l1clk),
    .io_clk(rvclkhdr_274_io_clk),
    .io_en(rvclkhdr_274_io_en),
    .io_scan_mode(rvclkhdr_274_io_scan_mode)
  );
  rvclkhdr rvclkhdr_275 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_275_io_l1clk),
    .io_clk(rvclkhdr_275_io_clk),
    .io_en(rvclkhdr_275_io_en),
    .io_scan_mode(rvclkhdr_275_io_scan_mode)
  );
  rvclkhdr rvclkhdr_276 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_276_io_l1clk),
    .io_clk(rvclkhdr_276_io_clk),
    .io_en(rvclkhdr_276_io_en),
    .io_scan_mode(rvclkhdr_276_io_scan_mode)
  );
  rvclkhdr rvclkhdr_277 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_277_io_l1clk),
    .io_clk(rvclkhdr_277_io_clk),
    .io_en(rvclkhdr_277_io_en),
    .io_scan_mode(rvclkhdr_277_io_scan_mode)
  );
  rvclkhdr rvclkhdr_278 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_278_io_l1clk),
    .io_clk(rvclkhdr_278_io_clk),
    .io_en(rvclkhdr_278_io_en),
    .io_scan_mode(rvclkhdr_278_io_scan_mode)
  );
  rvclkhdr rvclkhdr_279 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_279_io_l1clk),
    .io_clk(rvclkhdr_279_io_clk),
    .io_en(rvclkhdr_279_io_en),
    .io_scan_mode(rvclkhdr_279_io_scan_mode)
  );
  rvclkhdr rvclkhdr_280 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_280_io_l1clk),
    .io_clk(rvclkhdr_280_io_clk),
    .io_en(rvclkhdr_280_io_en),
    .io_scan_mode(rvclkhdr_280_io_scan_mode)
  );
  rvclkhdr rvclkhdr_281 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_281_io_l1clk),
    .io_clk(rvclkhdr_281_io_clk),
    .io_en(rvclkhdr_281_io_en),
    .io_scan_mode(rvclkhdr_281_io_scan_mode)
  );
  rvclkhdr rvclkhdr_282 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_282_io_l1clk),
    .io_clk(rvclkhdr_282_io_clk),
    .io_en(rvclkhdr_282_io_en),
    .io_scan_mode(rvclkhdr_282_io_scan_mode)
  );
  rvclkhdr rvclkhdr_283 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_283_io_l1clk),
    .io_clk(rvclkhdr_283_io_clk),
    .io_en(rvclkhdr_283_io_en),
    .io_scan_mode(rvclkhdr_283_io_scan_mode)
  );
  rvclkhdr rvclkhdr_284 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_284_io_l1clk),
    .io_clk(rvclkhdr_284_io_clk),
    .io_en(rvclkhdr_284_io_en),
    .io_scan_mode(rvclkhdr_284_io_scan_mode)
  );
  rvclkhdr rvclkhdr_285 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_285_io_l1clk),
    .io_clk(rvclkhdr_285_io_clk),
    .io_en(rvclkhdr_285_io_en),
    .io_scan_mode(rvclkhdr_285_io_scan_mode)
  );
  rvclkhdr rvclkhdr_286 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_286_io_l1clk),
    .io_clk(rvclkhdr_286_io_clk),
    .io_en(rvclkhdr_286_io_en),
    .io_scan_mode(rvclkhdr_286_io_scan_mode)
  );
  rvclkhdr rvclkhdr_287 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_287_io_l1clk),
    .io_clk(rvclkhdr_287_io_clk),
    .io_en(rvclkhdr_287_io_en),
    .io_scan_mode(rvclkhdr_287_io_scan_mode)
  );
  rvclkhdr rvclkhdr_288 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_288_io_l1clk),
    .io_clk(rvclkhdr_288_io_clk),
    .io_en(rvclkhdr_288_io_en),
    .io_scan_mode(rvclkhdr_288_io_scan_mode)
  );
  rvclkhdr rvclkhdr_289 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_289_io_l1clk),
    .io_clk(rvclkhdr_289_io_clk),
    .io_en(rvclkhdr_289_io_en),
    .io_scan_mode(rvclkhdr_289_io_scan_mode)
  );
  rvclkhdr rvclkhdr_290 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_290_io_l1clk),
    .io_clk(rvclkhdr_290_io_clk),
    .io_en(rvclkhdr_290_io_en),
    .io_scan_mode(rvclkhdr_290_io_scan_mode)
  );
  rvclkhdr rvclkhdr_291 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_291_io_l1clk),
    .io_clk(rvclkhdr_291_io_clk),
    .io_en(rvclkhdr_291_io_en),
    .io_scan_mode(rvclkhdr_291_io_scan_mode)
  );
  rvclkhdr rvclkhdr_292 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_292_io_l1clk),
    .io_clk(rvclkhdr_292_io_clk),
    .io_en(rvclkhdr_292_io_en),
    .io_scan_mode(rvclkhdr_292_io_scan_mode)
  );
  rvclkhdr rvclkhdr_293 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_293_io_l1clk),
    .io_clk(rvclkhdr_293_io_clk),
    .io_en(rvclkhdr_293_io_en),
    .io_scan_mode(rvclkhdr_293_io_scan_mode)
  );
  rvclkhdr rvclkhdr_294 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_294_io_l1clk),
    .io_clk(rvclkhdr_294_io_clk),
    .io_en(rvclkhdr_294_io_en),
    .io_scan_mode(rvclkhdr_294_io_scan_mode)
  );
  rvclkhdr rvclkhdr_295 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_295_io_l1clk),
    .io_clk(rvclkhdr_295_io_clk),
    .io_en(rvclkhdr_295_io_en),
    .io_scan_mode(rvclkhdr_295_io_scan_mode)
  );
  rvclkhdr rvclkhdr_296 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_296_io_l1clk),
    .io_clk(rvclkhdr_296_io_clk),
    .io_en(rvclkhdr_296_io_en),
    .io_scan_mode(rvclkhdr_296_io_scan_mode)
  );
  rvclkhdr rvclkhdr_297 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_297_io_l1clk),
    .io_clk(rvclkhdr_297_io_clk),
    .io_en(rvclkhdr_297_io_en),
    .io_scan_mode(rvclkhdr_297_io_scan_mode)
  );
  rvclkhdr rvclkhdr_298 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_298_io_l1clk),
    .io_clk(rvclkhdr_298_io_clk),
    .io_en(rvclkhdr_298_io_en),
    .io_scan_mode(rvclkhdr_298_io_scan_mode)
  );
  rvclkhdr rvclkhdr_299 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_299_io_l1clk),
    .io_clk(rvclkhdr_299_io_clk),
    .io_en(rvclkhdr_299_io_en),
    .io_scan_mode(rvclkhdr_299_io_scan_mode)
  );
  rvclkhdr rvclkhdr_300 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_300_io_l1clk),
    .io_clk(rvclkhdr_300_io_clk),
    .io_en(rvclkhdr_300_io_en),
    .io_scan_mode(rvclkhdr_300_io_scan_mode)
  );
  rvclkhdr rvclkhdr_301 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_301_io_l1clk),
    .io_clk(rvclkhdr_301_io_clk),
    .io_en(rvclkhdr_301_io_en),
    .io_scan_mode(rvclkhdr_301_io_scan_mode)
  );
  rvclkhdr rvclkhdr_302 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_302_io_l1clk),
    .io_clk(rvclkhdr_302_io_clk),
    .io_en(rvclkhdr_302_io_en),
    .io_scan_mode(rvclkhdr_302_io_scan_mode)
  );
  rvclkhdr rvclkhdr_303 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_303_io_l1clk),
    .io_clk(rvclkhdr_303_io_clk),
    .io_en(rvclkhdr_303_io_en),
    .io_scan_mode(rvclkhdr_303_io_scan_mode)
  );
  rvclkhdr rvclkhdr_304 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_304_io_l1clk),
    .io_clk(rvclkhdr_304_io_clk),
    .io_en(rvclkhdr_304_io_en),
    .io_scan_mode(rvclkhdr_304_io_scan_mode)
  );
  rvclkhdr rvclkhdr_305 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_305_io_l1clk),
    .io_clk(rvclkhdr_305_io_clk),
    .io_en(rvclkhdr_305_io_en),
    .io_scan_mode(rvclkhdr_305_io_scan_mode)
  );
  rvclkhdr rvclkhdr_306 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_306_io_l1clk),
    .io_clk(rvclkhdr_306_io_clk),
    .io_en(rvclkhdr_306_io_en),
    .io_scan_mode(rvclkhdr_306_io_scan_mode)
  );
  rvclkhdr rvclkhdr_307 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_307_io_l1clk),
    .io_clk(rvclkhdr_307_io_clk),
    .io_en(rvclkhdr_307_io_en),
    .io_scan_mode(rvclkhdr_307_io_scan_mode)
  );
  rvclkhdr rvclkhdr_308 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_308_io_l1clk),
    .io_clk(rvclkhdr_308_io_clk),
    .io_en(rvclkhdr_308_io_en),
    .io_scan_mode(rvclkhdr_308_io_scan_mode)
  );
  rvclkhdr rvclkhdr_309 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_309_io_l1clk),
    .io_clk(rvclkhdr_309_io_clk),
    .io_en(rvclkhdr_309_io_en),
    .io_scan_mode(rvclkhdr_309_io_scan_mode)
  );
  rvclkhdr rvclkhdr_310 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_310_io_l1clk),
    .io_clk(rvclkhdr_310_io_clk),
    .io_en(rvclkhdr_310_io_en),
    .io_scan_mode(rvclkhdr_310_io_scan_mode)
  );
  rvclkhdr rvclkhdr_311 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_311_io_l1clk),
    .io_clk(rvclkhdr_311_io_clk),
    .io_en(rvclkhdr_311_io_en),
    .io_scan_mode(rvclkhdr_311_io_scan_mode)
  );
  rvclkhdr rvclkhdr_312 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_312_io_l1clk),
    .io_clk(rvclkhdr_312_io_clk),
    .io_en(rvclkhdr_312_io_en),
    .io_scan_mode(rvclkhdr_312_io_scan_mode)
  );
  rvclkhdr rvclkhdr_313 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_313_io_l1clk),
    .io_clk(rvclkhdr_313_io_clk),
    .io_en(rvclkhdr_313_io_en),
    .io_scan_mode(rvclkhdr_313_io_scan_mode)
  );
  rvclkhdr rvclkhdr_314 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_314_io_l1clk),
    .io_clk(rvclkhdr_314_io_clk),
    .io_en(rvclkhdr_314_io_en),
    .io_scan_mode(rvclkhdr_314_io_scan_mode)
  );
  rvclkhdr rvclkhdr_315 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_315_io_l1clk),
    .io_clk(rvclkhdr_315_io_clk),
    .io_en(rvclkhdr_315_io_en),
    .io_scan_mode(rvclkhdr_315_io_scan_mode)
  );
  rvclkhdr rvclkhdr_316 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_316_io_l1clk),
    .io_clk(rvclkhdr_316_io_clk),
    .io_en(rvclkhdr_316_io_en),
    .io_scan_mode(rvclkhdr_316_io_scan_mode)
  );
  rvclkhdr rvclkhdr_317 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_317_io_l1clk),
    .io_clk(rvclkhdr_317_io_clk),
    .io_en(rvclkhdr_317_io_en),
    .io_scan_mode(rvclkhdr_317_io_scan_mode)
  );
  rvclkhdr rvclkhdr_318 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_318_io_l1clk),
    .io_clk(rvclkhdr_318_io_clk),
    .io_en(rvclkhdr_318_io_en),
    .io_scan_mode(rvclkhdr_318_io_scan_mode)
  );
  rvclkhdr rvclkhdr_319 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_319_io_l1clk),
    .io_clk(rvclkhdr_319_io_clk),
    .io_en(rvclkhdr_319_io_en),
    .io_scan_mode(rvclkhdr_319_io_scan_mode)
  );
  rvclkhdr rvclkhdr_320 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_320_io_l1clk),
    .io_clk(rvclkhdr_320_io_clk),
    .io_en(rvclkhdr_320_io_en),
    .io_scan_mode(rvclkhdr_320_io_scan_mode)
  );
  rvclkhdr rvclkhdr_321 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_321_io_l1clk),
    .io_clk(rvclkhdr_321_io_clk),
    .io_en(rvclkhdr_321_io_en),
    .io_scan_mode(rvclkhdr_321_io_scan_mode)
  );
  rvclkhdr rvclkhdr_322 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_322_io_l1clk),
    .io_clk(rvclkhdr_322_io_clk),
    .io_en(rvclkhdr_322_io_en),
    .io_scan_mode(rvclkhdr_322_io_scan_mode)
  );
  rvclkhdr rvclkhdr_323 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_323_io_l1clk),
    .io_clk(rvclkhdr_323_io_clk),
    .io_en(rvclkhdr_323_io_en),
    .io_scan_mode(rvclkhdr_323_io_scan_mode)
  );
  rvclkhdr rvclkhdr_324 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_324_io_l1clk),
    .io_clk(rvclkhdr_324_io_clk),
    .io_en(rvclkhdr_324_io_en),
    .io_scan_mode(rvclkhdr_324_io_scan_mode)
  );
  rvclkhdr rvclkhdr_325 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_325_io_l1clk),
    .io_clk(rvclkhdr_325_io_clk),
    .io_en(rvclkhdr_325_io_en),
    .io_scan_mode(rvclkhdr_325_io_scan_mode)
  );
  rvclkhdr rvclkhdr_326 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_326_io_l1clk),
    .io_clk(rvclkhdr_326_io_clk),
    .io_en(rvclkhdr_326_io_en),
    .io_scan_mode(rvclkhdr_326_io_scan_mode)
  );
  rvclkhdr rvclkhdr_327 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_327_io_l1clk),
    .io_clk(rvclkhdr_327_io_clk),
    .io_en(rvclkhdr_327_io_en),
    .io_scan_mode(rvclkhdr_327_io_scan_mode)
  );
  rvclkhdr rvclkhdr_328 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_328_io_l1clk),
    .io_clk(rvclkhdr_328_io_clk),
    .io_en(rvclkhdr_328_io_en),
    .io_scan_mode(rvclkhdr_328_io_scan_mode)
  );
  rvclkhdr rvclkhdr_329 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_329_io_l1clk),
    .io_clk(rvclkhdr_329_io_clk),
    .io_en(rvclkhdr_329_io_en),
    .io_scan_mode(rvclkhdr_329_io_scan_mode)
  );
  rvclkhdr rvclkhdr_330 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_330_io_l1clk),
    .io_clk(rvclkhdr_330_io_clk),
    .io_en(rvclkhdr_330_io_en),
    .io_scan_mode(rvclkhdr_330_io_scan_mode)
  );
  rvclkhdr rvclkhdr_331 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_331_io_l1clk),
    .io_clk(rvclkhdr_331_io_clk),
    .io_en(rvclkhdr_331_io_en),
    .io_scan_mode(rvclkhdr_331_io_scan_mode)
  );
  rvclkhdr rvclkhdr_332 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_332_io_l1clk),
    .io_clk(rvclkhdr_332_io_clk),
    .io_en(rvclkhdr_332_io_en),
    .io_scan_mode(rvclkhdr_332_io_scan_mode)
  );
  rvclkhdr rvclkhdr_333 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_333_io_l1clk),
    .io_clk(rvclkhdr_333_io_clk),
    .io_en(rvclkhdr_333_io_en),
    .io_scan_mode(rvclkhdr_333_io_scan_mode)
  );
  rvclkhdr rvclkhdr_334 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_334_io_l1clk),
    .io_clk(rvclkhdr_334_io_clk),
    .io_en(rvclkhdr_334_io_en),
    .io_scan_mode(rvclkhdr_334_io_scan_mode)
  );
  rvclkhdr rvclkhdr_335 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_335_io_l1clk),
    .io_clk(rvclkhdr_335_io_clk),
    .io_en(rvclkhdr_335_io_en),
    .io_scan_mode(rvclkhdr_335_io_scan_mode)
  );
  rvclkhdr rvclkhdr_336 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_336_io_l1clk),
    .io_clk(rvclkhdr_336_io_clk),
    .io_en(rvclkhdr_336_io_en),
    .io_scan_mode(rvclkhdr_336_io_scan_mode)
  );
  rvclkhdr rvclkhdr_337 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_337_io_l1clk),
    .io_clk(rvclkhdr_337_io_clk),
    .io_en(rvclkhdr_337_io_en),
    .io_scan_mode(rvclkhdr_337_io_scan_mode)
  );
  rvclkhdr rvclkhdr_338 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_338_io_l1clk),
    .io_clk(rvclkhdr_338_io_clk),
    .io_en(rvclkhdr_338_io_en),
    .io_scan_mode(rvclkhdr_338_io_scan_mode)
  );
  rvclkhdr rvclkhdr_339 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_339_io_l1clk),
    .io_clk(rvclkhdr_339_io_clk),
    .io_en(rvclkhdr_339_io_en),
    .io_scan_mode(rvclkhdr_339_io_scan_mode)
  );
  rvclkhdr rvclkhdr_340 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_340_io_l1clk),
    .io_clk(rvclkhdr_340_io_clk),
    .io_en(rvclkhdr_340_io_en),
    .io_scan_mode(rvclkhdr_340_io_scan_mode)
  );
  rvclkhdr rvclkhdr_341 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_341_io_l1clk),
    .io_clk(rvclkhdr_341_io_clk),
    .io_en(rvclkhdr_341_io_en),
    .io_scan_mode(rvclkhdr_341_io_scan_mode)
  );
  rvclkhdr rvclkhdr_342 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_342_io_l1clk),
    .io_clk(rvclkhdr_342_io_clk),
    .io_en(rvclkhdr_342_io_en),
    .io_scan_mode(rvclkhdr_342_io_scan_mode)
  );
  rvclkhdr rvclkhdr_343 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_343_io_l1clk),
    .io_clk(rvclkhdr_343_io_clk),
    .io_en(rvclkhdr_343_io_en),
    .io_scan_mode(rvclkhdr_343_io_scan_mode)
  );
  rvclkhdr rvclkhdr_344 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_344_io_l1clk),
    .io_clk(rvclkhdr_344_io_clk),
    .io_en(rvclkhdr_344_io_en),
    .io_scan_mode(rvclkhdr_344_io_scan_mode)
  );
  rvclkhdr rvclkhdr_345 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_345_io_l1clk),
    .io_clk(rvclkhdr_345_io_clk),
    .io_en(rvclkhdr_345_io_en),
    .io_scan_mode(rvclkhdr_345_io_scan_mode)
  );
  rvclkhdr rvclkhdr_346 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_346_io_l1clk),
    .io_clk(rvclkhdr_346_io_clk),
    .io_en(rvclkhdr_346_io_en),
    .io_scan_mode(rvclkhdr_346_io_scan_mode)
  );
  rvclkhdr rvclkhdr_347 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_347_io_l1clk),
    .io_clk(rvclkhdr_347_io_clk),
    .io_en(rvclkhdr_347_io_en),
    .io_scan_mode(rvclkhdr_347_io_scan_mode)
  );
  rvclkhdr rvclkhdr_348 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_348_io_l1clk),
    .io_clk(rvclkhdr_348_io_clk),
    .io_en(rvclkhdr_348_io_en),
    .io_scan_mode(rvclkhdr_348_io_scan_mode)
  );
  rvclkhdr rvclkhdr_349 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_349_io_l1clk),
    .io_clk(rvclkhdr_349_io_clk),
    .io_en(rvclkhdr_349_io_en),
    .io_scan_mode(rvclkhdr_349_io_scan_mode)
  );
  rvclkhdr rvclkhdr_350 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_350_io_l1clk),
    .io_clk(rvclkhdr_350_io_clk),
    .io_en(rvclkhdr_350_io_en),
    .io_scan_mode(rvclkhdr_350_io_scan_mode)
  );
  rvclkhdr rvclkhdr_351 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_351_io_l1clk),
    .io_clk(rvclkhdr_351_io_clk),
    .io_en(rvclkhdr_351_io_en),
    .io_scan_mode(rvclkhdr_351_io_scan_mode)
  );
  rvclkhdr rvclkhdr_352 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_352_io_l1clk),
    .io_clk(rvclkhdr_352_io_clk),
    .io_en(rvclkhdr_352_io_en),
    .io_scan_mode(rvclkhdr_352_io_scan_mode)
  );
  rvclkhdr rvclkhdr_353 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_353_io_l1clk),
    .io_clk(rvclkhdr_353_io_clk),
    .io_en(rvclkhdr_353_io_en),
    .io_scan_mode(rvclkhdr_353_io_scan_mode)
  );
  rvclkhdr rvclkhdr_354 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_354_io_l1clk),
    .io_clk(rvclkhdr_354_io_clk),
    .io_en(rvclkhdr_354_io_en),
    .io_scan_mode(rvclkhdr_354_io_scan_mode)
  );
  rvclkhdr rvclkhdr_355 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_355_io_l1clk),
    .io_clk(rvclkhdr_355_io_clk),
    .io_en(rvclkhdr_355_io_en),
    .io_scan_mode(rvclkhdr_355_io_scan_mode)
  );
  rvclkhdr rvclkhdr_356 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_356_io_l1clk),
    .io_clk(rvclkhdr_356_io_clk),
    .io_en(rvclkhdr_356_io_en),
    .io_scan_mode(rvclkhdr_356_io_scan_mode)
  );
  rvclkhdr rvclkhdr_357 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_357_io_l1clk),
    .io_clk(rvclkhdr_357_io_clk),
    .io_en(rvclkhdr_357_io_en),
    .io_scan_mode(rvclkhdr_357_io_scan_mode)
  );
  rvclkhdr rvclkhdr_358 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_358_io_l1clk),
    .io_clk(rvclkhdr_358_io_clk),
    .io_en(rvclkhdr_358_io_en),
    .io_scan_mode(rvclkhdr_358_io_scan_mode)
  );
  rvclkhdr rvclkhdr_359 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_359_io_l1clk),
    .io_clk(rvclkhdr_359_io_clk),
    .io_en(rvclkhdr_359_io_en),
    .io_scan_mode(rvclkhdr_359_io_scan_mode)
  );
  rvclkhdr rvclkhdr_360 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_360_io_l1clk),
    .io_clk(rvclkhdr_360_io_clk),
    .io_en(rvclkhdr_360_io_en),
    .io_scan_mode(rvclkhdr_360_io_scan_mode)
  );
  rvclkhdr rvclkhdr_361 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_361_io_l1clk),
    .io_clk(rvclkhdr_361_io_clk),
    .io_en(rvclkhdr_361_io_en),
    .io_scan_mode(rvclkhdr_361_io_scan_mode)
  );
  rvclkhdr rvclkhdr_362 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_362_io_l1clk),
    .io_clk(rvclkhdr_362_io_clk),
    .io_en(rvclkhdr_362_io_en),
    .io_scan_mode(rvclkhdr_362_io_scan_mode)
  );
  rvclkhdr rvclkhdr_363 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_363_io_l1clk),
    .io_clk(rvclkhdr_363_io_clk),
    .io_en(rvclkhdr_363_io_en),
    .io_scan_mode(rvclkhdr_363_io_scan_mode)
  );
  rvclkhdr rvclkhdr_364 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_364_io_l1clk),
    .io_clk(rvclkhdr_364_io_clk),
    .io_en(rvclkhdr_364_io_en),
    .io_scan_mode(rvclkhdr_364_io_scan_mode)
  );
  rvclkhdr rvclkhdr_365 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_365_io_l1clk),
    .io_clk(rvclkhdr_365_io_clk),
    .io_en(rvclkhdr_365_io_en),
    .io_scan_mode(rvclkhdr_365_io_scan_mode)
  );
  rvclkhdr rvclkhdr_366 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_366_io_l1clk),
    .io_clk(rvclkhdr_366_io_clk),
    .io_en(rvclkhdr_366_io_en),
    .io_scan_mode(rvclkhdr_366_io_scan_mode)
  );
  rvclkhdr rvclkhdr_367 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_367_io_l1clk),
    .io_clk(rvclkhdr_367_io_clk),
    .io_en(rvclkhdr_367_io_en),
    .io_scan_mode(rvclkhdr_367_io_scan_mode)
  );
  rvclkhdr rvclkhdr_368 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_368_io_l1clk),
    .io_clk(rvclkhdr_368_io_clk),
    .io_en(rvclkhdr_368_io_en),
    .io_scan_mode(rvclkhdr_368_io_scan_mode)
  );
  rvclkhdr rvclkhdr_369 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_369_io_l1clk),
    .io_clk(rvclkhdr_369_io_clk),
    .io_en(rvclkhdr_369_io_en),
    .io_scan_mode(rvclkhdr_369_io_scan_mode)
  );
  rvclkhdr rvclkhdr_370 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_370_io_l1clk),
    .io_clk(rvclkhdr_370_io_clk),
    .io_en(rvclkhdr_370_io_en),
    .io_scan_mode(rvclkhdr_370_io_scan_mode)
  );
  rvclkhdr rvclkhdr_371 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_371_io_l1clk),
    .io_clk(rvclkhdr_371_io_clk),
    .io_en(rvclkhdr_371_io_en),
    .io_scan_mode(rvclkhdr_371_io_scan_mode)
  );
  rvclkhdr rvclkhdr_372 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_372_io_l1clk),
    .io_clk(rvclkhdr_372_io_clk),
    .io_en(rvclkhdr_372_io_en),
    .io_scan_mode(rvclkhdr_372_io_scan_mode)
  );
  rvclkhdr rvclkhdr_373 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_373_io_l1clk),
    .io_clk(rvclkhdr_373_io_clk),
    .io_en(rvclkhdr_373_io_en),
    .io_scan_mode(rvclkhdr_373_io_scan_mode)
  );
  rvclkhdr rvclkhdr_374 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_374_io_l1clk),
    .io_clk(rvclkhdr_374_io_clk),
    .io_en(rvclkhdr_374_io_en),
    .io_scan_mode(rvclkhdr_374_io_scan_mode)
  );
  rvclkhdr rvclkhdr_375 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_375_io_l1clk),
    .io_clk(rvclkhdr_375_io_clk),
    .io_en(rvclkhdr_375_io_en),
    .io_scan_mode(rvclkhdr_375_io_scan_mode)
  );
  rvclkhdr rvclkhdr_376 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_376_io_l1clk),
    .io_clk(rvclkhdr_376_io_clk),
    .io_en(rvclkhdr_376_io_en),
    .io_scan_mode(rvclkhdr_376_io_scan_mode)
  );
  rvclkhdr rvclkhdr_377 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_377_io_l1clk),
    .io_clk(rvclkhdr_377_io_clk),
    .io_en(rvclkhdr_377_io_en),
    .io_scan_mode(rvclkhdr_377_io_scan_mode)
  );
  rvclkhdr rvclkhdr_378 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_378_io_l1clk),
    .io_clk(rvclkhdr_378_io_clk),
    .io_en(rvclkhdr_378_io_en),
    .io_scan_mode(rvclkhdr_378_io_scan_mode)
  );
  rvclkhdr rvclkhdr_379 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_379_io_l1clk),
    .io_clk(rvclkhdr_379_io_clk),
    .io_en(rvclkhdr_379_io_en),
    .io_scan_mode(rvclkhdr_379_io_scan_mode)
  );
  rvclkhdr rvclkhdr_380 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_380_io_l1clk),
    .io_clk(rvclkhdr_380_io_clk),
    .io_en(rvclkhdr_380_io_en),
    .io_scan_mode(rvclkhdr_380_io_scan_mode)
  );
  rvclkhdr rvclkhdr_381 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_381_io_l1clk),
    .io_clk(rvclkhdr_381_io_clk),
    .io_en(rvclkhdr_381_io_en),
    .io_scan_mode(rvclkhdr_381_io_scan_mode)
  );
  rvclkhdr rvclkhdr_382 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_382_io_l1clk),
    .io_clk(rvclkhdr_382_io_clk),
    .io_en(rvclkhdr_382_io_en),
    .io_scan_mode(rvclkhdr_382_io_scan_mode)
  );
  rvclkhdr rvclkhdr_383 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_383_io_l1clk),
    .io_clk(rvclkhdr_383_io_clk),
    .io_en(rvclkhdr_383_io_en),
    .io_scan_mode(rvclkhdr_383_io_scan_mode)
  );
  rvclkhdr rvclkhdr_384 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_384_io_l1clk),
    .io_clk(rvclkhdr_384_io_clk),
    .io_en(rvclkhdr_384_io_en),
    .io_scan_mode(rvclkhdr_384_io_scan_mode)
  );
  rvclkhdr rvclkhdr_385 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_385_io_l1clk),
    .io_clk(rvclkhdr_385_io_clk),
    .io_en(rvclkhdr_385_io_en),
    .io_scan_mode(rvclkhdr_385_io_scan_mode)
  );
  rvclkhdr rvclkhdr_386 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_386_io_l1clk),
    .io_clk(rvclkhdr_386_io_clk),
    .io_en(rvclkhdr_386_io_en),
    .io_scan_mode(rvclkhdr_386_io_scan_mode)
  );
  rvclkhdr rvclkhdr_387 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_387_io_l1clk),
    .io_clk(rvclkhdr_387_io_clk),
    .io_en(rvclkhdr_387_io_en),
    .io_scan_mode(rvclkhdr_387_io_scan_mode)
  );
  rvclkhdr rvclkhdr_388 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_388_io_l1clk),
    .io_clk(rvclkhdr_388_io_clk),
    .io_en(rvclkhdr_388_io_en),
    .io_scan_mode(rvclkhdr_388_io_scan_mode)
  );
  rvclkhdr rvclkhdr_389 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_389_io_l1clk),
    .io_clk(rvclkhdr_389_io_clk),
    .io_en(rvclkhdr_389_io_en),
    .io_scan_mode(rvclkhdr_389_io_scan_mode)
  );
  rvclkhdr rvclkhdr_390 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_390_io_l1clk),
    .io_clk(rvclkhdr_390_io_clk),
    .io_en(rvclkhdr_390_io_en),
    .io_scan_mode(rvclkhdr_390_io_scan_mode)
  );
  rvclkhdr rvclkhdr_391 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_391_io_l1clk),
    .io_clk(rvclkhdr_391_io_clk),
    .io_en(rvclkhdr_391_io_en),
    .io_scan_mode(rvclkhdr_391_io_scan_mode)
  );
  rvclkhdr rvclkhdr_392 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_392_io_l1clk),
    .io_clk(rvclkhdr_392_io_clk),
    .io_en(rvclkhdr_392_io_en),
    .io_scan_mode(rvclkhdr_392_io_scan_mode)
  );
  rvclkhdr rvclkhdr_393 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_393_io_l1clk),
    .io_clk(rvclkhdr_393_io_clk),
    .io_en(rvclkhdr_393_io_en),
    .io_scan_mode(rvclkhdr_393_io_scan_mode)
  );
  rvclkhdr rvclkhdr_394 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_394_io_l1clk),
    .io_clk(rvclkhdr_394_io_clk),
    .io_en(rvclkhdr_394_io_en),
    .io_scan_mode(rvclkhdr_394_io_scan_mode)
  );
  rvclkhdr rvclkhdr_395 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_395_io_l1clk),
    .io_clk(rvclkhdr_395_io_clk),
    .io_en(rvclkhdr_395_io_en),
    .io_scan_mode(rvclkhdr_395_io_scan_mode)
  );
  rvclkhdr rvclkhdr_396 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_396_io_l1clk),
    .io_clk(rvclkhdr_396_io_clk),
    .io_en(rvclkhdr_396_io_en),
    .io_scan_mode(rvclkhdr_396_io_scan_mode)
  );
  rvclkhdr rvclkhdr_397 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_397_io_l1clk),
    .io_clk(rvclkhdr_397_io_clk),
    .io_en(rvclkhdr_397_io_en),
    .io_scan_mode(rvclkhdr_397_io_scan_mode)
  );
  rvclkhdr rvclkhdr_398 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_398_io_l1clk),
    .io_clk(rvclkhdr_398_io_clk),
    .io_en(rvclkhdr_398_io_en),
    .io_scan_mode(rvclkhdr_398_io_scan_mode)
  );
  rvclkhdr rvclkhdr_399 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_399_io_l1clk),
    .io_clk(rvclkhdr_399_io_clk),
    .io_en(rvclkhdr_399_io_en),
    .io_scan_mode(rvclkhdr_399_io_scan_mode)
  );
  rvclkhdr rvclkhdr_400 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_400_io_l1clk),
    .io_clk(rvclkhdr_400_io_clk),
    .io_en(rvclkhdr_400_io_en),
    .io_scan_mode(rvclkhdr_400_io_scan_mode)
  );
  rvclkhdr rvclkhdr_401 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_401_io_l1clk),
    .io_clk(rvclkhdr_401_io_clk),
    .io_en(rvclkhdr_401_io_en),
    .io_scan_mode(rvclkhdr_401_io_scan_mode)
  );
  rvclkhdr rvclkhdr_402 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_402_io_l1clk),
    .io_clk(rvclkhdr_402_io_clk),
    .io_en(rvclkhdr_402_io_en),
    .io_scan_mode(rvclkhdr_402_io_scan_mode)
  );
  rvclkhdr rvclkhdr_403 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_403_io_l1clk),
    .io_clk(rvclkhdr_403_io_clk),
    .io_en(rvclkhdr_403_io_en),
    .io_scan_mode(rvclkhdr_403_io_scan_mode)
  );
  rvclkhdr rvclkhdr_404 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_404_io_l1clk),
    .io_clk(rvclkhdr_404_io_clk),
    .io_en(rvclkhdr_404_io_en),
    .io_scan_mode(rvclkhdr_404_io_scan_mode)
  );
  rvclkhdr rvclkhdr_405 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_405_io_l1clk),
    .io_clk(rvclkhdr_405_io_clk),
    .io_en(rvclkhdr_405_io_en),
    .io_scan_mode(rvclkhdr_405_io_scan_mode)
  );
  rvclkhdr rvclkhdr_406 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_406_io_l1clk),
    .io_clk(rvclkhdr_406_io_clk),
    .io_en(rvclkhdr_406_io_en),
    .io_scan_mode(rvclkhdr_406_io_scan_mode)
  );
  rvclkhdr rvclkhdr_407 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_407_io_l1clk),
    .io_clk(rvclkhdr_407_io_clk),
    .io_en(rvclkhdr_407_io_en),
    .io_scan_mode(rvclkhdr_407_io_scan_mode)
  );
  rvclkhdr rvclkhdr_408 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_408_io_l1clk),
    .io_clk(rvclkhdr_408_io_clk),
    .io_en(rvclkhdr_408_io_en),
    .io_scan_mode(rvclkhdr_408_io_scan_mode)
  );
  rvclkhdr rvclkhdr_409 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_409_io_l1clk),
    .io_clk(rvclkhdr_409_io_clk),
    .io_en(rvclkhdr_409_io_en),
    .io_scan_mode(rvclkhdr_409_io_scan_mode)
  );
  rvclkhdr rvclkhdr_410 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_410_io_l1clk),
    .io_clk(rvclkhdr_410_io_clk),
    .io_en(rvclkhdr_410_io_en),
    .io_scan_mode(rvclkhdr_410_io_scan_mode)
  );
  rvclkhdr rvclkhdr_411 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_411_io_l1clk),
    .io_clk(rvclkhdr_411_io_clk),
    .io_en(rvclkhdr_411_io_en),
    .io_scan_mode(rvclkhdr_411_io_scan_mode)
  );
  rvclkhdr rvclkhdr_412 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_412_io_l1clk),
    .io_clk(rvclkhdr_412_io_clk),
    .io_en(rvclkhdr_412_io_en),
    .io_scan_mode(rvclkhdr_412_io_scan_mode)
  );
  rvclkhdr rvclkhdr_413 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_413_io_l1clk),
    .io_clk(rvclkhdr_413_io_clk),
    .io_en(rvclkhdr_413_io_en),
    .io_scan_mode(rvclkhdr_413_io_scan_mode)
  );
  rvclkhdr rvclkhdr_414 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_414_io_l1clk),
    .io_clk(rvclkhdr_414_io_clk),
    .io_en(rvclkhdr_414_io_en),
    .io_scan_mode(rvclkhdr_414_io_scan_mode)
  );
  rvclkhdr rvclkhdr_415 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_415_io_l1clk),
    .io_clk(rvclkhdr_415_io_clk),
    .io_en(rvclkhdr_415_io_en),
    .io_scan_mode(rvclkhdr_415_io_scan_mode)
  );
  rvclkhdr rvclkhdr_416 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_416_io_l1clk),
    .io_clk(rvclkhdr_416_io_clk),
    .io_en(rvclkhdr_416_io_en),
    .io_scan_mode(rvclkhdr_416_io_scan_mode)
  );
  rvclkhdr rvclkhdr_417 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_417_io_l1clk),
    .io_clk(rvclkhdr_417_io_clk),
    .io_en(rvclkhdr_417_io_en),
    .io_scan_mode(rvclkhdr_417_io_scan_mode)
  );
  rvclkhdr rvclkhdr_418 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_418_io_l1clk),
    .io_clk(rvclkhdr_418_io_clk),
    .io_en(rvclkhdr_418_io_en),
    .io_scan_mode(rvclkhdr_418_io_scan_mode)
  );
  rvclkhdr rvclkhdr_419 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_419_io_l1clk),
    .io_clk(rvclkhdr_419_io_clk),
    .io_en(rvclkhdr_419_io_en),
    .io_scan_mode(rvclkhdr_419_io_scan_mode)
  );
  rvclkhdr rvclkhdr_420 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_420_io_l1clk),
    .io_clk(rvclkhdr_420_io_clk),
    .io_en(rvclkhdr_420_io_en),
    .io_scan_mode(rvclkhdr_420_io_scan_mode)
  );
  rvclkhdr rvclkhdr_421 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_421_io_l1clk),
    .io_clk(rvclkhdr_421_io_clk),
    .io_en(rvclkhdr_421_io_en),
    .io_scan_mode(rvclkhdr_421_io_scan_mode)
  );
  rvclkhdr rvclkhdr_422 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_422_io_l1clk),
    .io_clk(rvclkhdr_422_io_clk),
    .io_en(rvclkhdr_422_io_en),
    .io_scan_mode(rvclkhdr_422_io_scan_mode)
  );
  rvclkhdr rvclkhdr_423 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_423_io_l1clk),
    .io_clk(rvclkhdr_423_io_clk),
    .io_en(rvclkhdr_423_io_en),
    .io_scan_mode(rvclkhdr_423_io_scan_mode)
  );
  rvclkhdr rvclkhdr_424 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_424_io_l1clk),
    .io_clk(rvclkhdr_424_io_clk),
    .io_en(rvclkhdr_424_io_en),
    .io_scan_mode(rvclkhdr_424_io_scan_mode)
  );
  rvclkhdr rvclkhdr_425 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_425_io_l1clk),
    .io_clk(rvclkhdr_425_io_clk),
    .io_en(rvclkhdr_425_io_en),
    .io_scan_mode(rvclkhdr_425_io_scan_mode)
  );
  rvclkhdr rvclkhdr_426 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_426_io_l1clk),
    .io_clk(rvclkhdr_426_io_clk),
    .io_en(rvclkhdr_426_io_en),
    .io_scan_mode(rvclkhdr_426_io_scan_mode)
  );
  rvclkhdr rvclkhdr_427 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_427_io_l1clk),
    .io_clk(rvclkhdr_427_io_clk),
    .io_en(rvclkhdr_427_io_en),
    .io_scan_mode(rvclkhdr_427_io_scan_mode)
  );
  rvclkhdr rvclkhdr_428 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_428_io_l1clk),
    .io_clk(rvclkhdr_428_io_clk),
    .io_en(rvclkhdr_428_io_en),
    .io_scan_mode(rvclkhdr_428_io_scan_mode)
  );
  rvclkhdr rvclkhdr_429 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_429_io_l1clk),
    .io_clk(rvclkhdr_429_io_clk),
    .io_en(rvclkhdr_429_io_en),
    .io_scan_mode(rvclkhdr_429_io_scan_mode)
  );
  rvclkhdr rvclkhdr_430 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_430_io_l1clk),
    .io_clk(rvclkhdr_430_io_clk),
    .io_en(rvclkhdr_430_io_en),
    .io_scan_mode(rvclkhdr_430_io_scan_mode)
  );
  rvclkhdr rvclkhdr_431 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_431_io_l1clk),
    .io_clk(rvclkhdr_431_io_clk),
    .io_en(rvclkhdr_431_io_en),
    .io_scan_mode(rvclkhdr_431_io_scan_mode)
  );
  rvclkhdr rvclkhdr_432 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_432_io_l1clk),
    .io_clk(rvclkhdr_432_io_clk),
    .io_en(rvclkhdr_432_io_en),
    .io_scan_mode(rvclkhdr_432_io_scan_mode)
  );
  rvclkhdr rvclkhdr_433 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_433_io_l1clk),
    .io_clk(rvclkhdr_433_io_clk),
    .io_en(rvclkhdr_433_io_en),
    .io_scan_mode(rvclkhdr_433_io_scan_mode)
  );
  rvclkhdr rvclkhdr_434 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_434_io_l1clk),
    .io_clk(rvclkhdr_434_io_clk),
    .io_en(rvclkhdr_434_io_en),
    .io_scan_mode(rvclkhdr_434_io_scan_mode)
  );
  rvclkhdr rvclkhdr_435 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_435_io_l1clk),
    .io_clk(rvclkhdr_435_io_clk),
    .io_en(rvclkhdr_435_io_en),
    .io_scan_mode(rvclkhdr_435_io_scan_mode)
  );
  rvclkhdr rvclkhdr_436 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_436_io_l1clk),
    .io_clk(rvclkhdr_436_io_clk),
    .io_en(rvclkhdr_436_io_en),
    .io_scan_mode(rvclkhdr_436_io_scan_mode)
  );
  rvclkhdr rvclkhdr_437 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_437_io_l1clk),
    .io_clk(rvclkhdr_437_io_clk),
    .io_en(rvclkhdr_437_io_en),
    .io_scan_mode(rvclkhdr_437_io_scan_mode)
  );
  rvclkhdr rvclkhdr_438 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_438_io_l1clk),
    .io_clk(rvclkhdr_438_io_clk),
    .io_en(rvclkhdr_438_io_en),
    .io_scan_mode(rvclkhdr_438_io_scan_mode)
  );
  rvclkhdr rvclkhdr_439 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_439_io_l1clk),
    .io_clk(rvclkhdr_439_io_clk),
    .io_en(rvclkhdr_439_io_en),
    .io_scan_mode(rvclkhdr_439_io_scan_mode)
  );
  rvclkhdr rvclkhdr_440 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_440_io_l1clk),
    .io_clk(rvclkhdr_440_io_clk),
    .io_en(rvclkhdr_440_io_en),
    .io_scan_mode(rvclkhdr_440_io_scan_mode)
  );
  rvclkhdr rvclkhdr_441 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_441_io_l1clk),
    .io_clk(rvclkhdr_441_io_clk),
    .io_en(rvclkhdr_441_io_en),
    .io_scan_mode(rvclkhdr_441_io_scan_mode)
  );
  rvclkhdr rvclkhdr_442 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_442_io_l1clk),
    .io_clk(rvclkhdr_442_io_clk),
    .io_en(rvclkhdr_442_io_en),
    .io_scan_mode(rvclkhdr_442_io_scan_mode)
  );
  rvclkhdr rvclkhdr_443 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_443_io_l1clk),
    .io_clk(rvclkhdr_443_io_clk),
    .io_en(rvclkhdr_443_io_en),
    .io_scan_mode(rvclkhdr_443_io_scan_mode)
  );
  rvclkhdr rvclkhdr_444 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_444_io_l1clk),
    .io_clk(rvclkhdr_444_io_clk),
    .io_en(rvclkhdr_444_io_en),
    .io_scan_mode(rvclkhdr_444_io_scan_mode)
  );
  rvclkhdr rvclkhdr_445 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_445_io_l1clk),
    .io_clk(rvclkhdr_445_io_clk),
    .io_en(rvclkhdr_445_io_en),
    .io_scan_mode(rvclkhdr_445_io_scan_mode)
  );
  rvclkhdr rvclkhdr_446 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_446_io_l1clk),
    .io_clk(rvclkhdr_446_io_clk),
    .io_en(rvclkhdr_446_io_en),
    .io_scan_mode(rvclkhdr_446_io_scan_mode)
  );
  rvclkhdr rvclkhdr_447 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_447_io_l1clk),
    .io_clk(rvclkhdr_447_io_clk),
    .io_en(rvclkhdr_447_io_en),
    .io_scan_mode(rvclkhdr_447_io_scan_mode)
  );
  rvclkhdr rvclkhdr_448 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_448_io_l1clk),
    .io_clk(rvclkhdr_448_io_clk),
    .io_en(rvclkhdr_448_io_en),
    .io_scan_mode(rvclkhdr_448_io_scan_mode)
  );
  rvclkhdr rvclkhdr_449 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_449_io_l1clk),
    .io_clk(rvclkhdr_449_io_clk),
    .io_en(rvclkhdr_449_io_en),
    .io_scan_mode(rvclkhdr_449_io_scan_mode)
  );
  rvclkhdr rvclkhdr_450 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_450_io_l1clk),
    .io_clk(rvclkhdr_450_io_clk),
    .io_en(rvclkhdr_450_io_en),
    .io_scan_mode(rvclkhdr_450_io_scan_mode)
  );
  rvclkhdr rvclkhdr_451 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_451_io_l1clk),
    .io_clk(rvclkhdr_451_io_clk),
    .io_en(rvclkhdr_451_io_en),
    .io_scan_mode(rvclkhdr_451_io_scan_mode)
  );
  rvclkhdr rvclkhdr_452 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_452_io_l1clk),
    .io_clk(rvclkhdr_452_io_clk),
    .io_en(rvclkhdr_452_io_en),
    .io_scan_mode(rvclkhdr_452_io_scan_mode)
  );
  rvclkhdr rvclkhdr_453 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_453_io_l1clk),
    .io_clk(rvclkhdr_453_io_clk),
    .io_en(rvclkhdr_453_io_en),
    .io_scan_mode(rvclkhdr_453_io_scan_mode)
  );
  rvclkhdr rvclkhdr_454 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_454_io_l1clk),
    .io_clk(rvclkhdr_454_io_clk),
    .io_en(rvclkhdr_454_io_en),
    .io_scan_mode(rvclkhdr_454_io_scan_mode)
  );
  rvclkhdr rvclkhdr_455 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_455_io_l1clk),
    .io_clk(rvclkhdr_455_io_clk),
    .io_en(rvclkhdr_455_io_en),
    .io_scan_mode(rvclkhdr_455_io_scan_mode)
  );
  rvclkhdr rvclkhdr_456 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_456_io_l1clk),
    .io_clk(rvclkhdr_456_io_clk),
    .io_en(rvclkhdr_456_io_en),
    .io_scan_mode(rvclkhdr_456_io_scan_mode)
  );
  rvclkhdr rvclkhdr_457 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_457_io_l1clk),
    .io_clk(rvclkhdr_457_io_clk),
    .io_en(rvclkhdr_457_io_en),
    .io_scan_mode(rvclkhdr_457_io_scan_mode)
  );
  rvclkhdr rvclkhdr_458 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_458_io_l1clk),
    .io_clk(rvclkhdr_458_io_clk),
    .io_en(rvclkhdr_458_io_en),
    .io_scan_mode(rvclkhdr_458_io_scan_mode)
  );
  rvclkhdr rvclkhdr_459 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_459_io_l1clk),
    .io_clk(rvclkhdr_459_io_clk),
    .io_en(rvclkhdr_459_io_en),
    .io_scan_mode(rvclkhdr_459_io_scan_mode)
  );
  rvclkhdr rvclkhdr_460 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_460_io_l1clk),
    .io_clk(rvclkhdr_460_io_clk),
    .io_en(rvclkhdr_460_io_en),
    .io_scan_mode(rvclkhdr_460_io_scan_mode)
  );
  rvclkhdr rvclkhdr_461 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_461_io_l1clk),
    .io_clk(rvclkhdr_461_io_clk),
    .io_en(rvclkhdr_461_io_en),
    .io_scan_mode(rvclkhdr_461_io_scan_mode)
  );
  rvclkhdr rvclkhdr_462 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_462_io_l1clk),
    .io_clk(rvclkhdr_462_io_clk),
    .io_en(rvclkhdr_462_io_en),
    .io_scan_mode(rvclkhdr_462_io_scan_mode)
  );
  rvclkhdr rvclkhdr_463 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_463_io_l1clk),
    .io_clk(rvclkhdr_463_io_clk),
    .io_en(rvclkhdr_463_io_en),
    .io_scan_mode(rvclkhdr_463_io_scan_mode)
  );
  rvclkhdr rvclkhdr_464 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_464_io_l1clk),
    .io_clk(rvclkhdr_464_io_clk),
    .io_en(rvclkhdr_464_io_en),
    .io_scan_mode(rvclkhdr_464_io_scan_mode)
  );
  rvclkhdr rvclkhdr_465 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_465_io_l1clk),
    .io_clk(rvclkhdr_465_io_clk),
    .io_en(rvclkhdr_465_io_en),
    .io_scan_mode(rvclkhdr_465_io_scan_mode)
  );
  rvclkhdr rvclkhdr_466 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_466_io_l1clk),
    .io_clk(rvclkhdr_466_io_clk),
    .io_en(rvclkhdr_466_io_en),
    .io_scan_mode(rvclkhdr_466_io_scan_mode)
  );
  rvclkhdr rvclkhdr_467 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_467_io_l1clk),
    .io_clk(rvclkhdr_467_io_clk),
    .io_en(rvclkhdr_467_io_en),
    .io_scan_mode(rvclkhdr_467_io_scan_mode)
  );
  rvclkhdr rvclkhdr_468 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_468_io_l1clk),
    .io_clk(rvclkhdr_468_io_clk),
    .io_en(rvclkhdr_468_io_en),
    .io_scan_mode(rvclkhdr_468_io_scan_mode)
  );
  rvclkhdr rvclkhdr_469 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_469_io_l1clk),
    .io_clk(rvclkhdr_469_io_clk),
    .io_en(rvclkhdr_469_io_en),
    .io_scan_mode(rvclkhdr_469_io_scan_mode)
  );
  rvclkhdr rvclkhdr_470 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_470_io_l1clk),
    .io_clk(rvclkhdr_470_io_clk),
    .io_en(rvclkhdr_470_io_en),
    .io_scan_mode(rvclkhdr_470_io_scan_mode)
  );
  rvclkhdr rvclkhdr_471 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_471_io_l1clk),
    .io_clk(rvclkhdr_471_io_clk),
    .io_en(rvclkhdr_471_io_en),
    .io_scan_mode(rvclkhdr_471_io_scan_mode)
  );
  rvclkhdr rvclkhdr_472 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_472_io_l1clk),
    .io_clk(rvclkhdr_472_io_clk),
    .io_en(rvclkhdr_472_io_en),
    .io_scan_mode(rvclkhdr_472_io_scan_mode)
  );
  rvclkhdr rvclkhdr_473 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_473_io_l1clk),
    .io_clk(rvclkhdr_473_io_clk),
    .io_en(rvclkhdr_473_io_en),
    .io_scan_mode(rvclkhdr_473_io_scan_mode)
  );
  rvclkhdr rvclkhdr_474 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_474_io_l1clk),
    .io_clk(rvclkhdr_474_io_clk),
    .io_en(rvclkhdr_474_io_en),
    .io_scan_mode(rvclkhdr_474_io_scan_mode)
  );
  rvclkhdr rvclkhdr_475 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_475_io_l1clk),
    .io_clk(rvclkhdr_475_io_clk),
    .io_en(rvclkhdr_475_io_en),
    .io_scan_mode(rvclkhdr_475_io_scan_mode)
  );
  rvclkhdr rvclkhdr_476 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_476_io_l1clk),
    .io_clk(rvclkhdr_476_io_clk),
    .io_en(rvclkhdr_476_io_en),
    .io_scan_mode(rvclkhdr_476_io_scan_mode)
  );
  rvclkhdr rvclkhdr_477 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_477_io_l1clk),
    .io_clk(rvclkhdr_477_io_clk),
    .io_en(rvclkhdr_477_io_en),
    .io_scan_mode(rvclkhdr_477_io_scan_mode)
  );
  rvclkhdr rvclkhdr_478 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_478_io_l1clk),
    .io_clk(rvclkhdr_478_io_clk),
    .io_en(rvclkhdr_478_io_en),
    .io_scan_mode(rvclkhdr_478_io_scan_mode)
  );
  rvclkhdr rvclkhdr_479 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_479_io_l1clk),
    .io_clk(rvclkhdr_479_io_clk),
    .io_en(rvclkhdr_479_io_en),
    .io_scan_mode(rvclkhdr_479_io_scan_mode)
  );
  rvclkhdr rvclkhdr_480 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_480_io_l1clk),
    .io_clk(rvclkhdr_480_io_clk),
    .io_en(rvclkhdr_480_io_en),
    .io_scan_mode(rvclkhdr_480_io_scan_mode)
  );
  rvclkhdr rvclkhdr_481 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_481_io_l1clk),
    .io_clk(rvclkhdr_481_io_clk),
    .io_en(rvclkhdr_481_io_en),
    .io_scan_mode(rvclkhdr_481_io_scan_mode)
  );
  rvclkhdr rvclkhdr_482 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_482_io_l1clk),
    .io_clk(rvclkhdr_482_io_clk),
    .io_en(rvclkhdr_482_io_en),
    .io_scan_mode(rvclkhdr_482_io_scan_mode)
  );
  rvclkhdr rvclkhdr_483 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_483_io_l1clk),
    .io_clk(rvclkhdr_483_io_clk),
    .io_en(rvclkhdr_483_io_en),
    .io_scan_mode(rvclkhdr_483_io_scan_mode)
  );
  rvclkhdr rvclkhdr_484 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_484_io_l1clk),
    .io_clk(rvclkhdr_484_io_clk),
    .io_en(rvclkhdr_484_io_en),
    .io_scan_mode(rvclkhdr_484_io_scan_mode)
  );
  rvclkhdr rvclkhdr_485 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_485_io_l1clk),
    .io_clk(rvclkhdr_485_io_clk),
    .io_en(rvclkhdr_485_io_en),
    .io_scan_mode(rvclkhdr_485_io_scan_mode)
  );
  rvclkhdr rvclkhdr_486 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_486_io_l1clk),
    .io_clk(rvclkhdr_486_io_clk),
    .io_en(rvclkhdr_486_io_en),
    .io_scan_mode(rvclkhdr_486_io_scan_mode)
  );
  rvclkhdr rvclkhdr_487 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_487_io_l1clk),
    .io_clk(rvclkhdr_487_io_clk),
    .io_en(rvclkhdr_487_io_en),
    .io_scan_mode(rvclkhdr_487_io_scan_mode)
  );
  rvclkhdr rvclkhdr_488 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_488_io_l1clk),
    .io_clk(rvclkhdr_488_io_clk),
    .io_en(rvclkhdr_488_io_en),
    .io_scan_mode(rvclkhdr_488_io_scan_mode)
  );
  rvclkhdr rvclkhdr_489 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_489_io_l1clk),
    .io_clk(rvclkhdr_489_io_clk),
    .io_en(rvclkhdr_489_io_en),
    .io_scan_mode(rvclkhdr_489_io_scan_mode)
  );
  rvclkhdr rvclkhdr_490 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_490_io_l1clk),
    .io_clk(rvclkhdr_490_io_clk),
    .io_en(rvclkhdr_490_io_en),
    .io_scan_mode(rvclkhdr_490_io_scan_mode)
  );
  rvclkhdr rvclkhdr_491 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_491_io_l1clk),
    .io_clk(rvclkhdr_491_io_clk),
    .io_en(rvclkhdr_491_io_en),
    .io_scan_mode(rvclkhdr_491_io_scan_mode)
  );
  rvclkhdr rvclkhdr_492 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_492_io_l1clk),
    .io_clk(rvclkhdr_492_io_clk),
    .io_en(rvclkhdr_492_io_en),
    .io_scan_mode(rvclkhdr_492_io_scan_mode)
  );
  rvclkhdr rvclkhdr_493 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_493_io_l1clk),
    .io_clk(rvclkhdr_493_io_clk),
    .io_en(rvclkhdr_493_io_en),
    .io_scan_mode(rvclkhdr_493_io_scan_mode)
  );
  rvclkhdr rvclkhdr_494 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_494_io_l1clk),
    .io_clk(rvclkhdr_494_io_clk),
    .io_en(rvclkhdr_494_io_en),
    .io_scan_mode(rvclkhdr_494_io_scan_mode)
  );
  rvclkhdr rvclkhdr_495 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_495_io_l1clk),
    .io_clk(rvclkhdr_495_io_clk),
    .io_en(rvclkhdr_495_io_en),
    .io_scan_mode(rvclkhdr_495_io_scan_mode)
  );
  rvclkhdr rvclkhdr_496 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_496_io_l1clk),
    .io_clk(rvclkhdr_496_io_clk),
    .io_en(rvclkhdr_496_io_en),
    .io_scan_mode(rvclkhdr_496_io_scan_mode)
  );
  rvclkhdr rvclkhdr_497 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_497_io_l1clk),
    .io_clk(rvclkhdr_497_io_clk),
    .io_en(rvclkhdr_497_io_en),
    .io_scan_mode(rvclkhdr_497_io_scan_mode)
  );
  rvclkhdr rvclkhdr_498 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_498_io_l1clk),
    .io_clk(rvclkhdr_498_io_clk),
    .io_en(rvclkhdr_498_io_en),
    .io_scan_mode(rvclkhdr_498_io_scan_mode)
  );
  rvclkhdr rvclkhdr_499 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_499_io_l1clk),
    .io_clk(rvclkhdr_499_io_clk),
    .io_en(rvclkhdr_499_io_en),
    .io_scan_mode(rvclkhdr_499_io_scan_mode)
  );
  rvclkhdr rvclkhdr_500 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_500_io_l1clk),
    .io_clk(rvclkhdr_500_io_clk),
    .io_en(rvclkhdr_500_io_en),
    .io_scan_mode(rvclkhdr_500_io_scan_mode)
  );
  rvclkhdr rvclkhdr_501 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_501_io_l1clk),
    .io_clk(rvclkhdr_501_io_clk),
    .io_en(rvclkhdr_501_io_en),
    .io_scan_mode(rvclkhdr_501_io_scan_mode)
  );
  rvclkhdr rvclkhdr_502 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_502_io_l1clk),
    .io_clk(rvclkhdr_502_io_clk),
    .io_en(rvclkhdr_502_io_en),
    .io_scan_mode(rvclkhdr_502_io_scan_mode)
  );
  rvclkhdr rvclkhdr_503 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_503_io_l1clk),
    .io_clk(rvclkhdr_503_io_clk),
    .io_en(rvclkhdr_503_io_en),
    .io_scan_mode(rvclkhdr_503_io_scan_mode)
  );
  rvclkhdr rvclkhdr_504 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_504_io_l1clk),
    .io_clk(rvclkhdr_504_io_clk),
    .io_en(rvclkhdr_504_io_en),
    .io_scan_mode(rvclkhdr_504_io_scan_mode)
  );
  rvclkhdr rvclkhdr_505 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_505_io_l1clk),
    .io_clk(rvclkhdr_505_io_clk),
    .io_en(rvclkhdr_505_io_en),
    .io_scan_mode(rvclkhdr_505_io_scan_mode)
  );
  rvclkhdr rvclkhdr_506 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_506_io_l1clk),
    .io_clk(rvclkhdr_506_io_clk),
    .io_en(rvclkhdr_506_io_en),
    .io_scan_mode(rvclkhdr_506_io_scan_mode)
  );
  rvclkhdr rvclkhdr_507 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_507_io_l1clk),
    .io_clk(rvclkhdr_507_io_clk),
    .io_en(rvclkhdr_507_io_en),
    .io_scan_mode(rvclkhdr_507_io_scan_mode)
  );
  rvclkhdr rvclkhdr_508 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_508_io_l1clk),
    .io_clk(rvclkhdr_508_io_clk),
    .io_en(rvclkhdr_508_io_en),
    .io_scan_mode(rvclkhdr_508_io_scan_mode)
  );
  rvclkhdr rvclkhdr_509 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_509_io_l1clk),
    .io_clk(rvclkhdr_509_io_clk),
    .io_en(rvclkhdr_509_io_en),
    .io_scan_mode(rvclkhdr_509_io_scan_mode)
  );
  rvclkhdr rvclkhdr_510 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_510_io_l1clk),
    .io_clk(rvclkhdr_510_io_clk),
    .io_en(rvclkhdr_510_io_en),
    .io_scan_mode(rvclkhdr_510_io_scan_mode)
  );
  rvclkhdr rvclkhdr_511 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_511_io_l1clk),
    .io_clk(rvclkhdr_511_io_clk),
    .io_en(rvclkhdr_511_io_en),
    .io_scan_mode(rvclkhdr_511_io_scan_mode)
  );
  rvclkhdr rvclkhdr_512 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_512_io_l1clk),
    .io_clk(rvclkhdr_512_io_clk),
    .io_en(rvclkhdr_512_io_en),
    .io_scan_mode(rvclkhdr_512_io_scan_mode)
  );
  rvclkhdr rvclkhdr_513 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_513_io_l1clk),
    .io_clk(rvclkhdr_513_io_clk),
    .io_en(rvclkhdr_513_io_en),
    .io_scan_mode(rvclkhdr_513_io_scan_mode)
  );
  rvclkhdr rvclkhdr_514 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_514_io_l1clk),
    .io_clk(rvclkhdr_514_io_clk),
    .io_en(rvclkhdr_514_io_en),
    .io_scan_mode(rvclkhdr_514_io_scan_mode)
  );
  rvclkhdr rvclkhdr_515 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_515_io_l1clk),
    .io_clk(rvclkhdr_515_io_clk),
    .io_en(rvclkhdr_515_io_en),
    .io_scan_mode(rvclkhdr_515_io_scan_mode)
  );
  rvclkhdr rvclkhdr_516 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_516_io_l1clk),
    .io_clk(rvclkhdr_516_io_clk),
    .io_en(rvclkhdr_516_io_en),
    .io_scan_mode(rvclkhdr_516_io_scan_mode)
  );
  rvclkhdr rvclkhdr_517 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_517_io_l1clk),
    .io_clk(rvclkhdr_517_io_clk),
    .io_en(rvclkhdr_517_io_en),
    .io_scan_mode(rvclkhdr_517_io_scan_mode)
  );
  rvclkhdr rvclkhdr_518 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_518_io_l1clk),
    .io_clk(rvclkhdr_518_io_clk),
    .io_en(rvclkhdr_518_io_en),
    .io_scan_mode(rvclkhdr_518_io_scan_mode)
  );
  rvclkhdr rvclkhdr_519 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_519_io_l1clk),
    .io_clk(rvclkhdr_519_io_clk),
    .io_en(rvclkhdr_519_io_en),
    .io_scan_mode(rvclkhdr_519_io_scan_mode)
  );
  rvclkhdr rvclkhdr_520 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_520_io_l1clk),
    .io_clk(rvclkhdr_520_io_clk),
    .io_en(rvclkhdr_520_io_en),
    .io_scan_mode(rvclkhdr_520_io_scan_mode)
  );
  rvclkhdr rvclkhdr_521 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_521_io_l1clk),
    .io_clk(rvclkhdr_521_io_clk),
    .io_en(rvclkhdr_521_io_en),
    .io_scan_mode(rvclkhdr_521_io_scan_mode)
  );
  rvclkhdr rvclkhdr_522 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_522_io_l1clk),
    .io_clk(rvclkhdr_522_io_clk),
    .io_en(rvclkhdr_522_io_en),
    .io_scan_mode(rvclkhdr_522_io_scan_mode)
  );
  rvclkhdr rvclkhdr_523 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_523_io_l1clk),
    .io_clk(rvclkhdr_523_io_clk),
    .io_en(rvclkhdr_523_io_en),
    .io_scan_mode(rvclkhdr_523_io_scan_mode)
  );
  rvclkhdr rvclkhdr_524 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_524_io_l1clk),
    .io_clk(rvclkhdr_524_io_clk),
    .io_en(rvclkhdr_524_io_en),
    .io_scan_mode(rvclkhdr_524_io_scan_mode)
  );
  rvclkhdr rvclkhdr_525 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_525_io_l1clk),
    .io_clk(rvclkhdr_525_io_clk),
    .io_en(rvclkhdr_525_io_en),
    .io_scan_mode(rvclkhdr_525_io_scan_mode)
  );
  rvclkhdr rvclkhdr_526 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_526_io_l1clk),
    .io_clk(rvclkhdr_526_io_clk),
    .io_en(rvclkhdr_526_io_en),
    .io_scan_mode(rvclkhdr_526_io_scan_mode)
  );
  rvclkhdr rvclkhdr_527 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_527_io_l1clk),
    .io_clk(rvclkhdr_527_io_clk),
    .io_en(rvclkhdr_527_io_en),
    .io_scan_mode(rvclkhdr_527_io_scan_mode)
  );
  rvclkhdr rvclkhdr_528 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_528_io_l1clk),
    .io_clk(rvclkhdr_528_io_clk),
    .io_en(rvclkhdr_528_io_en),
    .io_scan_mode(rvclkhdr_528_io_scan_mode)
  );
  rvclkhdr rvclkhdr_529 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_529_io_l1clk),
    .io_clk(rvclkhdr_529_io_clk),
    .io_en(rvclkhdr_529_io_en),
    .io_scan_mode(rvclkhdr_529_io_scan_mode)
  );
  rvclkhdr rvclkhdr_530 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_530_io_l1clk),
    .io_clk(rvclkhdr_530_io_clk),
    .io_en(rvclkhdr_530_io_en),
    .io_scan_mode(rvclkhdr_530_io_scan_mode)
  );
  rvclkhdr rvclkhdr_531 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_531_io_l1clk),
    .io_clk(rvclkhdr_531_io_clk),
    .io_en(rvclkhdr_531_io_en),
    .io_scan_mode(rvclkhdr_531_io_scan_mode)
  );
  rvclkhdr rvclkhdr_532 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_532_io_l1clk),
    .io_clk(rvclkhdr_532_io_clk),
    .io_en(rvclkhdr_532_io_en),
    .io_scan_mode(rvclkhdr_532_io_scan_mode)
  );
  rvclkhdr rvclkhdr_533 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_533_io_l1clk),
    .io_clk(rvclkhdr_533_io_clk),
    .io_en(rvclkhdr_533_io_en),
    .io_scan_mode(rvclkhdr_533_io_scan_mode)
  );
  rvclkhdr rvclkhdr_534 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_534_io_l1clk),
    .io_clk(rvclkhdr_534_io_clk),
    .io_en(rvclkhdr_534_io_en),
    .io_scan_mode(rvclkhdr_534_io_scan_mode)
  );
  rvclkhdr rvclkhdr_535 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_535_io_l1clk),
    .io_clk(rvclkhdr_535_io_clk),
    .io_en(rvclkhdr_535_io_en),
    .io_scan_mode(rvclkhdr_535_io_scan_mode)
  );
  rvclkhdr rvclkhdr_536 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_536_io_l1clk),
    .io_clk(rvclkhdr_536_io_clk),
    .io_en(rvclkhdr_536_io_en),
    .io_scan_mode(rvclkhdr_536_io_scan_mode)
  );
  rvclkhdr rvclkhdr_537 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_537_io_l1clk),
    .io_clk(rvclkhdr_537_io_clk),
    .io_en(rvclkhdr_537_io_en),
    .io_scan_mode(rvclkhdr_537_io_scan_mode)
  );
  rvclkhdr rvclkhdr_538 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_538_io_l1clk),
    .io_clk(rvclkhdr_538_io_clk),
    .io_en(rvclkhdr_538_io_en),
    .io_scan_mode(rvclkhdr_538_io_scan_mode)
  );
  rvclkhdr rvclkhdr_539 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_539_io_l1clk),
    .io_clk(rvclkhdr_539_io_clk),
    .io_en(rvclkhdr_539_io_en),
    .io_scan_mode(rvclkhdr_539_io_scan_mode)
  );
  rvclkhdr rvclkhdr_540 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_540_io_l1clk),
    .io_clk(rvclkhdr_540_io_clk),
    .io_en(rvclkhdr_540_io_en),
    .io_scan_mode(rvclkhdr_540_io_scan_mode)
  );
  rvclkhdr rvclkhdr_541 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_541_io_l1clk),
    .io_clk(rvclkhdr_541_io_clk),
    .io_en(rvclkhdr_541_io_en),
    .io_scan_mode(rvclkhdr_541_io_scan_mode)
  );
  rvclkhdr rvclkhdr_542 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_542_io_l1clk),
    .io_clk(rvclkhdr_542_io_clk),
    .io_en(rvclkhdr_542_io_en),
    .io_scan_mode(rvclkhdr_542_io_scan_mode)
  );
  rvclkhdr rvclkhdr_543 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_543_io_l1clk),
    .io_clk(rvclkhdr_543_io_clk),
    .io_en(rvclkhdr_543_io_en),
    .io_scan_mode(rvclkhdr_543_io_scan_mode)
  );
  rvclkhdr rvclkhdr_544 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_544_io_l1clk),
    .io_clk(rvclkhdr_544_io_clk),
    .io_en(rvclkhdr_544_io_en),
    .io_scan_mode(rvclkhdr_544_io_scan_mode)
  );
  rvclkhdr rvclkhdr_545 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_545_io_l1clk),
    .io_clk(rvclkhdr_545_io_clk),
    .io_en(rvclkhdr_545_io_en),
    .io_scan_mode(rvclkhdr_545_io_scan_mode)
  );
  rvclkhdr rvclkhdr_546 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_546_io_l1clk),
    .io_clk(rvclkhdr_546_io_clk),
    .io_en(rvclkhdr_546_io_en),
    .io_scan_mode(rvclkhdr_546_io_scan_mode)
  );
  rvclkhdr rvclkhdr_547 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_547_io_l1clk),
    .io_clk(rvclkhdr_547_io_clk),
    .io_en(rvclkhdr_547_io_en),
    .io_scan_mode(rvclkhdr_547_io_scan_mode)
  );
  rvclkhdr rvclkhdr_548 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_548_io_l1clk),
    .io_clk(rvclkhdr_548_io_clk),
    .io_en(rvclkhdr_548_io_en),
    .io_scan_mode(rvclkhdr_548_io_scan_mode)
  );
  rvclkhdr rvclkhdr_549 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_549_io_l1clk),
    .io_clk(rvclkhdr_549_io_clk),
    .io_en(rvclkhdr_549_io_en),
    .io_scan_mode(rvclkhdr_549_io_scan_mode)
  );
  rvclkhdr rvclkhdr_550 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_550_io_l1clk),
    .io_clk(rvclkhdr_550_io_clk),
    .io_en(rvclkhdr_550_io_en),
    .io_scan_mode(rvclkhdr_550_io_scan_mode)
  );
  rvclkhdr rvclkhdr_551 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_551_io_l1clk),
    .io_clk(rvclkhdr_551_io_clk),
    .io_en(rvclkhdr_551_io_en),
    .io_scan_mode(rvclkhdr_551_io_scan_mode)
  );
  rvclkhdr rvclkhdr_552 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_552_io_l1clk),
    .io_clk(rvclkhdr_552_io_clk),
    .io_en(rvclkhdr_552_io_en),
    .io_scan_mode(rvclkhdr_552_io_scan_mode)
  );
  rvclkhdr rvclkhdr_553 ( // @[lib.scala 343:22]
    .io_l1clk(rvclkhdr_553_io_l1clk),
    .io_clk(rvclkhdr_553_io_clk),
    .io_en(rvclkhdr_553_io_en),
    .io_scan_mode(rvclkhdr_553_io_scan_mode)
  );
  assign io_ifu_bp_hit_taken_f = _T_238 & _T_239; // @[ifu_bp_ctl.scala 261:25]
  assign io_ifu_bp_btb_target_f = _T_429 ? rets_out_0[31:1] : bp_btb_target_adder_f[31:1]; // @[ifu_bp_ctl.scala 357:26]
  assign io_ifu_bp_inst_mask_f = _T_275 | _T_276; // @[ifu_bp_ctl.scala 285:25]
  assign io_ifu_bp_fghr_f = fghr; // @[ifu_bp_ctl.scala 325:20]
  assign io_ifu_bp_way_f = tag_match_vway1_expanded_f | _T_213; // @[ifu_bp_ctl.scala 235:19]
  assign io_ifu_bp_ret_f = {_T_295,_T_301}; // @[ifu_bp_ctl.scala 331:19]
  assign io_ifu_bp_hist1_f = bht_force_taken_f | _T_280; // @[ifu_bp_ctl.scala 326:21]
  assign io_ifu_bp_hist0_f = {bht_vbank1_rd_data_f[0],bht_vbank0_rd_data_f[0]}; // @[ifu_bp_ctl.scala 327:21]
  assign io_ifu_bp_pc4_f = {_T_286,_T_289}; // @[ifu_bp_ctl.scala 328:19]
  assign io_ifu_bp_valid_f = bht_valid_f & _T_345; // @[ifu_bp_ctl.scala 330:21]
  assign io_ifu_bp_poffset_f = btb_sel_data_f[15:4]; // @[ifu_bp_ctl.scala 344:23]
  assign rvclkhdr_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_io_en = io_ifc_fetch_req_f | exu_mp_valid; // @[lib.scala 371:17]
  assign rvclkhdr_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_1_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_1_io_en = _T_376 & io_ic_hit_f; // @[lib.scala 371:17]
  assign rvclkhdr_1_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_2_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_2_io_en = ~rs_hold; // @[lib.scala 371:17]
  assign rvclkhdr_2_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_3_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_3_io_en = rs_push | rs_pop; // @[lib.scala 371:17]
  assign rvclkhdr_3_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_4_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_4_io_en = rs_push | rs_pop; // @[lib.scala 371:17]
  assign rvclkhdr_4_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_5_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_5_io_en = rs_push | rs_pop; // @[lib.scala 371:17]
  assign rvclkhdr_5_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_6_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_6_io_en = rs_push | rs_pop; // @[lib.scala 371:17]
  assign rvclkhdr_6_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_7_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_7_io_en = rs_push | rs_pop; // @[lib.scala 371:17]
  assign rvclkhdr_7_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_8_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_8_io_en = rs_push | rs_pop; // @[lib.scala 371:17]
  assign rvclkhdr_8_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_9_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_9_io_en = _T_473 & io_ifu_bp_hit_taken_f; // @[lib.scala 371:17]
  assign rvclkhdr_9_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_10_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_10_io_en = _T_576 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_10_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_11_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_11_io_en = _T_579 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_11_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_12_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_12_io_en = _T_582 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_12_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_13_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_13_io_en = _T_585 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_13_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_14_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_14_io_en = _T_588 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_14_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_15_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_15_io_en = _T_591 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_15_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_16_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_16_io_en = _T_594 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_16_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_17_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_17_io_en = _T_597 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_17_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_18_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_18_io_en = _T_600 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_18_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_19_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_19_io_en = _T_603 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_19_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_20_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_20_io_en = _T_606 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_20_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_21_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_21_io_en = _T_609 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_21_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_22_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_22_io_en = _T_612 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_22_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_23_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_23_io_en = _T_615 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_23_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_24_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_24_io_en = _T_618 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_24_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_25_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_25_io_en = _T_621 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_25_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_26_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_26_io_en = _T_624 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_26_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_27_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_27_io_en = _T_627 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_27_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_28_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_28_io_en = _T_630 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_28_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_29_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_29_io_en = _T_633 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_29_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_30_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_30_io_en = _T_636 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_30_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_31_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_31_io_en = _T_639 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_31_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_32_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_32_io_en = _T_642 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_32_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_33_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_33_io_en = _T_645 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_33_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_34_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_34_io_en = _T_648 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_34_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_35_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_35_io_en = _T_651 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_35_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_36_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_36_io_en = _T_654 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_36_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_37_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_37_io_en = _T_657 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_37_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_38_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_38_io_en = _T_660 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_38_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_39_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_39_io_en = _T_663 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_39_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_40_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_40_io_en = _T_666 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_40_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_41_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_41_io_en = _T_669 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_41_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_42_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_42_io_en = _T_672 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_42_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_43_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_43_io_en = _T_675 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_43_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_44_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_44_io_en = _T_678 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_44_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_45_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_45_io_en = _T_681 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_45_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_46_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_46_io_en = _T_684 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_46_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_47_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_47_io_en = _T_687 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_47_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_48_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_48_io_en = _T_690 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_48_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_49_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_49_io_en = _T_693 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_49_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_50_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_50_io_en = _T_696 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_50_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_51_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_51_io_en = _T_699 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_51_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_52_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_52_io_en = _T_702 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_52_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_53_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_53_io_en = _T_705 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_53_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_54_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_54_io_en = _T_708 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_54_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_55_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_55_io_en = _T_711 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_55_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_56_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_56_io_en = _T_714 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_56_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_57_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_57_io_en = _T_717 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_57_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_58_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_58_io_en = _T_720 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_58_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_59_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_59_io_en = _T_723 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_59_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_60_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_60_io_en = _T_726 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_60_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_61_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_61_io_en = _T_729 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_61_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_62_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_62_io_en = _T_732 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_62_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_63_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_63_io_en = _T_735 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_63_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_64_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_64_io_en = _T_738 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_64_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_65_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_65_io_en = _T_741 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_65_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_66_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_66_io_en = _T_744 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_66_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_67_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_67_io_en = _T_747 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_67_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_68_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_68_io_en = _T_750 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_68_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_69_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_69_io_en = _T_753 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_69_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_70_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_70_io_en = _T_756 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_70_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_71_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_71_io_en = _T_759 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_71_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_72_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_72_io_en = _T_762 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_72_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_73_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_73_io_en = _T_765 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_73_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_74_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_74_io_en = _T_768 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_74_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_75_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_75_io_en = _T_771 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_75_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_76_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_76_io_en = _T_774 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_76_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_77_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_77_io_en = _T_777 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_77_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_78_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_78_io_en = _T_780 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_78_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_79_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_79_io_en = _T_783 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_79_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_80_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_80_io_en = _T_786 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_80_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_81_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_81_io_en = _T_789 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_81_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_82_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_82_io_en = _T_792 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_82_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_83_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_83_io_en = _T_795 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_83_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_84_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_84_io_en = _T_798 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_84_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_85_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_85_io_en = _T_801 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_85_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_86_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_86_io_en = _T_804 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_86_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_87_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_87_io_en = _T_807 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_87_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_88_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_88_io_en = _T_810 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_88_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_89_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_89_io_en = _T_813 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_89_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_90_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_90_io_en = _T_816 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_90_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_91_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_91_io_en = _T_819 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_91_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_92_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_92_io_en = _T_822 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_92_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_93_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_93_io_en = _T_825 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_93_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_94_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_94_io_en = _T_828 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_94_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_95_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_95_io_en = _T_831 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_95_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_96_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_96_io_en = _T_834 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_96_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_97_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_97_io_en = _T_837 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_97_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_98_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_98_io_en = _T_840 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_98_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_99_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_99_io_en = _T_843 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_99_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_100_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_100_io_en = _T_846 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_100_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_101_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_101_io_en = _T_849 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_101_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_102_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_102_io_en = _T_852 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_102_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_103_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_103_io_en = _T_855 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_103_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_104_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_104_io_en = _T_858 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_104_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_105_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_105_io_en = _T_861 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_105_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_106_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_106_io_en = _T_864 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_106_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_107_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_107_io_en = _T_867 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_107_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_108_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_108_io_en = _T_870 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_108_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_109_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_109_io_en = _T_873 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_109_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_110_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_110_io_en = _T_876 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_110_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_111_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_111_io_en = _T_879 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_111_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_112_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_112_io_en = _T_882 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_112_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_113_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_113_io_en = _T_885 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_113_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_114_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_114_io_en = _T_888 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_114_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_115_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_115_io_en = _T_891 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_115_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_116_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_116_io_en = _T_894 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_116_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_117_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_117_io_en = _T_897 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_117_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_118_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_118_io_en = _T_900 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_118_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_119_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_119_io_en = _T_903 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_119_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_120_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_120_io_en = _T_906 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_120_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_121_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_121_io_en = _T_909 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_121_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_122_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_122_io_en = _T_912 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_122_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_123_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_123_io_en = _T_915 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_123_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_124_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_124_io_en = _T_918 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_124_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_125_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_125_io_en = _T_921 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_125_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_126_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_126_io_en = _T_924 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_126_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_127_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_127_io_en = _T_927 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_127_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_128_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_128_io_en = _T_930 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_128_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_129_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_129_io_en = _T_933 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_129_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_130_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_130_io_en = _T_936 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_130_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_131_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_131_io_en = _T_939 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_131_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_132_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_132_io_en = _T_942 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_132_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_133_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_133_io_en = _T_945 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_133_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_134_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_134_io_en = _T_948 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_134_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_135_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_135_io_en = _T_951 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_135_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_136_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_136_io_en = _T_954 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_136_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_137_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_137_io_en = _T_957 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_137_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_138_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_138_io_en = _T_960 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_138_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_139_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_139_io_en = _T_963 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_139_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_140_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_140_io_en = _T_966 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_140_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_141_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_141_io_en = _T_969 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_141_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_142_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_142_io_en = _T_972 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_142_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_143_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_143_io_en = _T_975 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_143_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_144_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_144_io_en = _T_978 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_144_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_145_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_145_io_en = _T_981 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_145_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_146_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_146_io_en = _T_984 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_146_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_147_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_147_io_en = _T_987 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_147_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_148_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_148_io_en = _T_990 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_148_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_149_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_149_io_en = _T_993 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_149_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_150_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_150_io_en = _T_996 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_150_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_151_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_151_io_en = _T_999 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_151_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_152_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_152_io_en = _T_1002 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_152_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_153_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_153_io_en = _T_1005 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_153_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_154_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_154_io_en = _T_1008 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_154_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_155_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_155_io_en = _T_1011 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_155_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_156_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_156_io_en = _T_1014 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_156_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_157_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_157_io_en = _T_1017 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_157_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_158_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_158_io_en = _T_1020 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_158_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_159_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_159_io_en = _T_1023 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_159_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_160_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_160_io_en = _T_1026 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_160_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_161_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_161_io_en = _T_1029 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_161_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_162_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_162_io_en = _T_1032 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_162_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_163_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_163_io_en = _T_1035 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_163_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_164_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_164_io_en = _T_1038 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_164_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_165_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_165_io_en = _T_1041 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_165_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_166_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_166_io_en = _T_1044 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_166_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_167_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_167_io_en = _T_1047 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_167_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_168_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_168_io_en = _T_1050 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_168_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_169_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_169_io_en = _T_1053 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_169_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_170_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_170_io_en = _T_1056 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_170_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_171_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_171_io_en = _T_1059 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_171_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_172_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_172_io_en = _T_1062 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_172_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_173_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_173_io_en = _T_1065 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_173_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_174_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_174_io_en = _T_1068 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_174_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_175_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_175_io_en = _T_1071 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_175_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_176_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_176_io_en = _T_1074 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_176_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_177_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_177_io_en = _T_1077 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_177_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_178_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_178_io_en = _T_1080 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_178_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_179_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_179_io_en = _T_1083 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_179_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_180_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_180_io_en = _T_1086 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_180_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_181_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_181_io_en = _T_1089 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_181_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_182_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_182_io_en = _T_1092 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_182_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_183_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_183_io_en = _T_1095 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_183_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_184_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_184_io_en = _T_1098 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_184_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_185_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_185_io_en = _T_1101 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_185_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_186_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_186_io_en = _T_1104 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_186_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_187_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_187_io_en = _T_1107 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_187_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_188_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_188_io_en = _T_1110 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_188_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_189_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_189_io_en = _T_1113 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_189_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_190_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_190_io_en = _T_1116 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_190_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_191_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_191_io_en = _T_1119 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_191_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_192_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_192_io_en = _T_1122 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_192_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_193_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_193_io_en = _T_1125 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_193_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_194_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_194_io_en = _T_1128 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_194_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_195_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_195_io_en = _T_1131 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_195_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_196_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_196_io_en = _T_1134 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_196_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_197_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_197_io_en = _T_1137 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_197_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_198_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_198_io_en = _T_1140 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_198_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_199_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_199_io_en = _T_1143 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_199_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_200_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_200_io_en = _T_1146 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_200_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_201_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_201_io_en = _T_1149 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_201_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_202_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_202_io_en = _T_1152 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_202_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_203_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_203_io_en = _T_1155 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_203_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_204_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_204_io_en = _T_1158 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_204_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_205_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_205_io_en = _T_1161 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_205_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_206_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_206_io_en = _T_1164 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_206_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_207_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_207_io_en = _T_1167 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_207_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_208_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_208_io_en = _T_1170 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_208_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_209_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_209_io_en = _T_1173 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_209_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_210_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_210_io_en = _T_1176 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_210_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_211_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_211_io_en = _T_1179 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_211_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_212_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_212_io_en = _T_1182 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_212_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_213_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_213_io_en = _T_1185 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_213_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_214_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_214_io_en = _T_1188 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_214_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_215_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_215_io_en = _T_1191 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_215_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_216_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_216_io_en = _T_1194 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_216_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_217_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_217_io_en = _T_1197 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_217_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_218_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_218_io_en = _T_1200 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_218_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_219_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_219_io_en = _T_1203 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_219_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_220_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_220_io_en = _T_1206 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_220_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_221_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_221_io_en = _T_1209 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_221_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_222_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_222_io_en = _T_1212 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_222_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_223_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_223_io_en = _T_1215 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_223_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_224_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_224_io_en = _T_1218 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_224_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_225_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_225_io_en = _T_1221 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_225_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_226_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_226_io_en = _T_1224 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_226_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_227_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_227_io_en = _T_1227 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_227_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_228_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_228_io_en = _T_1230 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_228_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_229_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_229_io_en = _T_1233 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_229_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_230_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_230_io_en = _T_1236 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_230_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_231_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_231_io_en = _T_1239 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_231_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_232_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_232_io_en = _T_1242 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_232_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_233_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_233_io_en = _T_1245 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_233_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_234_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_234_io_en = _T_1248 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_234_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_235_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_235_io_en = _T_1251 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_235_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_236_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_236_io_en = _T_1254 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_236_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_237_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_237_io_en = _T_1257 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_237_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_238_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_238_io_en = _T_1260 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_238_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_239_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_239_io_en = _T_1263 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_239_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_240_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_240_io_en = _T_1266 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_240_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_241_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_241_io_en = _T_1269 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_241_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_242_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_242_io_en = _T_1272 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_242_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_243_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_243_io_en = _T_1275 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_243_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_244_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_244_io_en = _T_1278 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_244_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_245_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_245_io_en = _T_1281 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_245_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_246_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_246_io_en = _T_1284 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_246_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_247_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_247_io_en = _T_1287 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_247_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_248_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_248_io_en = _T_1290 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_248_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_249_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_249_io_en = _T_1293 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_249_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_250_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_250_io_en = _T_1296 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_250_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_251_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_251_io_en = _T_1299 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_251_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_252_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_252_io_en = _T_1302 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_252_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_253_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_253_io_en = _T_1305 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_253_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_254_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_254_io_en = _T_1308 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_254_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_255_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_255_io_en = _T_1311 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_255_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_256_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_256_io_en = _T_1314 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_256_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_257_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_257_io_en = _T_1317 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_257_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_258_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_258_io_en = _T_1320 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_258_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_259_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_259_io_en = _T_1323 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_259_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_260_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_260_io_en = _T_1326 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_260_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_261_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_261_io_en = _T_1329 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_261_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_262_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_262_io_en = _T_1332 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_262_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_263_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_263_io_en = _T_1335 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_263_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_264_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_264_io_en = _T_1338 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_264_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_265_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_265_io_en = _T_1341 & btb_wr_en_way0; // @[lib.scala 371:17]
  assign rvclkhdr_265_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_266_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_266_io_en = _T_576 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_266_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_267_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_267_io_en = _T_579 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_267_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_268_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_268_io_en = _T_582 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_268_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_269_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_269_io_en = _T_585 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_269_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_270_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_270_io_en = _T_588 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_270_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_271_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_271_io_en = _T_591 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_271_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_272_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_272_io_en = _T_594 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_272_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_273_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_273_io_en = _T_597 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_273_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_274_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_274_io_en = _T_600 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_274_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_275_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_275_io_en = _T_603 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_275_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_276_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_276_io_en = _T_606 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_276_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_277_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_277_io_en = _T_609 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_277_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_278_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_278_io_en = _T_612 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_278_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_279_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_279_io_en = _T_615 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_279_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_280_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_280_io_en = _T_618 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_280_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_281_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_281_io_en = _T_621 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_281_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_282_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_282_io_en = _T_624 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_282_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_283_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_283_io_en = _T_627 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_283_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_284_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_284_io_en = _T_630 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_284_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_285_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_285_io_en = _T_633 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_285_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_286_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_286_io_en = _T_636 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_286_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_287_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_287_io_en = _T_639 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_287_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_288_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_288_io_en = _T_642 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_288_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_289_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_289_io_en = _T_645 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_289_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_290_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_290_io_en = _T_648 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_290_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_291_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_291_io_en = _T_651 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_291_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_292_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_292_io_en = _T_654 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_292_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_293_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_293_io_en = _T_657 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_293_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_294_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_294_io_en = _T_660 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_294_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_295_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_295_io_en = _T_663 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_295_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_296_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_296_io_en = _T_666 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_296_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_297_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_297_io_en = _T_669 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_297_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_298_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_298_io_en = _T_672 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_298_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_299_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_299_io_en = _T_675 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_299_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_300_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_300_io_en = _T_678 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_300_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_301_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_301_io_en = _T_681 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_301_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_302_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_302_io_en = _T_684 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_302_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_303_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_303_io_en = _T_687 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_303_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_304_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_304_io_en = _T_690 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_304_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_305_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_305_io_en = _T_693 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_305_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_306_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_306_io_en = _T_696 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_306_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_307_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_307_io_en = _T_699 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_307_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_308_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_308_io_en = _T_702 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_308_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_309_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_309_io_en = _T_705 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_309_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_310_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_310_io_en = _T_708 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_310_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_311_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_311_io_en = _T_711 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_311_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_312_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_312_io_en = _T_714 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_312_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_313_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_313_io_en = _T_717 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_313_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_314_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_314_io_en = _T_720 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_314_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_315_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_315_io_en = _T_723 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_315_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_316_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_316_io_en = _T_726 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_316_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_317_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_317_io_en = _T_729 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_317_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_318_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_318_io_en = _T_732 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_318_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_319_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_319_io_en = _T_735 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_319_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_320_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_320_io_en = _T_738 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_320_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_321_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_321_io_en = _T_741 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_321_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_322_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_322_io_en = _T_744 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_322_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_323_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_323_io_en = _T_747 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_323_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_324_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_324_io_en = _T_750 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_324_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_325_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_325_io_en = _T_753 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_325_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_326_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_326_io_en = _T_756 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_326_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_327_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_327_io_en = _T_759 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_327_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_328_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_328_io_en = _T_762 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_328_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_329_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_329_io_en = _T_765 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_329_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_330_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_330_io_en = _T_768 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_330_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_331_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_331_io_en = _T_771 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_331_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_332_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_332_io_en = _T_774 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_332_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_333_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_333_io_en = _T_777 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_333_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_334_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_334_io_en = _T_780 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_334_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_335_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_335_io_en = _T_783 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_335_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_336_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_336_io_en = _T_786 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_336_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_337_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_337_io_en = _T_789 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_337_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_338_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_338_io_en = _T_792 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_338_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_339_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_339_io_en = _T_795 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_339_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_340_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_340_io_en = _T_798 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_340_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_341_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_341_io_en = _T_801 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_341_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_342_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_342_io_en = _T_804 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_342_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_343_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_343_io_en = _T_807 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_343_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_344_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_344_io_en = _T_810 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_344_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_345_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_345_io_en = _T_813 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_345_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_346_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_346_io_en = _T_816 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_346_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_347_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_347_io_en = _T_819 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_347_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_348_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_348_io_en = _T_822 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_348_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_349_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_349_io_en = _T_825 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_349_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_350_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_350_io_en = _T_828 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_350_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_351_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_351_io_en = _T_831 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_351_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_352_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_352_io_en = _T_834 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_352_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_353_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_353_io_en = _T_837 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_353_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_354_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_354_io_en = _T_840 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_354_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_355_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_355_io_en = _T_843 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_355_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_356_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_356_io_en = _T_846 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_356_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_357_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_357_io_en = _T_849 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_357_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_358_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_358_io_en = _T_852 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_358_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_359_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_359_io_en = _T_855 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_359_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_360_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_360_io_en = _T_858 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_360_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_361_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_361_io_en = _T_861 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_361_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_362_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_362_io_en = _T_864 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_362_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_363_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_363_io_en = _T_867 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_363_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_364_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_364_io_en = _T_870 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_364_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_365_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_365_io_en = _T_873 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_365_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_366_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_366_io_en = _T_876 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_366_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_367_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_367_io_en = _T_879 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_367_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_368_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_368_io_en = _T_882 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_368_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_369_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_369_io_en = _T_885 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_369_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_370_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_370_io_en = _T_888 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_370_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_371_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_371_io_en = _T_891 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_371_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_372_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_372_io_en = _T_894 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_372_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_373_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_373_io_en = _T_897 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_373_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_374_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_374_io_en = _T_900 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_374_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_375_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_375_io_en = _T_903 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_375_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_376_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_376_io_en = _T_906 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_376_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_377_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_377_io_en = _T_909 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_377_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_378_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_378_io_en = _T_912 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_378_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_379_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_379_io_en = _T_915 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_379_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_380_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_380_io_en = _T_918 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_380_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_381_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_381_io_en = _T_921 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_381_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_382_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_382_io_en = _T_924 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_382_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_383_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_383_io_en = _T_927 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_383_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_384_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_384_io_en = _T_930 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_384_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_385_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_385_io_en = _T_933 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_385_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_386_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_386_io_en = _T_936 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_386_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_387_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_387_io_en = _T_939 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_387_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_388_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_388_io_en = _T_942 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_388_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_389_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_389_io_en = _T_945 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_389_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_390_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_390_io_en = _T_948 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_390_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_391_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_391_io_en = _T_951 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_391_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_392_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_392_io_en = _T_954 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_392_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_393_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_393_io_en = _T_957 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_393_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_394_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_394_io_en = _T_960 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_394_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_395_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_395_io_en = _T_963 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_395_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_396_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_396_io_en = _T_966 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_396_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_397_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_397_io_en = _T_969 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_397_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_398_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_398_io_en = _T_972 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_398_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_399_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_399_io_en = _T_975 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_399_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_400_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_400_io_en = _T_978 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_400_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_401_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_401_io_en = _T_981 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_401_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_402_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_402_io_en = _T_984 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_402_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_403_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_403_io_en = _T_987 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_403_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_404_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_404_io_en = _T_990 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_404_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_405_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_405_io_en = _T_993 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_405_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_406_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_406_io_en = _T_996 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_406_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_407_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_407_io_en = _T_999 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_407_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_408_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_408_io_en = _T_1002 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_408_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_409_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_409_io_en = _T_1005 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_409_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_410_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_410_io_en = _T_1008 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_410_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_411_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_411_io_en = _T_1011 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_411_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_412_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_412_io_en = _T_1014 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_412_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_413_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_413_io_en = _T_1017 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_413_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_414_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_414_io_en = _T_1020 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_414_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_415_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_415_io_en = _T_1023 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_415_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_416_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_416_io_en = _T_1026 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_416_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_417_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_417_io_en = _T_1029 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_417_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_418_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_418_io_en = _T_1032 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_418_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_419_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_419_io_en = _T_1035 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_419_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_420_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_420_io_en = _T_1038 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_420_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_421_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_421_io_en = _T_1041 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_421_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_422_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_422_io_en = _T_1044 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_422_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_423_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_423_io_en = _T_1047 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_423_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_424_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_424_io_en = _T_1050 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_424_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_425_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_425_io_en = _T_1053 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_425_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_426_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_426_io_en = _T_1056 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_426_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_427_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_427_io_en = _T_1059 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_427_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_428_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_428_io_en = _T_1062 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_428_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_429_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_429_io_en = _T_1065 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_429_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_430_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_430_io_en = _T_1068 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_430_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_431_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_431_io_en = _T_1071 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_431_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_432_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_432_io_en = _T_1074 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_432_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_433_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_433_io_en = _T_1077 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_433_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_434_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_434_io_en = _T_1080 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_434_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_435_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_435_io_en = _T_1083 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_435_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_436_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_436_io_en = _T_1086 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_436_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_437_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_437_io_en = _T_1089 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_437_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_438_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_438_io_en = _T_1092 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_438_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_439_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_439_io_en = _T_1095 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_439_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_440_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_440_io_en = _T_1098 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_440_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_441_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_441_io_en = _T_1101 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_441_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_442_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_442_io_en = _T_1104 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_442_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_443_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_443_io_en = _T_1107 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_443_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_444_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_444_io_en = _T_1110 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_444_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_445_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_445_io_en = _T_1113 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_445_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_446_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_446_io_en = _T_1116 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_446_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_447_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_447_io_en = _T_1119 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_447_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_448_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_448_io_en = _T_1122 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_448_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_449_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_449_io_en = _T_1125 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_449_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_450_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_450_io_en = _T_1128 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_450_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_451_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_451_io_en = _T_1131 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_451_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_452_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_452_io_en = _T_1134 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_452_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_453_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_453_io_en = _T_1137 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_453_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_454_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_454_io_en = _T_1140 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_454_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_455_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_455_io_en = _T_1143 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_455_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_456_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_456_io_en = _T_1146 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_456_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_457_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_457_io_en = _T_1149 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_457_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_458_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_458_io_en = _T_1152 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_458_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_459_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_459_io_en = _T_1155 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_459_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_460_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_460_io_en = _T_1158 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_460_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_461_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_461_io_en = _T_1161 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_461_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_462_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_462_io_en = _T_1164 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_462_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_463_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_463_io_en = _T_1167 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_463_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_464_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_464_io_en = _T_1170 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_464_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_465_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_465_io_en = _T_1173 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_465_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_466_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_466_io_en = _T_1176 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_466_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_467_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_467_io_en = _T_1179 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_467_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_468_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_468_io_en = _T_1182 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_468_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_469_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_469_io_en = _T_1185 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_469_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_470_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_470_io_en = _T_1188 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_470_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_471_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_471_io_en = _T_1191 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_471_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_472_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_472_io_en = _T_1194 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_472_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_473_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_473_io_en = _T_1197 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_473_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_474_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_474_io_en = _T_1200 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_474_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_475_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_475_io_en = _T_1203 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_475_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_476_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_476_io_en = _T_1206 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_476_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_477_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_477_io_en = _T_1209 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_477_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_478_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_478_io_en = _T_1212 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_478_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_479_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_479_io_en = _T_1215 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_479_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_480_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_480_io_en = _T_1218 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_480_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_481_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_481_io_en = _T_1221 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_481_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_482_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_482_io_en = _T_1224 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_482_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_483_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_483_io_en = _T_1227 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_483_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_484_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_484_io_en = _T_1230 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_484_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_485_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_485_io_en = _T_1233 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_485_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_486_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_486_io_en = _T_1236 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_486_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_487_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_487_io_en = _T_1239 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_487_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_488_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_488_io_en = _T_1242 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_488_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_489_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_489_io_en = _T_1245 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_489_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_490_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_490_io_en = _T_1248 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_490_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_491_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_491_io_en = _T_1251 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_491_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_492_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_492_io_en = _T_1254 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_492_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_493_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_493_io_en = _T_1257 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_493_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_494_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_494_io_en = _T_1260 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_494_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_495_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_495_io_en = _T_1263 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_495_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_496_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_496_io_en = _T_1266 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_496_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_497_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_497_io_en = _T_1269 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_497_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_498_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_498_io_en = _T_1272 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_498_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_499_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_499_io_en = _T_1275 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_499_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_500_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_500_io_en = _T_1278 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_500_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_501_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_501_io_en = _T_1281 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_501_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_502_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_502_io_en = _T_1284 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_502_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_503_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_503_io_en = _T_1287 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_503_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_504_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_504_io_en = _T_1290 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_504_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_505_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_505_io_en = _T_1293 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_505_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_506_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_506_io_en = _T_1296 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_506_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_507_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_507_io_en = _T_1299 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_507_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_508_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_508_io_en = _T_1302 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_508_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_509_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_509_io_en = _T_1305 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_509_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_510_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_510_io_en = _T_1308 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_510_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_511_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_511_io_en = _T_1311 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_511_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_512_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_512_io_en = _T_1314 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_512_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_513_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_513_io_en = _T_1317 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_513_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_514_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_514_io_en = _T_1320 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_514_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_515_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_515_io_en = _T_1323 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_515_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_516_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_516_io_en = _T_1326 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_516_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_517_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_517_io_en = _T_1329 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_517_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_518_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_518_io_en = _T_1332 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_518_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_519_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_519_io_en = _T_1335 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_519_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_520_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_520_io_en = _T_1338 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_520_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_521_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_521_io_en = _T_1341 & btb_wr_en_way1; // @[lib.scala 371:17]
  assign rvclkhdr_521_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_522_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_522_io_en = _T_6212 | _T_6217; // @[lib.scala 345:16]
  assign rvclkhdr_522_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_523_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_523_io_en = _T_6223 | _T_6228; // @[lib.scala 345:16]
  assign rvclkhdr_523_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_524_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_524_io_en = _T_6234 | _T_6239; // @[lib.scala 345:16]
  assign rvclkhdr_524_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_525_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_525_io_en = _T_6245 | _T_6250; // @[lib.scala 345:16]
  assign rvclkhdr_525_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_526_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_526_io_en = _T_6256 | _T_6261; // @[lib.scala 345:16]
  assign rvclkhdr_526_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_527_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_527_io_en = _T_6267 | _T_6272; // @[lib.scala 345:16]
  assign rvclkhdr_527_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_528_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_528_io_en = _T_6278 | _T_6283; // @[lib.scala 345:16]
  assign rvclkhdr_528_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_529_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_529_io_en = _T_6289 | _T_6294; // @[lib.scala 345:16]
  assign rvclkhdr_529_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_530_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_530_io_en = _T_6300 | _T_6305; // @[lib.scala 345:16]
  assign rvclkhdr_530_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_531_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_531_io_en = _T_6311 | _T_6316; // @[lib.scala 345:16]
  assign rvclkhdr_531_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_532_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_532_io_en = _T_6322 | _T_6327; // @[lib.scala 345:16]
  assign rvclkhdr_532_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_533_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_533_io_en = _T_6333 | _T_6338; // @[lib.scala 345:16]
  assign rvclkhdr_533_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_534_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_534_io_en = _T_6344 | _T_6349; // @[lib.scala 345:16]
  assign rvclkhdr_534_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_535_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_535_io_en = _T_6355 | _T_6360; // @[lib.scala 345:16]
  assign rvclkhdr_535_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_536_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_536_io_en = _T_6366 | _T_6371; // @[lib.scala 345:16]
  assign rvclkhdr_536_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_537_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_537_io_en = _T_6377 | _T_6382; // @[lib.scala 345:16]
  assign rvclkhdr_537_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_538_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_538_io_en = _T_6388 | _T_6393; // @[lib.scala 345:16]
  assign rvclkhdr_538_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_539_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_539_io_en = _T_6399 | _T_6404; // @[lib.scala 345:16]
  assign rvclkhdr_539_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_540_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_540_io_en = _T_6410 | _T_6415; // @[lib.scala 345:16]
  assign rvclkhdr_540_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_541_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_541_io_en = _T_6421 | _T_6426; // @[lib.scala 345:16]
  assign rvclkhdr_541_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_542_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_542_io_en = _T_6432 | _T_6437; // @[lib.scala 345:16]
  assign rvclkhdr_542_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_543_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_543_io_en = _T_6443 | _T_6448; // @[lib.scala 345:16]
  assign rvclkhdr_543_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_544_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_544_io_en = _T_6454 | _T_6459; // @[lib.scala 345:16]
  assign rvclkhdr_544_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_545_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_545_io_en = _T_6465 | _T_6470; // @[lib.scala 345:16]
  assign rvclkhdr_545_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_546_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_546_io_en = _T_6476 | _T_6481; // @[lib.scala 345:16]
  assign rvclkhdr_546_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_547_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_547_io_en = _T_6487 | _T_6492; // @[lib.scala 345:16]
  assign rvclkhdr_547_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_548_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_548_io_en = _T_6498 | _T_6503; // @[lib.scala 345:16]
  assign rvclkhdr_548_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_549_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_549_io_en = _T_6509 | _T_6514; // @[lib.scala 345:16]
  assign rvclkhdr_549_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_550_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_550_io_en = _T_6520 | _T_6525; // @[lib.scala 345:16]
  assign rvclkhdr_550_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_551_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_551_io_en = _T_6531 | _T_6536; // @[lib.scala 345:16]
  assign rvclkhdr_551_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_552_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_552_io_en = _T_6542 | _T_6547; // @[lib.scala 345:16]
  assign rvclkhdr_552_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
  assign rvclkhdr_553_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_553_io_en = _T_6553 | _T_6558; // @[lib.scala 345:16]
  assign rvclkhdr_553_io_scan_mode = io_scan_mode; // @[lib.scala 346:23]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  leak_one_f_d1 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_0 = _RAND_1[21:0];
  _RAND_2 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_1 = _RAND_2[21:0];
  _RAND_3 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_2 = _RAND_3[21:0];
  _RAND_4 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_3 = _RAND_4[21:0];
  _RAND_5 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_4 = _RAND_5[21:0];
  _RAND_6 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_5 = _RAND_6[21:0];
  _RAND_7 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_6 = _RAND_7[21:0];
  _RAND_8 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_7 = _RAND_8[21:0];
  _RAND_9 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_8 = _RAND_9[21:0];
  _RAND_10 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_9 = _RAND_10[21:0];
  _RAND_11 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_10 = _RAND_11[21:0];
  _RAND_12 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_11 = _RAND_12[21:0];
  _RAND_13 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_12 = _RAND_13[21:0];
  _RAND_14 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_13 = _RAND_14[21:0];
  _RAND_15 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_14 = _RAND_15[21:0];
  _RAND_16 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_15 = _RAND_16[21:0];
  _RAND_17 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_16 = _RAND_17[21:0];
  _RAND_18 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_17 = _RAND_18[21:0];
  _RAND_19 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_18 = _RAND_19[21:0];
  _RAND_20 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_19 = _RAND_20[21:0];
  _RAND_21 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_20 = _RAND_21[21:0];
  _RAND_22 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_21 = _RAND_22[21:0];
  _RAND_23 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_22 = _RAND_23[21:0];
  _RAND_24 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_23 = _RAND_24[21:0];
  _RAND_25 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_24 = _RAND_25[21:0];
  _RAND_26 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_25 = _RAND_26[21:0];
  _RAND_27 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_26 = _RAND_27[21:0];
  _RAND_28 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_27 = _RAND_28[21:0];
  _RAND_29 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_28 = _RAND_29[21:0];
  _RAND_30 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_29 = _RAND_30[21:0];
  _RAND_31 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_30 = _RAND_31[21:0];
  _RAND_32 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_31 = _RAND_32[21:0];
  _RAND_33 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_32 = _RAND_33[21:0];
  _RAND_34 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_33 = _RAND_34[21:0];
  _RAND_35 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_34 = _RAND_35[21:0];
  _RAND_36 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_35 = _RAND_36[21:0];
  _RAND_37 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_36 = _RAND_37[21:0];
  _RAND_38 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_37 = _RAND_38[21:0];
  _RAND_39 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_38 = _RAND_39[21:0];
  _RAND_40 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_39 = _RAND_40[21:0];
  _RAND_41 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_40 = _RAND_41[21:0];
  _RAND_42 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_41 = _RAND_42[21:0];
  _RAND_43 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_42 = _RAND_43[21:0];
  _RAND_44 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_43 = _RAND_44[21:0];
  _RAND_45 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_44 = _RAND_45[21:0];
  _RAND_46 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_45 = _RAND_46[21:0];
  _RAND_47 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_46 = _RAND_47[21:0];
  _RAND_48 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_47 = _RAND_48[21:0];
  _RAND_49 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_48 = _RAND_49[21:0];
  _RAND_50 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_49 = _RAND_50[21:0];
  _RAND_51 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_50 = _RAND_51[21:0];
  _RAND_52 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_51 = _RAND_52[21:0];
  _RAND_53 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_52 = _RAND_53[21:0];
  _RAND_54 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_53 = _RAND_54[21:0];
  _RAND_55 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_54 = _RAND_55[21:0];
  _RAND_56 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_55 = _RAND_56[21:0];
  _RAND_57 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_56 = _RAND_57[21:0];
  _RAND_58 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_57 = _RAND_58[21:0];
  _RAND_59 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_58 = _RAND_59[21:0];
  _RAND_60 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_59 = _RAND_60[21:0];
  _RAND_61 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_60 = _RAND_61[21:0];
  _RAND_62 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_61 = _RAND_62[21:0];
  _RAND_63 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_62 = _RAND_63[21:0];
  _RAND_64 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_63 = _RAND_64[21:0];
  _RAND_65 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_64 = _RAND_65[21:0];
  _RAND_66 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_65 = _RAND_66[21:0];
  _RAND_67 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_66 = _RAND_67[21:0];
  _RAND_68 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_67 = _RAND_68[21:0];
  _RAND_69 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_68 = _RAND_69[21:0];
  _RAND_70 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_69 = _RAND_70[21:0];
  _RAND_71 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_70 = _RAND_71[21:0];
  _RAND_72 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_71 = _RAND_72[21:0];
  _RAND_73 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_72 = _RAND_73[21:0];
  _RAND_74 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_73 = _RAND_74[21:0];
  _RAND_75 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_74 = _RAND_75[21:0];
  _RAND_76 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_75 = _RAND_76[21:0];
  _RAND_77 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_76 = _RAND_77[21:0];
  _RAND_78 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_77 = _RAND_78[21:0];
  _RAND_79 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_78 = _RAND_79[21:0];
  _RAND_80 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_79 = _RAND_80[21:0];
  _RAND_81 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_80 = _RAND_81[21:0];
  _RAND_82 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_81 = _RAND_82[21:0];
  _RAND_83 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_82 = _RAND_83[21:0];
  _RAND_84 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_83 = _RAND_84[21:0];
  _RAND_85 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_84 = _RAND_85[21:0];
  _RAND_86 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_85 = _RAND_86[21:0];
  _RAND_87 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_86 = _RAND_87[21:0];
  _RAND_88 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_87 = _RAND_88[21:0];
  _RAND_89 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_88 = _RAND_89[21:0];
  _RAND_90 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_89 = _RAND_90[21:0];
  _RAND_91 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_90 = _RAND_91[21:0];
  _RAND_92 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_91 = _RAND_92[21:0];
  _RAND_93 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_92 = _RAND_93[21:0];
  _RAND_94 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_93 = _RAND_94[21:0];
  _RAND_95 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_94 = _RAND_95[21:0];
  _RAND_96 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_95 = _RAND_96[21:0];
  _RAND_97 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_96 = _RAND_97[21:0];
  _RAND_98 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_97 = _RAND_98[21:0];
  _RAND_99 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_98 = _RAND_99[21:0];
  _RAND_100 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_99 = _RAND_100[21:0];
  _RAND_101 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_100 = _RAND_101[21:0];
  _RAND_102 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_101 = _RAND_102[21:0];
  _RAND_103 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_102 = _RAND_103[21:0];
  _RAND_104 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_103 = _RAND_104[21:0];
  _RAND_105 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_104 = _RAND_105[21:0];
  _RAND_106 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_105 = _RAND_106[21:0];
  _RAND_107 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_106 = _RAND_107[21:0];
  _RAND_108 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_107 = _RAND_108[21:0];
  _RAND_109 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_108 = _RAND_109[21:0];
  _RAND_110 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_109 = _RAND_110[21:0];
  _RAND_111 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_110 = _RAND_111[21:0];
  _RAND_112 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_111 = _RAND_112[21:0];
  _RAND_113 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_112 = _RAND_113[21:0];
  _RAND_114 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_113 = _RAND_114[21:0];
  _RAND_115 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_114 = _RAND_115[21:0];
  _RAND_116 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_115 = _RAND_116[21:0];
  _RAND_117 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_116 = _RAND_117[21:0];
  _RAND_118 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_117 = _RAND_118[21:0];
  _RAND_119 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_118 = _RAND_119[21:0];
  _RAND_120 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_119 = _RAND_120[21:0];
  _RAND_121 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_120 = _RAND_121[21:0];
  _RAND_122 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_121 = _RAND_122[21:0];
  _RAND_123 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_122 = _RAND_123[21:0];
  _RAND_124 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_123 = _RAND_124[21:0];
  _RAND_125 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_124 = _RAND_125[21:0];
  _RAND_126 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_125 = _RAND_126[21:0];
  _RAND_127 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_126 = _RAND_127[21:0];
  _RAND_128 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_127 = _RAND_128[21:0];
  _RAND_129 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_128 = _RAND_129[21:0];
  _RAND_130 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_129 = _RAND_130[21:0];
  _RAND_131 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_130 = _RAND_131[21:0];
  _RAND_132 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_131 = _RAND_132[21:0];
  _RAND_133 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_132 = _RAND_133[21:0];
  _RAND_134 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_133 = _RAND_134[21:0];
  _RAND_135 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_134 = _RAND_135[21:0];
  _RAND_136 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_135 = _RAND_136[21:0];
  _RAND_137 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_136 = _RAND_137[21:0];
  _RAND_138 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_137 = _RAND_138[21:0];
  _RAND_139 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_138 = _RAND_139[21:0];
  _RAND_140 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_139 = _RAND_140[21:0];
  _RAND_141 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_140 = _RAND_141[21:0];
  _RAND_142 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_141 = _RAND_142[21:0];
  _RAND_143 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_142 = _RAND_143[21:0];
  _RAND_144 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_143 = _RAND_144[21:0];
  _RAND_145 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_144 = _RAND_145[21:0];
  _RAND_146 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_145 = _RAND_146[21:0];
  _RAND_147 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_146 = _RAND_147[21:0];
  _RAND_148 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_147 = _RAND_148[21:0];
  _RAND_149 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_148 = _RAND_149[21:0];
  _RAND_150 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_149 = _RAND_150[21:0];
  _RAND_151 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_150 = _RAND_151[21:0];
  _RAND_152 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_151 = _RAND_152[21:0];
  _RAND_153 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_152 = _RAND_153[21:0];
  _RAND_154 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_153 = _RAND_154[21:0];
  _RAND_155 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_154 = _RAND_155[21:0];
  _RAND_156 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_155 = _RAND_156[21:0];
  _RAND_157 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_156 = _RAND_157[21:0];
  _RAND_158 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_157 = _RAND_158[21:0];
  _RAND_159 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_158 = _RAND_159[21:0];
  _RAND_160 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_159 = _RAND_160[21:0];
  _RAND_161 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_160 = _RAND_161[21:0];
  _RAND_162 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_161 = _RAND_162[21:0];
  _RAND_163 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_162 = _RAND_163[21:0];
  _RAND_164 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_163 = _RAND_164[21:0];
  _RAND_165 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_164 = _RAND_165[21:0];
  _RAND_166 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_165 = _RAND_166[21:0];
  _RAND_167 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_166 = _RAND_167[21:0];
  _RAND_168 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_167 = _RAND_168[21:0];
  _RAND_169 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_168 = _RAND_169[21:0];
  _RAND_170 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_169 = _RAND_170[21:0];
  _RAND_171 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_170 = _RAND_171[21:0];
  _RAND_172 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_171 = _RAND_172[21:0];
  _RAND_173 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_172 = _RAND_173[21:0];
  _RAND_174 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_173 = _RAND_174[21:0];
  _RAND_175 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_174 = _RAND_175[21:0];
  _RAND_176 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_175 = _RAND_176[21:0];
  _RAND_177 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_176 = _RAND_177[21:0];
  _RAND_178 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_177 = _RAND_178[21:0];
  _RAND_179 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_178 = _RAND_179[21:0];
  _RAND_180 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_179 = _RAND_180[21:0];
  _RAND_181 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_180 = _RAND_181[21:0];
  _RAND_182 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_181 = _RAND_182[21:0];
  _RAND_183 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_182 = _RAND_183[21:0];
  _RAND_184 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_183 = _RAND_184[21:0];
  _RAND_185 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_184 = _RAND_185[21:0];
  _RAND_186 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_185 = _RAND_186[21:0];
  _RAND_187 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_186 = _RAND_187[21:0];
  _RAND_188 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_187 = _RAND_188[21:0];
  _RAND_189 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_188 = _RAND_189[21:0];
  _RAND_190 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_189 = _RAND_190[21:0];
  _RAND_191 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_190 = _RAND_191[21:0];
  _RAND_192 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_191 = _RAND_192[21:0];
  _RAND_193 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_192 = _RAND_193[21:0];
  _RAND_194 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_193 = _RAND_194[21:0];
  _RAND_195 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_194 = _RAND_195[21:0];
  _RAND_196 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_195 = _RAND_196[21:0];
  _RAND_197 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_196 = _RAND_197[21:0];
  _RAND_198 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_197 = _RAND_198[21:0];
  _RAND_199 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_198 = _RAND_199[21:0];
  _RAND_200 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_199 = _RAND_200[21:0];
  _RAND_201 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_200 = _RAND_201[21:0];
  _RAND_202 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_201 = _RAND_202[21:0];
  _RAND_203 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_202 = _RAND_203[21:0];
  _RAND_204 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_203 = _RAND_204[21:0];
  _RAND_205 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_204 = _RAND_205[21:0];
  _RAND_206 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_205 = _RAND_206[21:0];
  _RAND_207 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_206 = _RAND_207[21:0];
  _RAND_208 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_207 = _RAND_208[21:0];
  _RAND_209 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_208 = _RAND_209[21:0];
  _RAND_210 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_209 = _RAND_210[21:0];
  _RAND_211 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_210 = _RAND_211[21:0];
  _RAND_212 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_211 = _RAND_212[21:0];
  _RAND_213 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_212 = _RAND_213[21:0];
  _RAND_214 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_213 = _RAND_214[21:0];
  _RAND_215 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_214 = _RAND_215[21:0];
  _RAND_216 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_215 = _RAND_216[21:0];
  _RAND_217 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_216 = _RAND_217[21:0];
  _RAND_218 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_217 = _RAND_218[21:0];
  _RAND_219 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_218 = _RAND_219[21:0];
  _RAND_220 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_219 = _RAND_220[21:0];
  _RAND_221 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_220 = _RAND_221[21:0];
  _RAND_222 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_221 = _RAND_222[21:0];
  _RAND_223 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_222 = _RAND_223[21:0];
  _RAND_224 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_223 = _RAND_224[21:0];
  _RAND_225 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_224 = _RAND_225[21:0];
  _RAND_226 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_225 = _RAND_226[21:0];
  _RAND_227 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_226 = _RAND_227[21:0];
  _RAND_228 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_227 = _RAND_228[21:0];
  _RAND_229 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_228 = _RAND_229[21:0];
  _RAND_230 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_229 = _RAND_230[21:0];
  _RAND_231 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_230 = _RAND_231[21:0];
  _RAND_232 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_231 = _RAND_232[21:0];
  _RAND_233 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_232 = _RAND_233[21:0];
  _RAND_234 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_233 = _RAND_234[21:0];
  _RAND_235 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_234 = _RAND_235[21:0];
  _RAND_236 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_235 = _RAND_236[21:0];
  _RAND_237 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_236 = _RAND_237[21:0];
  _RAND_238 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_237 = _RAND_238[21:0];
  _RAND_239 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_238 = _RAND_239[21:0];
  _RAND_240 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_239 = _RAND_240[21:0];
  _RAND_241 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_240 = _RAND_241[21:0];
  _RAND_242 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_241 = _RAND_242[21:0];
  _RAND_243 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_242 = _RAND_243[21:0];
  _RAND_244 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_243 = _RAND_244[21:0];
  _RAND_245 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_244 = _RAND_245[21:0];
  _RAND_246 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_245 = _RAND_246[21:0];
  _RAND_247 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_246 = _RAND_247[21:0];
  _RAND_248 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_247 = _RAND_248[21:0];
  _RAND_249 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_248 = _RAND_249[21:0];
  _RAND_250 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_249 = _RAND_250[21:0];
  _RAND_251 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_250 = _RAND_251[21:0];
  _RAND_252 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_251 = _RAND_252[21:0];
  _RAND_253 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_252 = _RAND_253[21:0];
  _RAND_254 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_253 = _RAND_254[21:0];
  _RAND_255 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_254 = _RAND_255[21:0];
  _RAND_256 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_255 = _RAND_256[21:0];
  _RAND_257 = {1{`RANDOM}};
  dec_tlu_way_wb_f = _RAND_257[0:0];
  _RAND_258 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_0 = _RAND_258[21:0];
  _RAND_259 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_1 = _RAND_259[21:0];
  _RAND_260 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_2 = _RAND_260[21:0];
  _RAND_261 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_3 = _RAND_261[21:0];
  _RAND_262 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_4 = _RAND_262[21:0];
  _RAND_263 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_5 = _RAND_263[21:0];
  _RAND_264 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_6 = _RAND_264[21:0];
  _RAND_265 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_7 = _RAND_265[21:0];
  _RAND_266 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_8 = _RAND_266[21:0];
  _RAND_267 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_9 = _RAND_267[21:0];
  _RAND_268 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_10 = _RAND_268[21:0];
  _RAND_269 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_11 = _RAND_269[21:0];
  _RAND_270 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_12 = _RAND_270[21:0];
  _RAND_271 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_13 = _RAND_271[21:0];
  _RAND_272 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_14 = _RAND_272[21:0];
  _RAND_273 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_15 = _RAND_273[21:0];
  _RAND_274 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_16 = _RAND_274[21:0];
  _RAND_275 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_17 = _RAND_275[21:0];
  _RAND_276 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_18 = _RAND_276[21:0];
  _RAND_277 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_19 = _RAND_277[21:0];
  _RAND_278 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_20 = _RAND_278[21:0];
  _RAND_279 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_21 = _RAND_279[21:0];
  _RAND_280 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_22 = _RAND_280[21:0];
  _RAND_281 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_23 = _RAND_281[21:0];
  _RAND_282 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_24 = _RAND_282[21:0];
  _RAND_283 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_25 = _RAND_283[21:0];
  _RAND_284 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_26 = _RAND_284[21:0];
  _RAND_285 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_27 = _RAND_285[21:0];
  _RAND_286 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_28 = _RAND_286[21:0];
  _RAND_287 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_29 = _RAND_287[21:0];
  _RAND_288 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_30 = _RAND_288[21:0];
  _RAND_289 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_31 = _RAND_289[21:0];
  _RAND_290 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_32 = _RAND_290[21:0];
  _RAND_291 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_33 = _RAND_291[21:0];
  _RAND_292 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_34 = _RAND_292[21:0];
  _RAND_293 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_35 = _RAND_293[21:0];
  _RAND_294 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_36 = _RAND_294[21:0];
  _RAND_295 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_37 = _RAND_295[21:0];
  _RAND_296 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_38 = _RAND_296[21:0];
  _RAND_297 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_39 = _RAND_297[21:0];
  _RAND_298 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_40 = _RAND_298[21:0];
  _RAND_299 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_41 = _RAND_299[21:0];
  _RAND_300 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_42 = _RAND_300[21:0];
  _RAND_301 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_43 = _RAND_301[21:0];
  _RAND_302 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_44 = _RAND_302[21:0];
  _RAND_303 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_45 = _RAND_303[21:0];
  _RAND_304 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_46 = _RAND_304[21:0];
  _RAND_305 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_47 = _RAND_305[21:0];
  _RAND_306 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_48 = _RAND_306[21:0];
  _RAND_307 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_49 = _RAND_307[21:0];
  _RAND_308 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_50 = _RAND_308[21:0];
  _RAND_309 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_51 = _RAND_309[21:0];
  _RAND_310 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_52 = _RAND_310[21:0];
  _RAND_311 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_53 = _RAND_311[21:0];
  _RAND_312 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_54 = _RAND_312[21:0];
  _RAND_313 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_55 = _RAND_313[21:0];
  _RAND_314 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_56 = _RAND_314[21:0];
  _RAND_315 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_57 = _RAND_315[21:0];
  _RAND_316 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_58 = _RAND_316[21:0];
  _RAND_317 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_59 = _RAND_317[21:0];
  _RAND_318 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_60 = _RAND_318[21:0];
  _RAND_319 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_61 = _RAND_319[21:0];
  _RAND_320 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_62 = _RAND_320[21:0];
  _RAND_321 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_63 = _RAND_321[21:0];
  _RAND_322 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_64 = _RAND_322[21:0];
  _RAND_323 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_65 = _RAND_323[21:0];
  _RAND_324 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_66 = _RAND_324[21:0];
  _RAND_325 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_67 = _RAND_325[21:0];
  _RAND_326 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_68 = _RAND_326[21:0];
  _RAND_327 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_69 = _RAND_327[21:0];
  _RAND_328 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_70 = _RAND_328[21:0];
  _RAND_329 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_71 = _RAND_329[21:0];
  _RAND_330 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_72 = _RAND_330[21:0];
  _RAND_331 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_73 = _RAND_331[21:0];
  _RAND_332 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_74 = _RAND_332[21:0];
  _RAND_333 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_75 = _RAND_333[21:0];
  _RAND_334 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_76 = _RAND_334[21:0];
  _RAND_335 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_77 = _RAND_335[21:0];
  _RAND_336 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_78 = _RAND_336[21:0];
  _RAND_337 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_79 = _RAND_337[21:0];
  _RAND_338 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_80 = _RAND_338[21:0];
  _RAND_339 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_81 = _RAND_339[21:0];
  _RAND_340 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_82 = _RAND_340[21:0];
  _RAND_341 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_83 = _RAND_341[21:0];
  _RAND_342 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_84 = _RAND_342[21:0];
  _RAND_343 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_85 = _RAND_343[21:0];
  _RAND_344 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_86 = _RAND_344[21:0];
  _RAND_345 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_87 = _RAND_345[21:0];
  _RAND_346 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_88 = _RAND_346[21:0];
  _RAND_347 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_89 = _RAND_347[21:0];
  _RAND_348 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_90 = _RAND_348[21:0];
  _RAND_349 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_91 = _RAND_349[21:0];
  _RAND_350 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_92 = _RAND_350[21:0];
  _RAND_351 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_93 = _RAND_351[21:0];
  _RAND_352 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_94 = _RAND_352[21:0];
  _RAND_353 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_95 = _RAND_353[21:0];
  _RAND_354 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_96 = _RAND_354[21:0];
  _RAND_355 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_97 = _RAND_355[21:0];
  _RAND_356 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_98 = _RAND_356[21:0];
  _RAND_357 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_99 = _RAND_357[21:0];
  _RAND_358 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_100 = _RAND_358[21:0];
  _RAND_359 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_101 = _RAND_359[21:0];
  _RAND_360 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_102 = _RAND_360[21:0];
  _RAND_361 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_103 = _RAND_361[21:0];
  _RAND_362 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_104 = _RAND_362[21:0];
  _RAND_363 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_105 = _RAND_363[21:0];
  _RAND_364 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_106 = _RAND_364[21:0];
  _RAND_365 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_107 = _RAND_365[21:0];
  _RAND_366 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_108 = _RAND_366[21:0];
  _RAND_367 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_109 = _RAND_367[21:0];
  _RAND_368 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_110 = _RAND_368[21:0];
  _RAND_369 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_111 = _RAND_369[21:0];
  _RAND_370 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_112 = _RAND_370[21:0];
  _RAND_371 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_113 = _RAND_371[21:0];
  _RAND_372 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_114 = _RAND_372[21:0];
  _RAND_373 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_115 = _RAND_373[21:0];
  _RAND_374 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_116 = _RAND_374[21:0];
  _RAND_375 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_117 = _RAND_375[21:0];
  _RAND_376 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_118 = _RAND_376[21:0];
  _RAND_377 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_119 = _RAND_377[21:0];
  _RAND_378 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_120 = _RAND_378[21:0];
  _RAND_379 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_121 = _RAND_379[21:0];
  _RAND_380 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_122 = _RAND_380[21:0];
  _RAND_381 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_123 = _RAND_381[21:0];
  _RAND_382 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_124 = _RAND_382[21:0];
  _RAND_383 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_125 = _RAND_383[21:0];
  _RAND_384 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_126 = _RAND_384[21:0];
  _RAND_385 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_127 = _RAND_385[21:0];
  _RAND_386 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_128 = _RAND_386[21:0];
  _RAND_387 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_129 = _RAND_387[21:0];
  _RAND_388 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_130 = _RAND_388[21:0];
  _RAND_389 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_131 = _RAND_389[21:0];
  _RAND_390 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_132 = _RAND_390[21:0];
  _RAND_391 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_133 = _RAND_391[21:0];
  _RAND_392 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_134 = _RAND_392[21:0];
  _RAND_393 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_135 = _RAND_393[21:0];
  _RAND_394 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_136 = _RAND_394[21:0];
  _RAND_395 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_137 = _RAND_395[21:0];
  _RAND_396 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_138 = _RAND_396[21:0];
  _RAND_397 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_139 = _RAND_397[21:0];
  _RAND_398 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_140 = _RAND_398[21:0];
  _RAND_399 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_141 = _RAND_399[21:0];
  _RAND_400 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_142 = _RAND_400[21:0];
  _RAND_401 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_143 = _RAND_401[21:0];
  _RAND_402 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_144 = _RAND_402[21:0];
  _RAND_403 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_145 = _RAND_403[21:0];
  _RAND_404 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_146 = _RAND_404[21:0];
  _RAND_405 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_147 = _RAND_405[21:0];
  _RAND_406 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_148 = _RAND_406[21:0];
  _RAND_407 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_149 = _RAND_407[21:0];
  _RAND_408 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_150 = _RAND_408[21:0];
  _RAND_409 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_151 = _RAND_409[21:0];
  _RAND_410 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_152 = _RAND_410[21:0];
  _RAND_411 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_153 = _RAND_411[21:0];
  _RAND_412 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_154 = _RAND_412[21:0];
  _RAND_413 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_155 = _RAND_413[21:0];
  _RAND_414 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_156 = _RAND_414[21:0];
  _RAND_415 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_157 = _RAND_415[21:0];
  _RAND_416 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_158 = _RAND_416[21:0];
  _RAND_417 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_159 = _RAND_417[21:0];
  _RAND_418 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_160 = _RAND_418[21:0];
  _RAND_419 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_161 = _RAND_419[21:0];
  _RAND_420 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_162 = _RAND_420[21:0];
  _RAND_421 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_163 = _RAND_421[21:0];
  _RAND_422 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_164 = _RAND_422[21:0];
  _RAND_423 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_165 = _RAND_423[21:0];
  _RAND_424 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_166 = _RAND_424[21:0];
  _RAND_425 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_167 = _RAND_425[21:0];
  _RAND_426 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_168 = _RAND_426[21:0];
  _RAND_427 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_169 = _RAND_427[21:0];
  _RAND_428 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_170 = _RAND_428[21:0];
  _RAND_429 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_171 = _RAND_429[21:0];
  _RAND_430 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_172 = _RAND_430[21:0];
  _RAND_431 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_173 = _RAND_431[21:0];
  _RAND_432 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_174 = _RAND_432[21:0];
  _RAND_433 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_175 = _RAND_433[21:0];
  _RAND_434 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_176 = _RAND_434[21:0];
  _RAND_435 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_177 = _RAND_435[21:0];
  _RAND_436 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_178 = _RAND_436[21:0];
  _RAND_437 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_179 = _RAND_437[21:0];
  _RAND_438 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_180 = _RAND_438[21:0];
  _RAND_439 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_181 = _RAND_439[21:0];
  _RAND_440 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_182 = _RAND_440[21:0];
  _RAND_441 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_183 = _RAND_441[21:0];
  _RAND_442 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_184 = _RAND_442[21:0];
  _RAND_443 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_185 = _RAND_443[21:0];
  _RAND_444 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_186 = _RAND_444[21:0];
  _RAND_445 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_187 = _RAND_445[21:0];
  _RAND_446 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_188 = _RAND_446[21:0];
  _RAND_447 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_189 = _RAND_447[21:0];
  _RAND_448 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_190 = _RAND_448[21:0];
  _RAND_449 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_191 = _RAND_449[21:0];
  _RAND_450 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_192 = _RAND_450[21:0];
  _RAND_451 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_193 = _RAND_451[21:0];
  _RAND_452 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_194 = _RAND_452[21:0];
  _RAND_453 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_195 = _RAND_453[21:0];
  _RAND_454 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_196 = _RAND_454[21:0];
  _RAND_455 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_197 = _RAND_455[21:0];
  _RAND_456 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_198 = _RAND_456[21:0];
  _RAND_457 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_199 = _RAND_457[21:0];
  _RAND_458 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_200 = _RAND_458[21:0];
  _RAND_459 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_201 = _RAND_459[21:0];
  _RAND_460 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_202 = _RAND_460[21:0];
  _RAND_461 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_203 = _RAND_461[21:0];
  _RAND_462 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_204 = _RAND_462[21:0];
  _RAND_463 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_205 = _RAND_463[21:0];
  _RAND_464 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_206 = _RAND_464[21:0];
  _RAND_465 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_207 = _RAND_465[21:0];
  _RAND_466 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_208 = _RAND_466[21:0];
  _RAND_467 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_209 = _RAND_467[21:0];
  _RAND_468 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_210 = _RAND_468[21:0];
  _RAND_469 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_211 = _RAND_469[21:0];
  _RAND_470 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_212 = _RAND_470[21:0];
  _RAND_471 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_213 = _RAND_471[21:0];
  _RAND_472 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_214 = _RAND_472[21:0];
  _RAND_473 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_215 = _RAND_473[21:0];
  _RAND_474 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_216 = _RAND_474[21:0];
  _RAND_475 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_217 = _RAND_475[21:0];
  _RAND_476 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_218 = _RAND_476[21:0];
  _RAND_477 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_219 = _RAND_477[21:0];
  _RAND_478 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_220 = _RAND_478[21:0];
  _RAND_479 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_221 = _RAND_479[21:0];
  _RAND_480 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_222 = _RAND_480[21:0];
  _RAND_481 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_223 = _RAND_481[21:0];
  _RAND_482 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_224 = _RAND_482[21:0];
  _RAND_483 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_225 = _RAND_483[21:0];
  _RAND_484 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_226 = _RAND_484[21:0];
  _RAND_485 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_227 = _RAND_485[21:0];
  _RAND_486 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_228 = _RAND_486[21:0];
  _RAND_487 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_229 = _RAND_487[21:0];
  _RAND_488 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_230 = _RAND_488[21:0];
  _RAND_489 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_231 = _RAND_489[21:0];
  _RAND_490 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_232 = _RAND_490[21:0];
  _RAND_491 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_233 = _RAND_491[21:0];
  _RAND_492 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_234 = _RAND_492[21:0];
  _RAND_493 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_235 = _RAND_493[21:0];
  _RAND_494 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_236 = _RAND_494[21:0];
  _RAND_495 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_237 = _RAND_495[21:0];
  _RAND_496 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_238 = _RAND_496[21:0];
  _RAND_497 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_239 = _RAND_497[21:0];
  _RAND_498 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_240 = _RAND_498[21:0];
  _RAND_499 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_241 = _RAND_499[21:0];
  _RAND_500 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_242 = _RAND_500[21:0];
  _RAND_501 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_243 = _RAND_501[21:0];
  _RAND_502 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_244 = _RAND_502[21:0];
  _RAND_503 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_245 = _RAND_503[21:0];
  _RAND_504 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_246 = _RAND_504[21:0];
  _RAND_505 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_247 = _RAND_505[21:0];
  _RAND_506 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_248 = _RAND_506[21:0];
  _RAND_507 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_249 = _RAND_507[21:0];
  _RAND_508 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_250 = _RAND_508[21:0];
  _RAND_509 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_251 = _RAND_509[21:0];
  _RAND_510 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_252 = _RAND_510[21:0];
  _RAND_511 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_253 = _RAND_511[21:0];
  _RAND_512 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_254 = _RAND_512[21:0];
  _RAND_513 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_255 = _RAND_513[21:0];
  _RAND_514 = {1{`RANDOM}};
  fghr = _RAND_514[7:0];
  _RAND_515 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_0 = _RAND_515[1:0];
  _RAND_516 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_1 = _RAND_516[1:0];
  _RAND_517 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_2 = _RAND_517[1:0];
  _RAND_518 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_3 = _RAND_518[1:0];
  _RAND_519 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_4 = _RAND_519[1:0];
  _RAND_520 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_5 = _RAND_520[1:0];
  _RAND_521 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_6 = _RAND_521[1:0];
  _RAND_522 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_7 = _RAND_522[1:0];
  _RAND_523 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_8 = _RAND_523[1:0];
  _RAND_524 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_9 = _RAND_524[1:0];
  _RAND_525 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_10 = _RAND_525[1:0];
  _RAND_526 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_11 = _RAND_526[1:0];
  _RAND_527 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_12 = _RAND_527[1:0];
  _RAND_528 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_13 = _RAND_528[1:0];
  _RAND_529 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_14 = _RAND_529[1:0];
  _RAND_530 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_15 = _RAND_530[1:0];
  _RAND_531 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_16 = _RAND_531[1:0];
  _RAND_532 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_17 = _RAND_532[1:0];
  _RAND_533 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_18 = _RAND_533[1:0];
  _RAND_534 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_19 = _RAND_534[1:0];
  _RAND_535 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_20 = _RAND_535[1:0];
  _RAND_536 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_21 = _RAND_536[1:0];
  _RAND_537 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_22 = _RAND_537[1:0];
  _RAND_538 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_23 = _RAND_538[1:0];
  _RAND_539 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_24 = _RAND_539[1:0];
  _RAND_540 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_25 = _RAND_540[1:0];
  _RAND_541 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_26 = _RAND_541[1:0];
  _RAND_542 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_27 = _RAND_542[1:0];
  _RAND_543 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_28 = _RAND_543[1:0];
  _RAND_544 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_29 = _RAND_544[1:0];
  _RAND_545 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_30 = _RAND_545[1:0];
  _RAND_546 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_31 = _RAND_546[1:0];
  _RAND_547 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_32 = _RAND_547[1:0];
  _RAND_548 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_33 = _RAND_548[1:0];
  _RAND_549 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_34 = _RAND_549[1:0];
  _RAND_550 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_35 = _RAND_550[1:0];
  _RAND_551 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_36 = _RAND_551[1:0];
  _RAND_552 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_37 = _RAND_552[1:0];
  _RAND_553 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_38 = _RAND_553[1:0];
  _RAND_554 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_39 = _RAND_554[1:0];
  _RAND_555 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_40 = _RAND_555[1:0];
  _RAND_556 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_41 = _RAND_556[1:0];
  _RAND_557 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_42 = _RAND_557[1:0];
  _RAND_558 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_43 = _RAND_558[1:0];
  _RAND_559 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_44 = _RAND_559[1:0];
  _RAND_560 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_45 = _RAND_560[1:0];
  _RAND_561 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_46 = _RAND_561[1:0];
  _RAND_562 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_47 = _RAND_562[1:0];
  _RAND_563 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_48 = _RAND_563[1:0];
  _RAND_564 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_49 = _RAND_564[1:0];
  _RAND_565 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_50 = _RAND_565[1:0];
  _RAND_566 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_51 = _RAND_566[1:0];
  _RAND_567 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_52 = _RAND_567[1:0];
  _RAND_568 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_53 = _RAND_568[1:0];
  _RAND_569 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_54 = _RAND_569[1:0];
  _RAND_570 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_55 = _RAND_570[1:0];
  _RAND_571 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_56 = _RAND_571[1:0];
  _RAND_572 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_57 = _RAND_572[1:0];
  _RAND_573 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_58 = _RAND_573[1:0];
  _RAND_574 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_59 = _RAND_574[1:0];
  _RAND_575 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_60 = _RAND_575[1:0];
  _RAND_576 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_61 = _RAND_576[1:0];
  _RAND_577 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_62 = _RAND_577[1:0];
  _RAND_578 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_63 = _RAND_578[1:0];
  _RAND_579 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_64 = _RAND_579[1:0];
  _RAND_580 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_65 = _RAND_580[1:0];
  _RAND_581 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_66 = _RAND_581[1:0];
  _RAND_582 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_67 = _RAND_582[1:0];
  _RAND_583 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_68 = _RAND_583[1:0];
  _RAND_584 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_69 = _RAND_584[1:0];
  _RAND_585 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_70 = _RAND_585[1:0];
  _RAND_586 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_71 = _RAND_586[1:0];
  _RAND_587 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_72 = _RAND_587[1:0];
  _RAND_588 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_73 = _RAND_588[1:0];
  _RAND_589 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_74 = _RAND_589[1:0];
  _RAND_590 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_75 = _RAND_590[1:0];
  _RAND_591 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_76 = _RAND_591[1:0];
  _RAND_592 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_77 = _RAND_592[1:0];
  _RAND_593 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_78 = _RAND_593[1:0];
  _RAND_594 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_79 = _RAND_594[1:0];
  _RAND_595 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_80 = _RAND_595[1:0];
  _RAND_596 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_81 = _RAND_596[1:0];
  _RAND_597 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_82 = _RAND_597[1:0];
  _RAND_598 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_83 = _RAND_598[1:0];
  _RAND_599 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_84 = _RAND_599[1:0];
  _RAND_600 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_85 = _RAND_600[1:0];
  _RAND_601 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_86 = _RAND_601[1:0];
  _RAND_602 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_87 = _RAND_602[1:0];
  _RAND_603 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_88 = _RAND_603[1:0];
  _RAND_604 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_89 = _RAND_604[1:0];
  _RAND_605 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_90 = _RAND_605[1:0];
  _RAND_606 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_91 = _RAND_606[1:0];
  _RAND_607 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_92 = _RAND_607[1:0];
  _RAND_608 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_93 = _RAND_608[1:0];
  _RAND_609 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_94 = _RAND_609[1:0];
  _RAND_610 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_95 = _RAND_610[1:0];
  _RAND_611 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_96 = _RAND_611[1:0];
  _RAND_612 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_97 = _RAND_612[1:0];
  _RAND_613 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_98 = _RAND_613[1:0];
  _RAND_614 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_99 = _RAND_614[1:0];
  _RAND_615 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_100 = _RAND_615[1:0];
  _RAND_616 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_101 = _RAND_616[1:0];
  _RAND_617 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_102 = _RAND_617[1:0];
  _RAND_618 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_103 = _RAND_618[1:0];
  _RAND_619 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_104 = _RAND_619[1:0];
  _RAND_620 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_105 = _RAND_620[1:0];
  _RAND_621 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_106 = _RAND_621[1:0];
  _RAND_622 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_107 = _RAND_622[1:0];
  _RAND_623 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_108 = _RAND_623[1:0];
  _RAND_624 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_109 = _RAND_624[1:0];
  _RAND_625 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_110 = _RAND_625[1:0];
  _RAND_626 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_111 = _RAND_626[1:0];
  _RAND_627 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_112 = _RAND_627[1:0];
  _RAND_628 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_113 = _RAND_628[1:0];
  _RAND_629 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_114 = _RAND_629[1:0];
  _RAND_630 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_115 = _RAND_630[1:0];
  _RAND_631 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_116 = _RAND_631[1:0];
  _RAND_632 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_117 = _RAND_632[1:0];
  _RAND_633 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_118 = _RAND_633[1:0];
  _RAND_634 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_119 = _RAND_634[1:0];
  _RAND_635 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_120 = _RAND_635[1:0];
  _RAND_636 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_121 = _RAND_636[1:0];
  _RAND_637 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_122 = _RAND_637[1:0];
  _RAND_638 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_123 = _RAND_638[1:0];
  _RAND_639 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_124 = _RAND_639[1:0];
  _RAND_640 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_125 = _RAND_640[1:0];
  _RAND_641 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_126 = _RAND_641[1:0];
  _RAND_642 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_127 = _RAND_642[1:0];
  _RAND_643 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_128 = _RAND_643[1:0];
  _RAND_644 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_129 = _RAND_644[1:0];
  _RAND_645 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_130 = _RAND_645[1:0];
  _RAND_646 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_131 = _RAND_646[1:0];
  _RAND_647 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_132 = _RAND_647[1:0];
  _RAND_648 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_133 = _RAND_648[1:0];
  _RAND_649 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_134 = _RAND_649[1:0];
  _RAND_650 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_135 = _RAND_650[1:0];
  _RAND_651 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_136 = _RAND_651[1:0];
  _RAND_652 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_137 = _RAND_652[1:0];
  _RAND_653 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_138 = _RAND_653[1:0];
  _RAND_654 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_139 = _RAND_654[1:0];
  _RAND_655 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_140 = _RAND_655[1:0];
  _RAND_656 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_141 = _RAND_656[1:0];
  _RAND_657 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_142 = _RAND_657[1:0];
  _RAND_658 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_143 = _RAND_658[1:0];
  _RAND_659 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_144 = _RAND_659[1:0];
  _RAND_660 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_145 = _RAND_660[1:0];
  _RAND_661 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_146 = _RAND_661[1:0];
  _RAND_662 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_147 = _RAND_662[1:0];
  _RAND_663 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_148 = _RAND_663[1:0];
  _RAND_664 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_149 = _RAND_664[1:0];
  _RAND_665 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_150 = _RAND_665[1:0];
  _RAND_666 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_151 = _RAND_666[1:0];
  _RAND_667 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_152 = _RAND_667[1:0];
  _RAND_668 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_153 = _RAND_668[1:0];
  _RAND_669 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_154 = _RAND_669[1:0];
  _RAND_670 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_155 = _RAND_670[1:0];
  _RAND_671 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_156 = _RAND_671[1:0];
  _RAND_672 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_157 = _RAND_672[1:0];
  _RAND_673 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_158 = _RAND_673[1:0];
  _RAND_674 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_159 = _RAND_674[1:0];
  _RAND_675 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_160 = _RAND_675[1:0];
  _RAND_676 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_161 = _RAND_676[1:0];
  _RAND_677 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_162 = _RAND_677[1:0];
  _RAND_678 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_163 = _RAND_678[1:0];
  _RAND_679 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_164 = _RAND_679[1:0];
  _RAND_680 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_165 = _RAND_680[1:0];
  _RAND_681 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_166 = _RAND_681[1:0];
  _RAND_682 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_167 = _RAND_682[1:0];
  _RAND_683 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_168 = _RAND_683[1:0];
  _RAND_684 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_169 = _RAND_684[1:0];
  _RAND_685 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_170 = _RAND_685[1:0];
  _RAND_686 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_171 = _RAND_686[1:0];
  _RAND_687 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_172 = _RAND_687[1:0];
  _RAND_688 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_173 = _RAND_688[1:0];
  _RAND_689 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_174 = _RAND_689[1:0];
  _RAND_690 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_175 = _RAND_690[1:0];
  _RAND_691 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_176 = _RAND_691[1:0];
  _RAND_692 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_177 = _RAND_692[1:0];
  _RAND_693 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_178 = _RAND_693[1:0];
  _RAND_694 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_179 = _RAND_694[1:0];
  _RAND_695 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_180 = _RAND_695[1:0];
  _RAND_696 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_181 = _RAND_696[1:0];
  _RAND_697 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_182 = _RAND_697[1:0];
  _RAND_698 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_183 = _RAND_698[1:0];
  _RAND_699 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_184 = _RAND_699[1:0];
  _RAND_700 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_185 = _RAND_700[1:0];
  _RAND_701 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_186 = _RAND_701[1:0];
  _RAND_702 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_187 = _RAND_702[1:0];
  _RAND_703 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_188 = _RAND_703[1:0];
  _RAND_704 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_189 = _RAND_704[1:0];
  _RAND_705 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_190 = _RAND_705[1:0];
  _RAND_706 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_191 = _RAND_706[1:0];
  _RAND_707 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_192 = _RAND_707[1:0];
  _RAND_708 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_193 = _RAND_708[1:0];
  _RAND_709 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_194 = _RAND_709[1:0];
  _RAND_710 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_195 = _RAND_710[1:0];
  _RAND_711 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_196 = _RAND_711[1:0];
  _RAND_712 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_197 = _RAND_712[1:0];
  _RAND_713 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_198 = _RAND_713[1:0];
  _RAND_714 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_199 = _RAND_714[1:0];
  _RAND_715 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_200 = _RAND_715[1:0];
  _RAND_716 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_201 = _RAND_716[1:0];
  _RAND_717 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_202 = _RAND_717[1:0];
  _RAND_718 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_203 = _RAND_718[1:0];
  _RAND_719 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_204 = _RAND_719[1:0];
  _RAND_720 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_205 = _RAND_720[1:0];
  _RAND_721 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_206 = _RAND_721[1:0];
  _RAND_722 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_207 = _RAND_722[1:0];
  _RAND_723 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_208 = _RAND_723[1:0];
  _RAND_724 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_209 = _RAND_724[1:0];
  _RAND_725 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_210 = _RAND_725[1:0];
  _RAND_726 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_211 = _RAND_726[1:0];
  _RAND_727 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_212 = _RAND_727[1:0];
  _RAND_728 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_213 = _RAND_728[1:0];
  _RAND_729 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_214 = _RAND_729[1:0];
  _RAND_730 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_215 = _RAND_730[1:0];
  _RAND_731 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_216 = _RAND_731[1:0];
  _RAND_732 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_217 = _RAND_732[1:0];
  _RAND_733 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_218 = _RAND_733[1:0];
  _RAND_734 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_219 = _RAND_734[1:0];
  _RAND_735 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_220 = _RAND_735[1:0];
  _RAND_736 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_221 = _RAND_736[1:0];
  _RAND_737 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_222 = _RAND_737[1:0];
  _RAND_738 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_223 = _RAND_738[1:0];
  _RAND_739 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_224 = _RAND_739[1:0];
  _RAND_740 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_225 = _RAND_740[1:0];
  _RAND_741 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_226 = _RAND_741[1:0];
  _RAND_742 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_227 = _RAND_742[1:0];
  _RAND_743 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_228 = _RAND_743[1:0];
  _RAND_744 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_229 = _RAND_744[1:0];
  _RAND_745 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_230 = _RAND_745[1:0];
  _RAND_746 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_231 = _RAND_746[1:0];
  _RAND_747 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_232 = _RAND_747[1:0];
  _RAND_748 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_233 = _RAND_748[1:0];
  _RAND_749 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_234 = _RAND_749[1:0];
  _RAND_750 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_235 = _RAND_750[1:0];
  _RAND_751 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_236 = _RAND_751[1:0];
  _RAND_752 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_237 = _RAND_752[1:0];
  _RAND_753 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_238 = _RAND_753[1:0];
  _RAND_754 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_239 = _RAND_754[1:0];
  _RAND_755 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_240 = _RAND_755[1:0];
  _RAND_756 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_241 = _RAND_756[1:0];
  _RAND_757 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_242 = _RAND_757[1:0];
  _RAND_758 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_243 = _RAND_758[1:0];
  _RAND_759 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_244 = _RAND_759[1:0];
  _RAND_760 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_245 = _RAND_760[1:0];
  _RAND_761 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_246 = _RAND_761[1:0];
  _RAND_762 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_247 = _RAND_762[1:0];
  _RAND_763 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_248 = _RAND_763[1:0];
  _RAND_764 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_249 = _RAND_764[1:0];
  _RAND_765 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_250 = _RAND_765[1:0];
  _RAND_766 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_251 = _RAND_766[1:0];
  _RAND_767 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_252 = _RAND_767[1:0];
  _RAND_768 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_253 = _RAND_768[1:0];
  _RAND_769 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_254 = _RAND_769[1:0];
  _RAND_770 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_255 = _RAND_770[1:0];
  _RAND_771 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_0 = _RAND_771[1:0];
  _RAND_772 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_1 = _RAND_772[1:0];
  _RAND_773 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_2 = _RAND_773[1:0];
  _RAND_774 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_3 = _RAND_774[1:0];
  _RAND_775 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_4 = _RAND_775[1:0];
  _RAND_776 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_5 = _RAND_776[1:0];
  _RAND_777 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_6 = _RAND_777[1:0];
  _RAND_778 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_7 = _RAND_778[1:0];
  _RAND_779 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_8 = _RAND_779[1:0];
  _RAND_780 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_9 = _RAND_780[1:0];
  _RAND_781 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_10 = _RAND_781[1:0];
  _RAND_782 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_11 = _RAND_782[1:0];
  _RAND_783 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_12 = _RAND_783[1:0];
  _RAND_784 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_13 = _RAND_784[1:0];
  _RAND_785 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_14 = _RAND_785[1:0];
  _RAND_786 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_15 = _RAND_786[1:0];
  _RAND_787 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_16 = _RAND_787[1:0];
  _RAND_788 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_17 = _RAND_788[1:0];
  _RAND_789 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_18 = _RAND_789[1:0];
  _RAND_790 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_19 = _RAND_790[1:0];
  _RAND_791 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_20 = _RAND_791[1:0];
  _RAND_792 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_21 = _RAND_792[1:0];
  _RAND_793 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_22 = _RAND_793[1:0];
  _RAND_794 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_23 = _RAND_794[1:0];
  _RAND_795 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_24 = _RAND_795[1:0];
  _RAND_796 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_25 = _RAND_796[1:0];
  _RAND_797 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_26 = _RAND_797[1:0];
  _RAND_798 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_27 = _RAND_798[1:0];
  _RAND_799 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_28 = _RAND_799[1:0];
  _RAND_800 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_29 = _RAND_800[1:0];
  _RAND_801 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_30 = _RAND_801[1:0];
  _RAND_802 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_31 = _RAND_802[1:0];
  _RAND_803 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_32 = _RAND_803[1:0];
  _RAND_804 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_33 = _RAND_804[1:0];
  _RAND_805 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_34 = _RAND_805[1:0];
  _RAND_806 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_35 = _RAND_806[1:0];
  _RAND_807 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_36 = _RAND_807[1:0];
  _RAND_808 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_37 = _RAND_808[1:0];
  _RAND_809 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_38 = _RAND_809[1:0];
  _RAND_810 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_39 = _RAND_810[1:0];
  _RAND_811 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_40 = _RAND_811[1:0];
  _RAND_812 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_41 = _RAND_812[1:0];
  _RAND_813 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_42 = _RAND_813[1:0];
  _RAND_814 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_43 = _RAND_814[1:0];
  _RAND_815 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_44 = _RAND_815[1:0];
  _RAND_816 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_45 = _RAND_816[1:0];
  _RAND_817 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_46 = _RAND_817[1:0];
  _RAND_818 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_47 = _RAND_818[1:0];
  _RAND_819 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_48 = _RAND_819[1:0];
  _RAND_820 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_49 = _RAND_820[1:0];
  _RAND_821 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_50 = _RAND_821[1:0];
  _RAND_822 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_51 = _RAND_822[1:0];
  _RAND_823 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_52 = _RAND_823[1:0];
  _RAND_824 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_53 = _RAND_824[1:0];
  _RAND_825 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_54 = _RAND_825[1:0];
  _RAND_826 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_55 = _RAND_826[1:0];
  _RAND_827 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_56 = _RAND_827[1:0];
  _RAND_828 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_57 = _RAND_828[1:0];
  _RAND_829 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_58 = _RAND_829[1:0];
  _RAND_830 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_59 = _RAND_830[1:0];
  _RAND_831 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_60 = _RAND_831[1:0];
  _RAND_832 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_61 = _RAND_832[1:0];
  _RAND_833 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_62 = _RAND_833[1:0];
  _RAND_834 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_63 = _RAND_834[1:0];
  _RAND_835 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_64 = _RAND_835[1:0];
  _RAND_836 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_65 = _RAND_836[1:0];
  _RAND_837 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_66 = _RAND_837[1:0];
  _RAND_838 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_67 = _RAND_838[1:0];
  _RAND_839 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_68 = _RAND_839[1:0];
  _RAND_840 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_69 = _RAND_840[1:0];
  _RAND_841 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_70 = _RAND_841[1:0];
  _RAND_842 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_71 = _RAND_842[1:0];
  _RAND_843 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_72 = _RAND_843[1:0];
  _RAND_844 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_73 = _RAND_844[1:0];
  _RAND_845 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_74 = _RAND_845[1:0];
  _RAND_846 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_75 = _RAND_846[1:0];
  _RAND_847 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_76 = _RAND_847[1:0];
  _RAND_848 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_77 = _RAND_848[1:0];
  _RAND_849 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_78 = _RAND_849[1:0];
  _RAND_850 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_79 = _RAND_850[1:0];
  _RAND_851 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_80 = _RAND_851[1:0];
  _RAND_852 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_81 = _RAND_852[1:0];
  _RAND_853 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_82 = _RAND_853[1:0];
  _RAND_854 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_83 = _RAND_854[1:0];
  _RAND_855 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_84 = _RAND_855[1:0];
  _RAND_856 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_85 = _RAND_856[1:0];
  _RAND_857 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_86 = _RAND_857[1:0];
  _RAND_858 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_87 = _RAND_858[1:0];
  _RAND_859 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_88 = _RAND_859[1:0];
  _RAND_860 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_89 = _RAND_860[1:0];
  _RAND_861 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_90 = _RAND_861[1:0];
  _RAND_862 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_91 = _RAND_862[1:0];
  _RAND_863 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_92 = _RAND_863[1:0];
  _RAND_864 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_93 = _RAND_864[1:0];
  _RAND_865 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_94 = _RAND_865[1:0];
  _RAND_866 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_95 = _RAND_866[1:0];
  _RAND_867 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_96 = _RAND_867[1:0];
  _RAND_868 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_97 = _RAND_868[1:0];
  _RAND_869 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_98 = _RAND_869[1:0];
  _RAND_870 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_99 = _RAND_870[1:0];
  _RAND_871 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_100 = _RAND_871[1:0];
  _RAND_872 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_101 = _RAND_872[1:0];
  _RAND_873 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_102 = _RAND_873[1:0];
  _RAND_874 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_103 = _RAND_874[1:0];
  _RAND_875 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_104 = _RAND_875[1:0];
  _RAND_876 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_105 = _RAND_876[1:0];
  _RAND_877 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_106 = _RAND_877[1:0];
  _RAND_878 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_107 = _RAND_878[1:0];
  _RAND_879 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_108 = _RAND_879[1:0];
  _RAND_880 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_109 = _RAND_880[1:0];
  _RAND_881 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_110 = _RAND_881[1:0];
  _RAND_882 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_111 = _RAND_882[1:0];
  _RAND_883 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_112 = _RAND_883[1:0];
  _RAND_884 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_113 = _RAND_884[1:0];
  _RAND_885 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_114 = _RAND_885[1:0];
  _RAND_886 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_115 = _RAND_886[1:0];
  _RAND_887 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_116 = _RAND_887[1:0];
  _RAND_888 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_117 = _RAND_888[1:0];
  _RAND_889 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_118 = _RAND_889[1:0];
  _RAND_890 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_119 = _RAND_890[1:0];
  _RAND_891 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_120 = _RAND_891[1:0];
  _RAND_892 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_121 = _RAND_892[1:0];
  _RAND_893 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_122 = _RAND_893[1:0];
  _RAND_894 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_123 = _RAND_894[1:0];
  _RAND_895 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_124 = _RAND_895[1:0];
  _RAND_896 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_125 = _RAND_896[1:0];
  _RAND_897 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_126 = _RAND_897[1:0];
  _RAND_898 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_127 = _RAND_898[1:0];
  _RAND_899 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_128 = _RAND_899[1:0];
  _RAND_900 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_129 = _RAND_900[1:0];
  _RAND_901 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_130 = _RAND_901[1:0];
  _RAND_902 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_131 = _RAND_902[1:0];
  _RAND_903 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_132 = _RAND_903[1:0];
  _RAND_904 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_133 = _RAND_904[1:0];
  _RAND_905 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_134 = _RAND_905[1:0];
  _RAND_906 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_135 = _RAND_906[1:0];
  _RAND_907 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_136 = _RAND_907[1:0];
  _RAND_908 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_137 = _RAND_908[1:0];
  _RAND_909 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_138 = _RAND_909[1:0];
  _RAND_910 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_139 = _RAND_910[1:0];
  _RAND_911 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_140 = _RAND_911[1:0];
  _RAND_912 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_141 = _RAND_912[1:0];
  _RAND_913 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_142 = _RAND_913[1:0];
  _RAND_914 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_143 = _RAND_914[1:0];
  _RAND_915 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_144 = _RAND_915[1:0];
  _RAND_916 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_145 = _RAND_916[1:0];
  _RAND_917 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_146 = _RAND_917[1:0];
  _RAND_918 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_147 = _RAND_918[1:0];
  _RAND_919 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_148 = _RAND_919[1:0];
  _RAND_920 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_149 = _RAND_920[1:0];
  _RAND_921 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_150 = _RAND_921[1:0];
  _RAND_922 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_151 = _RAND_922[1:0];
  _RAND_923 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_152 = _RAND_923[1:0];
  _RAND_924 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_153 = _RAND_924[1:0];
  _RAND_925 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_154 = _RAND_925[1:0];
  _RAND_926 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_155 = _RAND_926[1:0];
  _RAND_927 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_156 = _RAND_927[1:0];
  _RAND_928 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_157 = _RAND_928[1:0];
  _RAND_929 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_158 = _RAND_929[1:0];
  _RAND_930 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_159 = _RAND_930[1:0];
  _RAND_931 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_160 = _RAND_931[1:0];
  _RAND_932 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_161 = _RAND_932[1:0];
  _RAND_933 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_162 = _RAND_933[1:0];
  _RAND_934 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_163 = _RAND_934[1:0];
  _RAND_935 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_164 = _RAND_935[1:0];
  _RAND_936 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_165 = _RAND_936[1:0];
  _RAND_937 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_166 = _RAND_937[1:0];
  _RAND_938 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_167 = _RAND_938[1:0];
  _RAND_939 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_168 = _RAND_939[1:0];
  _RAND_940 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_169 = _RAND_940[1:0];
  _RAND_941 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_170 = _RAND_941[1:0];
  _RAND_942 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_171 = _RAND_942[1:0];
  _RAND_943 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_172 = _RAND_943[1:0];
  _RAND_944 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_173 = _RAND_944[1:0];
  _RAND_945 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_174 = _RAND_945[1:0];
  _RAND_946 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_175 = _RAND_946[1:0];
  _RAND_947 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_176 = _RAND_947[1:0];
  _RAND_948 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_177 = _RAND_948[1:0];
  _RAND_949 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_178 = _RAND_949[1:0];
  _RAND_950 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_179 = _RAND_950[1:0];
  _RAND_951 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_180 = _RAND_951[1:0];
  _RAND_952 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_181 = _RAND_952[1:0];
  _RAND_953 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_182 = _RAND_953[1:0];
  _RAND_954 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_183 = _RAND_954[1:0];
  _RAND_955 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_184 = _RAND_955[1:0];
  _RAND_956 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_185 = _RAND_956[1:0];
  _RAND_957 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_186 = _RAND_957[1:0];
  _RAND_958 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_187 = _RAND_958[1:0];
  _RAND_959 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_188 = _RAND_959[1:0];
  _RAND_960 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_189 = _RAND_960[1:0];
  _RAND_961 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_190 = _RAND_961[1:0];
  _RAND_962 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_191 = _RAND_962[1:0];
  _RAND_963 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_192 = _RAND_963[1:0];
  _RAND_964 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_193 = _RAND_964[1:0];
  _RAND_965 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_194 = _RAND_965[1:0];
  _RAND_966 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_195 = _RAND_966[1:0];
  _RAND_967 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_196 = _RAND_967[1:0];
  _RAND_968 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_197 = _RAND_968[1:0];
  _RAND_969 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_198 = _RAND_969[1:0];
  _RAND_970 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_199 = _RAND_970[1:0];
  _RAND_971 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_200 = _RAND_971[1:0];
  _RAND_972 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_201 = _RAND_972[1:0];
  _RAND_973 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_202 = _RAND_973[1:0];
  _RAND_974 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_203 = _RAND_974[1:0];
  _RAND_975 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_204 = _RAND_975[1:0];
  _RAND_976 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_205 = _RAND_976[1:0];
  _RAND_977 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_206 = _RAND_977[1:0];
  _RAND_978 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_207 = _RAND_978[1:0];
  _RAND_979 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_208 = _RAND_979[1:0];
  _RAND_980 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_209 = _RAND_980[1:0];
  _RAND_981 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_210 = _RAND_981[1:0];
  _RAND_982 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_211 = _RAND_982[1:0];
  _RAND_983 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_212 = _RAND_983[1:0];
  _RAND_984 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_213 = _RAND_984[1:0];
  _RAND_985 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_214 = _RAND_985[1:0];
  _RAND_986 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_215 = _RAND_986[1:0];
  _RAND_987 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_216 = _RAND_987[1:0];
  _RAND_988 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_217 = _RAND_988[1:0];
  _RAND_989 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_218 = _RAND_989[1:0];
  _RAND_990 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_219 = _RAND_990[1:0];
  _RAND_991 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_220 = _RAND_991[1:0];
  _RAND_992 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_221 = _RAND_992[1:0];
  _RAND_993 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_222 = _RAND_993[1:0];
  _RAND_994 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_223 = _RAND_994[1:0];
  _RAND_995 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_224 = _RAND_995[1:0];
  _RAND_996 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_225 = _RAND_996[1:0];
  _RAND_997 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_226 = _RAND_997[1:0];
  _RAND_998 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_227 = _RAND_998[1:0];
  _RAND_999 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_228 = _RAND_999[1:0];
  _RAND_1000 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_229 = _RAND_1000[1:0];
  _RAND_1001 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_230 = _RAND_1001[1:0];
  _RAND_1002 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_231 = _RAND_1002[1:0];
  _RAND_1003 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_232 = _RAND_1003[1:0];
  _RAND_1004 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_233 = _RAND_1004[1:0];
  _RAND_1005 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_234 = _RAND_1005[1:0];
  _RAND_1006 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_235 = _RAND_1006[1:0];
  _RAND_1007 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_236 = _RAND_1007[1:0];
  _RAND_1008 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_237 = _RAND_1008[1:0];
  _RAND_1009 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_238 = _RAND_1009[1:0];
  _RAND_1010 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_239 = _RAND_1010[1:0];
  _RAND_1011 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_240 = _RAND_1011[1:0];
  _RAND_1012 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_241 = _RAND_1012[1:0];
  _RAND_1013 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_242 = _RAND_1013[1:0];
  _RAND_1014 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_243 = _RAND_1014[1:0];
  _RAND_1015 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_244 = _RAND_1015[1:0];
  _RAND_1016 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_245 = _RAND_1016[1:0];
  _RAND_1017 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_246 = _RAND_1017[1:0];
  _RAND_1018 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_247 = _RAND_1018[1:0];
  _RAND_1019 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_248 = _RAND_1019[1:0];
  _RAND_1020 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_249 = _RAND_1020[1:0];
  _RAND_1021 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_250 = _RAND_1021[1:0];
  _RAND_1022 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_251 = _RAND_1022[1:0];
  _RAND_1023 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_252 = _RAND_1023[1:0];
  _RAND_1024 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_253 = _RAND_1024[1:0];
  _RAND_1025 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_254 = _RAND_1025[1:0];
  _RAND_1026 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_255 = _RAND_1026[1:0];
  _RAND_1027 = {1{`RANDOM}};
  exu_mp_way_f = _RAND_1027[0:0];
  _RAND_1028 = {1{`RANDOM}};
  exu_flush_final_d1 = _RAND_1028[0:0];
  _RAND_1029 = {8{`RANDOM}};
  btb_lru_b0_f = _RAND_1029[255:0];
  _RAND_1030 = {1{`RANDOM}};
  ifc_fetch_adder_prior = _RAND_1030[29:0];
  _RAND_1031 = {1{`RANDOM}};
  rets_out_0 = _RAND_1031[31:0];
  _RAND_1032 = {1{`RANDOM}};
  rets_out_1 = _RAND_1032[31:0];
  _RAND_1033 = {1{`RANDOM}};
  rets_out_2 = _RAND_1033[31:0];
  _RAND_1034 = {1{`RANDOM}};
  rets_out_3 = _RAND_1034[31:0];
  _RAND_1035 = {1{`RANDOM}};
  rets_out_4 = _RAND_1035[31:0];
  _RAND_1036 = {1{`RANDOM}};
  rets_out_5 = _RAND_1036[31:0];
  _RAND_1037 = {1{`RANDOM}};
  rets_out_6 = _RAND_1037[31:0];
  _RAND_1038 = {1{`RANDOM}};
  rets_out_7 = _RAND_1038[31:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    leak_one_f_d1 = 1'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_0 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_1 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_2 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_3 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_4 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_5 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_6 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_7 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_8 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_9 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_10 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_11 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_12 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_13 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_14 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_15 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_16 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_17 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_18 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_19 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_20 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_21 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_22 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_23 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_24 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_25 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_26 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_27 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_28 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_29 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_30 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_31 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_32 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_33 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_34 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_35 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_36 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_37 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_38 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_39 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_40 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_41 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_42 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_43 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_44 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_45 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_46 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_47 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_48 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_49 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_50 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_51 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_52 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_53 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_54 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_55 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_56 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_57 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_58 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_59 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_60 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_61 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_62 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_63 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_64 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_65 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_66 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_67 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_68 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_69 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_70 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_71 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_72 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_73 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_74 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_75 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_76 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_77 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_78 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_79 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_80 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_81 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_82 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_83 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_84 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_85 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_86 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_87 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_88 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_89 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_90 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_91 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_92 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_93 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_94 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_95 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_96 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_97 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_98 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_99 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_100 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_101 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_102 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_103 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_104 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_105 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_106 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_107 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_108 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_109 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_110 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_111 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_112 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_113 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_114 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_115 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_116 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_117 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_118 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_119 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_120 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_121 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_122 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_123 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_124 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_125 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_126 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_127 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_128 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_129 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_130 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_131 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_132 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_133 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_134 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_135 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_136 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_137 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_138 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_139 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_140 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_141 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_142 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_143 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_144 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_145 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_146 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_147 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_148 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_149 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_150 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_151 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_152 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_153 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_154 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_155 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_156 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_157 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_158 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_159 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_160 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_161 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_162 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_163 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_164 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_165 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_166 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_167 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_168 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_169 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_170 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_171 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_172 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_173 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_174 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_175 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_176 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_177 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_178 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_179 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_180 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_181 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_182 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_183 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_184 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_185 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_186 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_187 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_188 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_189 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_190 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_191 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_192 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_193 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_194 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_195 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_196 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_197 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_198 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_199 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_200 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_201 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_202 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_203 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_204 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_205 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_206 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_207 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_208 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_209 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_210 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_211 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_212 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_213 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_214 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_215 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_216 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_217 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_218 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_219 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_220 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_221 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_222 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_223 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_224 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_225 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_226 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_227 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_228 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_229 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_230 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_231 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_232 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_233 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_234 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_235 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_236 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_237 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_238 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_239 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_240 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_241 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_242 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_243 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_244 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_245 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_246 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_247 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_248 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_249 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_250 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_251 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_252 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_253 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_254 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_255 = 22'h0;
  end
  if (reset) begin
    dec_tlu_way_wb_f = 1'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_0 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_1 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_2 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_3 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_4 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_5 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_6 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_7 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_8 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_9 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_10 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_11 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_12 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_13 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_14 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_15 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_16 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_17 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_18 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_19 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_20 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_21 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_22 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_23 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_24 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_25 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_26 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_27 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_28 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_29 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_30 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_31 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_32 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_33 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_34 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_35 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_36 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_37 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_38 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_39 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_40 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_41 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_42 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_43 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_44 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_45 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_46 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_47 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_48 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_49 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_50 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_51 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_52 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_53 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_54 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_55 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_56 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_57 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_58 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_59 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_60 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_61 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_62 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_63 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_64 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_65 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_66 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_67 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_68 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_69 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_70 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_71 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_72 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_73 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_74 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_75 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_76 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_77 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_78 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_79 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_80 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_81 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_82 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_83 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_84 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_85 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_86 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_87 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_88 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_89 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_90 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_91 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_92 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_93 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_94 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_95 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_96 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_97 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_98 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_99 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_100 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_101 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_102 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_103 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_104 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_105 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_106 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_107 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_108 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_109 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_110 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_111 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_112 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_113 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_114 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_115 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_116 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_117 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_118 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_119 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_120 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_121 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_122 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_123 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_124 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_125 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_126 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_127 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_128 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_129 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_130 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_131 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_132 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_133 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_134 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_135 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_136 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_137 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_138 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_139 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_140 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_141 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_142 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_143 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_144 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_145 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_146 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_147 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_148 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_149 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_150 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_151 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_152 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_153 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_154 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_155 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_156 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_157 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_158 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_159 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_160 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_161 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_162 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_163 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_164 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_165 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_166 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_167 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_168 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_169 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_170 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_171 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_172 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_173 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_174 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_175 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_176 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_177 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_178 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_179 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_180 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_181 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_182 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_183 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_184 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_185 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_186 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_187 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_188 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_189 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_190 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_191 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_192 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_193 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_194 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_195 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_196 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_197 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_198 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_199 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_200 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_201 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_202 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_203 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_204 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_205 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_206 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_207 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_208 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_209 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_210 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_211 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_212 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_213 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_214 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_215 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_216 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_217 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_218 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_219 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_220 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_221 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_222 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_223 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_224 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_225 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_226 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_227 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_228 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_229 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_230 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_231 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_232 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_233 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_234 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_235 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_236 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_237 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_238 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_239 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_240 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_241 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_242 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_243 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_244 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_245 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_246 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_247 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_248 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_249 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_250 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_251 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_252 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_253 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_254 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_255 = 22'h0;
  end
  if (reset) begin
    fghr = 8'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_0 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_1 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_2 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_3 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_4 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_5 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_6 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_7 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_8 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_9 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_10 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_11 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_12 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_13 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_14 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_15 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_16 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_17 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_18 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_19 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_20 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_21 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_22 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_23 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_24 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_25 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_26 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_27 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_28 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_29 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_30 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_31 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_32 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_33 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_34 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_35 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_36 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_37 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_38 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_39 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_40 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_41 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_42 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_43 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_44 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_45 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_46 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_47 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_48 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_49 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_50 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_51 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_52 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_53 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_54 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_55 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_56 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_57 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_58 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_59 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_60 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_61 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_62 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_63 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_64 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_65 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_66 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_67 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_68 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_69 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_70 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_71 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_72 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_73 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_74 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_75 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_76 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_77 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_78 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_79 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_80 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_81 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_82 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_83 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_84 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_85 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_86 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_87 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_88 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_89 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_90 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_91 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_92 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_93 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_94 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_95 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_96 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_97 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_98 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_99 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_100 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_101 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_102 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_103 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_104 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_105 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_106 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_107 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_108 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_109 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_110 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_111 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_112 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_113 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_114 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_115 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_116 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_117 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_118 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_119 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_120 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_121 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_122 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_123 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_124 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_125 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_126 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_127 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_128 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_129 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_130 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_131 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_132 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_133 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_134 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_135 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_136 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_137 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_138 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_139 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_140 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_141 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_142 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_143 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_144 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_145 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_146 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_147 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_148 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_149 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_150 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_151 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_152 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_153 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_154 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_155 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_156 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_157 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_158 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_159 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_160 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_161 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_162 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_163 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_164 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_165 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_166 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_167 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_168 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_169 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_170 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_171 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_172 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_173 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_174 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_175 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_176 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_177 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_178 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_179 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_180 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_181 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_182 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_183 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_184 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_185 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_186 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_187 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_188 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_189 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_190 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_191 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_192 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_193 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_194 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_195 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_196 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_197 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_198 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_199 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_200 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_201 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_202 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_203 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_204 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_205 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_206 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_207 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_208 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_209 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_210 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_211 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_212 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_213 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_214 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_215 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_216 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_217 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_218 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_219 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_220 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_221 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_222 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_223 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_224 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_225 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_226 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_227 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_228 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_229 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_230 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_231 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_232 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_233 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_234 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_235 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_236 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_237 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_238 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_239 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_240 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_241 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_242 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_243 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_244 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_245 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_246 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_247 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_248 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_249 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_250 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_251 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_252 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_253 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_254 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_255 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_0 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_1 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_2 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_3 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_4 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_5 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_6 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_7 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_8 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_9 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_10 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_11 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_12 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_13 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_14 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_15 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_16 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_17 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_18 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_19 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_20 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_21 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_22 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_23 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_24 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_25 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_26 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_27 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_28 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_29 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_30 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_31 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_32 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_33 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_34 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_35 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_36 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_37 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_38 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_39 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_40 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_41 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_42 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_43 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_44 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_45 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_46 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_47 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_48 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_49 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_50 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_51 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_52 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_53 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_54 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_55 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_56 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_57 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_58 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_59 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_60 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_61 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_62 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_63 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_64 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_65 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_66 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_67 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_68 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_69 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_70 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_71 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_72 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_73 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_74 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_75 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_76 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_77 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_78 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_79 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_80 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_81 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_82 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_83 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_84 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_85 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_86 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_87 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_88 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_89 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_90 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_91 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_92 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_93 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_94 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_95 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_96 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_97 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_98 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_99 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_100 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_101 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_102 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_103 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_104 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_105 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_106 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_107 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_108 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_109 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_110 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_111 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_112 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_113 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_114 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_115 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_116 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_117 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_118 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_119 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_120 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_121 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_122 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_123 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_124 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_125 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_126 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_127 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_128 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_129 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_130 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_131 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_132 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_133 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_134 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_135 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_136 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_137 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_138 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_139 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_140 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_141 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_142 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_143 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_144 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_145 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_146 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_147 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_148 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_149 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_150 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_151 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_152 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_153 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_154 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_155 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_156 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_157 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_158 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_159 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_160 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_161 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_162 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_163 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_164 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_165 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_166 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_167 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_168 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_169 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_170 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_171 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_172 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_173 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_174 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_175 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_176 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_177 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_178 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_179 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_180 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_181 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_182 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_183 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_184 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_185 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_186 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_187 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_188 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_189 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_190 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_191 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_192 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_193 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_194 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_195 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_196 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_197 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_198 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_199 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_200 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_201 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_202 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_203 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_204 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_205 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_206 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_207 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_208 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_209 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_210 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_211 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_212 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_213 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_214 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_215 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_216 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_217 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_218 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_219 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_220 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_221 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_222 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_223 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_224 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_225 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_226 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_227 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_228 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_229 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_230 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_231 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_232 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_233 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_234 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_235 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_236 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_237 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_238 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_239 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_240 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_241 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_242 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_243 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_244 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_245 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_246 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_247 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_248 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_249 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_250 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_251 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_252 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_253 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_254 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_255 = 2'h0;
  end
  if (reset) begin
    exu_mp_way_f = 1'h0;
  end
  if (reset) begin
    exu_flush_final_d1 = 1'h0;
  end
  if (reset) begin
    btb_lru_b0_f = 256'h0;
  end
  if (reset) begin
    ifc_fetch_adder_prior = 30'h0;
  end
  if (reset) begin
    rets_out_0 = 32'h0;
  end
  if (reset) begin
    rets_out_1 = 32'h0;
  end
  if (reset) begin
    rets_out_2 = 32'h0;
  end
  if (reset) begin
    rets_out_3 = 32'h0;
  end
  if (reset) begin
    rets_out_4 = 32'h0;
  end
  if (reset) begin
    rets_out_5 = 32'h0;
  end
  if (reset) begin
    rets_out_6 = 32'h0;
  end
  if (reset) begin
    rets_out_7 = 32'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      leak_one_f_d1 <= 1'h0;
    end else begin
      leak_one_f_d1 <= _T_40 | _T_42;
    end
  end
  always @(posedge rvclkhdr_10_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_0 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_0 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_11_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_1 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_1 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_12_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_2 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_2 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_13_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_3 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_3 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_14_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_4 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_4 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_15_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_5 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_5 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_16_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_6 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_6 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_17_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_7 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_7 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_18_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_8 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_8 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_19_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_9 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_9 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_20_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_10 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_10 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_21_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_11 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_11 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_22_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_12 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_12 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_23_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_13 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_13 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_24_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_14 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_14 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_25_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_15 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_15 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_26_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_16 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_16 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_27_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_17 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_17 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_28_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_18 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_18 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_29_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_19 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_19 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_30_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_20 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_20 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_31_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_21 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_21 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_32_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_22 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_22 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_33_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_23 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_23 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_34_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_24 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_24 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_35_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_25 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_25 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_36_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_26 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_26 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_37_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_27 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_27 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_38_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_28 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_28 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_39_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_29 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_29 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_40_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_30 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_30 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_41_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_31 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_31 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_42_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_32 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_32 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_43_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_33 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_33 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_44_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_34 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_34 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_45_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_35 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_35 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_46_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_36 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_36 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_47_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_37 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_37 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_48_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_38 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_38 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_49_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_39 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_39 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_50_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_40 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_40 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_51_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_41 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_41 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_52_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_42 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_42 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_53_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_43 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_43 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_54_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_44 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_44 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_55_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_45 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_45 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_56_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_46 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_46 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_57_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_47 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_47 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_58_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_48 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_48 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_59_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_49 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_49 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_60_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_50 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_50 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_61_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_51 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_51 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_62_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_52 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_52 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_63_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_53 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_53 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_64_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_54 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_54 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_65_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_55 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_55 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_66_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_56 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_56 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_67_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_57 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_57 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_68_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_58 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_58 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_69_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_59 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_59 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_70_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_60 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_60 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_71_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_61 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_61 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_72_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_62 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_62 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_73_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_63 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_63 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_74_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_64 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_64 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_75_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_65 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_65 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_76_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_66 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_66 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_77_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_67 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_67 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_78_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_68 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_68 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_79_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_69 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_69 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_80_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_70 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_70 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_81_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_71 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_71 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_82_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_72 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_72 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_83_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_73 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_73 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_84_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_74 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_74 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_85_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_75 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_75 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_76 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_76 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_77 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_77 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_78 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_78 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_79 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_79 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_80 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_80 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_81 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_81 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_82 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_82 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_83 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_83 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_94_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_84 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_84 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_95_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_85 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_85 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_96_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_86 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_86 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_97_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_87 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_87 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_98_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_88 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_88 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_99_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_89 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_89 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_100_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_90 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_90 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_101_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_91 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_91 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_102_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_92 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_92 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_103_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_93 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_93 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_104_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_94 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_94 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_105_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_95 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_95 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_106_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_96 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_96 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_107_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_97 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_97 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_108_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_98 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_98 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_109_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_99 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_99 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_110_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_100 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_100 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_111_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_101 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_101 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_112_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_102 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_102 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_113_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_103 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_103 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_114_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_104 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_104 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_115_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_105 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_105 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_116_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_106 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_106 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_117_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_107 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_107 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_118_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_108 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_108 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_119_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_109 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_109 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_120_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_110 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_110 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_121_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_111 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_111 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_122_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_112 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_112 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_123_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_113 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_113 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_124_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_114 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_114 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_125_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_115 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_115 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_126_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_116 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_116 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_127_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_117 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_117 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_128_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_118 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_118 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_129_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_119 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_119 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_130_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_120 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_120 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_131_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_121 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_121 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_132_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_122 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_122 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_133_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_123 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_123 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_134_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_124 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_124 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_135_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_125 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_125 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_136_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_126 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_126 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_137_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_127 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_127 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_138_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_128 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_128 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_139_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_129 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_129 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_140_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_130 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_130 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_141_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_131 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_131 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_142_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_132 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_132 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_143_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_133 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_133 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_144_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_134 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_134 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_145_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_135 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_135 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_146_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_136 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_136 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_147_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_137 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_137 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_148_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_138 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_138 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_149_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_139 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_139 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_150_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_140 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_140 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_151_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_141 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_141 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_152_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_142 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_142 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_153_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_143 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_143 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_154_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_144 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_144 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_155_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_145 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_145 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_156_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_146 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_146 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_157_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_147 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_147 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_158_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_148 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_148 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_159_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_149 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_149 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_160_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_150 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_150 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_161_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_151 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_151 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_162_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_152 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_152 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_163_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_153 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_153 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_164_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_154 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_154 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_165_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_155 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_155 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_166_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_156 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_156 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_167_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_157 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_157 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_168_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_158 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_158 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_169_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_159 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_159 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_170_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_160 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_160 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_171_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_161 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_161 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_172_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_162 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_162 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_173_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_163 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_163 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_174_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_164 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_164 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_175_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_165 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_165 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_176_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_166 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_166 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_177_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_167 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_167 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_178_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_168 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_168 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_179_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_169 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_169 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_180_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_170 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_170 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_181_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_171 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_171 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_182_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_172 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_172 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_183_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_173 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_173 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_184_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_174 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_174 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_185_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_175 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_175 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_186_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_176 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_176 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_187_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_177 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_177 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_188_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_178 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_178 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_189_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_179 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_179 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_190_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_180 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_180 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_191_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_181 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_181 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_192_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_182 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_182 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_193_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_183 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_183 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_194_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_184 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_184 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_195_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_185 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_185 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_196_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_186 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_186 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_197_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_187 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_187 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_198_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_188 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_188 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_199_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_189 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_189 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_200_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_190 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_190 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_201_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_191 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_191 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_202_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_192 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_192 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_203_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_193 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_193 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_204_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_194 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_194 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_205_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_195 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_195 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_206_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_196 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_196 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_207_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_197 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_197 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_208_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_198 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_198 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_209_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_199 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_199 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_210_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_200 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_200 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_211_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_201 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_201 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_212_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_202 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_202 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_213_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_203 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_203 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_214_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_204 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_204 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_215_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_205 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_205 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_216_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_206 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_206 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_217_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_207 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_207 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_218_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_208 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_208 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_219_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_209 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_209 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_220_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_210 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_210 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_221_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_211 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_211 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_222_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_212 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_212 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_223_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_213 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_213 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_224_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_214 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_214 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_225_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_215 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_215 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_226_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_216 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_216 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_227_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_217 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_217 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_228_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_218 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_218 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_229_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_219 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_219 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_230_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_220 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_220 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_231_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_221 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_221 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_232_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_222 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_222 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_233_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_223 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_223 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_234_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_224 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_224 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_235_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_225 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_225 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_236_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_226 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_226 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_237_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_227 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_227 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_238_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_228 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_228 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_239_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_229 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_229 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_240_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_230 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_230 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_241_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_231 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_231 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_242_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_232 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_232 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_243_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_233 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_233 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_244_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_234 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_234 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_245_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_235 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_235 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_246_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_236 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_236 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_247_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_237 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_237 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_248_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_238 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_238 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_249_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_239 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_239 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_250_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_240 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_240 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_251_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_241 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_241 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_252_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_242 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_242 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_253_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_243 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_243 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_254_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_244 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_244 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_255_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_245 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_245 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_256_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_246 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_246 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_257_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_247 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_247 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_258_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_248 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_248 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_259_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_249 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_249 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_260_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_250 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_250 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_261_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_251 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_251 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_262_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_252 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_252 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_263_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_253 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_253 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_264_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_254 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_254 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_265_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_255 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way0_out_255 <= {_T_538,_T_535};
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      dec_tlu_way_wb_f <= 1'h0;
    end else begin
      dec_tlu_way_wb_f <= io_dec_bp_dec_tlu_br0_r_pkt_bits_way;
    end
  end
  always @(posedge rvclkhdr_266_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_0 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_0 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_267_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_1 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_1 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_268_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_2 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_2 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_269_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_3 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_3 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_270_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_4 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_4 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_271_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_5 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_5 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_272_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_6 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_6 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_273_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_7 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_7 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_274_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_8 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_8 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_275_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_9 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_9 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_276_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_10 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_10 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_277_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_11 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_11 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_278_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_12 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_12 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_279_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_13 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_13 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_280_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_14 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_14 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_281_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_15 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_15 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_282_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_16 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_16 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_283_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_17 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_17 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_284_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_18 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_18 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_285_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_19 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_19 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_286_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_20 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_20 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_287_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_21 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_21 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_288_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_22 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_22 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_289_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_23 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_23 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_290_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_24 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_24 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_291_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_25 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_25 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_292_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_26 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_26 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_293_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_27 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_27 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_294_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_28 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_28 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_295_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_29 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_29 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_296_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_30 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_30 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_297_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_31 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_31 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_298_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_32 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_32 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_299_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_33 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_33 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_300_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_34 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_34 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_301_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_35 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_35 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_302_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_36 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_36 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_303_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_37 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_37 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_304_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_38 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_38 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_305_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_39 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_39 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_306_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_40 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_40 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_307_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_41 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_41 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_308_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_42 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_42 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_309_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_43 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_43 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_310_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_44 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_44 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_311_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_45 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_45 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_312_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_46 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_46 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_313_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_47 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_47 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_314_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_48 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_48 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_315_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_49 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_49 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_316_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_50 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_50 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_317_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_51 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_51 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_318_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_52 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_52 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_319_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_53 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_53 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_320_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_54 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_54 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_321_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_55 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_55 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_322_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_56 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_56 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_323_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_57 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_57 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_324_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_58 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_58 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_325_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_59 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_59 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_326_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_60 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_60 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_327_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_61 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_61 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_328_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_62 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_62 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_329_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_63 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_63 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_330_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_64 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_64 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_331_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_65 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_65 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_332_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_66 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_66 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_333_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_67 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_67 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_334_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_68 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_68 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_335_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_69 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_69 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_336_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_70 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_70 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_337_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_71 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_71 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_338_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_72 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_72 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_339_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_73 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_73 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_340_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_74 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_74 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_341_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_75 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_75 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_342_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_76 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_76 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_343_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_77 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_77 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_344_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_78 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_78 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_345_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_79 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_79 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_346_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_80 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_80 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_347_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_81 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_81 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_348_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_82 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_82 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_349_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_83 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_83 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_350_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_84 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_84 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_351_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_85 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_85 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_352_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_86 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_86 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_353_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_87 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_87 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_354_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_88 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_88 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_355_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_89 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_89 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_356_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_90 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_90 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_357_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_91 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_91 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_358_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_92 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_92 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_359_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_93 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_93 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_360_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_94 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_94 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_361_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_95 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_95 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_362_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_96 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_96 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_363_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_97 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_97 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_364_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_98 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_98 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_365_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_99 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_99 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_366_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_100 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_100 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_367_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_101 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_101 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_368_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_102 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_102 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_369_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_103 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_103 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_370_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_104 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_104 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_371_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_105 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_105 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_372_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_106 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_106 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_373_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_107 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_107 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_374_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_108 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_108 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_375_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_109 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_109 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_376_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_110 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_110 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_377_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_111 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_111 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_378_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_112 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_112 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_379_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_113 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_113 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_380_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_114 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_114 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_381_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_115 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_115 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_382_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_116 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_116 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_383_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_117 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_117 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_384_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_118 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_118 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_385_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_119 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_119 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_386_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_120 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_120 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_387_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_121 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_121 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_388_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_122 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_122 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_389_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_123 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_123 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_390_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_124 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_124 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_391_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_125 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_125 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_392_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_126 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_126 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_393_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_127 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_127 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_394_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_128 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_128 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_395_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_129 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_129 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_396_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_130 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_130 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_397_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_131 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_131 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_398_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_132 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_132 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_399_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_133 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_133 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_400_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_134 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_134 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_401_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_135 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_135 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_402_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_136 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_136 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_403_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_137 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_137 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_404_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_138 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_138 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_405_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_139 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_139 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_406_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_140 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_140 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_407_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_141 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_141 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_408_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_142 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_142 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_409_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_143 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_143 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_410_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_144 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_144 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_411_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_145 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_145 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_412_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_146 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_146 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_413_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_147 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_147 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_414_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_148 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_148 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_415_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_149 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_149 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_416_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_150 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_150 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_417_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_151 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_151 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_418_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_152 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_152 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_419_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_153 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_153 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_420_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_154 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_154 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_421_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_155 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_155 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_422_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_156 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_156 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_423_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_157 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_157 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_424_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_158 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_158 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_425_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_159 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_159 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_426_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_160 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_160 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_427_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_161 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_161 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_428_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_162 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_162 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_429_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_163 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_163 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_430_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_164 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_164 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_431_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_165 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_165 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_432_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_166 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_166 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_433_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_167 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_167 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_434_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_168 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_168 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_435_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_169 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_169 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_436_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_170 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_170 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_437_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_171 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_171 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_438_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_172 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_172 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_439_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_173 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_173 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_440_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_174 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_174 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_441_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_175 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_175 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_442_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_176 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_176 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_443_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_177 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_177 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_444_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_178 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_178 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_445_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_179 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_179 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_446_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_180 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_180 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_447_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_181 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_181 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_448_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_182 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_182 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_449_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_183 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_183 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_450_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_184 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_184 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_451_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_185 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_185 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_452_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_186 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_186 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_453_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_187 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_187 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_454_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_188 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_188 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_455_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_189 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_189 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_456_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_190 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_190 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_457_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_191 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_191 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_458_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_192 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_192 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_459_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_193 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_193 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_460_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_194 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_194 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_461_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_195 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_195 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_462_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_196 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_196 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_463_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_197 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_197 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_464_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_198 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_198 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_465_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_199 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_199 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_466_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_200 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_200 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_467_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_201 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_201 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_468_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_202 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_202 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_469_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_203 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_203 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_470_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_204 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_204 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_471_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_205 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_205 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_472_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_206 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_206 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_473_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_207 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_207 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_474_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_208 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_208 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_475_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_209 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_209 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_476_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_210 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_210 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_477_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_211 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_211 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_478_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_212 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_212 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_479_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_213 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_213 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_480_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_214 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_214 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_481_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_215 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_215 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_482_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_216 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_216 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_483_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_217 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_217 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_484_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_218 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_218 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_485_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_219 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_219 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_486_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_220 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_220 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_487_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_221 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_221 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_488_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_222 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_222 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_489_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_223 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_223 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_490_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_224 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_224 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_491_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_225 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_225 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_492_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_226 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_226 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_493_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_227 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_227 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_494_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_228 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_228 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_495_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_229 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_229 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_496_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_230 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_230 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_497_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_231 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_231 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_498_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_232 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_232 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_499_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_233 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_233 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_500_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_234 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_234 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_501_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_235 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_235 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_502_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_236 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_236 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_503_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_237 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_237 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_504_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_238 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_238 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_505_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_239 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_239 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_506_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_240 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_240 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_507_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_241 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_241 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_508_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_242 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_242 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_509_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_243 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_243 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_510_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_244 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_244 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_511_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_245 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_245 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_512_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_246 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_246 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_513_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_247 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_247 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_514_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_248 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_248 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_515_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_249 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_249 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_516_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_250 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_250 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_517_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_251 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_251 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_518_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_252 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_252 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_519_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_253 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_253 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_520_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_254 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_254 <= {_T_538,_T_535};
    end
  end
  always @(posedge rvclkhdr_521_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_255 <= 22'h0;
    end else begin
      btb_bank0_rd_data_way1_out_255 <= {_T_538,_T_535};
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      fghr <= 8'h0;
    end else begin
      fghr <= _T_339 | _T_338;
    end
  end
  always @(posedge rvclkhdr_538_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_0 <= 2'h0;
    end else if (bht_bank_sel_1_0_0) begin
      if (_T_8870) begin
        bht_bank_rd_data_out_1_0 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_0 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_538_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_1 <= 2'h0;
    end else if (bht_bank_sel_1_0_1) begin
      if (_T_8879) begin
        bht_bank_rd_data_out_1_1 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_1 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_538_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_2 <= 2'h0;
    end else if (bht_bank_sel_1_0_2) begin
      if (_T_8888) begin
        bht_bank_rd_data_out_1_2 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_2 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_538_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_3 <= 2'h0;
    end else if (bht_bank_sel_1_0_3) begin
      if (_T_8897) begin
        bht_bank_rd_data_out_1_3 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_3 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_538_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_4 <= 2'h0;
    end else if (bht_bank_sel_1_0_4) begin
      if (_T_8906) begin
        bht_bank_rd_data_out_1_4 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_4 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_538_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_5 <= 2'h0;
    end else if (bht_bank_sel_1_0_5) begin
      if (_T_8915) begin
        bht_bank_rd_data_out_1_5 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_5 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_538_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_6 <= 2'h0;
    end else if (bht_bank_sel_1_0_6) begin
      if (_T_8924) begin
        bht_bank_rd_data_out_1_6 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_6 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_538_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_7 <= 2'h0;
    end else if (bht_bank_sel_1_0_7) begin
      if (_T_8933) begin
        bht_bank_rd_data_out_1_7 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_7 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_538_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_8 <= 2'h0;
    end else if (bht_bank_sel_1_0_8) begin
      if (_T_8942) begin
        bht_bank_rd_data_out_1_8 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_8 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_538_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_9 <= 2'h0;
    end else if (bht_bank_sel_1_0_9) begin
      if (_T_8951) begin
        bht_bank_rd_data_out_1_9 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_9 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_538_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_10 <= 2'h0;
    end else if (bht_bank_sel_1_0_10) begin
      if (_T_8960) begin
        bht_bank_rd_data_out_1_10 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_10 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_538_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_11 <= 2'h0;
    end else if (bht_bank_sel_1_0_11) begin
      if (_T_8969) begin
        bht_bank_rd_data_out_1_11 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_11 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_538_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_12 <= 2'h0;
    end else if (bht_bank_sel_1_0_12) begin
      if (_T_8978) begin
        bht_bank_rd_data_out_1_12 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_12 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_538_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_13 <= 2'h0;
    end else if (bht_bank_sel_1_0_13) begin
      if (_T_8987) begin
        bht_bank_rd_data_out_1_13 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_13 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_538_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_14 <= 2'h0;
    end else if (bht_bank_sel_1_0_14) begin
      if (_T_8996) begin
        bht_bank_rd_data_out_1_14 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_14 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_538_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_15 <= 2'h0;
    end else if (bht_bank_sel_1_0_15) begin
      if (_T_9005) begin
        bht_bank_rd_data_out_1_15 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_15 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_539_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_16 <= 2'h0;
    end else if (bht_bank_sel_1_1_0) begin
      if (_T_9014) begin
        bht_bank_rd_data_out_1_16 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_16 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_539_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_17 <= 2'h0;
    end else if (bht_bank_sel_1_1_1) begin
      if (_T_9023) begin
        bht_bank_rd_data_out_1_17 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_17 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_539_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_18 <= 2'h0;
    end else if (bht_bank_sel_1_1_2) begin
      if (_T_9032) begin
        bht_bank_rd_data_out_1_18 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_18 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_539_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_19 <= 2'h0;
    end else if (bht_bank_sel_1_1_3) begin
      if (_T_9041) begin
        bht_bank_rd_data_out_1_19 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_19 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_539_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_20 <= 2'h0;
    end else if (bht_bank_sel_1_1_4) begin
      if (_T_9050) begin
        bht_bank_rd_data_out_1_20 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_20 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_539_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_21 <= 2'h0;
    end else if (bht_bank_sel_1_1_5) begin
      if (_T_9059) begin
        bht_bank_rd_data_out_1_21 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_21 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_539_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_22 <= 2'h0;
    end else if (bht_bank_sel_1_1_6) begin
      if (_T_9068) begin
        bht_bank_rd_data_out_1_22 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_22 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_539_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_23 <= 2'h0;
    end else if (bht_bank_sel_1_1_7) begin
      if (_T_9077) begin
        bht_bank_rd_data_out_1_23 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_23 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_539_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_24 <= 2'h0;
    end else if (bht_bank_sel_1_1_8) begin
      if (_T_9086) begin
        bht_bank_rd_data_out_1_24 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_24 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_539_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_25 <= 2'h0;
    end else if (bht_bank_sel_1_1_9) begin
      if (_T_9095) begin
        bht_bank_rd_data_out_1_25 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_25 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_539_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_26 <= 2'h0;
    end else if (bht_bank_sel_1_1_10) begin
      if (_T_9104) begin
        bht_bank_rd_data_out_1_26 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_26 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_539_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_27 <= 2'h0;
    end else if (bht_bank_sel_1_1_11) begin
      if (_T_9113) begin
        bht_bank_rd_data_out_1_27 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_27 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_539_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_28 <= 2'h0;
    end else if (bht_bank_sel_1_1_12) begin
      if (_T_9122) begin
        bht_bank_rd_data_out_1_28 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_28 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_539_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_29 <= 2'h0;
    end else if (bht_bank_sel_1_1_13) begin
      if (_T_9131) begin
        bht_bank_rd_data_out_1_29 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_29 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_539_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_30 <= 2'h0;
    end else if (bht_bank_sel_1_1_14) begin
      if (_T_9140) begin
        bht_bank_rd_data_out_1_30 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_30 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_539_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_31 <= 2'h0;
    end else if (bht_bank_sel_1_1_15) begin
      if (_T_9149) begin
        bht_bank_rd_data_out_1_31 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_31 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_540_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_32 <= 2'h0;
    end else if (bht_bank_sel_1_2_0) begin
      if (_T_9158) begin
        bht_bank_rd_data_out_1_32 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_32 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_540_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_33 <= 2'h0;
    end else if (bht_bank_sel_1_2_1) begin
      if (_T_9167) begin
        bht_bank_rd_data_out_1_33 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_33 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_540_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_34 <= 2'h0;
    end else if (bht_bank_sel_1_2_2) begin
      if (_T_9176) begin
        bht_bank_rd_data_out_1_34 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_34 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_540_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_35 <= 2'h0;
    end else if (bht_bank_sel_1_2_3) begin
      if (_T_9185) begin
        bht_bank_rd_data_out_1_35 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_35 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_540_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_36 <= 2'h0;
    end else if (bht_bank_sel_1_2_4) begin
      if (_T_9194) begin
        bht_bank_rd_data_out_1_36 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_36 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_540_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_37 <= 2'h0;
    end else if (bht_bank_sel_1_2_5) begin
      if (_T_9203) begin
        bht_bank_rd_data_out_1_37 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_37 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_540_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_38 <= 2'h0;
    end else if (bht_bank_sel_1_2_6) begin
      if (_T_9212) begin
        bht_bank_rd_data_out_1_38 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_38 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_540_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_39 <= 2'h0;
    end else if (bht_bank_sel_1_2_7) begin
      if (_T_9221) begin
        bht_bank_rd_data_out_1_39 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_39 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_540_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_40 <= 2'h0;
    end else if (bht_bank_sel_1_2_8) begin
      if (_T_9230) begin
        bht_bank_rd_data_out_1_40 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_40 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_540_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_41 <= 2'h0;
    end else if (bht_bank_sel_1_2_9) begin
      if (_T_9239) begin
        bht_bank_rd_data_out_1_41 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_41 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_540_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_42 <= 2'h0;
    end else if (bht_bank_sel_1_2_10) begin
      if (_T_9248) begin
        bht_bank_rd_data_out_1_42 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_42 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_540_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_43 <= 2'h0;
    end else if (bht_bank_sel_1_2_11) begin
      if (_T_9257) begin
        bht_bank_rd_data_out_1_43 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_43 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_540_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_44 <= 2'h0;
    end else if (bht_bank_sel_1_2_12) begin
      if (_T_9266) begin
        bht_bank_rd_data_out_1_44 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_44 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_540_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_45 <= 2'h0;
    end else if (bht_bank_sel_1_2_13) begin
      if (_T_9275) begin
        bht_bank_rd_data_out_1_45 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_45 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_540_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_46 <= 2'h0;
    end else if (bht_bank_sel_1_2_14) begin
      if (_T_9284) begin
        bht_bank_rd_data_out_1_46 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_46 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_540_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_47 <= 2'h0;
    end else if (bht_bank_sel_1_2_15) begin
      if (_T_9293) begin
        bht_bank_rd_data_out_1_47 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_47 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_541_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_48 <= 2'h0;
    end else if (bht_bank_sel_1_3_0) begin
      if (_T_9302) begin
        bht_bank_rd_data_out_1_48 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_48 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_541_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_49 <= 2'h0;
    end else if (bht_bank_sel_1_3_1) begin
      if (_T_9311) begin
        bht_bank_rd_data_out_1_49 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_49 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_541_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_50 <= 2'h0;
    end else if (bht_bank_sel_1_3_2) begin
      if (_T_9320) begin
        bht_bank_rd_data_out_1_50 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_50 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_541_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_51 <= 2'h0;
    end else if (bht_bank_sel_1_3_3) begin
      if (_T_9329) begin
        bht_bank_rd_data_out_1_51 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_51 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_541_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_52 <= 2'h0;
    end else if (bht_bank_sel_1_3_4) begin
      if (_T_9338) begin
        bht_bank_rd_data_out_1_52 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_52 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_541_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_53 <= 2'h0;
    end else if (bht_bank_sel_1_3_5) begin
      if (_T_9347) begin
        bht_bank_rd_data_out_1_53 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_53 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_541_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_54 <= 2'h0;
    end else if (bht_bank_sel_1_3_6) begin
      if (_T_9356) begin
        bht_bank_rd_data_out_1_54 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_54 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_541_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_55 <= 2'h0;
    end else if (bht_bank_sel_1_3_7) begin
      if (_T_9365) begin
        bht_bank_rd_data_out_1_55 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_55 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_541_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_56 <= 2'h0;
    end else if (bht_bank_sel_1_3_8) begin
      if (_T_9374) begin
        bht_bank_rd_data_out_1_56 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_56 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_541_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_57 <= 2'h0;
    end else if (bht_bank_sel_1_3_9) begin
      if (_T_9383) begin
        bht_bank_rd_data_out_1_57 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_57 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_541_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_58 <= 2'h0;
    end else if (bht_bank_sel_1_3_10) begin
      if (_T_9392) begin
        bht_bank_rd_data_out_1_58 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_58 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_541_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_59 <= 2'h0;
    end else if (bht_bank_sel_1_3_11) begin
      if (_T_9401) begin
        bht_bank_rd_data_out_1_59 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_59 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_541_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_60 <= 2'h0;
    end else if (bht_bank_sel_1_3_12) begin
      if (_T_9410) begin
        bht_bank_rd_data_out_1_60 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_60 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_541_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_61 <= 2'h0;
    end else if (bht_bank_sel_1_3_13) begin
      if (_T_9419) begin
        bht_bank_rd_data_out_1_61 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_61 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_541_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_62 <= 2'h0;
    end else if (bht_bank_sel_1_3_14) begin
      if (_T_9428) begin
        bht_bank_rd_data_out_1_62 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_62 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_541_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_63 <= 2'h0;
    end else if (bht_bank_sel_1_3_15) begin
      if (_T_9437) begin
        bht_bank_rd_data_out_1_63 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_63 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_542_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_64 <= 2'h0;
    end else if (bht_bank_sel_1_4_0) begin
      if (_T_9446) begin
        bht_bank_rd_data_out_1_64 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_64 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_542_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_65 <= 2'h0;
    end else if (bht_bank_sel_1_4_1) begin
      if (_T_9455) begin
        bht_bank_rd_data_out_1_65 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_65 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_542_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_66 <= 2'h0;
    end else if (bht_bank_sel_1_4_2) begin
      if (_T_9464) begin
        bht_bank_rd_data_out_1_66 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_66 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_542_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_67 <= 2'h0;
    end else if (bht_bank_sel_1_4_3) begin
      if (_T_9473) begin
        bht_bank_rd_data_out_1_67 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_67 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_542_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_68 <= 2'h0;
    end else if (bht_bank_sel_1_4_4) begin
      if (_T_9482) begin
        bht_bank_rd_data_out_1_68 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_68 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_542_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_69 <= 2'h0;
    end else if (bht_bank_sel_1_4_5) begin
      if (_T_9491) begin
        bht_bank_rd_data_out_1_69 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_69 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_542_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_70 <= 2'h0;
    end else if (bht_bank_sel_1_4_6) begin
      if (_T_9500) begin
        bht_bank_rd_data_out_1_70 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_70 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_542_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_71 <= 2'h0;
    end else if (bht_bank_sel_1_4_7) begin
      if (_T_9509) begin
        bht_bank_rd_data_out_1_71 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_71 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_542_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_72 <= 2'h0;
    end else if (bht_bank_sel_1_4_8) begin
      if (_T_9518) begin
        bht_bank_rd_data_out_1_72 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_72 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_542_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_73 <= 2'h0;
    end else if (bht_bank_sel_1_4_9) begin
      if (_T_9527) begin
        bht_bank_rd_data_out_1_73 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_73 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_542_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_74 <= 2'h0;
    end else if (bht_bank_sel_1_4_10) begin
      if (_T_9536) begin
        bht_bank_rd_data_out_1_74 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_74 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_542_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_75 <= 2'h0;
    end else if (bht_bank_sel_1_4_11) begin
      if (_T_9545) begin
        bht_bank_rd_data_out_1_75 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_75 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_542_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_76 <= 2'h0;
    end else if (bht_bank_sel_1_4_12) begin
      if (_T_9554) begin
        bht_bank_rd_data_out_1_76 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_76 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_542_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_77 <= 2'h0;
    end else if (bht_bank_sel_1_4_13) begin
      if (_T_9563) begin
        bht_bank_rd_data_out_1_77 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_77 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_542_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_78 <= 2'h0;
    end else if (bht_bank_sel_1_4_14) begin
      if (_T_9572) begin
        bht_bank_rd_data_out_1_78 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_78 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_542_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_79 <= 2'h0;
    end else if (bht_bank_sel_1_4_15) begin
      if (_T_9581) begin
        bht_bank_rd_data_out_1_79 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_79 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_543_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_80 <= 2'h0;
    end else if (bht_bank_sel_1_5_0) begin
      if (_T_9590) begin
        bht_bank_rd_data_out_1_80 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_80 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_543_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_81 <= 2'h0;
    end else if (bht_bank_sel_1_5_1) begin
      if (_T_9599) begin
        bht_bank_rd_data_out_1_81 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_81 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_543_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_82 <= 2'h0;
    end else if (bht_bank_sel_1_5_2) begin
      if (_T_9608) begin
        bht_bank_rd_data_out_1_82 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_82 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_543_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_83 <= 2'h0;
    end else if (bht_bank_sel_1_5_3) begin
      if (_T_9617) begin
        bht_bank_rd_data_out_1_83 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_83 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_543_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_84 <= 2'h0;
    end else if (bht_bank_sel_1_5_4) begin
      if (_T_9626) begin
        bht_bank_rd_data_out_1_84 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_84 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_543_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_85 <= 2'h0;
    end else if (bht_bank_sel_1_5_5) begin
      if (_T_9635) begin
        bht_bank_rd_data_out_1_85 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_85 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_543_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_86 <= 2'h0;
    end else if (bht_bank_sel_1_5_6) begin
      if (_T_9644) begin
        bht_bank_rd_data_out_1_86 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_86 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_543_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_87 <= 2'h0;
    end else if (bht_bank_sel_1_5_7) begin
      if (_T_9653) begin
        bht_bank_rd_data_out_1_87 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_87 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_543_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_88 <= 2'h0;
    end else if (bht_bank_sel_1_5_8) begin
      if (_T_9662) begin
        bht_bank_rd_data_out_1_88 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_88 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_543_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_89 <= 2'h0;
    end else if (bht_bank_sel_1_5_9) begin
      if (_T_9671) begin
        bht_bank_rd_data_out_1_89 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_89 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_543_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_90 <= 2'h0;
    end else if (bht_bank_sel_1_5_10) begin
      if (_T_9680) begin
        bht_bank_rd_data_out_1_90 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_90 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_543_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_91 <= 2'h0;
    end else if (bht_bank_sel_1_5_11) begin
      if (_T_9689) begin
        bht_bank_rd_data_out_1_91 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_91 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_543_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_92 <= 2'h0;
    end else if (bht_bank_sel_1_5_12) begin
      if (_T_9698) begin
        bht_bank_rd_data_out_1_92 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_92 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_543_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_93 <= 2'h0;
    end else if (bht_bank_sel_1_5_13) begin
      if (_T_9707) begin
        bht_bank_rd_data_out_1_93 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_93 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_543_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_94 <= 2'h0;
    end else if (bht_bank_sel_1_5_14) begin
      if (_T_9716) begin
        bht_bank_rd_data_out_1_94 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_94 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_543_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_95 <= 2'h0;
    end else if (bht_bank_sel_1_5_15) begin
      if (_T_9725) begin
        bht_bank_rd_data_out_1_95 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_95 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_544_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_96 <= 2'h0;
    end else if (bht_bank_sel_1_6_0) begin
      if (_T_9734) begin
        bht_bank_rd_data_out_1_96 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_96 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_544_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_97 <= 2'h0;
    end else if (bht_bank_sel_1_6_1) begin
      if (_T_9743) begin
        bht_bank_rd_data_out_1_97 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_97 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_544_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_98 <= 2'h0;
    end else if (bht_bank_sel_1_6_2) begin
      if (_T_9752) begin
        bht_bank_rd_data_out_1_98 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_98 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_544_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_99 <= 2'h0;
    end else if (bht_bank_sel_1_6_3) begin
      if (_T_9761) begin
        bht_bank_rd_data_out_1_99 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_99 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_544_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_100 <= 2'h0;
    end else if (bht_bank_sel_1_6_4) begin
      if (_T_9770) begin
        bht_bank_rd_data_out_1_100 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_100 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_544_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_101 <= 2'h0;
    end else if (bht_bank_sel_1_6_5) begin
      if (_T_9779) begin
        bht_bank_rd_data_out_1_101 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_101 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_544_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_102 <= 2'h0;
    end else if (bht_bank_sel_1_6_6) begin
      if (_T_9788) begin
        bht_bank_rd_data_out_1_102 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_102 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_544_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_103 <= 2'h0;
    end else if (bht_bank_sel_1_6_7) begin
      if (_T_9797) begin
        bht_bank_rd_data_out_1_103 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_103 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_544_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_104 <= 2'h0;
    end else if (bht_bank_sel_1_6_8) begin
      if (_T_9806) begin
        bht_bank_rd_data_out_1_104 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_104 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_544_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_105 <= 2'h0;
    end else if (bht_bank_sel_1_6_9) begin
      if (_T_9815) begin
        bht_bank_rd_data_out_1_105 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_105 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_544_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_106 <= 2'h0;
    end else if (bht_bank_sel_1_6_10) begin
      if (_T_9824) begin
        bht_bank_rd_data_out_1_106 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_106 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_544_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_107 <= 2'h0;
    end else if (bht_bank_sel_1_6_11) begin
      if (_T_9833) begin
        bht_bank_rd_data_out_1_107 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_107 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_544_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_108 <= 2'h0;
    end else if (bht_bank_sel_1_6_12) begin
      if (_T_9842) begin
        bht_bank_rd_data_out_1_108 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_108 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_544_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_109 <= 2'h0;
    end else if (bht_bank_sel_1_6_13) begin
      if (_T_9851) begin
        bht_bank_rd_data_out_1_109 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_109 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_544_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_110 <= 2'h0;
    end else if (bht_bank_sel_1_6_14) begin
      if (_T_9860) begin
        bht_bank_rd_data_out_1_110 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_110 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_544_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_111 <= 2'h0;
    end else if (bht_bank_sel_1_6_15) begin
      if (_T_9869) begin
        bht_bank_rd_data_out_1_111 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_111 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_545_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_112 <= 2'h0;
    end else if (bht_bank_sel_1_7_0) begin
      if (_T_9878) begin
        bht_bank_rd_data_out_1_112 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_112 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_545_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_113 <= 2'h0;
    end else if (bht_bank_sel_1_7_1) begin
      if (_T_9887) begin
        bht_bank_rd_data_out_1_113 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_113 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_545_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_114 <= 2'h0;
    end else if (bht_bank_sel_1_7_2) begin
      if (_T_9896) begin
        bht_bank_rd_data_out_1_114 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_114 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_545_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_115 <= 2'h0;
    end else if (bht_bank_sel_1_7_3) begin
      if (_T_9905) begin
        bht_bank_rd_data_out_1_115 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_115 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_545_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_116 <= 2'h0;
    end else if (bht_bank_sel_1_7_4) begin
      if (_T_9914) begin
        bht_bank_rd_data_out_1_116 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_116 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_545_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_117 <= 2'h0;
    end else if (bht_bank_sel_1_7_5) begin
      if (_T_9923) begin
        bht_bank_rd_data_out_1_117 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_117 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_545_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_118 <= 2'h0;
    end else if (bht_bank_sel_1_7_6) begin
      if (_T_9932) begin
        bht_bank_rd_data_out_1_118 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_118 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_545_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_119 <= 2'h0;
    end else if (bht_bank_sel_1_7_7) begin
      if (_T_9941) begin
        bht_bank_rd_data_out_1_119 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_119 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_545_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_120 <= 2'h0;
    end else if (bht_bank_sel_1_7_8) begin
      if (_T_9950) begin
        bht_bank_rd_data_out_1_120 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_120 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_545_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_121 <= 2'h0;
    end else if (bht_bank_sel_1_7_9) begin
      if (_T_9959) begin
        bht_bank_rd_data_out_1_121 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_121 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_545_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_122 <= 2'h0;
    end else if (bht_bank_sel_1_7_10) begin
      if (_T_9968) begin
        bht_bank_rd_data_out_1_122 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_122 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_545_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_123 <= 2'h0;
    end else if (bht_bank_sel_1_7_11) begin
      if (_T_9977) begin
        bht_bank_rd_data_out_1_123 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_123 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_545_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_124 <= 2'h0;
    end else if (bht_bank_sel_1_7_12) begin
      if (_T_9986) begin
        bht_bank_rd_data_out_1_124 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_124 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_545_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_125 <= 2'h0;
    end else if (bht_bank_sel_1_7_13) begin
      if (_T_9995) begin
        bht_bank_rd_data_out_1_125 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_125 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_545_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_126 <= 2'h0;
    end else if (bht_bank_sel_1_7_14) begin
      if (_T_10004) begin
        bht_bank_rd_data_out_1_126 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_126 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_545_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_127 <= 2'h0;
    end else if (bht_bank_sel_1_7_15) begin
      if (_T_10013) begin
        bht_bank_rd_data_out_1_127 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_127 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_546_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_128 <= 2'h0;
    end else if (bht_bank_sel_1_8_0) begin
      if (_T_10022) begin
        bht_bank_rd_data_out_1_128 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_128 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_546_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_129 <= 2'h0;
    end else if (bht_bank_sel_1_8_1) begin
      if (_T_10031) begin
        bht_bank_rd_data_out_1_129 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_129 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_546_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_130 <= 2'h0;
    end else if (bht_bank_sel_1_8_2) begin
      if (_T_10040) begin
        bht_bank_rd_data_out_1_130 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_130 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_546_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_131 <= 2'h0;
    end else if (bht_bank_sel_1_8_3) begin
      if (_T_10049) begin
        bht_bank_rd_data_out_1_131 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_131 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_546_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_132 <= 2'h0;
    end else if (bht_bank_sel_1_8_4) begin
      if (_T_10058) begin
        bht_bank_rd_data_out_1_132 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_132 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_546_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_133 <= 2'h0;
    end else if (bht_bank_sel_1_8_5) begin
      if (_T_10067) begin
        bht_bank_rd_data_out_1_133 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_133 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_546_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_134 <= 2'h0;
    end else if (bht_bank_sel_1_8_6) begin
      if (_T_10076) begin
        bht_bank_rd_data_out_1_134 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_134 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_546_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_135 <= 2'h0;
    end else if (bht_bank_sel_1_8_7) begin
      if (_T_10085) begin
        bht_bank_rd_data_out_1_135 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_135 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_546_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_136 <= 2'h0;
    end else if (bht_bank_sel_1_8_8) begin
      if (_T_10094) begin
        bht_bank_rd_data_out_1_136 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_136 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_546_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_137 <= 2'h0;
    end else if (bht_bank_sel_1_8_9) begin
      if (_T_10103) begin
        bht_bank_rd_data_out_1_137 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_137 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_546_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_138 <= 2'h0;
    end else if (bht_bank_sel_1_8_10) begin
      if (_T_10112) begin
        bht_bank_rd_data_out_1_138 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_138 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_546_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_139 <= 2'h0;
    end else if (bht_bank_sel_1_8_11) begin
      if (_T_10121) begin
        bht_bank_rd_data_out_1_139 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_139 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_546_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_140 <= 2'h0;
    end else if (bht_bank_sel_1_8_12) begin
      if (_T_10130) begin
        bht_bank_rd_data_out_1_140 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_140 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_546_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_141 <= 2'h0;
    end else if (bht_bank_sel_1_8_13) begin
      if (_T_10139) begin
        bht_bank_rd_data_out_1_141 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_141 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_546_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_142 <= 2'h0;
    end else if (bht_bank_sel_1_8_14) begin
      if (_T_10148) begin
        bht_bank_rd_data_out_1_142 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_142 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_546_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_143 <= 2'h0;
    end else if (bht_bank_sel_1_8_15) begin
      if (_T_10157) begin
        bht_bank_rd_data_out_1_143 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_143 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_547_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_144 <= 2'h0;
    end else if (bht_bank_sel_1_9_0) begin
      if (_T_10166) begin
        bht_bank_rd_data_out_1_144 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_144 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_547_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_145 <= 2'h0;
    end else if (bht_bank_sel_1_9_1) begin
      if (_T_10175) begin
        bht_bank_rd_data_out_1_145 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_145 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_547_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_146 <= 2'h0;
    end else if (bht_bank_sel_1_9_2) begin
      if (_T_10184) begin
        bht_bank_rd_data_out_1_146 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_146 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_547_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_147 <= 2'h0;
    end else if (bht_bank_sel_1_9_3) begin
      if (_T_10193) begin
        bht_bank_rd_data_out_1_147 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_147 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_547_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_148 <= 2'h0;
    end else if (bht_bank_sel_1_9_4) begin
      if (_T_10202) begin
        bht_bank_rd_data_out_1_148 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_148 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_547_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_149 <= 2'h0;
    end else if (bht_bank_sel_1_9_5) begin
      if (_T_10211) begin
        bht_bank_rd_data_out_1_149 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_149 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_547_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_150 <= 2'h0;
    end else if (bht_bank_sel_1_9_6) begin
      if (_T_10220) begin
        bht_bank_rd_data_out_1_150 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_150 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_547_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_151 <= 2'h0;
    end else if (bht_bank_sel_1_9_7) begin
      if (_T_10229) begin
        bht_bank_rd_data_out_1_151 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_151 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_547_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_152 <= 2'h0;
    end else if (bht_bank_sel_1_9_8) begin
      if (_T_10238) begin
        bht_bank_rd_data_out_1_152 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_152 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_547_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_153 <= 2'h0;
    end else if (bht_bank_sel_1_9_9) begin
      if (_T_10247) begin
        bht_bank_rd_data_out_1_153 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_153 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_547_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_154 <= 2'h0;
    end else if (bht_bank_sel_1_9_10) begin
      if (_T_10256) begin
        bht_bank_rd_data_out_1_154 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_154 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_547_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_155 <= 2'h0;
    end else if (bht_bank_sel_1_9_11) begin
      if (_T_10265) begin
        bht_bank_rd_data_out_1_155 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_155 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_547_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_156 <= 2'h0;
    end else if (bht_bank_sel_1_9_12) begin
      if (_T_10274) begin
        bht_bank_rd_data_out_1_156 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_156 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_547_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_157 <= 2'h0;
    end else if (bht_bank_sel_1_9_13) begin
      if (_T_10283) begin
        bht_bank_rd_data_out_1_157 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_157 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_547_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_158 <= 2'h0;
    end else if (bht_bank_sel_1_9_14) begin
      if (_T_10292) begin
        bht_bank_rd_data_out_1_158 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_158 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_547_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_159 <= 2'h0;
    end else if (bht_bank_sel_1_9_15) begin
      if (_T_10301) begin
        bht_bank_rd_data_out_1_159 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_159 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_548_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_160 <= 2'h0;
    end else if (bht_bank_sel_1_10_0) begin
      if (_T_10310) begin
        bht_bank_rd_data_out_1_160 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_160 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_548_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_161 <= 2'h0;
    end else if (bht_bank_sel_1_10_1) begin
      if (_T_10319) begin
        bht_bank_rd_data_out_1_161 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_161 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_548_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_162 <= 2'h0;
    end else if (bht_bank_sel_1_10_2) begin
      if (_T_10328) begin
        bht_bank_rd_data_out_1_162 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_162 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_548_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_163 <= 2'h0;
    end else if (bht_bank_sel_1_10_3) begin
      if (_T_10337) begin
        bht_bank_rd_data_out_1_163 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_163 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_548_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_164 <= 2'h0;
    end else if (bht_bank_sel_1_10_4) begin
      if (_T_10346) begin
        bht_bank_rd_data_out_1_164 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_164 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_548_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_165 <= 2'h0;
    end else if (bht_bank_sel_1_10_5) begin
      if (_T_10355) begin
        bht_bank_rd_data_out_1_165 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_165 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_548_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_166 <= 2'h0;
    end else if (bht_bank_sel_1_10_6) begin
      if (_T_10364) begin
        bht_bank_rd_data_out_1_166 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_166 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_548_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_167 <= 2'h0;
    end else if (bht_bank_sel_1_10_7) begin
      if (_T_10373) begin
        bht_bank_rd_data_out_1_167 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_167 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_548_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_168 <= 2'h0;
    end else if (bht_bank_sel_1_10_8) begin
      if (_T_10382) begin
        bht_bank_rd_data_out_1_168 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_168 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_548_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_169 <= 2'h0;
    end else if (bht_bank_sel_1_10_9) begin
      if (_T_10391) begin
        bht_bank_rd_data_out_1_169 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_169 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_548_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_170 <= 2'h0;
    end else if (bht_bank_sel_1_10_10) begin
      if (_T_10400) begin
        bht_bank_rd_data_out_1_170 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_170 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_548_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_171 <= 2'h0;
    end else if (bht_bank_sel_1_10_11) begin
      if (_T_10409) begin
        bht_bank_rd_data_out_1_171 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_171 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_548_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_172 <= 2'h0;
    end else if (bht_bank_sel_1_10_12) begin
      if (_T_10418) begin
        bht_bank_rd_data_out_1_172 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_172 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_548_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_173 <= 2'h0;
    end else if (bht_bank_sel_1_10_13) begin
      if (_T_10427) begin
        bht_bank_rd_data_out_1_173 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_173 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_548_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_174 <= 2'h0;
    end else if (bht_bank_sel_1_10_14) begin
      if (_T_10436) begin
        bht_bank_rd_data_out_1_174 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_174 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_548_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_175 <= 2'h0;
    end else if (bht_bank_sel_1_10_15) begin
      if (_T_10445) begin
        bht_bank_rd_data_out_1_175 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_175 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_549_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_176 <= 2'h0;
    end else if (bht_bank_sel_1_11_0) begin
      if (_T_10454) begin
        bht_bank_rd_data_out_1_176 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_176 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_549_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_177 <= 2'h0;
    end else if (bht_bank_sel_1_11_1) begin
      if (_T_10463) begin
        bht_bank_rd_data_out_1_177 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_177 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_549_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_178 <= 2'h0;
    end else if (bht_bank_sel_1_11_2) begin
      if (_T_10472) begin
        bht_bank_rd_data_out_1_178 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_178 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_549_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_179 <= 2'h0;
    end else if (bht_bank_sel_1_11_3) begin
      if (_T_10481) begin
        bht_bank_rd_data_out_1_179 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_179 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_549_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_180 <= 2'h0;
    end else if (bht_bank_sel_1_11_4) begin
      if (_T_10490) begin
        bht_bank_rd_data_out_1_180 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_180 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_549_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_181 <= 2'h0;
    end else if (bht_bank_sel_1_11_5) begin
      if (_T_10499) begin
        bht_bank_rd_data_out_1_181 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_181 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_549_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_182 <= 2'h0;
    end else if (bht_bank_sel_1_11_6) begin
      if (_T_10508) begin
        bht_bank_rd_data_out_1_182 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_182 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_549_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_183 <= 2'h0;
    end else if (bht_bank_sel_1_11_7) begin
      if (_T_10517) begin
        bht_bank_rd_data_out_1_183 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_183 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_549_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_184 <= 2'h0;
    end else if (bht_bank_sel_1_11_8) begin
      if (_T_10526) begin
        bht_bank_rd_data_out_1_184 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_184 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_549_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_185 <= 2'h0;
    end else if (bht_bank_sel_1_11_9) begin
      if (_T_10535) begin
        bht_bank_rd_data_out_1_185 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_185 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_549_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_186 <= 2'h0;
    end else if (bht_bank_sel_1_11_10) begin
      if (_T_10544) begin
        bht_bank_rd_data_out_1_186 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_186 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_549_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_187 <= 2'h0;
    end else if (bht_bank_sel_1_11_11) begin
      if (_T_10553) begin
        bht_bank_rd_data_out_1_187 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_187 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_549_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_188 <= 2'h0;
    end else if (bht_bank_sel_1_11_12) begin
      if (_T_10562) begin
        bht_bank_rd_data_out_1_188 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_188 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_549_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_189 <= 2'h0;
    end else if (bht_bank_sel_1_11_13) begin
      if (_T_10571) begin
        bht_bank_rd_data_out_1_189 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_189 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_549_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_190 <= 2'h0;
    end else if (bht_bank_sel_1_11_14) begin
      if (_T_10580) begin
        bht_bank_rd_data_out_1_190 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_190 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_549_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_191 <= 2'h0;
    end else if (bht_bank_sel_1_11_15) begin
      if (_T_10589) begin
        bht_bank_rd_data_out_1_191 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_191 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_550_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_192 <= 2'h0;
    end else if (bht_bank_sel_1_12_0) begin
      if (_T_10598) begin
        bht_bank_rd_data_out_1_192 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_192 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_550_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_193 <= 2'h0;
    end else if (bht_bank_sel_1_12_1) begin
      if (_T_10607) begin
        bht_bank_rd_data_out_1_193 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_193 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_550_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_194 <= 2'h0;
    end else if (bht_bank_sel_1_12_2) begin
      if (_T_10616) begin
        bht_bank_rd_data_out_1_194 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_194 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_550_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_195 <= 2'h0;
    end else if (bht_bank_sel_1_12_3) begin
      if (_T_10625) begin
        bht_bank_rd_data_out_1_195 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_195 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_550_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_196 <= 2'h0;
    end else if (bht_bank_sel_1_12_4) begin
      if (_T_10634) begin
        bht_bank_rd_data_out_1_196 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_196 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_550_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_197 <= 2'h0;
    end else if (bht_bank_sel_1_12_5) begin
      if (_T_10643) begin
        bht_bank_rd_data_out_1_197 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_197 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_550_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_198 <= 2'h0;
    end else if (bht_bank_sel_1_12_6) begin
      if (_T_10652) begin
        bht_bank_rd_data_out_1_198 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_198 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_550_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_199 <= 2'h0;
    end else if (bht_bank_sel_1_12_7) begin
      if (_T_10661) begin
        bht_bank_rd_data_out_1_199 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_199 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_550_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_200 <= 2'h0;
    end else if (bht_bank_sel_1_12_8) begin
      if (_T_10670) begin
        bht_bank_rd_data_out_1_200 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_200 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_550_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_201 <= 2'h0;
    end else if (bht_bank_sel_1_12_9) begin
      if (_T_10679) begin
        bht_bank_rd_data_out_1_201 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_201 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_550_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_202 <= 2'h0;
    end else if (bht_bank_sel_1_12_10) begin
      if (_T_10688) begin
        bht_bank_rd_data_out_1_202 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_202 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_550_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_203 <= 2'h0;
    end else if (bht_bank_sel_1_12_11) begin
      if (_T_10697) begin
        bht_bank_rd_data_out_1_203 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_203 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_550_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_204 <= 2'h0;
    end else if (bht_bank_sel_1_12_12) begin
      if (_T_10706) begin
        bht_bank_rd_data_out_1_204 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_204 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_550_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_205 <= 2'h0;
    end else if (bht_bank_sel_1_12_13) begin
      if (_T_10715) begin
        bht_bank_rd_data_out_1_205 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_205 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_550_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_206 <= 2'h0;
    end else if (bht_bank_sel_1_12_14) begin
      if (_T_10724) begin
        bht_bank_rd_data_out_1_206 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_206 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_550_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_207 <= 2'h0;
    end else if (bht_bank_sel_1_12_15) begin
      if (_T_10733) begin
        bht_bank_rd_data_out_1_207 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_207 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_551_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_208 <= 2'h0;
    end else if (bht_bank_sel_1_13_0) begin
      if (_T_10742) begin
        bht_bank_rd_data_out_1_208 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_208 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_551_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_209 <= 2'h0;
    end else if (bht_bank_sel_1_13_1) begin
      if (_T_10751) begin
        bht_bank_rd_data_out_1_209 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_209 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_551_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_210 <= 2'h0;
    end else if (bht_bank_sel_1_13_2) begin
      if (_T_10760) begin
        bht_bank_rd_data_out_1_210 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_210 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_551_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_211 <= 2'h0;
    end else if (bht_bank_sel_1_13_3) begin
      if (_T_10769) begin
        bht_bank_rd_data_out_1_211 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_211 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_551_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_212 <= 2'h0;
    end else if (bht_bank_sel_1_13_4) begin
      if (_T_10778) begin
        bht_bank_rd_data_out_1_212 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_212 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_551_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_213 <= 2'h0;
    end else if (bht_bank_sel_1_13_5) begin
      if (_T_10787) begin
        bht_bank_rd_data_out_1_213 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_213 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_551_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_214 <= 2'h0;
    end else if (bht_bank_sel_1_13_6) begin
      if (_T_10796) begin
        bht_bank_rd_data_out_1_214 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_214 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_551_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_215 <= 2'h0;
    end else if (bht_bank_sel_1_13_7) begin
      if (_T_10805) begin
        bht_bank_rd_data_out_1_215 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_215 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_551_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_216 <= 2'h0;
    end else if (bht_bank_sel_1_13_8) begin
      if (_T_10814) begin
        bht_bank_rd_data_out_1_216 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_216 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_551_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_217 <= 2'h0;
    end else if (bht_bank_sel_1_13_9) begin
      if (_T_10823) begin
        bht_bank_rd_data_out_1_217 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_217 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_551_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_218 <= 2'h0;
    end else if (bht_bank_sel_1_13_10) begin
      if (_T_10832) begin
        bht_bank_rd_data_out_1_218 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_218 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_551_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_219 <= 2'h0;
    end else if (bht_bank_sel_1_13_11) begin
      if (_T_10841) begin
        bht_bank_rd_data_out_1_219 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_219 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_551_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_220 <= 2'h0;
    end else if (bht_bank_sel_1_13_12) begin
      if (_T_10850) begin
        bht_bank_rd_data_out_1_220 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_220 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_551_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_221 <= 2'h0;
    end else if (bht_bank_sel_1_13_13) begin
      if (_T_10859) begin
        bht_bank_rd_data_out_1_221 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_221 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_551_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_222 <= 2'h0;
    end else if (bht_bank_sel_1_13_14) begin
      if (_T_10868) begin
        bht_bank_rd_data_out_1_222 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_222 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_551_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_223 <= 2'h0;
    end else if (bht_bank_sel_1_13_15) begin
      if (_T_10877) begin
        bht_bank_rd_data_out_1_223 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_223 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_552_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_224 <= 2'h0;
    end else if (bht_bank_sel_1_14_0) begin
      if (_T_10886) begin
        bht_bank_rd_data_out_1_224 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_224 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_552_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_225 <= 2'h0;
    end else if (bht_bank_sel_1_14_1) begin
      if (_T_10895) begin
        bht_bank_rd_data_out_1_225 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_225 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_552_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_226 <= 2'h0;
    end else if (bht_bank_sel_1_14_2) begin
      if (_T_10904) begin
        bht_bank_rd_data_out_1_226 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_226 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_552_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_227 <= 2'h0;
    end else if (bht_bank_sel_1_14_3) begin
      if (_T_10913) begin
        bht_bank_rd_data_out_1_227 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_227 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_552_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_228 <= 2'h0;
    end else if (bht_bank_sel_1_14_4) begin
      if (_T_10922) begin
        bht_bank_rd_data_out_1_228 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_228 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_552_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_229 <= 2'h0;
    end else if (bht_bank_sel_1_14_5) begin
      if (_T_10931) begin
        bht_bank_rd_data_out_1_229 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_229 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_552_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_230 <= 2'h0;
    end else if (bht_bank_sel_1_14_6) begin
      if (_T_10940) begin
        bht_bank_rd_data_out_1_230 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_230 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_552_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_231 <= 2'h0;
    end else if (bht_bank_sel_1_14_7) begin
      if (_T_10949) begin
        bht_bank_rd_data_out_1_231 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_231 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_552_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_232 <= 2'h0;
    end else if (bht_bank_sel_1_14_8) begin
      if (_T_10958) begin
        bht_bank_rd_data_out_1_232 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_232 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_552_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_233 <= 2'h0;
    end else if (bht_bank_sel_1_14_9) begin
      if (_T_10967) begin
        bht_bank_rd_data_out_1_233 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_233 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_552_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_234 <= 2'h0;
    end else if (bht_bank_sel_1_14_10) begin
      if (_T_10976) begin
        bht_bank_rd_data_out_1_234 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_234 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_552_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_235 <= 2'h0;
    end else if (bht_bank_sel_1_14_11) begin
      if (_T_10985) begin
        bht_bank_rd_data_out_1_235 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_235 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_552_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_236 <= 2'h0;
    end else if (bht_bank_sel_1_14_12) begin
      if (_T_10994) begin
        bht_bank_rd_data_out_1_236 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_236 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_552_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_237 <= 2'h0;
    end else if (bht_bank_sel_1_14_13) begin
      if (_T_11003) begin
        bht_bank_rd_data_out_1_237 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_237 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_552_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_238 <= 2'h0;
    end else if (bht_bank_sel_1_14_14) begin
      if (_T_11012) begin
        bht_bank_rd_data_out_1_238 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_238 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_552_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_239 <= 2'h0;
    end else if (bht_bank_sel_1_14_15) begin
      if (_T_11021) begin
        bht_bank_rd_data_out_1_239 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_239 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_553_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_240 <= 2'h0;
    end else if (bht_bank_sel_1_15_0) begin
      if (_T_11030) begin
        bht_bank_rd_data_out_1_240 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_240 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_553_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_241 <= 2'h0;
    end else if (bht_bank_sel_1_15_1) begin
      if (_T_11039) begin
        bht_bank_rd_data_out_1_241 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_241 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_553_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_242 <= 2'h0;
    end else if (bht_bank_sel_1_15_2) begin
      if (_T_11048) begin
        bht_bank_rd_data_out_1_242 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_242 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_553_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_243 <= 2'h0;
    end else if (bht_bank_sel_1_15_3) begin
      if (_T_11057) begin
        bht_bank_rd_data_out_1_243 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_243 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_553_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_244 <= 2'h0;
    end else if (bht_bank_sel_1_15_4) begin
      if (_T_11066) begin
        bht_bank_rd_data_out_1_244 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_244 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_553_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_245 <= 2'h0;
    end else if (bht_bank_sel_1_15_5) begin
      if (_T_11075) begin
        bht_bank_rd_data_out_1_245 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_245 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_553_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_246 <= 2'h0;
    end else if (bht_bank_sel_1_15_6) begin
      if (_T_11084) begin
        bht_bank_rd_data_out_1_246 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_246 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_553_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_247 <= 2'h0;
    end else if (bht_bank_sel_1_15_7) begin
      if (_T_11093) begin
        bht_bank_rd_data_out_1_247 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_247 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_553_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_248 <= 2'h0;
    end else if (bht_bank_sel_1_15_8) begin
      if (_T_11102) begin
        bht_bank_rd_data_out_1_248 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_248 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_553_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_249 <= 2'h0;
    end else if (bht_bank_sel_1_15_9) begin
      if (_T_11111) begin
        bht_bank_rd_data_out_1_249 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_249 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_553_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_250 <= 2'h0;
    end else if (bht_bank_sel_1_15_10) begin
      if (_T_11120) begin
        bht_bank_rd_data_out_1_250 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_250 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_553_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_251 <= 2'h0;
    end else if (bht_bank_sel_1_15_11) begin
      if (_T_11129) begin
        bht_bank_rd_data_out_1_251 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_251 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_553_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_252 <= 2'h0;
    end else if (bht_bank_sel_1_15_12) begin
      if (_T_11138) begin
        bht_bank_rd_data_out_1_252 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_252 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_553_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_253 <= 2'h0;
    end else if (bht_bank_sel_1_15_13) begin
      if (_T_11147) begin
        bht_bank_rd_data_out_1_253 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_253 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_553_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_254 <= 2'h0;
    end else if (bht_bank_sel_1_15_14) begin
      if (_T_11156) begin
        bht_bank_rd_data_out_1_254 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_254 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_553_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_255 <= 2'h0;
    end else if (bht_bank_sel_1_15_15) begin
      if (_T_11165) begin
        bht_bank_rd_data_out_1_255 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_255 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_522_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_0 <= 2'h0;
    end else if (bht_bank_sel_0_0_0) begin
      if (_T_6566) begin
        bht_bank_rd_data_out_0_0 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_0 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_522_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_1 <= 2'h0;
    end else if (bht_bank_sel_0_0_1) begin
      if (_T_6575) begin
        bht_bank_rd_data_out_0_1 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_1 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_522_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_2 <= 2'h0;
    end else if (bht_bank_sel_0_0_2) begin
      if (_T_6584) begin
        bht_bank_rd_data_out_0_2 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_2 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_522_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_3 <= 2'h0;
    end else if (bht_bank_sel_0_0_3) begin
      if (_T_6593) begin
        bht_bank_rd_data_out_0_3 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_3 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_522_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_4 <= 2'h0;
    end else if (bht_bank_sel_0_0_4) begin
      if (_T_6602) begin
        bht_bank_rd_data_out_0_4 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_4 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_522_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_5 <= 2'h0;
    end else if (bht_bank_sel_0_0_5) begin
      if (_T_6611) begin
        bht_bank_rd_data_out_0_5 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_5 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_522_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_6 <= 2'h0;
    end else if (bht_bank_sel_0_0_6) begin
      if (_T_6620) begin
        bht_bank_rd_data_out_0_6 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_6 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_522_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_7 <= 2'h0;
    end else if (bht_bank_sel_0_0_7) begin
      if (_T_6629) begin
        bht_bank_rd_data_out_0_7 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_7 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_522_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_8 <= 2'h0;
    end else if (bht_bank_sel_0_0_8) begin
      if (_T_6638) begin
        bht_bank_rd_data_out_0_8 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_8 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_522_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_9 <= 2'h0;
    end else if (bht_bank_sel_0_0_9) begin
      if (_T_6647) begin
        bht_bank_rd_data_out_0_9 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_9 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_522_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_10 <= 2'h0;
    end else if (bht_bank_sel_0_0_10) begin
      if (_T_6656) begin
        bht_bank_rd_data_out_0_10 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_10 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_522_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_11 <= 2'h0;
    end else if (bht_bank_sel_0_0_11) begin
      if (_T_6665) begin
        bht_bank_rd_data_out_0_11 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_11 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_522_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_12 <= 2'h0;
    end else if (bht_bank_sel_0_0_12) begin
      if (_T_6674) begin
        bht_bank_rd_data_out_0_12 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_12 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_522_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_13 <= 2'h0;
    end else if (bht_bank_sel_0_0_13) begin
      if (_T_6683) begin
        bht_bank_rd_data_out_0_13 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_13 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_522_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_14 <= 2'h0;
    end else if (bht_bank_sel_0_0_14) begin
      if (_T_6692) begin
        bht_bank_rd_data_out_0_14 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_14 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_522_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_15 <= 2'h0;
    end else if (bht_bank_sel_0_0_15) begin
      if (_T_6701) begin
        bht_bank_rd_data_out_0_15 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_15 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_523_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_16 <= 2'h0;
    end else if (bht_bank_sel_0_1_0) begin
      if (_T_6710) begin
        bht_bank_rd_data_out_0_16 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_16 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_523_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_17 <= 2'h0;
    end else if (bht_bank_sel_0_1_1) begin
      if (_T_6719) begin
        bht_bank_rd_data_out_0_17 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_17 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_523_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_18 <= 2'h0;
    end else if (bht_bank_sel_0_1_2) begin
      if (_T_6728) begin
        bht_bank_rd_data_out_0_18 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_18 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_523_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_19 <= 2'h0;
    end else if (bht_bank_sel_0_1_3) begin
      if (_T_6737) begin
        bht_bank_rd_data_out_0_19 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_19 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_523_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_20 <= 2'h0;
    end else if (bht_bank_sel_0_1_4) begin
      if (_T_6746) begin
        bht_bank_rd_data_out_0_20 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_20 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_523_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_21 <= 2'h0;
    end else if (bht_bank_sel_0_1_5) begin
      if (_T_6755) begin
        bht_bank_rd_data_out_0_21 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_21 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_523_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_22 <= 2'h0;
    end else if (bht_bank_sel_0_1_6) begin
      if (_T_6764) begin
        bht_bank_rd_data_out_0_22 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_22 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_523_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_23 <= 2'h0;
    end else if (bht_bank_sel_0_1_7) begin
      if (_T_6773) begin
        bht_bank_rd_data_out_0_23 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_23 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_523_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_24 <= 2'h0;
    end else if (bht_bank_sel_0_1_8) begin
      if (_T_6782) begin
        bht_bank_rd_data_out_0_24 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_24 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_523_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_25 <= 2'h0;
    end else if (bht_bank_sel_0_1_9) begin
      if (_T_6791) begin
        bht_bank_rd_data_out_0_25 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_25 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_523_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_26 <= 2'h0;
    end else if (bht_bank_sel_0_1_10) begin
      if (_T_6800) begin
        bht_bank_rd_data_out_0_26 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_26 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_523_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_27 <= 2'h0;
    end else if (bht_bank_sel_0_1_11) begin
      if (_T_6809) begin
        bht_bank_rd_data_out_0_27 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_27 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_523_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_28 <= 2'h0;
    end else if (bht_bank_sel_0_1_12) begin
      if (_T_6818) begin
        bht_bank_rd_data_out_0_28 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_28 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_523_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_29 <= 2'h0;
    end else if (bht_bank_sel_0_1_13) begin
      if (_T_6827) begin
        bht_bank_rd_data_out_0_29 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_29 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_523_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_30 <= 2'h0;
    end else if (bht_bank_sel_0_1_14) begin
      if (_T_6836) begin
        bht_bank_rd_data_out_0_30 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_30 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_523_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_31 <= 2'h0;
    end else if (bht_bank_sel_0_1_15) begin
      if (_T_6845) begin
        bht_bank_rd_data_out_0_31 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_31 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_524_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_32 <= 2'h0;
    end else if (bht_bank_sel_0_2_0) begin
      if (_T_6854) begin
        bht_bank_rd_data_out_0_32 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_32 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_524_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_33 <= 2'h0;
    end else if (bht_bank_sel_0_2_1) begin
      if (_T_6863) begin
        bht_bank_rd_data_out_0_33 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_33 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_524_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_34 <= 2'h0;
    end else if (bht_bank_sel_0_2_2) begin
      if (_T_6872) begin
        bht_bank_rd_data_out_0_34 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_34 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_524_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_35 <= 2'h0;
    end else if (bht_bank_sel_0_2_3) begin
      if (_T_6881) begin
        bht_bank_rd_data_out_0_35 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_35 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_524_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_36 <= 2'h0;
    end else if (bht_bank_sel_0_2_4) begin
      if (_T_6890) begin
        bht_bank_rd_data_out_0_36 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_36 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_524_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_37 <= 2'h0;
    end else if (bht_bank_sel_0_2_5) begin
      if (_T_6899) begin
        bht_bank_rd_data_out_0_37 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_37 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_524_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_38 <= 2'h0;
    end else if (bht_bank_sel_0_2_6) begin
      if (_T_6908) begin
        bht_bank_rd_data_out_0_38 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_38 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_524_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_39 <= 2'h0;
    end else if (bht_bank_sel_0_2_7) begin
      if (_T_6917) begin
        bht_bank_rd_data_out_0_39 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_39 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_524_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_40 <= 2'h0;
    end else if (bht_bank_sel_0_2_8) begin
      if (_T_6926) begin
        bht_bank_rd_data_out_0_40 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_40 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_524_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_41 <= 2'h0;
    end else if (bht_bank_sel_0_2_9) begin
      if (_T_6935) begin
        bht_bank_rd_data_out_0_41 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_41 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_524_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_42 <= 2'h0;
    end else if (bht_bank_sel_0_2_10) begin
      if (_T_6944) begin
        bht_bank_rd_data_out_0_42 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_42 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_524_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_43 <= 2'h0;
    end else if (bht_bank_sel_0_2_11) begin
      if (_T_6953) begin
        bht_bank_rd_data_out_0_43 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_43 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_524_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_44 <= 2'h0;
    end else if (bht_bank_sel_0_2_12) begin
      if (_T_6962) begin
        bht_bank_rd_data_out_0_44 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_44 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_524_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_45 <= 2'h0;
    end else if (bht_bank_sel_0_2_13) begin
      if (_T_6971) begin
        bht_bank_rd_data_out_0_45 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_45 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_524_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_46 <= 2'h0;
    end else if (bht_bank_sel_0_2_14) begin
      if (_T_6980) begin
        bht_bank_rd_data_out_0_46 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_46 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_524_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_47 <= 2'h0;
    end else if (bht_bank_sel_0_2_15) begin
      if (_T_6989) begin
        bht_bank_rd_data_out_0_47 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_47 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_525_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_48 <= 2'h0;
    end else if (bht_bank_sel_0_3_0) begin
      if (_T_6998) begin
        bht_bank_rd_data_out_0_48 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_48 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_525_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_49 <= 2'h0;
    end else if (bht_bank_sel_0_3_1) begin
      if (_T_7007) begin
        bht_bank_rd_data_out_0_49 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_49 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_525_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_50 <= 2'h0;
    end else if (bht_bank_sel_0_3_2) begin
      if (_T_7016) begin
        bht_bank_rd_data_out_0_50 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_50 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_525_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_51 <= 2'h0;
    end else if (bht_bank_sel_0_3_3) begin
      if (_T_7025) begin
        bht_bank_rd_data_out_0_51 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_51 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_525_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_52 <= 2'h0;
    end else if (bht_bank_sel_0_3_4) begin
      if (_T_7034) begin
        bht_bank_rd_data_out_0_52 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_52 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_525_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_53 <= 2'h0;
    end else if (bht_bank_sel_0_3_5) begin
      if (_T_7043) begin
        bht_bank_rd_data_out_0_53 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_53 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_525_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_54 <= 2'h0;
    end else if (bht_bank_sel_0_3_6) begin
      if (_T_7052) begin
        bht_bank_rd_data_out_0_54 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_54 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_525_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_55 <= 2'h0;
    end else if (bht_bank_sel_0_3_7) begin
      if (_T_7061) begin
        bht_bank_rd_data_out_0_55 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_55 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_525_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_56 <= 2'h0;
    end else if (bht_bank_sel_0_3_8) begin
      if (_T_7070) begin
        bht_bank_rd_data_out_0_56 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_56 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_525_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_57 <= 2'h0;
    end else if (bht_bank_sel_0_3_9) begin
      if (_T_7079) begin
        bht_bank_rd_data_out_0_57 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_57 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_525_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_58 <= 2'h0;
    end else if (bht_bank_sel_0_3_10) begin
      if (_T_7088) begin
        bht_bank_rd_data_out_0_58 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_58 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_525_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_59 <= 2'h0;
    end else if (bht_bank_sel_0_3_11) begin
      if (_T_7097) begin
        bht_bank_rd_data_out_0_59 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_59 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_525_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_60 <= 2'h0;
    end else if (bht_bank_sel_0_3_12) begin
      if (_T_7106) begin
        bht_bank_rd_data_out_0_60 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_60 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_525_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_61 <= 2'h0;
    end else if (bht_bank_sel_0_3_13) begin
      if (_T_7115) begin
        bht_bank_rd_data_out_0_61 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_61 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_525_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_62 <= 2'h0;
    end else if (bht_bank_sel_0_3_14) begin
      if (_T_7124) begin
        bht_bank_rd_data_out_0_62 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_62 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_525_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_63 <= 2'h0;
    end else if (bht_bank_sel_0_3_15) begin
      if (_T_7133) begin
        bht_bank_rd_data_out_0_63 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_63 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_526_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_64 <= 2'h0;
    end else if (bht_bank_sel_0_4_0) begin
      if (_T_7142) begin
        bht_bank_rd_data_out_0_64 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_64 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_526_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_65 <= 2'h0;
    end else if (bht_bank_sel_0_4_1) begin
      if (_T_7151) begin
        bht_bank_rd_data_out_0_65 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_65 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_526_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_66 <= 2'h0;
    end else if (bht_bank_sel_0_4_2) begin
      if (_T_7160) begin
        bht_bank_rd_data_out_0_66 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_66 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_526_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_67 <= 2'h0;
    end else if (bht_bank_sel_0_4_3) begin
      if (_T_7169) begin
        bht_bank_rd_data_out_0_67 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_67 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_526_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_68 <= 2'h0;
    end else if (bht_bank_sel_0_4_4) begin
      if (_T_7178) begin
        bht_bank_rd_data_out_0_68 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_68 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_526_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_69 <= 2'h0;
    end else if (bht_bank_sel_0_4_5) begin
      if (_T_7187) begin
        bht_bank_rd_data_out_0_69 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_69 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_526_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_70 <= 2'h0;
    end else if (bht_bank_sel_0_4_6) begin
      if (_T_7196) begin
        bht_bank_rd_data_out_0_70 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_70 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_526_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_71 <= 2'h0;
    end else if (bht_bank_sel_0_4_7) begin
      if (_T_7205) begin
        bht_bank_rd_data_out_0_71 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_71 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_526_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_72 <= 2'h0;
    end else if (bht_bank_sel_0_4_8) begin
      if (_T_7214) begin
        bht_bank_rd_data_out_0_72 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_72 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_526_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_73 <= 2'h0;
    end else if (bht_bank_sel_0_4_9) begin
      if (_T_7223) begin
        bht_bank_rd_data_out_0_73 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_73 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_526_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_74 <= 2'h0;
    end else if (bht_bank_sel_0_4_10) begin
      if (_T_7232) begin
        bht_bank_rd_data_out_0_74 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_74 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_526_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_75 <= 2'h0;
    end else if (bht_bank_sel_0_4_11) begin
      if (_T_7241) begin
        bht_bank_rd_data_out_0_75 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_75 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_526_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_76 <= 2'h0;
    end else if (bht_bank_sel_0_4_12) begin
      if (_T_7250) begin
        bht_bank_rd_data_out_0_76 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_76 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_526_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_77 <= 2'h0;
    end else if (bht_bank_sel_0_4_13) begin
      if (_T_7259) begin
        bht_bank_rd_data_out_0_77 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_77 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_526_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_78 <= 2'h0;
    end else if (bht_bank_sel_0_4_14) begin
      if (_T_7268) begin
        bht_bank_rd_data_out_0_78 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_78 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_526_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_79 <= 2'h0;
    end else if (bht_bank_sel_0_4_15) begin
      if (_T_7277) begin
        bht_bank_rd_data_out_0_79 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_79 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_527_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_80 <= 2'h0;
    end else if (bht_bank_sel_0_5_0) begin
      if (_T_7286) begin
        bht_bank_rd_data_out_0_80 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_80 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_527_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_81 <= 2'h0;
    end else if (bht_bank_sel_0_5_1) begin
      if (_T_7295) begin
        bht_bank_rd_data_out_0_81 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_81 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_527_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_82 <= 2'h0;
    end else if (bht_bank_sel_0_5_2) begin
      if (_T_7304) begin
        bht_bank_rd_data_out_0_82 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_82 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_527_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_83 <= 2'h0;
    end else if (bht_bank_sel_0_5_3) begin
      if (_T_7313) begin
        bht_bank_rd_data_out_0_83 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_83 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_527_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_84 <= 2'h0;
    end else if (bht_bank_sel_0_5_4) begin
      if (_T_7322) begin
        bht_bank_rd_data_out_0_84 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_84 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_527_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_85 <= 2'h0;
    end else if (bht_bank_sel_0_5_5) begin
      if (_T_7331) begin
        bht_bank_rd_data_out_0_85 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_85 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_527_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_86 <= 2'h0;
    end else if (bht_bank_sel_0_5_6) begin
      if (_T_7340) begin
        bht_bank_rd_data_out_0_86 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_86 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_527_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_87 <= 2'h0;
    end else if (bht_bank_sel_0_5_7) begin
      if (_T_7349) begin
        bht_bank_rd_data_out_0_87 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_87 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_527_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_88 <= 2'h0;
    end else if (bht_bank_sel_0_5_8) begin
      if (_T_7358) begin
        bht_bank_rd_data_out_0_88 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_88 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_527_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_89 <= 2'h0;
    end else if (bht_bank_sel_0_5_9) begin
      if (_T_7367) begin
        bht_bank_rd_data_out_0_89 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_89 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_527_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_90 <= 2'h0;
    end else if (bht_bank_sel_0_5_10) begin
      if (_T_7376) begin
        bht_bank_rd_data_out_0_90 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_90 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_527_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_91 <= 2'h0;
    end else if (bht_bank_sel_0_5_11) begin
      if (_T_7385) begin
        bht_bank_rd_data_out_0_91 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_91 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_527_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_92 <= 2'h0;
    end else if (bht_bank_sel_0_5_12) begin
      if (_T_7394) begin
        bht_bank_rd_data_out_0_92 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_92 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_527_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_93 <= 2'h0;
    end else if (bht_bank_sel_0_5_13) begin
      if (_T_7403) begin
        bht_bank_rd_data_out_0_93 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_93 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_527_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_94 <= 2'h0;
    end else if (bht_bank_sel_0_5_14) begin
      if (_T_7412) begin
        bht_bank_rd_data_out_0_94 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_94 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_527_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_95 <= 2'h0;
    end else if (bht_bank_sel_0_5_15) begin
      if (_T_7421) begin
        bht_bank_rd_data_out_0_95 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_95 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_528_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_96 <= 2'h0;
    end else if (bht_bank_sel_0_6_0) begin
      if (_T_7430) begin
        bht_bank_rd_data_out_0_96 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_96 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_528_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_97 <= 2'h0;
    end else if (bht_bank_sel_0_6_1) begin
      if (_T_7439) begin
        bht_bank_rd_data_out_0_97 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_97 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_528_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_98 <= 2'h0;
    end else if (bht_bank_sel_0_6_2) begin
      if (_T_7448) begin
        bht_bank_rd_data_out_0_98 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_98 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_528_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_99 <= 2'h0;
    end else if (bht_bank_sel_0_6_3) begin
      if (_T_7457) begin
        bht_bank_rd_data_out_0_99 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_99 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_528_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_100 <= 2'h0;
    end else if (bht_bank_sel_0_6_4) begin
      if (_T_7466) begin
        bht_bank_rd_data_out_0_100 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_100 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_528_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_101 <= 2'h0;
    end else if (bht_bank_sel_0_6_5) begin
      if (_T_7475) begin
        bht_bank_rd_data_out_0_101 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_101 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_528_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_102 <= 2'h0;
    end else if (bht_bank_sel_0_6_6) begin
      if (_T_7484) begin
        bht_bank_rd_data_out_0_102 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_102 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_528_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_103 <= 2'h0;
    end else if (bht_bank_sel_0_6_7) begin
      if (_T_7493) begin
        bht_bank_rd_data_out_0_103 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_103 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_528_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_104 <= 2'h0;
    end else if (bht_bank_sel_0_6_8) begin
      if (_T_7502) begin
        bht_bank_rd_data_out_0_104 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_104 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_528_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_105 <= 2'h0;
    end else if (bht_bank_sel_0_6_9) begin
      if (_T_7511) begin
        bht_bank_rd_data_out_0_105 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_105 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_528_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_106 <= 2'h0;
    end else if (bht_bank_sel_0_6_10) begin
      if (_T_7520) begin
        bht_bank_rd_data_out_0_106 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_106 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_528_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_107 <= 2'h0;
    end else if (bht_bank_sel_0_6_11) begin
      if (_T_7529) begin
        bht_bank_rd_data_out_0_107 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_107 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_528_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_108 <= 2'h0;
    end else if (bht_bank_sel_0_6_12) begin
      if (_T_7538) begin
        bht_bank_rd_data_out_0_108 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_108 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_528_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_109 <= 2'h0;
    end else if (bht_bank_sel_0_6_13) begin
      if (_T_7547) begin
        bht_bank_rd_data_out_0_109 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_109 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_528_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_110 <= 2'h0;
    end else if (bht_bank_sel_0_6_14) begin
      if (_T_7556) begin
        bht_bank_rd_data_out_0_110 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_110 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_528_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_111 <= 2'h0;
    end else if (bht_bank_sel_0_6_15) begin
      if (_T_7565) begin
        bht_bank_rd_data_out_0_111 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_111 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_529_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_112 <= 2'h0;
    end else if (bht_bank_sel_0_7_0) begin
      if (_T_7574) begin
        bht_bank_rd_data_out_0_112 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_112 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_529_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_113 <= 2'h0;
    end else if (bht_bank_sel_0_7_1) begin
      if (_T_7583) begin
        bht_bank_rd_data_out_0_113 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_113 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_529_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_114 <= 2'h0;
    end else if (bht_bank_sel_0_7_2) begin
      if (_T_7592) begin
        bht_bank_rd_data_out_0_114 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_114 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_529_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_115 <= 2'h0;
    end else if (bht_bank_sel_0_7_3) begin
      if (_T_7601) begin
        bht_bank_rd_data_out_0_115 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_115 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_529_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_116 <= 2'h0;
    end else if (bht_bank_sel_0_7_4) begin
      if (_T_7610) begin
        bht_bank_rd_data_out_0_116 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_116 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_529_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_117 <= 2'h0;
    end else if (bht_bank_sel_0_7_5) begin
      if (_T_7619) begin
        bht_bank_rd_data_out_0_117 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_117 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_529_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_118 <= 2'h0;
    end else if (bht_bank_sel_0_7_6) begin
      if (_T_7628) begin
        bht_bank_rd_data_out_0_118 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_118 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_529_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_119 <= 2'h0;
    end else if (bht_bank_sel_0_7_7) begin
      if (_T_7637) begin
        bht_bank_rd_data_out_0_119 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_119 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_529_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_120 <= 2'h0;
    end else if (bht_bank_sel_0_7_8) begin
      if (_T_7646) begin
        bht_bank_rd_data_out_0_120 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_120 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_529_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_121 <= 2'h0;
    end else if (bht_bank_sel_0_7_9) begin
      if (_T_7655) begin
        bht_bank_rd_data_out_0_121 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_121 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_529_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_122 <= 2'h0;
    end else if (bht_bank_sel_0_7_10) begin
      if (_T_7664) begin
        bht_bank_rd_data_out_0_122 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_122 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_529_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_123 <= 2'h0;
    end else if (bht_bank_sel_0_7_11) begin
      if (_T_7673) begin
        bht_bank_rd_data_out_0_123 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_123 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_529_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_124 <= 2'h0;
    end else if (bht_bank_sel_0_7_12) begin
      if (_T_7682) begin
        bht_bank_rd_data_out_0_124 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_124 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_529_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_125 <= 2'h0;
    end else if (bht_bank_sel_0_7_13) begin
      if (_T_7691) begin
        bht_bank_rd_data_out_0_125 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_125 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_529_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_126 <= 2'h0;
    end else if (bht_bank_sel_0_7_14) begin
      if (_T_7700) begin
        bht_bank_rd_data_out_0_126 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_126 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_529_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_127 <= 2'h0;
    end else if (bht_bank_sel_0_7_15) begin
      if (_T_7709) begin
        bht_bank_rd_data_out_0_127 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_127 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_530_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_128 <= 2'h0;
    end else if (bht_bank_sel_0_8_0) begin
      if (_T_7718) begin
        bht_bank_rd_data_out_0_128 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_128 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_530_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_129 <= 2'h0;
    end else if (bht_bank_sel_0_8_1) begin
      if (_T_7727) begin
        bht_bank_rd_data_out_0_129 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_129 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_530_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_130 <= 2'h0;
    end else if (bht_bank_sel_0_8_2) begin
      if (_T_7736) begin
        bht_bank_rd_data_out_0_130 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_130 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_530_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_131 <= 2'h0;
    end else if (bht_bank_sel_0_8_3) begin
      if (_T_7745) begin
        bht_bank_rd_data_out_0_131 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_131 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_530_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_132 <= 2'h0;
    end else if (bht_bank_sel_0_8_4) begin
      if (_T_7754) begin
        bht_bank_rd_data_out_0_132 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_132 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_530_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_133 <= 2'h0;
    end else if (bht_bank_sel_0_8_5) begin
      if (_T_7763) begin
        bht_bank_rd_data_out_0_133 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_133 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_530_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_134 <= 2'h0;
    end else if (bht_bank_sel_0_8_6) begin
      if (_T_7772) begin
        bht_bank_rd_data_out_0_134 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_134 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_530_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_135 <= 2'h0;
    end else if (bht_bank_sel_0_8_7) begin
      if (_T_7781) begin
        bht_bank_rd_data_out_0_135 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_135 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_530_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_136 <= 2'h0;
    end else if (bht_bank_sel_0_8_8) begin
      if (_T_7790) begin
        bht_bank_rd_data_out_0_136 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_136 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_530_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_137 <= 2'h0;
    end else if (bht_bank_sel_0_8_9) begin
      if (_T_7799) begin
        bht_bank_rd_data_out_0_137 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_137 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_530_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_138 <= 2'h0;
    end else if (bht_bank_sel_0_8_10) begin
      if (_T_7808) begin
        bht_bank_rd_data_out_0_138 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_138 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_530_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_139 <= 2'h0;
    end else if (bht_bank_sel_0_8_11) begin
      if (_T_7817) begin
        bht_bank_rd_data_out_0_139 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_139 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_530_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_140 <= 2'h0;
    end else if (bht_bank_sel_0_8_12) begin
      if (_T_7826) begin
        bht_bank_rd_data_out_0_140 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_140 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_530_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_141 <= 2'h0;
    end else if (bht_bank_sel_0_8_13) begin
      if (_T_7835) begin
        bht_bank_rd_data_out_0_141 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_141 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_530_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_142 <= 2'h0;
    end else if (bht_bank_sel_0_8_14) begin
      if (_T_7844) begin
        bht_bank_rd_data_out_0_142 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_142 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_530_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_143 <= 2'h0;
    end else if (bht_bank_sel_0_8_15) begin
      if (_T_7853) begin
        bht_bank_rd_data_out_0_143 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_143 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_531_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_144 <= 2'h0;
    end else if (bht_bank_sel_0_9_0) begin
      if (_T_7862) begin
        bht_bank_rd_data_out_0_144 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_144 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_531_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_145 <= 2'h0;
    end else if (bht_bank_sel_0_9_1) begin
      if (_T_7871) begin
        bht_bank_rd_data_out_0_145 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_145 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_531_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_146 <= 2'h0;
    end else if (bht_bank_sel_0_9_2) begin
      if (_T_7880) begin
        bht_bank_rd_data_out_0_146 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_146 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_531_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_147 <= 2'h0;
    end else if (bht_bank_sel_0_9_3) begin
      if (_T_7889) begin
        bht_bank_rd_data_out_0_147 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_147 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_531_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_148 <= 2'h0;
    end else if (bht_bank_sel_0_9_4) begin
      if (_T_7898) begin
        bht_bank_rd_data_out_0_148 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_148 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_531_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_149 <= 2'h0;
    end else if (bht_bank_sel_0_9_5) begin
      if (_T_7907) begin
        bht_bank_rd_data_out_0_149 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_149 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_531_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_150 <= 2'h0;
    end else if (bht_bank_sel_0_9_6) begin
      if (_T_7916) begin
        bht_bank_rd_data_out_0_150 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_150 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_531_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_151 <= 2'h0;
    end else if (bht_bank_sel_0_9_7) begin
      if (_T_7925) begin
        bht_bank_rd_data_out_0_151 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_151 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_531_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_152 <= 2'h0;
    end else if (bht_bank_sel_0_9_8) begin
      if (_T_7934) begin
        bht_bank_rd_data_out_0_152 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_152 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_531_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_153 <= 2'h0;
    end else if (bht_bank_sel_0_9_9) begin
      if (_T_7943) begin
        bht_bank_rd_data_out_0_153 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_153 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_531_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_154 <= 2'h0;
    end else if (bht_bank_sel_0_9_10) begin
      if (_T_7952) begin
        bht_bank_rd_data_out_0_154 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_154 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_531_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_155 <= 2'h0;
    end else if (bht_bank_sel_0_9_11) begin
      if (_T_7961) begin
        bht_bank_rd_data_out_0_155 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_155 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_531_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_156 <= 2'h0;
    end else if (bht_bank_sel_0_9_12) begin
      if (_T_7970) begin
        bht_bank_rd_data_out_0_156 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_156 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_531_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_157 <= 2'h0;
    end else if (bht_bank_sel_0_9_13) begin
      if (_T_7979) begin
        bht_bank_rd_data_out_0_157 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_157 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_531_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_158 <= 2'h0;
    end else if (bht_bank_sel_0_9_14) begin
      if (_T_7988) begin
        bht_bank_rd_data_out_0_158 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_158 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_531_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_159 <= 2'h0;
    end else if (bht_bank_sel_0_9_15) begin
      if (_T_7997) begin
        bht_bank_rd_data_out_0_159 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_159 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_532_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_160 <= 2'h0;
    end else if (bht_bank_sel_0_10_0) begin
      if (_T_8006) begin
        bht_bank_rd_data_out_0_160 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_160 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_532_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_161 <= 2'h0;
    end else if (bht_bank_sel_0_10_1) begin
      if (_T_8015) begin
        bht_bank_rd_data_out_0_161 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_161 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_532_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_162 <= 2'h0;
    end else if (bht_bank_sel_0_10_2) begin
      if (_T_8024) begin
        bht_bank_rd_data_out_0_162 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_162 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_532_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_163 <= 2'h0;
    end else if (bht_bank_sel_0_10_3) begin
      if (_T_8033) begin
        bht_bank_rd_data_out_0_163 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_163 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_532_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_164 <= 2'h0;
    end else if (bht_bank_sel_0_10_4) begin
      if (_T_8042) begin
        bht_bank_rd_data_out_0_164 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_164 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_532_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_165 <= 2'h0;
    end else if (bht_bank_sel_0_10_5) begin
      if (_T_8051) begin
        bht_bank_rd_data_out_0_165 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_165 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_532_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_166 <= 2'h0;
    end else if (bht_bank_sel_0_10_6) begin
      if (_T_8060) begin
        bht_bank_rd_data_out_0_166 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_166 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_532_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_167 <= 2'h0;
    end else if (bht_bank_sel_0_10_7) begin
      if (_T_8069) begin
        bht_bank_rd_data_out_0_167 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_167 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_532_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_168 <= 2'h0;
    end else if (bht_bank_sel_0_10_8) begin
      if (_T_8078) begin
        bht_bank_rd_data_out_0_168 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_168 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_532_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_169 <= 2'h0;
    end else if (bht_bank_sel_0_10_9) begin
      if (_T_8087) begin
        bht_bank_rd_data_out_0_169 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_169 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_532_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_170 <= 2'h0;
    end else if (bht_bank_sel_0_10_10) begin
      if (_T_8096) begin
        bht_bank_rd_data_out_0_170 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_170 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_532_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_171 <= 2'h0;
    end else if (bht_bank_sel_0_10_11) begin
      if (_T_8105) begin
        bht_bank_rd_data_out_0_171 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_171 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_532_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_172 <= 2'h0;
    end else if (bht_bank_sel_0_10_12) begin
      if (_T_8114) begin
        bht_bank_rd_data_out_0_172 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_172 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_532_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_173 <= 2'h0;
    end else if (bht_bank_sel_0_10_13) begin
      if (_T_8123) begin
        bht_bank_rd_data_out_0_173 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_173 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_532_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_174 <= 2'h0;
    end else if (bht_bank_sel_0_10_14) begin
      if (_T_8132) begin
        bht_bank_rd_data_out_0_174 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_174 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_532_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_175 <= 2'h0;
    end else if (bht_bank_sel_0_10_15) begin
      if (_T_8141) begin
        bht_bank_rd_data_out_0_175 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_175 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_533_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_176 <= 2'h0;
    end else if (bht_bank_sel_0_11_0) begin
      if (_T_8150) begin
        bht_bank_rd_data_out_0_176 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_176 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_533_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_177 <= 2'h0;
    end else if (bht_bank_sel_0_11_1) begin
      if (_T_8159) begin
        bht_bank_rd_data_out_0_177 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_177 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_533_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_178 <= 2'h0;
    end else if (bht_bank_sel_0_11_2) begin
      if (_T_8168) begin
        bht_bank_rd_data_out_0_178 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_178 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_533_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_179 <= 2'h0;
    end else if (bht_bank_sel_0_11_3) begin
      if (_T_8177) begin
        bht_bank_rd_data_out_0_179 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_179 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_533_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_180 <= 2'h0;
    end else if (bht_bank_sel_0_11_4) begin
      if (_T_8186) begin
        bht_bank_rd_data_out_0_180 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_180 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_533_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_181 <= 2'h0;
    end else if (bht_bank_sel_0_11_5) begin
      if (_T_8195) begin
        bht_bank_rd_data_out_0_181 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_181 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_533_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_182 <= 2'h0;
    end else if (bht_bank_sel_0_11_6) begin
      if (_T_8204) begin
        bht_bank_rd_data_out_0_182 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_182 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_533_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_183 <= 2'h0;
    end else if (bht_bank_sel_0_11_7) begin
      if (_T_8213) begin
        bht_bank_rd_data_out_0_183 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_183 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_533_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_184 <= 2'h0;
    end else if (bht_bank_sel_0_11_8) begin
      if (_T_8222) begin
        bht_bank_rd_data_out_0_184 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_184 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_533_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_185 <= 2'h0;
    end else if (bht_bank_sel_0_11_9) begin
      if (_T_8231) begin
        bht_bank_rd_data_out_0_185 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_185 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_533_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_186 <= 2'h0;
    end else if (bht_bank_sel_0_11_10) begin
      if (_T_8240) begin
        bht_bank_rd_data_out_0_186 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_186 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_533_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_187 <= 2'h0;
    end else if (bht_bank_sel_0_11_11) begin
      if (_T_8249) begin
        bht_bank_rd_data_out_0_187 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_187 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_533_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_188 <= 2'h0;
    end else if (bht_bank_sel_0_11_12) begin
      if (_T_8258) begin
        bht_bank_rd_data_out_0_188 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_188 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_533_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_189 <= 2'h0;
    end else if (bht_bank_sel_0_11_13) begin
      if (_T_8267) begin
        bht_bank_rd_data_out_0_189 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_189 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_533_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_190 <= 2'h0;
    end else if (bht_bank_sel_0_11_14) begin
      if (_T_8276) begin
        bht_bank_rd_data_out_0_190 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_190 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_533_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_191 <= 2'h0;
    end else if (bht_bank_sel_0_11_15) begin
      if (_T_8285) begin
        bht_bank_rd_data_out_0_191 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_191 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_534_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_192 <= 2'h0;
    end else if (bht_bank_sel_0_12_0) begin
      if (_T_8294) begin
        bht_bank_rd_data_out_0_192 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_192 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_534_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_193 <= 2'h0;
    end else if (bht_bank_sel_0_12_1) begin
      if (_T_8303) begin
        bht_bank_rd_data_out_0_193 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_193 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_534_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_194 <= 2'h0;
    end else if (bht_bank_sel_0_12_2) begin
      if (_T_8312) begin
        bht_bank_rd_data_out_0_194 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_194 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_534_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_195 <= 2'h0;
    end else if (bht_bank_sel_0_12_3) begin
      if (_T_8321) begin
        bht_bank_rd_data_out_0_195 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_195 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_534_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_196 <= 2'h0;
    end else if (bht_bank_sel_0_12_4) begin
      if (_T_8330) begin
        bht_bank_rd_data_out_0_196 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_196 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_534_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_197 <= 2'h0;
    end else if (bht_bank_sel_0_12_5) begin
      if (_T_8339) begin
        bht_bank_rd_data_out_0_197 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_197 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_534_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_198 <= 2'h0;
    end else if (bht_bank_sel_0_12_6) begin
      if (_T_8348) begin
        bht_bank_rd_data_out_0_198 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_198 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_534_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_199 <= 2'h0;
    end else if (bht_bank_sel_0_12_7) begin
      if (_T_8357) begin
        bht_bank_rd_data_out_0_199 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_199 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_534_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_200 <= 2'h0;
    end else if (bht_bank_sel_0_12_8) begin
      if (_T_8366) begin
        bht_bank_rd_data_out_0_200 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_200 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_534_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_201 <= 2'h0;
    end else if (bht_bank_sel_0_12_9) begin
      if (_T_8375) begin
        bht_bank_rd_data_out_0_201 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_201 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_534_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_202 <= 2'h0;
    end else if (bht_bank_sel_0_12_10) begin
      if (_T_8384) begin
        bht_bank_rd_data_out_0_202 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_202 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_534_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_203 <= 2'h0;
    end else if (bht_bank_sel_0_12_11) begin
      if (_T_8393) begin
        bht_bank_rd_data_out_0_203 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_203 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_534_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_204 <= 2'h0;
    end else if (bht_bank_sel_0_12_12) begin
      if (_T_8402) begin
        bht_bank_rd_data_out_0_204 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_204 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_534_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_205 <= 2'h0;
    end else if (bht_bank_sel_0_12_13) begin
      if (_T_8411) begin
        bht_bank_rd_data_out_0_205 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_205 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_534_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_206 <= 2'h0;
    end else if (bht_bank_sel_0_12_14) begin
      if (_T_8420) begin
        bht_bank_rd_data_out_0_206 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_206 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_534_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_207 <= 2'h0;
    end else if (bht_bank_sel_0_12_15) begin
      if (_T_8429) begin
        bht_bank_rd_data_out_0_207 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_207 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_535_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_208 <= 2'h0;
    end else if (bht_bank_sel_0_13_0) begin
      if (_T_8438) begin
        bht_bank_rd_data_out_0_208 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_208 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_535_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_209 <= 2'h0;
    end else if (bht_bank_sel_0_13_1) begin
      if (_T_8447) begin
        bht_bank_rd_data_out_0_209 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_209 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_535_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_210 <= 2'h0;
    end else if (bht_bank_sel_0_13_2) begin
      if (_T_8456) begin
        bht_bank_rd_data_out_0_210 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_210 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_535_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_211 <= 2'h0;
    end else if (bht_bank_sel_0_13_3) begin
      if (_T_8465) begin
        bht_bank_rd_data_out_0_211 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_211 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_535_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_212 <= 2'h0;
    end else if (bht_bank_sel_0_13_4) begin
      if (_T_8474) begin
        bht_bank_rd_data_out_0_212 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_212 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_535_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_213 <= 2'h0;
    end else if (bht_bank_sel_0_13_5) begin
      if (_T_8483) begin
        bht_bank_rd_data_out_0_213 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_213 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_535_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_214 <= 2'h0;
    end else if (bht_bank_sel_0_13_6) begin
      if (_T_8492) begin
        bht_bank_rd_data_out_0_214 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_214 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_535_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_215 <= 2'h0;
    end else if (bht_bank_sel_0_13_7) begin
      if (_T_8501) begin
        bht_bank_rd_data_out_0_215 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_215 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_535_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_216 <= 2'h0;
    end else if (bht_bank_sel_0_13_8) begin
      if (_T_8510) begin
        bht_bank_rd_data_out_0_216 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_216 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_535_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_217 <= 2'h0;
    end else if (bht_bank_sel_0_13_9) begin
      if (_T_8519) begin
        bht_bank_rd_data_out_0_217 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_217 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_535_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_218 <= 2'h0;
    end else if (bht_bank_sel_0_13_10) begin
      if (_T_8528) begin
        bht_bank_rd_data_out_0_218 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_218 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_535_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_219 <= 2'h0;
    end else if (bht_bank_sel_0_13_11) begin
      if (_T_8537) begin
        bht_bank_rd_data_out_0_219 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_219 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_535_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_220 <= 2'h0;
    end else if (bht_bank_sel_0_13_12) begin
      if (_T_8546) begin
        bht_bank_rd_data_out_0_220 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_220 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_535_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_221 <= 2'h0;
    end else if (bht_bank_sel_0_13_13) begin
      if (_T_8555) begin
        bht_bank_rd_data_out_0_221 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_221 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_535_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_222 <= 2'h0;
    end else if (bht_bank_sel_0_13_14) begin
      if (_T_8564) begin
        bht_bank_rd_data_out_0_222 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_222 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_535_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_223 <= 2'h0;
    end else if (bht_bank_sel_0_13_15) begin
      if (_T_8573) begin
        bht_bank_rd_data_out_0_223 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_223 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_536_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_224 <= 2'h0;
    end else if (bht_bank_sel_0_14_0) begin
      if (_T_8582) begin
        bht_bank_rd_data_out_0_224 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_224 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_536_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_225 <= 2'h0;
    end else if (bht_bank_sel_0_14_1) begin
      if (_T_8591) begin
        bht_bank_rd_data_out_0_225 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_225 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_536_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_226 <= 2'h0;
    end else if (bht_bank_sel_0_14_2) begin
      if (_T_8600) begin
        bht_bank_rd_data_out_0_226 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_226 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_536_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_227 <= 2'h0;
    end else if (bht_bank_sel_0_14_3) begin
      if (_T_8609) begin
        bht_bank_rd_data_out_0_227 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_227 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_536_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_228 <= 2'h0;
    end else if (bht_bank_sel_0_14_4) begin
      if (_T_8618) begin
        bht_bank_rd_data_out_0_228 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_228 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_536_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_229 <= 2'h0;
    end else if (bht_bank_sel_0_14_5) begin
      if (_T_8627) begin
        bht_bank_rd_data_out_0_229 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_229 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_536_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_230 <= 2'h0;
    end else if (bht_bank_sel_0_14_6) begin
      if (_T_8636) begin
        bht_bank_rd_data_out_0_230 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_230 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_536_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_231 <= 2'h0;
    end else if (bht_bank_sel_0_14_7) begin
      if (_T_8645) begin
        bht_bank_rd_data_out_0_231 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_231 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_536_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_232 <= 2'h0;
    end else if (bht_bank_sel_0_14_8) begin
      if (_T_8654) begin
        bht_bank_rd_data_out_0_232 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_232 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_536_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_233 <= 2'h0;
    end else if (bht_bank_sel_0_14_9) begin
      if (_T_8663) begin
        bht_bank_rd_data_out_0_233 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_233 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_536_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_234 <= 2'h0;
    end else if (bht_bank_sel_0_14_10) begin
      if (_T_8672) begin
        bht_bank_rd_data_out_0_234 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_234 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_536_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_235 <= 2'h0;
    end else if (bht_bank_sel_0_14_11) begin
      if (_T_8681) begin
        bht_bank_rd_data_out_0_235 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_235 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_536_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_236 <= 2'h0;
    end else if (bht_bank_sel_0_14_12) begin
      if (_T_8690) begin
        bht_bank_rd_data_out_0_236 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_236 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_536_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_237 <= 2'h0;
    end else if (bht_bank_sel_0_14_13) begin
      if (_T_8699) begin
        bht_bank_rd_data_out_0_237 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_237 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_536_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_238 <= 2'h0;
    end else if (bht_bank_sel_0_14_14) begin
      if (_T_8708) begin
        bht_bank_rd_data_out_0_238 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_238 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_536_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_239 <= 2'h0;
    end else if (bht_bank_sel_0_14_15) begin
      if (_T_8717) begin
        bht_bank_rd_data_out_0_239 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_239 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_537_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_240 <= 2'h0;
    end else if (bht_bank_sel_0_15_0) begin
      if (_T_8726) begin
        bht_bank_rd_data_out_0_240 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_240 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_537_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_241 <= 2'h0;
    end else if (bht_bank_sel_0_15_1) begin
      if (_T_8735) begin
        bht_bank_rd_data_out_0_241 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_241 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_537_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_242 <= 2'h0;
    end else if (bht_bank_sel_0_15_2) begin
      if (_T_8744) begin
        bht_bank_rd_data_out_0_242 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_242 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_537_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_243 <= 2'h0;
    end else if (bht_bank_sel_0_15_3) begin
      if (_T_8753) begin
        bht_bank_rd_data_out_0_243 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_243 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_537_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_244 <= 2'h0;
    end else if (bht_bank_sel_0_15_4) begin
      if (_T_8762) begin
        bht_bank_rd_data_out_0_244 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_244 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_537_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_245 <= 2'h0;
    end else if (bht_bank_sel_0_15_5) begin
      if (_T_8771) begin
        bht_bank_rd_data_out_0_245 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_245 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_537_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_246 <= 2'h0;
    end else if (bht_bank_sel_0_15_6) begin
      if (_T_8780) begin
        bht_bank_rd_data_out_0_246 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_246 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_537_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_247 <= 2'h0;
    end else if (bht_bank_sel_0_15_7) begin
      if (_T_8789) begin
        bht_bank_rd_data_out_0_247 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_247 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_537_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_248 <= 2'h0;
    end else if (bht_bank_sel_0_15_8) begin
      if (_T_8798) begin
        bht_bank_rd_data_out_0_248 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_248 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_537_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_249 <= 2'h0;
    end else if (bht_bank_sel_0_15_9) begin
      if (_T_8807) begin
        bht_bank_rd_data_out_0_249 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_249 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_537_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_250 <= 2'h0;
    end else if (bht_bank_sel_0_15_10) begin
      if (_T_8816) begin
        bht_bank_rd_data_out_0_250 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_250 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_537_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_251 <= 2'h0;
    end else if (bht_bank_sel_0_15_11) begin
      if (_T_8825) begin
        bht_bank_rd_data_out_0_251 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_251 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_537_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_252 <= 2'h0;
    end else if (bht_bank_sel_0_15_12) begin
      if (_T_8834) begin
        bht_bank_rd_data_out_0_252 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_252 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_537_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_253 <= 2'h0;
    end else if (bht_bank_sel_0_15_13) begin
      if (_T_8843) begin
        bht_bank_rd_data_out_0_253 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_253 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_537_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_254 <= 2'h0;
    end else if (bht_bank_sel_0_15_14) begin
      if (_T_8852) begin
        bht_bank_rd_data_out_0_254 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_254 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge rvclkhdr_537_io_l1clk or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_255 <= 2'h0;
    end else if (bht_bank_sel_0_15_15) begin
      if (_T_8861) begin
        bht_bank_rd_data_out_0_255 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_255 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      exu_mp_way_f <= 1'h0;
    end else begin
      exu_mp_way_f <= io_exu_bp_exu_mp_pkt_bits_way;
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      exu_flush_final_d1 <= 1'h0;
    end else begin
      exu_flush_final_d1 <= io_exu_flush_final;
    end
  end
  always @(posedge rvclkhdr_io_l1clk or posedge reset) begin
    if (reset) begin
      btb_lru_b0_f <= 256'h0;
    end else begin
      btb_lru_b0_f <= _T_183 | _T_185;
    end
  end
  always @(posedge rvclkhdr_1_io_l1clk or posedge reset) begin
    if (reset) begin
      ifc_fetch_adder_prior <= 30'h0;
    end else begin
      ifc_fetch_adder_prior <= io_ifc_fetch_addr_f[30:1];
    end
  end
  always @(posedge rvclkhdr_2_io_l1clk or posedge reset) begin
    if (reset) begin
      rets_out_0 <= 32'h0;
    end else begin
      rets_out_0 <= _T_482 | _T_483;
    end
  end
  always @(posedge rvclkhdr_3_io_l1clk or posedge reset) begin
    if (reset) begin
      rets_out_1 <= 32'h0;
    end else begin
      rets_out_1 <= _T_487 | _T_488;
    end
  end
  always @(posedge rvclkhdr_4_io_l1clk or posedge reset) begin
    if (reset) begin
      rets_out_2 <= 32'h0;
    end else begin
      rets_out_2 <= _T_492 | _T_493;
    end
  end
  always @(posedge rvclkhdr_5_io_l1clk or posedge reset) begin
    if (reset) begin
      rets_out_3 <= 32'h0;
    end else begin
      rets_out_3 <= _T_497 | _T_498;
    end
  end
  always @(posedge rvclkhdr_6_io_l1clk or posedge reset) begin
    if (reset) begin
      rets_out_4 <= 32'h0;
    end else begin
      rets_out_4 <= _T_502 | _T_503;
    end
  end
  always @(posedge rvclkhdr_7_io_l1clk or posedge reset) begin
    if (reset) begin
      rets_out_5 <= 32'h0;
    end else begin
      rets_out_5 <= _T_507 | _T_508;
    end
  end
  always @(posedge rvclkhdr_8_io_l1clk or posedge reset) begin
    if (reset) begin
      rets_out_6 <= 32'h0;
    end else begin
      rets_out_6 <= _T_512 | _T_513;
    end
  end
  always @(posedge rvclkhdr_9_io_l1clk or posedge reset) begin
    if (reset) begin
      rets_out_7 <= 32'h0;
    end else begin
      rets_out_7 <= rets_out_6;
    end
  end
endmodule
module ifu_compress_ctl(
  input  [15:0] io_din,
  output [31:0] io_dout
);
  wire  _T_2 = ~io_din[14]; // @[ifu_compress_ctl.scala 12:83]
  wire  _T_4 = ~io_din[13]; // @[ifu_compress_ctl.scala 12:83]
  wire  _T_7 = ~io_din[6]; // @[ifu_compress_ctl.scala 12:83]
  wire  _T_9 = ~io_din[5]; // @[ifu_compress_ctl.scala 12:83]
  wire  _T_11 = io_din[15] & _T_2; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_12 = _T_11 & _T_4; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_13 = _T_12 & io_din[10]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_14 = _T_13 & _T_7; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_15 = _T_14 & _T_9; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_16 = _T_15 & io_din[0]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_23 = ~io_din[11]; // @[ifu_compress_ctl.scala 12:83]
  wire  _T_28 = _T_12 & _T_23; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_29 = _T_28 & io_din[10]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_30 = _T_29 & io_din[0]; // @[ifu_compress_ctl.scala 12:110]
  wire  out_30 = _T_16 | _T_30; // @[ifu_compress_ctl.scala 17:53]
  wire  _T_38 = ~io_din[10]; // @[ifu_compress_ctl.scala 12:83]
  wire  _T_40 = ~io_din[9]; // @[ifu_compress_ctl.scala 12:83]
  wire  _T_42 = ~io_din[8]; // @[ifu_compress_ctl.scala 12:83]
  wire  _T_44 = ~io_din[7]; // @[ifu_compress_ctl.scala 12:83]
  wire  _T_50 = ~io_din[4]; // @[ifu_compress_ctl.scala 12:83]
  wire  _T_52 = ~io_din[3]; // @[ifu_compress_ctl.scala 12:83]
  wire  _T_54 = ~io_din[2]; // @[ifu_compress_ctl.scala 12:83]
  wire  _T_56 = _T_2 & io_din[12]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_57 = _T_56 & _T_23; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_58 = _T_57 & _T_38; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_59 = _T_58 & _T_40; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_60 = _T_59 & _T_42; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_61 = _T_60 & _T_44; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_62 = _T_61 & _T_7; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_63 = _T_62 & _T_9; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_64 = _T_63 & _T_50; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_65 = _T_64 & _T_52; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_66 = _T_65 & _T_54; // @[ifu_compress_ctl.scala 12:110]
  wire  out_20 = _T_66 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_79 = _T_28 & io_din[0]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_90 = _T_12 & _T_38; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_91 = _T_90 & io_din[0]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_92 = _T_79 | _T_91; // @[ifu_compress_ctl.scala 21:46]
  wire  _T_102 = _T_12 & io_din[6]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_103 = _T_102 & io_din[0]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_104 = _T_92 | _T_103; // @[ifu_compress_ctl.scala 21:80]
  wire  _T_114 = _T_12 & io_din[5]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_115 = _T_114 & io_din[0]; // @[ifu_compress_ctl.scala 12:110]
  wire  out_14 = _T_104 | _T_115; // @[ifu_compress_ctl.scala 21:113]
  wire  _T_128 = _T_12 & io_din[11]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_129 = _T_128 & _T_38; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_130 = _T_129 & io_din[0]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_142 = _T_128 & io_din[6]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_143 = _T_142 & io_din[0]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_144 = _T_130 | _T_143; // @[ifu_compress_ctl.scala 23:50]
  wire  _T_147 = ~io_din[0]; // @[ifu_compress_ctl.scala 23:101]
  wire  _T_148 = io_din[14] & _T_147; // @[ifu_compress_ctl.scala 23:99]
  wire  out_13 = _T_144 | _T_148; // @[ifu_compress_ctl.scala 23:86]
  wire  _T_161 = _T_102 & io_din[5]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_162 = _T_161 & io_din[0]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_175 = _T_162 | _T_79; // @[ifu_compress_ctl.scala 25:47]
  wire  _T_188 = _T_175 | _T_91; // @[ifu_compress_ctl.scala 25:81]
  wire  _T_190 = ~io_din[15]; // @[ifu_compress_ctl.scala 12:83]
  wire  _T_194 = _T_190 & _T_2; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_195 = _T_194 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_196 = _T_188 | _T_195; // @[ifu_compress_ctl.scala 25:115]
  wire  _T_200 = io_din[15] & io_din[14]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_201 = _T_200 & io_din[13]; // @[ifu_compress_ctl.scala 12:110]
  wire  out_12 = _T_196 | _T_201; // @[ifu_compress_ctl.scala 26:26]
  wire  _T_217 = _T_11 & _T_7; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_218 = _T_217 & _T_9; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_219 = _T_218 & _T_50; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_220 = _T_219 & _T_52; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_221 = _T_220 & _T_54; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_224 = _T_221 & _T_147; // @[ifu_compress_ctl.scala 28:53]
  wire  _T_228 = _T_2 & io_din[13]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_229 = _T_224 | _T_228; // @[ifu_compress_ctl.scala 28:67]
  wire  _T_234 = _T_200 & io_din[0]; // @[ifu_compress_ctl.scala 12:110]
  wire  out_6 = _T_229 | _T_234; // @[ifu_compress_ctl.scala 28:88]
  wire  _T_239 = io_din[15] & _T_147; // @[ifu_compress_ctl.scala 30:24]
  wire  _T_243 = io_din[15] & io_din[11]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_244 = _T_243 & io_din[10]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_245 = _T_239 | _T_244; // @[ifu_compress_ctl.scala 30:39]
  wire  _T_249 = io_din[13] & _T_42; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_250 = _T_245 | _T_249; // @[ifu_compress_ctl.scala 30:63]
  wire  _T_253 = io_din[13] & io_din[7]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_254 = _T_250 | _T_253; // @[ifu_compress_ctl.scala 30:83]
  wire  _T_257 = io_din[13] & io_din[9]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_258 = _T_254 | _T_257; // @[ifu_compress_ctl.scala 30:102]
  wire  _T_261 = io_din[13] & io_din[10]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_262 = _T_258 | _T_261; // @[ifu_compress_ctl.scala 31:22]
  wire  _T_265 = io_din[13] & io_din[11]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_266 = _T_262 | _T_265; // @[ifu_compress_ctl.scala 31:42]
  wire  _T_271 = _T_266 | _T_228; // @[ifu_compress_ctl.scala 31:62]
  wire  out_5 = _T_271 | _T_200; // @[ifu_compress_ctl.scala 31:83]
  wire  _T_288 = _T_2 & _T_23; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_289 = _T_288 & _T_38; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_290 = _T_289 & _T_40; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_291 = _T_290 & _T_42; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_292 = _T_291 & _T_44; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_295 = _T_292 & _T_147; // @[ifu_compress_ctl.scala 33:50]
  wire  _T_303 = _T_194 & _T_147; // @[ifu_compress_ctl.scala 33:87]
  wire  _T_304 = _T_295 | _T_303; // @[ifu_compress_ctl.scala 33:65]
  wire  _T_308 = _T_2 & io_din[6]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_311 = _T_308 & _T_147; // @[ifu_compress_ctl.scala 34:23]
  wire  _T_312 = _T_304 | _T_311; // @[ifu_compress_ctl.scala 33:102]
  wire  _T_317 = _T_190 & io_din[14]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_318 = _T_317 & io_din[0]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_319 = _T_312 | _T_318; // @[ifu_compress_ctl.scala 34:38]
  wire  _T_323 = _T_2 & io_din[5]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_326 = _T_323 & _T_147; // @[ifu_compress_ctl.scala 34:82]
  wire  _T_327 = _T_319 | _T_326; // @[ifu_compress_ctl.scala 34:62]
  wire  _T_331 = _T_2 & io_din[4]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_334 = _T_331 & _T_147; // @[ifu_compress_ctl.scala 35:23]
  wire  _T_335 = _T_327 | _T_334; // @[ifu_compress_ctl.scala 34:97]
  wire  _T_339 = _T_2 & io_din[3]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_342 = _T_339 & _T_147; // @[ifu_compress_ctl.scala 35:58]
  wire  _T_343 = _T_335 | _T_342; // @[ifu_compress_ctl.scala 35:38]
  wire  _T_347 = _T_2 & io_din[2]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_350 = _T_347 & _T_147; // @[ifu_compress_ctl.scala 35:93]
  wire  _T_351 = _T_343 | _T_350; // @[ifu_compress_ctl.scala 35:73]
  wire  _T_357 = _T_2 & _T_4; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_358 = _T_357 & io_din[0]; // @[ifu_compress_ctl.scala 12:110]
  wire  out_4 = _T_351 | _T_358; // @[ifu_compress_ctl.scala 35:108]
  wire  _T_380 = _T_56 & io_din[11]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_381 = _T_380 & _T_7; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_382 = _T_381 & _T_9; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_383 = _T_382 & _T_50; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_384 = _T_383 & _T_52; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_385 = _T_384 & _T_54; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_386 = _T_385 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_403 = _T_56 & io_din[10]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_404 = _T_403 & _T_7; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_405 = _T_404 & _T_9; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_406 = _T_405 & _T_50; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_407 = _T_406 & _T_52; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_408 = _T_407 & _T_54; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_409 = _T_408 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_410 = _T_386 | _T_409; // @[ifu_compress_ctl.scala 40:59]
  wire  _T_427 = _T_56 & io_din[9]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_428 = _T_427 & _T_7; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_429 = _T_428 & _T_9; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_430 = _T_429 & _T_50; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_431 = _T_430 & _T_52; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_432 = _T_431 & _T_54; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_433 = _T_432 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_434 = _T_410 | _T_433; // @[ifu_compress_ctl.scala 40:107]
  wire  _T_451 = _T_56 & io_din[8]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_452 = _T_451 & _T_7; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_453 = _T_452 & _T_9; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_454 = _T_453 & _T_50; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_455 = _T_454 & _T_52; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_456 = _T_455 & _T_54; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_457 = _T_456 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_458 = _T_434 | _T_457; // @[ifu_compress_ctl.scala 41:50]
  wire  _T_475 = _T_56 & io_din[7]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_476 = _T_475 & _T_7; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_477 = _T_476 & _T_9; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_478 = _T_477 & _T_50; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_479 = _T_478 & _T_52; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_480 = _T_479 & _T_54; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_481 = _T_480 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_482 = _T_458 | _T_481; // @[ifu_compress_ctl.scala 41:94]
  wire  _T_487 = ~io_din[12]; // @[ifu_compress_ctl.scala 12:83]
  wire  _T_499 = _T_11 & _T_487; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_500 = _T_499 & _T_7; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_501 = _T_500 & _T_9; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_502 = _T_501 & _T_50; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_503 = _T_502 & _T_52; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_504 = _T_503 & _T_54; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_507 = _T_504 & _T_147; // @[ifu_compress_ctl.scala 42:94]
  wire  _T_508 = _T_482 | _T_507; // @[ifu_compress_ctl.scala 42:49]
  wire  _T_514 = _T_190 & io_din[13]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_515 = _T_514 & _T_42; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_516 = _T_508 | _T_515; // @[ifu_compress_ctl.scala 42:109]
  wire  _T_522 = _T_514 & io_din[7]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_523 = _T_516 | _T_522; // @[ifu_compress_ctl.scala 43:26]
  wire  _T_529 = _T_514 & io_din[9]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_530 = _T_523 | _T_529; // @[ifu_compress_ctl.scala 43:48]
  wire  _T_536 = _T_514 & io_din[10]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_537 = _T_530 | _T_536; // @[ifu_compress_ctl.scala 43:70]
  wire  _T_543 = _T_514 & io_din[11]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_544 = _T_537 | _T_543; // @[ifu_compress_ctl.scala 43:93]
  wire  out_2 = _T_544 | _T_228; // @[ifu_compress_ctl.scala 44:26]
  wire [4:0] rs2d = io_din[6:2]; // @[ifu_compress_ctl.scala 50:20]
  wire [4:0] rdd = io_din[11:7]; // @[ifu_compress_ctl.scala 51:19]
  wire [4:0] rdpd = {2'h1,io_din[9:7]}; // @[Cat.scala 29:58]
  wire [4:0] rs2pd = {2'h1,io_din[4:2]}; // @[Cat.scala 29:58]
  wire  _T_557 = _T_308 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_564 = _T_317 & io_din[11]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_565 = _T_564 & io_din[0]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_566 = _T_557 | _T_565; // @[ifu_compress_ctl.scala 55:33]
  wire  _T_572 = _T_323 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_573 = _T_566 | _T_572; // @[ifu_compress_ctl.scala 55:58]
  wire  _T_580 = _T_317 & io_din[10]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_581 = _T_580 & io_din[0]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_582 = _T_573 | _T_581; // @[ifu_compress_ctl.scala 55:79]
  wire  _T_588 = _T_331 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_589 = _T_582 | _T_588; // @[ifu_compress_ctl.scala 55:104]
  wire  _T_596 = _T_317 & io_din[9]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_597 = _T_596 & io_din[0]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_598 = _T_589 | _T_597; // @[ifu_compress_ctl.scala 56:24]
  wire  _T_604 = _T_339 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_605 = _T_598 | _T_604; // @[ifu_compress_ctl.scala 56:48]
  wire  _T_613 = _T_317 & _T_42; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_614 = _T_613 & io_din[0]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_615 = _T_605 | _T_614; // @[ifu_compress_ctl.scala 56:69]
  wire  _T_621 = _T_347 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_622 = _T_615 | _T_621; // @[ifu_compress_ctl.scala 56:94]
  wire  _T_629 = _T_317 & io_din[7]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_630 = _T_629 & io_din[0]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_631 = _T_622 | _T_630; // @[ifu_compress_ctl.scala 57:22]
  wire  _T_635 = _T_190 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_636 = _T_631 | _T_635; // @[ifu_compress_ctl.scala 57:46]
  wire  _T_642 = _T_190 & _T_4; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_643 = _T_642 & io_din[0]; // @[ifu_compress_ctl.scala 12:110]
  wire  rdrd = _T_636 | _T_643; // @[ifu_compress_ctl.scala 57:65]
  wire  _T_651 = _T_380 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_659 = _T_403 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_660 = _T_651 | _T_659; // @[ifu_compress_ctl.scala 59:38]
  wire  _T_668 = _T_427 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_669 = _T_660 | _T_668; // @[ifu_compress_ctl.scala 59:63]
  wire  _T_677 = _T_451 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_678 = _T_669 | _T_677; // @[ifu_compress_ctl.scala 59:87]
  wire  _T_686 = _T_475 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_687 = _T_678 | _T_686; // @[ifu_compress_ctl.scala 60:27]
  wire  _T_703 = _T_2 & _T_487; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_704 = _T_703 & _T_7; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_705 = _T_704 & _T_9; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_706 = _T_705 & _T_50; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_707 = _T_706 & _T_52; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_708 = _T_707 & _T_54; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_709 = _T_708 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_710 = _T_687 | _T_709; // @[ifu_compress_ctl.scala 60:51]
  wire  _T_717 = _T_56 & io_din[6]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_718 = _T_717 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_719 = _T_710 | _T_718; // @[ifu_compress_ctl.scala 60:89]
  wire  _T_726 = _T_56 & io_din[5]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_727 = _T_726 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_728 = _T_719 | _T_727; // @[ifu_compress_ctl.scala 61:27]
  wire  _T_735 = _T_56 & io_din[4]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_736 = _T_735 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_737 = _T_728 | _T_736; // @[ifu_compress_ctl.scala 61:51]
  wire  _T_744 = _T_56 & io_din[3]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_745 = _T_744 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_746 = _T_737 | _T_745; // @[ifu_compress_ctl.scala 61:75]
  wire  _T_753 = _T_56 & io_din[2]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_754 = _T_753 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_755 = _T_746 | _T_754; // @[ifu_compress_ctl.scala 61:99]
  wire  _T_764 = _T_194 & _T_4; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_765 = _T_764 & io_din[0]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_766 = _T_755 | _T_765; // @[ifu_compress_ctl.scala 62:27]
  wire  rdrs1 = _T_766 | _T_195; // @[ifu_compress_ctl.scala 62:54]
  wire  _T_777 = io_din[15] & io_din[6]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_778 = _T_777 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_782 = io_din[15] & io_din[5]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_783 = _T_782 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_784 = _T_778 | _T_783; // @[ifu_compress_ctl.scala 64:34]
  wire  _T_788 = io_din[15] & io_din[4]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_789 = _T_788 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_790 = _T_784 | _T_789; // @[ifu_compress_ctl.scala 64:54]
  wire  _T_794 = io_din[15] & io_din[3]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_795 = _T_794 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_796 = _T_790 | _T_795; // @[ifu_compress_ctl.scala 64:74]
  wire  _T_800 = io_din[15] & io_din[2]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_801 = _T_800 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_802 = _T_796 | _T_801; // @[ifu_compress_ctl.scala 64:94]
  wire  _T_807 = _T_200 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  rs2rs2 = _T_802 | _T_807; // @[ifu_compress_ctl.scala 64:114]
  wire  rdprd = _T_12 & io_din[0]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_820 = io_din[15] & _T_4; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_821 = _T_820 & io_din[0]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_827 = _T_821 | _T_234; // @[ifu_compress_ctl.scala 68:36]
  wire  _T_830 = ~io_din[1]; // @[ifu_compress_ctl.scala 12:83]
  wire  _T_831 = io_din[14] & _T_830; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_834 = _T_831 & _T_147; // @[ifu_compress_ctl.scala 68:76]
  wire  rdprs1 = _T_827 | _T_834; // @[ifu_compress_ctl.scala 68:57]
  wire  _T_846 = _T_128 & io_din[10]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_847 = _T_846 & io_din[0]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_851 = io_din[15] & _T_830; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_854 = _T_851 & _T_147; // @[ifu_compress_ctl.scala 70:66]
  wire  rs2prs2 = _T_847 | _T_854; // @[ifu_compress_ctl.scala 70:47]
  wire  _T_859 = _T_190 & _T_830; // @[ifu_compress_ctl.scala 12:110]
  wire  rs2prd = _T_859 & _T_147; // @[ifu_compress_ctl.scala 72:33]
  wire  _T_866 = _T_2 & _T_830; // @[ifu_compress_ctl.scala 12:110]
  wire  uimm9_2 = _T_866 & _T_147; // @[ifu_compress_ctl.scala 74:34]
  wire  _T_875 = _T_317 & _T_830; // @[ifu_compress_ctl.scala 12:110]
  wire  ulwimm6_2 = _T_875 & _T_147; // @[ifu_compress_ctl.scala 76:39]
  wire  ulwspimm7_2 = _T_317 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_897 = _T_317 & io_din[13]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_898 = _T_897 & _T_23; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_899 = _T_898 & _T_38; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_900 = _T_899 & _T_40; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_901 = _T_900 & io_din[8]; // @[ifu_compress_ctl.scala 12:110]
  wire  rdeq2 = _T_901 & _T_44; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1027 = _T_194 & io_din[13]; // @[ifu_compress_ctl.scala 12:110]
  wire  rdeq1 = _T_482 | _T_1027; // @[ifu_compress_ctl.scala 84:42]
  wire  _T_1050 = io_din[14] & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1051 = rdeq2 | _T_1050; // @[ifu_compress_ctl.scala 86:53]
  wire  rs1eq2 = _T_1051 | uimm9_2; // @[ifu_compress_ctl.scala 86:71]
  wire  _T_1092 = _T_357 & io_din[11]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1093 = _T_1092 & _T_38; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1094 = _T_1093 & io_din[0]; // @[ifu_compress_ctl.scala 12:110]
  wire  simm5_0 = _T_1094 | _T_643; // @[ifu_compress_ctl.scala 92:45]
  wire  _T_1112 = _T_897 & io_din[7]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1121 = _T_897 & _T_42; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1122 = _T_1112 | _T_1121; // @[ifu_compress_ctl.scala 96:44]
  wire  _T_1130 = _T_897 & io_din[9]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1131 = _T_1122 | _T_1130; // @[ifu_compress_ctl.scala 96:70]
  wire  _T_1139 = _T_897 & io_din[10]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1140 = _T_1131 | _T_1139; // @[ifu_compress_ctl.scala 96:95]
  wire  _T_1148 = _T_897 & io_din[11]; // @[ifu_compress_ctl.scala 12:110]
  wire  sluimm17_12 = _T_1140 | _T_1148; // @[ifu_compress_ctl.scala 96:121]
  wire  uimm5_0 = _T_79 | _T_195; // @[ifu_compress_ctl.scala 98:45]
  wire [6:0] l1_6 = {out_6,out_5,out_4,_T_228,out_2,1'h1,1'h1}; // @[Cat.scala 29:58]
  wire [4:0] _T_1192 = rdrd ? rdd : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_1193 = rdprd ? rdpd : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_1194 = rs2prd ? rs2pd : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_1195 = rdeq1 ? 5'h1 : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_1196 = rdeq2 ? 5'h2 : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_1197 = _T_1192 | _T_1193; // @[Mux.scala 27:72]
  wire [4:0] _T_1198 = _T_1197 | _T_1194; // @[Mux.scala 27:72]
  wire [4:0] _T_1199 = _T_1198 | _T_1195; // @[Mux.scala 27:72]
  wire [4:0] l1_11 = _T_1199 | _T_1196; // @[Mux.scala 27:72]
  wire [4:0] _T_1210 = rdrs1 ? rdd : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_1211 = rdprs1 ? rdpd : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_1212 = rs1eq2 ? 5'h2 : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_1213 = _T_1210 | _T_1211; // @[Mux.scala 27:72]
  wire [4:0] l1_19 = _T_1213 | _T_1212; // @[Mux.scala 27:72]
  wire [4:0] _T_1219 = {3'h0,1'h0,out_20}; // @[Cat.scala 29:58]
  wire [4:0] _T_1222 = rs2rs2 ? rs2d : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_1223 = rs2prs2 ? rs2pd : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_1224 = _T_1222 | _T_1223; // @[Mux.scala 27:72]
  wire [4:0] l1_24 = _T_1219 | _T_1224; // @[ifu_compress_ctl.scala 114:67]
  wire [14:0] _T_1232 = {out_14,out_13,out_12,l1_11,l1_6}; // @[Cat.scala 29:58]
  wire [31:0] l1 = {1'h0,out_30,2'h0,3'h0,l1_24,l1_19,_T_1232}; // @[Cat.scala 29:58]
  wire [5:0] simm5d = {io_din[12],rs2d}; // @[Cat.scala 29:58]
  wire [5:0] simm9d = {io_din[12],io_din[4:3],io_din[5],io_din[2],io_din[6]}; // @[Cat.scala 29:58]
  wire [10:0] sjald_1 = {io_din[12],io_din[8],io_din[10:9],io_din[6],io_din[7],io_din[2],io_din[11],io_din[5:4],io_din[3]}; // @[Cat.scala 29:58]
  wire [19:0] sjald = {io_din[12],io_din[12],io_din[12],io_din[12],io_din[12],io_din[12],io_din[12],io_din[12],io_din[12],sjald_1}; // @[Cat.scala 29:58]
  wire [9:0] _T_1296 = {io_din[12],io_din[12],io_din[12],io_din[12],io_din[12],io_din[12],io_din[12],io_din[12],io_din[12],io_din[12]}; // @[Cat.scala 29:58]
  wire [19:0] sluimmd = {_T_1296,io_din[12],io_din[12],io_din[12],io_din[12],io_din[12],rs2d}; // @[Cat.scala 29:58]
  wire [11:0] _T_1314 = {simm5d[5],simm5d[5],simm5d[5],simm5d[5],simm5d[5],simm5d[5],simm5d[5],simm5d[4:0]}; // @[Cat.scala 29:58]
  wire [11:0] _T_1317 = {2'h0,io_din[10:7],io_din[12:11],io_din[5],io_din[6],2'h0}; // @[Cat.scala 29:58]
  wire [11:0] _T_1325 = {simm9d[5],simm9d[5],simm9d[5],simm9d[4:0],4'h0}; // @[Cat.scala 29:58]
  wire [11:0] _T_1328 = {5'h0,io_din[5],io_din[12:10],io_din[6],2'h0}; // @[Cat.scala 29:58]
  wire [11:0] _T_1331 = {4'h0,io_din[3:2],io_din[12],io_din[6:4],2'h0}; // @[Cat.scala 29:58]
  wire [11:0] _T_1333 = {6'h0,io_din[12],rs2d}; // @[Cat.scala 29:58]
  wire [11:0] _T_1339 = {sjald[19],sjald[9:0],sjald[10]}; // @[Cat.scala 29:58]
  wire [11:0] _T_1342 = simm5_0 ? _T_1314 : 12'h0; // @[Mux.scala 27:72]
  wire [11:0] _T_1343 = uimm9_2 ? _T_1317 : 12'h0; // @[Mux.scala 27:72]
  wire [11:0] _T_1344 = rdeq2 ? _T_1325 : 12'h0; // @[Mux.scala 27:72]
  wire [11:0] _T_1345 = ulwimm6_2 ? _T_1328 : 12'h0; // @[Mux.scala 27:72]
  wire [11:0] _T_1346 = ulwspimm7_2 ? _T_1331 : 12'h0; // @[Mux.scala 27:72]
  wire [11:0] _T_1347 = uimm5_0 ? _T_1333 : 12'h0; // @[Mux.scala 27:72]
  wire [11:0] _T_1348 = _T_228 ? _T_1339 : 12'h0; // @[Mux.scala 27:72]
  wire [11:0] _T_1349 = sluimm17_12 ? sluimmd[19:8] : 12'h0; // @[Mux.scala 27:72]
  wire [11:0] _T_1350 = _T_1342 | _T_1343; // @[Mux.scala 27:72]
  wire [11:0] _T_1351 = _T_1350 | _T_1344; // @[Mux.scala 27:72]
  wire [11:0] _T_1352 = _T_1351 | _T_1345; // @[Mux.scala 27:72]
  wire [11:0] _T_1353 = _T_1352 | _T_1346; // @[Mux.scala 27:72]
  wire [11:0] _T_1354 = _T_1353 | _T_1347; // @[Mux.scala 27:72]
  wire [11:0] _T_1355 = _T_1354 | _T_1348; // @[Mux.scala 27:72]
  wire [11:0] _T_1356 = _T_1355 | _T_1349; // @[Mux.scala 27:72]
  wire [11:0] l2_31 = l1[31:20] | _T_1356; // @[ifu_compress_ctl.scala 133:25]
  wire [7:0] _T_1363 = _T_228 ? sjald[19:12] : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_1364 = sluimm17_12 ? sluimmd[7:0] : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_1365 = _T_1363 | _T_1364; // @[Mux.scala 27:72]
  wire [7:0] l2_19 = l1[19:12] | _T_1365; // @[ifu_compress_ctl.scala 143:25]
  wire [31:0] l2 = {l2_31,l2_19,l1[11:0]}; // @[Cat.scala 29:58]
  wire [8:0] sbr8d = {io_din[12],io_din[6],io_din[5],io_din[2],io_din[11],io_din[10],io_din[4],io_din[3],1'h0}; // @[Cat.scala 29:58]
  wire [6:0] uswimm6d = {io_din[5],io_din[12:10],io_din[6],2'h0}; // @[Cat.scala 29:58]
  wire [7:0] uswspimm7d = {io_din[8:7],io_din[12:9],2'h0}; // @[Cat.scala 29:58]
  wire [6:0] _T_1400 = {sbr8d[8],sbr8d[8],sbr8d[8],sbr8d[8],sbr8d[7:5]}; // @[Cat.scala 29:58]
  wire [6:0] _T_1403 = {5'h0,uswimm6d[6:5]}; // @[Cat.scala 29:58]
  wire [6:0] _T_1406 = {4'h0,uswspimm7d[7:5]}; // @[Cat.scala 29:58]
  wire [6:0] _T_1407 = _T_234 ? _T_1400 : 7'h0; // @[Mux.scala 27:72]
  wire [6:0] _T_1408 = _T_854 ? _T_1403 : 7'h0; // @[Mux.scala 27:72]
  wire [6:0] _T_1409 = _T_807 ? _T_1406 : 7'h0; // @[Mux.scala 27:72]
  wire [6:0] _T_1410 = _T_1407 | _T_1408; // @[Mux.scala 27:72]
  wire [6:0] _T_1411 = _T_1410 | _T_1409; // @[Mux.scala 27:72]
  wire [6:0] l3_31 = l2[31:25] | _T_1411; // @[ifu_compress_ctl.scala 151:25]
  wire [12:0] l3_24 = l2[24:12]; // @[ifu_compress_ctl.scala 154:17]
  wire [4:0] _T_1417 = {sbr8d[4:1],sbr8d[8]}; // @[Cat.scala 29:58]
  wire [4:0] _T_1422 = _T_234 ? _T_1417 : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_1423 = _T_854 ? uswimm6d[4:0] : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_1424 = _T_807 ? uswspimm7d[4:0] : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_1425 = _T_1422 | _T_1423; // @[Mux.scala 27:72]
  wire [4:0] _T_1426 = _T_1425 | _T_1424; // @[Mux.scala 27:72]
  wire [4:0] l3_11 = l2[11:7] | _T_1426; // @[ifu_compress_ctl.scala 156:24]
  wire [31:0] l3 = {l3_31,l3_24,l3_11,l2[6:0]}; // @[Cat.scala 29:58]
  wire  _T_1437 = _T_4 & _T_487; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1438 = _T_1437 & io_din[11]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1439 = _T_1438 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1442 = _T_1439 & _T_147; // @[ifu_compress_ctl.scala 162:39]
  wire  _T_1450 = _T_1437 & io_din[6]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1451 = _T_1450 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1454 = _T_1451 & _T_147; // @[ifu_compress_ctl.scala 162:79]
  wire  _T_1455 = _T_1442 | _T_1454; // @[ifu_compress_ctl.scala 162:54]
  wire  _T_1464 = _T_642 & io_din[11]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1465 = _T_1464 & _T_830; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1466 = _T_1455 | _T_1465; // @[ifu_compress_ctl.scala 162:94]
  wire  _T_1474 = _T_1437 & io_din[5]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1475 = _T_1474 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1478 = _T_1475 & _T_147; // @[ifu_compress_ctl.scala 163:55]
  wire  _T_1479 = _T_1466 | _T_1478; // @[ifu_compress_ctl.scala 163:30]
  wire  _T_1487 = _T_1437 & io_din[10]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1488 = _T_1487 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1491 = _T_1488 & _T_147; // @[ifu_compress_ctl.scala 163:96]
  wire  _T_1492 = _T_1479 | _T_1491; // @[ifu_compress_ctl.scala 163:70]
  wire  _T_1501 = _T_642 & io_din[6]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1502 = _T_1501 & _T_830; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1503 = _T_1492 | _T_1502; // @[ifu_compress_ctl.scala 163:111]
  wire  _T_1510 = io_din[15] & _T_487; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1511 = _T_1510 & _T_830; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1512 = _T_1511 & io_din[0]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1513 = _T_1503 | _T_1512; // @[ifu_compress_ctl.scala 164:29]
  wire  _T_1521 = _T_1437 & io_din[9]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1522 = _T_1521 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1525 = _T_1522 & _T_147; // @[ifu_compress_ctl.scala 164:79]
  wire  _T_1526 = _T_1513 | _T_1525; // @[ifu_compress_ctl.scala 164:54]
  wire  _T_1533 = _T_487 & io_din[6]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1534 = _T_1533 & _T_830; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1535 = _T_1534 & io_din[0]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1536 = _T_1526 | _T_1535; // @[ifu_compress_ctl.scala 164:94]
  wire  _T_1545 = _T_642 & io_din[5]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1546 = _T_1545 & _T_830; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1547 = _T_1536 | _T_1546; // @[ifu_compress_ctl.scala 164:118]
  wire  _T_1555 = _T_1437 & io_din[8]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1556 = _T_1555 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1559 = _T_1556 & _T_147; // @[ifu_compress_ctl.scala 165:28]
  wire  _T_1560 = _T_1547 | _T_1559; // @[ifu_compress_ctl.scala 164:144]
  wire  _T_1567 = _T_487 & io_din[5]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1568 = _T_1567 & _T_830; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1569 = _T_1568 & io_din[0]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1570 = _T_1560 | _T_1569; // @[ifu_compress_ctl.scala 165:43]
  wire  _T_1579 = _T_642 & io_din[10]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1580 = _T_1579 & _T_830; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1581 = _T_1570 | _T_1580; // @[ifu_compress_ctl.scala 165:67]
  wire  _T_1589 = _T_1437 & io_din[7]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1590 = _T_1589 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1593 = _T_1590 & _T_147; // @[ifu_compress_ctl.scala 166:28]
  wire  _T_1594 = _T_1581 | _T_1593; // @[ifu_compress_ctl.scala 165:94]
  wire  _T_1602 = io_din[12] & io_din[11]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1603 = _T_1602 & _T_38; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1604 = _T_1603 & _T_830; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1605 = _T_1604 & io_din[0]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1606 = _T_1594 | _T_1605; // @[ifu_compress_ctl.scala 166:43]
  wire  _T_1615 = _T_642 & io_din[9]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1616 = _T_1615 & _T_830; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1617 = _T_1606 | _T_1616; // @[ifu_compress_ctl.scala 166:71]
  wire  _T_1625 = _T_1437 & io_din[4]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1626 = _T_1625 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1629 = _T_1626 & _T_147; // @[ifu_compress_ctl.scala 167:28]
  wire  _T_1630 = _T_1617 | _T_1629; // @[ifu_compress_ctl.scala 166:97]
  wire  _T_1636 = io_din[13] & io_din[12]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1637 = _T_1636 & _T_830; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1638 = _T_1637 & io_din[0]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1639 = _T_1630 | _T_1638; // @[ifu_compress_ctl.scala 167:43]
  wire  _T_1648 = _T_642 & io_din[8]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1649 = _T_1648 & _T_830; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1650 = _T_1639 | _T_1649; // @[ifu_compress_ctl.scala 167:67]
  wire  _T_1658 = _T_1437 & io_din[3]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1659 = _T_1658 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1662 = _T_1659 & _T_147; // @[ifu_compress_ctl.scala 168:28]
  wire  _T_1663 = _T_1650 | _T_1662; // @[ifu_compress_ctl.scala 167:93]
  wire  _T_1669 = io_din[13] & io_din[4]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1670 = _T_1669 & _T_830; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1671 = _T_1670 & io_din[0]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1672 = _T_1663 | _T_1671; // @[ifu_compress_ctl.scala 168:43]
  wire  _T_1680 = _T_1437 & io_din[2]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1681 = _T_1680 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1684 = _T_1681 & _T_147; // @[ifu_compress_ctl.scala 168:91]
  wire  _T_1685 = _T_1672 | _T_1684; // @[ifu_compress_ctl.scala 168:66]
  wire  _T_1694 = _T_642 & io_din[7]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1695 = _T_1694 & _T_830; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1696 = _T_1685 | _T_1695; // @[ifu_compress_ctl.scala 168:106]
  wire  _T_1702 = io_din[13] & io_din[3]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1703 = _T_1702 & _T_830; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1704 = _T_1703 & io_din[0]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1705 = _T_1696 | _T_1704; // @[ifu_compress_ctl.scala 169:29]
  wire  _T_1711 = io_din[13] & io_din[2]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1712 = _T_1711 & _T_830; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1713 = _T_1712 & io_din[0]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1714 = _T_1705 | _T_1713; // @[ifu_compress_ctl.scala 169:52]
  wire  _T_1720 = io_din[14] & _T_4; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1721 = _T_1720 & _T_830; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1722 = _T_1714 | _T_1721; // @[ifu_compress_ctl.scala 169:75]
  wire  _T_1731 = _T_703 & _T_830; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1732 = _T_1731 & io_din[0]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1733 = _T_1722 | _T_1732; // @[ifu_compress_ctl.scala 169:98]
  wire  _T_1740 = _T_820 & io_din[12]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1741 = _T_1740 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1744 = _T_1741 & _T_147; // @[ifu_compress_ctl.scala 170:54]
  wire  _T_1745 = _T_1733 | _T_1744; // @[ifu_compress_ctl.scala 170:29]
  wire  _T_1754 = _T_642 & _T_487; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1755 = _T_1754 & io_din[1]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1758 = _T_1755 & _T_147; // @[ifu_compress_ctl.scala 170:96]
  wire  _T_1759 = _T_1745 | _T_1758; // @[ifu_compress_ctl.scala 170:69]
  wire  _T_1768 = _T_642 & io_din[12]; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1769 = _T_1768 & _T_830; // @[ifu_compress_ctl.scala 12:110]
  wire  _T_1770 = _T_1759 | _T_1769; // @[ifu_compress_ctl.scala 170:111]
  wire  _T_1777 = _T_1720 & _T_147; // @[ifu_compress_ctl.scala 171:50]
  wire  legal = _T_1770 | _T_1777; // @[ifu_compress_ctl.scala 171:30]
  wire [9:0] _T_1787 = {legal,legal,legal,legal,legal,legal,legal,legal,legal,legal}; // @[Cat.scala 29:58]
  wire [18:0] _T_1796 = {_T_1787,legal,legal,legal,legal,legal,legal,legal,legal,legal}; // @[Cat.scala 29:58]
  wire [27:0] _T_1805 = {_T_1796,legal,legal,legal,legal,legal,legal,legal,legal,legal}; // @[Cat.scala 29:58]
  wire [31:0] _T_1809 = {_T_1805,legal,legal,legal,legal}; // @[Cat.scala 29:58]
  assign io_dout = l3 & _T_1809; // @[ifu_compress_ctl.scala 173:10]
endmodule
module ifu_aln_ctl(
  input         clock,
  input         reset,
  input         io_scan_mode,
  input         io_active_clk,
  input         io_ifu_async_error_start,
  input         io_iccm_rd_ecc_double_err,
  input         io_ic_access_fault_f,
  input  [1:0]  io_ic_access_fault_type_f,
  input  [7:0]  io_ifu_bp_fghr_f,
  input  [30:0] io_ifu_bp_btb_target_f,
  input  [11:0] io_ifu_bp_poffset_f,
  input  [1:0]  io_ifu_bp_hist0_f,
  input  [1:0]  io_ifu_bp_hist1_f,
  input  [1:0]  io_ifu_bp_pc4_f,
  input  [1:0]  io_ifu_bp_way_f,
  input  [1:0]  io_ifu_bp_valid_f,
  input  [1:0]  io_ifu_bp_ret_f,
  input         io_exu_flush_final,
  input         io_dec_aln_aln_dec_dec_i0_decode_d,
  output [15:0] io_dec_aln_aln_dec_ifu_i0_cinst,
  output        io_dec_aln_aln_ib_ifu_i0_icaf,
  output [1:0]  io_dec_aln_aln_ib_ifu_i0_icaf_type,
  output        io_dec_aln_aln_ib_ifu_i0_icaf_f1,
  output        io_dec_aln_aln_ib_ifu_i0_dbecc,
  output [7:0]  io_dec_aln_aln_ib_ifu_i0_bp_index,
  output [7:0]  io_dec_aln_aln_ib_ifu_i0_bp_fghr,
  output [4:0]  io_dec_aln_aln_ib_ifu_i0_bp_btag,
  output        io_dec_aln_aln_ib_ifu_i0_valid,
  output [31:0] io_dec_aln_aln_ib_ifu_i0_instr,
  output [30:0] io_dec_aln_aln_ib_ifu_i0_pc,
  output        io_dec_aln_aln_ib_ifu_i0_pc4,
  output        io_dec_aln_aln_ib_i0_brp_valid,
  output [11:0] io_dec_aln_aln_ib_i0_brp_bits_toffset,
  output [1:0]  io_dec_aln_aln_ib_i0_brp_bits_hist,
  output        io_dec_aln_aln_ib_i0_brp_bits_br_error,
  output        io_dec_aln_aln_ib_i0_brp_bits_br_start_error,
  output        io_dec_aln_aln_ib_i0_brp_bits_bank,
  output [30:0] io_dec_aln_aln_ib_i0_brp_bits_prett,
  output        io_dec_aln_aln_ib_i0_brp_bits_way,
  output        io_dec_aln_aln_ib_i0_brp_bits_ret,
  output        io_dec_aln_ifu_pmu_instr_aligned,
  input  [31:0] io_ifu_fetch_data_f,
  input  [1:0]  io_ifu_fetch_val,
  input  [30:0] io_ifu_fetch_pc,
  output        io_ifu_fb_consume1,
  output        io_ifu_fb_consume2
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
`endif // RANDOMIZE_REG_INIT
  wire  rvclkhdr_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_1_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_1_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_1_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_1_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_2_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_2_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_2_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_2_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_3_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_3_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_3_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_3_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_4_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_4_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_4_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_4_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_5_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_5_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_5_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_5_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_6_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_6_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_6_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_6_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_7_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_7_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_7_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_7_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_8_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_8_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_8_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_8_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_9_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_9_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_9_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_9_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_10_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_10_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_10_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_10_io_scan_mode; // @[lib.scala 368:23]
  wire  rvclkhdr_11_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_11_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_11_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_11_io_scan_mode; // @[lib.scala 368:23]
  wire [15:0] decompressed_io_din; // @[ifu_aln_ctl.scala 352:28]
  wire [31:0] decompressed_io_dout; // @[ifu_aln_ctl.scala 352:28]
  reg  error_stall; // @[ifu_aln_ctl.scala 102:51]
  wire  _T = error_stall | io_ifu_async_error_start; // @[ifu_aln_ctl.scala 99:34]
  wire  _T_1 = ~io_exu_flush_final; // @[ifu_aln_ctl.scala 99:64]
  reg [1:0] wrptr; // @[ifu_aln_ctl.scala 104:48]
  reg [1:0] rdptr; // @[ifu_aln_ctl.scala 106:48]
  reg [1:0] f2val; // @[ifu_aln_ctl.scala 108:48]
  reg [1:0] f1val; // @[ifu_aln_ctl.scala 109:48]
  reg [1:0] f0val; // @[ifu_aln_ctl.scala 110:48]
  reg  q2off; // @[ifu_aln_ctl.scala 112:48]
  reg  q1off; // @[ifu_aln_ctl.scala 113:48]
  reg  q0off; // @[ifu_aln_ctl.scala 114:48]
  wire  _T_785 = ~error_stall; // @[ifu_aln_ctl.scala 395:55]
  wire  i0_shift = io_dec_aln_aln_dec_dec_i0_decode_d & _T_785; // @[ifu_aln_ctl.scala 395:53]
  wire  _T_186 = rdptr == 2'h0; // @[ifu_aln_ctl.scala 169:31]
  wire  _T_189 = _T_186 & q0off; // @[Mux.scala 27:72]
  wire  _T_187 = rdptr == 2'h1; // @[ifu_aln_ctl.scala 170:11]
  wire  _T_190 = _T_187 & q1off; // @[Mux.scala 27:72]
  wire  _T_192 = _T_189 | _T_190; // @[Mux.scala 27:72]
  wire  _T_188 = rdptr == 2'h2; // @[ifu_aln_ctl.scala 171:11]
  wire  _T_191 = _T_188 & q2off; // @[Mux.scala 27:72]
  wire  q0ptr = _T_192 | _T_191; // @[Mux.scala 27:72]
  wire  _T_202 = ~q0ptr; // @[ifu_aln_ctl.scala 175:26]
  wire [1:0] q0sel = {q0ptr,_T_202}; // @[Cat.scala 29:58]
  wire [2:0] qren = {_T_188,_T_187,_T_186}; // @[Cat.scala 29:58]
  reg [31:0] q1; // @[lib.scala 374:16]
  reg [31:0] q0; // @[lib.scala 374:16]
  wire [63:0] _T_479 = {q1,q0}; // @[Cat.scala 29:58]
  wire [63:0] _T_486 = qren[0] ? _T_479 : 64'h0; // @[Mux.scala 27:72]
  reg [31:0] q2; // @[lib.scala 374:16]
  wire [63:0] _T_482 = {q2,q1}; // @[Cat.scala 29:58]
  wire [63:0] _T_487 = qren[1] ? _T_482 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_489 = _T_486 | _T_487; // @[Mux.scala 27:72]
  wire [63:0] _T_485 = {q0,q2}; // @[Cat.scala 29:58]
  wire [63:0] _T_488 = qren[2] ? _T_485 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] qeff = _T_489 | _T_488; // @[Mux.scala 27:72]
  wire [31:0] q0eff = qeff[31:0]; // @[ifu_aln_ctl.scala 294:42]
  wire [31:0] _T_496 = q0sel[0] ? q0eff : 32'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_497 = q0sel[1] ? q0eff[31:16] : 16'h0; // @[Mux.scala 27:72]
  wire [31:0] _GEN_0 = {{16'd0}, _T_497}; // @[Mux.scala 27:72]
  wire [31:0] q0final = _T_496 | _GEN_0; // @[Mux.scala 27:72]
  wire [31:0] _T_520 = f0val[1] ? q0final : 32'h0; // @[Mux.scala 27:72]
  wire  _T_513 = ~f0val[1]; // @[ifu_aln_ctl.scala 301:58]
  wire  _T_515 = _T_513 & f0val[0]; // @[ifu_aln_ctl.scala 301:68]
  wire  _T_197 = _T_186 & q1off; // @[Mux.scala 27:72]
  wire  _T_198 = _T_187 & q2off; // @[Mux.scala 27:72]
  wire  _T_200 = _T_197 | _T_198; // @[Mux.scala 27:72]
  wire  _T_199 = _T_188 & q0off; // @[Mux.scala 27:72]
  wire  q1ptr = _T_200 | _T_199; // @[Mux.scala 27:72]
  wire  _T_203 = ~q1ptr; // @[ifu_aln_ctl.scala 177:26]
  wire [1:0] q1sel = {q1ptr,_T_203}; // @[Cat.scala 29:58]
  wire [31:0] q1eff = qeff[63:32]; // @[ifu_aln_ctl.scala 294:29]
  wire [15:0] _T_506 = q1sel[0] ? q1eff[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_507 = q1sel[1] ? q1eff[31:16] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] q1final = _T_506 | _T_507; // @[Mux.scala 27:72]
  wire [31:0] _T_519 = {q1final,q0final[15:0]}; // @[Cat.scala 29:58]
  wire [31:0] _T_521 = _T_515 ? _T_519 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] aligndata = _T_520 | _T_521; // @[Mux.scala 27:72]
  wire  first4B = aligndata[1:0] == 2'h3; // @[ifu_aln_ctl.scala 334:29]
  wire  first2B = ~first4B; // @[ifu_aln_ctl.scala 336:17]
  wire  shift_2B = i0_shift & first2B; // @[ifu_aln_ctl.scala 399:24]
  wire [1:0] _T_443 = {1'h0,f0val[1]}; // @[Cat.scala 29:58]
  wire [1:0] _T_448 = shift_2B ? _T_443 : 2'h0; // @[Mux.scala 27:72]
  wire  _T_444 = ~shift_2B; // @[ifu_aln_ctl.scala 284:18]
  wire  shift_4B = i0_shift & first4B; // @[ifu_aln_ctl.scala 400:24]
  wire  _T_445 = ~shift_4B; // @[ifu_aln_ctl.scala 284:30]
  wire  _T_446 = _T_444 & _T_445; // @[ifu_aln_ctl.scala 284:28]
  wire [1:0] _T_449 = _T_446 ? f0val : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] sf0val = _T_448 | _T_449; // @[Mux.scala 27:72]
  wire  sf0_valid = sf0val[0]; // @[ifu_aln_ctl.scala 235:22]
  wire  _T_351 = ~sf0_valid; // @[ifu_aln_ctl.scala 256:26]
  wire  _T_802 = f0val[0] & _T_513; // @[ifu_aln_ctl.scala 403:28]
  wire  f1_shift_2B = _T_802 & shift_4B; // @[ifu_aln_ctl.scala 403:40]
  wire  _T_417 = f1_shift_2B & f1val[1]; // @[Mux.scala 27:72]
  wire  _T_416 = ~f1_shift_2B; // @[ifu_aln_ctl.scala 277:53]
  wire [1:0] _T_418 = _T_416 ? f1val : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _GEN_1 = {{1'd0}, _T_417}; // @[Mux.scala 27:72]
  wire [1:0] sf1val = _GEN_1 | _T_418; // @[Mux.scala 27:72]
  wire  sf1_valid = sf1val[0]; // @[ifu_aln_ctl.scala 234:22]
  wire  _T_352 = _T_351 & sf1_valid; // @[ifu_aln_ctl.scala 256:37]
  wire  f2_valid = f2val[0]; // @[ifu_aln_ctl.scala 233:20]
  wire  _T_353 = _T_352 & f2_valid; // @[ifu_aln_ctl.scala 256:50]
  wire  ifvalid = io_ifu_fetch_val[0]; // @[ifu_aln_ctl.scala 244:30]
  wire  _T_354 = _T_353 & ifvalid; // @[ifu_aln_ctl.scala 256:62]
  wire  _T_355 = sf0_valid & sf1_valid; // @[ifu_aln_ctl.scala 257:37]
  wire  _T_356 = ~f2_valid; // @[ifu_aln_ctl.scala 257:52]
  wire  _T_357 = _T_355 & _T_356; // @[ifu_aln_ctl.scala 257:50]
  wire  _T_358 = _T_357 & ifvalid; // @[ifu_aln_ctl.scala 257:62]
  wire  fetch_to_f2 = _T_354 | _T_358; // @[ifu_aln_ctl.scala 256:74]
  reg [30:0] f2pc; // @[lib.scala 374:16]
  wire  _T_335 = ~sf1_valid; // @[ifu_aln_ctl.scala 252:39]
  wire  _T_336 = _T_351 & _T_335; // @[ifu_aln_ctl.scala 252:37]
  wire  _T_337 = _T_336 & f2_valid; // @[ifu_aln_ctl.scala 252:50]
  wire  _T_338 = _T_337 & ifvalid; // @[ifu_aln_ctl.scala 252:62]
  wire  _T_342 = _T_352 & _T_356; // @[ifu_aln_ctl.scala 253:50]
  wire  _T_343 = _T_342 & ifvalid; // @[ifu_aln_ctl.scala 253:62]
  wire  _T_344 = _T_338 | _T_343; // @[ifu_aln_ctl.scala 252:74]
  wire  _T_346 = sf0_valid & _T_335; // @[ifu_aln_ctl.scala 254:37]
  wire  _T_348 = _T_346 & _T_356; // @[ifu_aln_ctl.scala 254:50]
  wire  _T_349 = _T_348 & ifvalid; // @[ifu_aln_ctl.scala 254:62]
  wire  fetch_to_f1 = _T_344 | _T_349; // @[ifu_aln_ctl.scala 253:74]
  wire  _T_25 = fetch_to_f1 | _T_353; // @[ifu_aln_ctl.scala 134:33]
  reg [30:0] f1pc; // @[lib.scala 374:16]
  wire  _T_332 = _T_336 & _T_356; // @[ifu_aln_ctl.scala 251:50]
  wire  fetch_to_f0 = _T_332 & ifvalid; // @[ifu_aln_ctl.scala 251:62]
  wire  _T_27 = fetch_to_f0 | _T_337; // @[ifu_aln_ctl.scala 135:33]
  wire  _T_28 = _T_27 | _T_352; // @[ifu_aln_ctl.scala 135:47]
  wire  _T_29 = _T_28 | shift_2B; // @[ifu_aln_ctl.scala 135:61]
  reg [30:0] f0pc; // @[lib.scala 374:16]
  wire  _T_35 = wrptr == 2'h2; // @[ifu_aln_ctl.scala 139:21]
  wire  _T_36 = _T_35 & ifvalid; // @[ifu_aln_ctl.scala 139:29]
  wire  _T_37 = wrptr == 2'h1; // @[ifu_aln_ctl.scala 139:46]
  wire  _T_38 = _T_37 & ifvalid; // @[ifu_aln_ctl.scala 139:54]
  wire  _T_39 = wrptr == 2'h0; // @[ifu_aln_ctl.scala 139:71]
  wire  _T_40 = _T_39 & ifvalid; // @[ifu_aln_ctl.scala 139:79]
  wire [2:0] qwen = {_T_36,_T_38,_T_40}; // @[Cat.scala 29:58]
  reg [11:0] brdata2; // @[lib.scala 374:16]
  reg [11:0] brdata1; // @[lib.scala 374:16]
  reg [11:0] brdata0; // @[lib.scala 374:16]
  reg [54:0] misc2; // @[lib.scala 374:16]
  reg [54:0] misc1; // @[lib.scala 374:16]
  reg [54:0] misc0; // @[lib.scala 374:16]
  wire  _T_44 = qren[0] & io_ifu_fb_consume1; // @[ifu_aln_ctl.scala 143:34]
  wire  _T_46 = _T_44 & _T_1; // @[ifu_aln_ctl.scala 143:55]
  wire  _T_49 = qren[1] & io_ifu_fb_consume1; // @[ifu_aln_ctl.scala 144:14]
  wire  _T_51 = _T_49 & _T_1; // @[ifu_aln_ctl.scala 144:35]
  wire  _T_59 = qren[0] & io_ifu_fb_consume2; // @[ifu_aln_ctl.scala 146:14]
  wire  _T_61 = _T_59 & _T_1; // @[ifu_aln_ctl.scala 146:35]
  wire  _T_69 = qren[2] & io_ifu_fb_consume2; // @[ifu_aln_ctl.scala 148:14]
  wire  _T_71 = _T_69 & _T_1; // @[ifu_aln_ctl.scala 148:35]
  wire  _T_73 = ~io_ifu_fb_consume1; // @[ifu_aln_ctl.scala 149:6]
  wire  _T_74 = ~io_ifu_fb_consume2; // @[ifu_aln_ctl.scala 149:28]
  wire  _T_75 = _T_73 & _T_74; // @[ifu_aln_ctl.scala 149:26]
  wire  _T_77 = _T_75 & _T_1; // @[ifu_aln_ctl.scala 149:48]
  wire [1:0] _T_80 = _T_51 ? 2'h2 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_82 = _T_61 ? 2'h2 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_85 = _T_77 ? rdptr : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _GEN_2 = {{1'd0}, _T_46}; // @[Mux.scala 27:72]
  wire [1:0] _T_86 = _GEN_2 | _T_80; // @[Mux.scala 27:72]
  wire [1:0] _T_88 = _T_86 | _T_82; // @[Mux.scala 27:72]
  wire [1:0] _GEN_3 = {{1'd0}, _T_71}; // @[Mux.scala 27:72]
  wire [1:0] _T_90 = _T_88 | _GEN_3; // @[Mux.scala 27:72]
  wire  _T_95 = qwen[0] & _T_1; // @[ifu_aln_ctl.scala 152:34]
  wire  _T_99 = qwen[1] & _T_1; // @[ifu_aln_ctl.scala 153:14]
  wire  _T_105 = ~ifvalid; // @[ifu_aln_ctl.scala 155:6]
  wire  _T_107 = _T_105 & _T_1; // @[ifu_aln_ctl.scala 155:15]
  wire [1:0] _T_110 = _T_99 ? 2'h2 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_112 = _T_107 ? wrptr : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _GEN_4 = {{1'd0}, _T_95}; // @[Mux.scala 27:72]
  wire [1:0] _T_113 = _GEN_4 | _T_110; // @[Mux.scala 27:72]
  wire  _T_118 = ~qwen[2]; // @[ifu_aln_ctl.scala 157:26]
  wire  _T_120 = _T_118 & _T_188; // @[ifu_aln_ctl.scala 157:35]
  wire  _T_795 = shift_2B & f0val[0]; // @[Mux.scala 27:72]
  wire  _T_796 = shift_4B & _T_802; // @[Mux.scala 27:72]
  wire  f0_shift_2B = _T_795 | _T_796; // @[Mux.scala 27:72]
  wire  _T_122 = q2off | f0_shift_2B; // @[ifu_aln_ctl.scala 157:74]
  wire  _T_126 = _T_118 & _T_187; // @[ifu_aln_ctl.scala 158:15]
  wire  _T_128 = q2off | f1_shift_2B; // @[ifu_aln_ctl.scala 158:54]
  wire  _T_132 = _T_118 & _T_186; // @[ifu_aln_ctl.scala 159:15]
  wire  _T_134 = _T_120 & _T_122; // @[Mux.scala 27:72]
  wire  _T_135 = _T_126 & _T_128; // @[Mux.scala 27:72]
  wire  _T_136 = _T_132 & q2off; // @[Mux.scala 27:72]
  wire  _T_137 = _T_134 | _T_135; // @[Mux.scala 27:72]
  wire  _T_141 = ~qwen[1]; // @[ifu_aln_ctl.scala 161:26]
  wire  _T_143 = _T_141 & _T_187; // @[ifu_aln_ctl.scala 161:35]
  wire  _T_145 = q1off | f0_shift_2B; // @[ifu_aln_ctl.scala 161:74]
  wire  _T_149 = _T_141 & _T_186; // @[ifu_aln_ctl.scala 162:15]
  wire  _T_151 = q1off | f1_shift_2B; // @[ifu_aln_ctl.scala 162:54]
  wire  _T_155 = _T_141 & _T_188; // @[ifu_aln_ctl.scala 163:15]
  wire  _T_157 = _T_143 & _T_145; // @[Mux.scala 27:72]
  wire  _T_158 = _T_149 & _T_151; // @[Mux.scala 27:72]
  wire  _T_159 = _T_155 & q1off; // @[Mux.scala 27:72]
  wire  _T_160 = _T_157 | _T_158; // @[Mux.scala 27:72]
  wire  _T_164 = ~qwen[0]; // @[ifu_aln_ctl.scala 165:26]
  wire  _T_166 = _T_164 & _T_186; // @[ifu_aln_ctl.scala 165:35]
  wire  _T_168 = q0off | f0_shift_2B; // @[ifu_aln_ctl.scala 165:76]
  wire  _T_172 = _T_164 & _T_188; // @[ifu_aln_ctl.scala 166:35]
  wire  _T_174 = q0off | f1_shift_2B; // @[ifu_aln_ctl.scala 166:76]
  wire  _T_178 = _T_164 & _T_187; // @[ifu_aln_ctl.scala 167:35]
  wire  _T_180 = _T_166 & _T_168; // @[Mux.scala 27:72]
  wire  _T_181 = _T_172 & _T_174; // @[Mux.scala 27:72]
  wire  _T_182 = _T_178 & q0off; // @[Mux.scala 27:72]
  wire  _T_183 = _T_180 | _T_181; // @[Mux.scala 27:72]
  wire [50:0] _T_205 = {io_ifu_bp_btb_target_f,io_ifu_bp_poffset_f,io_ifu_bp_fghr_f}; // @[Cat.scala 29:58]
  wire [3:0] _T_207 = {io_iccm_rd_ecc_double_err,io_ic_access_fault_f,io_ic_access_fault_type_f}; // @[Cat.scala 29:58]
  wire [109:0] _T_211 = {misc1,misc0}; // @[Cat.scala 29:58]
  wire [109:0] _T_214 = {misc2,misc1}; // @[Cat.scala 29:58]
  wire [109:0] _T_217 = {misc0,misc2}; // @[Cat.scala 29:58]
  wire [109:0] _T_218 = qren[0] ? _T_211 : 110'h0; // @[Mux.scala 27:72]
  wire [109:0] _T_219 = qren[1] ? _T_214 : 110'h0; // @[Mux.scala 27:72]
  wire [109:0] _T_220 = qren[2] ? _T_217 : 110'h0; // @[Mux.scala 27:72]
  wire [109:0] _T_221 = _T_218 | _T_219; // @[Mux.scala 27:72]
  wire [109:0] misceff = _T_221 | _T_220; // @[Mux.scala 27:72]
  wire [54:0] misc1eff = misceff[109:55]; // @[ifu_aln_ctl.scala 186:25]
  wire [54:0] misc0eff = misceff[54:0]; // @[ifu_aln_ctl.scala 187:25]
  wire  f1dbecc = misc1eff[54]; // @[ifu_aln_ctl.scala 190:25]
  wire  f1icaf = misc1eff[53]; // @[ifu_aln_ctl.scala 191:21]
  wire [1:0] f1ictype = misc1eff[52:51]; // @[ifu_aln_ctl.scala 192:26]
  wire [30:0] f1prett = misc1eff[50:20]; // @[ifu_aln_ctl.scala 193:25]
  wire [11:0] f1poffset = misc1eff[19:8]; // @[ifu_aln_ctl.scala 194:27]
  wire [7:0] f1fghr = misc1eff[7:0]; // @[ifu_aln_ctl.scala 195:24]
  wire  f0dbecc = misc0eff[54]; // @[ifu_aln_ctl.scala 197:25]
  wire  f0icaf = misc0eff[53]; // @[ifu_aln_ctl.scala 198:21]
  wire [1:0] f0ictype = misc0eff[52:51]; // @[ifu_aln_ctl.scala 199:26]
  wire [30:0] f0prett = misc0eff[50:20]; // @[ifu_aln_ctl.scala 200:25]
  wire [11:0] f0poffset = misc0eff[19:8]; // @[ifu_aln_ctl.scala 201:27]
  wire [7:0] f0fghr = misc0eff[7:0]; // @[ifu_aln_ctl.scala 202:24]
  wire [5:0] _T_241 = {io_ifu_bp_hist1_f[0],io_ifu_bp_hist0_f[0],io_ifu_bp_pc4_f[0],io_ifu_bp_way_f[0],io_ifu_bp_valid_f[0],io_ifu_bp_ret_f[0]}; // @[Cat.scala 29:58]
  wire [5:0] _T_246 = {io_ifu_bp_hist1_f[1],io_ifu_bp_hist0_f[1],io_ifu_bp_pc4_f[1],io_ifu_bp_way_f[1],io_ifu_bp_valid_f[1],io_ifu_bp_ret_f[1]}; // @[Cat.scala 29:58]
  wire [23:0] _T_250 = {brdata1,brdata0}; // @[Cat.scala 29:58]
  wire [23:0] _T_253 = {brdata2,brdata1}; // @[Cat.scala 29:58]
  wire [23:0] _T_256 = {brdata0,brdata2}; // @[Cat.scala 29:58]
  wire [23:0] _T_257 = qren[0] ? _T_250 : 24'h0; // @[Mux.scala 27:72]
  wire [23:0] _T_258 = qren[1] ? _T_253 : 24'h0; // @[Mux.scala 27:72]
  wire [23:0] _T_259 = qren[2] ? _T_256 : 24'h0; // @[Mux.scala 27:72]
  wire [23:0] _T_260 = _T_257 | _T_258; // @[Mux.scala 27:72]
  wire [23:0] brdataeff = _T_260 | _T_259; // @[Mux.scala 27:72]
  wire [11:0] brdata0eff = brdataeff[11:0]; // @[ifu_aln_ctl.scala 213:43]
  wire [11:0] brdata1eff = brdataeff[23:12]; // @[ifu_aln_ctl.scala 213:61]
  wire [11:0] _T_267 = q0sel[0] ? brdata0eff : 12'h0; // @[Mux.scala 27:72]
  wire [5:0] _T_268 = q0sel[1] ? brdata0eff[11:6] : 6'h0; // @[Mux.scala 27:72]
  wire [11:0] _GEN_5 = {{6'd0}, _T_268}; // @[Mux.scala 27:72]
  wire [11:0] brdata0final = _T_267 | _GEN_5; // @[Mux.scala 27:72]
  wire [11:0] _T_275 = q1sel[0] ? brdata1eff : 12'h0; // @[Mux.scala 27:72]
  wire [5:0] _T_276 = q1sel[1] ? brdata1eff[11:6] : 6'h0; // @[Mux.scala 27:72]
  wire [11:0] _GEN_6 = {{6'd0}, _T_276}; // @[Mux.scala 27:72]
  wire [11:0] brdata1final = _T_275 | _GEN_6; // @[Mux.scala 27:72]
  wire [1:0] f0ret = {brdata0final[6],brdata0final[0]}; // @[Cat.scala 29:58]
  wire [1:0] f0brend = {brdata0final[7],brdata0final[1]}; // @[Cat.scala 29:58]
  wire [1:0] f0way = {brdata0final[8],brdata0final[2]}; // @[Cat.scala 29:58]
  wire [1:0] f0pc4 = {brdata0final[9],brdata0final[3]}; // @[Cat.scala 29:58]
  wire [1:0] f0hist0 = {brdata0final[10],brdata0final[4]}; // @[Cat.scala 29:58]
  wire [1:0] f0hist1 = {brdata0final[11],brdata0final[5]}; // @[Cat.scala 29:58]
  wire [1:0] f1ret = {brdata1final[6],brdata1final[0]}; // @[Cat.scala 29:58]
  wire [1:0] f1brend = {brdata1final[7],brdata1final[1]}; // @[Cat.scala 29:58]
  wire [1:0] f1way = {brdata1final[8],brdata1final[2]}; // @[Cat.scala 29:58]
  wire [1:0] f1pc4 = {brdata1final[9],brdata1final[3]}; // @[Cat.scala 29:58]
  wire [1:0] f1hist0 = {brdata1final[10],brdata1final[4]}; // @[Cat.scala 29:58]
  wire [1:0] f1hist1 = {brdata1final[11],brdata1final[5]}; // @[Cat.scala 29:58]
  wire  consume_fb0 = _T_351 & f0val[0]; // @[ifu_aln_ctl.scala 237:32]
  wire  consume_fb1 = _T_335 & f1val[0]; // @[ifu_aln_ctl.scala 238:32]
  wire  _T_311 = ~consume_fb1; // @[ifu_aln_ctl.scala 241:39]
  wire  _T_312 = consume_fb0 & _T_311; // @[ifu_aln_ctl.scala 241:37]
  wire  _T_315 = consume_fb0 & consume_fb1; // @[ifu_aln_ctl.scala 242:37]
  wire [30:0] f0pc_plus1 = f0pc + 31'h1; // @[ifu_aln_ctl.scala 259:25]
  wire [30:0] f1pc_plus1 = f1pc + 31'h1; // @[ifu_aln_ctl.scala 261:25]
  wire [30:0] _T_363 = f1_shift_2B ? 31'h7fffffff : 31'h0; // @[Bitwise.scala 72:12]
  wire [30:0] _T_364 = _T_363 & f1pc_plus1; // @[ifu_aln_ctl.scala 263:38]
  wire [30:0] _T_367 = _T_416 ? 31'h7fffffff : 31'h0; // @[Bitwise.scala 72:12]
  wire [30:0] _T_368 = _T_367 & f1pc; // @[ifu_aln_ctl.scala 263:78]
  wire [30:0] sf1pc = _T_364 | _T_368; // @[ifu_aln_ctl.scala 263:52]
  wire  _T_371 = ~fetch_to_f1; // @[ifu_aln_ctl.scala 267:6]
  wire  _T_372 = ~_T_353; // @[ifu_aln_ctl.scala 267:21]
  wire  _T_373 = _T_371 & _T_372; // @[ifu_aln_ctl.scala 267:19]
  wire [30:0] _T_375 = fetch_to_f1 ? io_ifu_fetch_pc : 31'h0; // @[Mux.scala 27:72]
  wire [30:0] _T_376 = _T_353 ? f2pc : 31'h0; // @[Mux.scala 27:72]
  wire [30:0] _T_377 = _T_373 ? sf1pc : 31'h0; // @[Mux.scala 27:72]
  wire [30:0] _T_378 = _T_375 | _T_376; // @[Mux.scala 27:72]
  wire  _T_384 = ~fetch_to_f0; // @[ifu_aln_ctl.scala 272:24]
  wire  _T_385 = ~_T_337; // @[ifu_aln_ctl.scala 272:39]
  wire  _T_386 = _T_384 & _T_385; // @[ifu_aln_ctl.scala 272:37]
  wire  _T_387 = ~_T_352; // @[ifu_aln_ctl.scala 272:54]
  wire  _T_388 = _T_386 & _T_387; // @[ifu_aln_ctl.scala 272:52]
  wire [30:0] _T_390 = fetch_to_f0 ? io_ifu_fetch_pc : 31'h0; // @[Mux.scala 27:72]
  wire [30:0] _T_391 = _T_337 ? f2pc : 31'h0; // @[Mux.scala 27:72]
  wire [30:0] _T_392 = _T_352 ? sf1pc : 31'h0; // @[Mux.scala 27:72]
  wire [30:0] _T_393 = _T_388 ? f0pc_plus1 : 31'h0; // @[Mux.scala 27:72]
  wire [30:0] _T_394 = _T_390 | _T_391; // @[Mux.scala 27:72]
  wire [30:0] _T_395 = _T_394 | _T_392; // @[Mux.scala 27:72]
  wire  _T_399 = fetch_to_f2 & _T_1; // @[ifu_aln_ctl.scala 274:38]
  wire  _T_401 = ~fetch_to_f2; // @[ifu_aln_ctl.scala 275:25]
  wire  _T_403 = _T_401 & _T_372; // @[ifu_aln_ctl.scala 275:38]
  wire  _T_405 = _T_403 & _T_385; // @[ifu_aln_ctl.scala 275:53]
  wire  _T_407 = _T_405 & _T_1; // @[ifu_aln_ctl.scala 275:68]
  wire [1:0] _T_409 = _T_399 ? io_ifu_fetch_val : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_410 = _T_407 ? f2val : 2'h0; // @[Mux.scala 27:72]
  wire  _T_422 = fetch_to_f1 & _T_1; // @[ifu_aln_ctl.scala 279:39]
  wire  _T_425 = _T_353 & _T_1; // @[ifu_aln_ctl.scala 280:54]
  wire  _T_431 = _T_373 & _T_387; // @[ifu_aln_ctl.scala 281:54]
  wire  _T_433 = _T_431 & _T_1; // @[ifu_aln_ctl.scala 281:69]
  wire [1:0] _T_435 = _T_422 ? io_ifu_fetch_val : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_436 = _T_425 ? f2val : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_437 = _T_433 ? sf1val : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_438 = _T_435 | _T_436; // @[Mux.scala 27:72]
  wire  _T_453 = fetch_to_f0 & _T_1; // @[ifu_aln_ctl.scala 286:38]
  wire  _T_456 = _T_337 & _T_1; // @[ifu_aln_ctl.scala 287:54]
  wire  _T_459 = _T_352 & _T_1; // @[ifu_aln_ctl.scala 288:69]
  wire  _T_467 = _T_388 & _T_1; // @[ifu_aln_ctl.scala 289:69]
  wire [1:0] _T_469 = _T_453 ? io_ifu_fetch_val : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_470 = _T_456 ? f2val : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_471 = _T_459 ? sf1val : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_472 = _T_467 ? sf0val : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_473 = _T_469 | _T_470; // @[Mux.scala 27:72]
  wire [1:0] _T_474 = _T_473 | _T_471; // @[Mux.scala 27:72]
  wire [1:0] _T_530 = {f1val[0],1'h1}; // @[Cat.scala 29:58]
  wire [1:0] _T_531 = f0val[1] ? 2'h3 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_532 = _T_515 ? _T_530 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] alignval = _T_531 | _T_532; // @[Mux.scala 27:72]
  wire [1:0] _T_542 = {f1icaf,f0icaf}; // @[Cat.scala 29:58]
  wire  _T_543 = f0val[1] & f0icaf; // @[Mux.scala 27:72]
  wire [1:0] _T_544 = _T_515 ? _T_542 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _GEN_7 = {{1'd0}, _T_543}; // @[Mux.scala 27:72]
  wire [1:0] alignicaf = _GEN_7 | _T_544; // @[Mux.scala 27:72]
  wire [1:0] _T_549 = f0dbecc ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [1:0] _T_555 = {f1dbecc,f0dbecc}; // @[Cat.scala 29:58]
  wire [1:0] _T_556 = f0val[1] ? _T_549 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_557 = _T_515 ? _T_555 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] aligndbecc = _T_556 | _T_557; // @[Mux.scala 27:72]
  wire [1:0] _T_568 = {f1brend[0],f0brend[0]}; // @[Cat.scala 29:58]
  wire [1:0] _T_569 = f0val[1] ? f0brend : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_570 = _T_515 ? _T_568 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] alignbrend = _T_569 | _T_570; // @[Mux.scala 27:72]
  wire [1:0] _T_581 = {f1pc4[0],f0pc4[0]}; // @[Cat.scala 29:58]
  wire [1:0] _T_582 = f0val[1] ? f0pc4 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_583 = _T_515 ? _T_581 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] alignpc4 = _T_582 | _T_583; // @[Mux.scala 27:72]
  wire [1:0] _T_594 = {f1ret[0],f0ret[0]}; // @[Cat.scala 29:58]
  wire [1:0] _T_595 = f0val[1] ? f0ret : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_596 = _T_515 ? _T_594 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] alignret = _T_595 | _T_596; // @[Mux.scala 27:72]
  wire [1:0] _T_607 = {f1way[0],f0way[0]}; // @[Cat.scala 29:58]
  wire [1:0] _T_608 = f0val[1] ? f0way : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_609 = _T_515 ? _T_607 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] alignway = _T_608 | _T_609; // @[Mux.scala 27:72]
  wire [1:0] _T_620 = {f1hist1[0],f0hist1[0]}; // @[Cat.scala 29:58]
  wire [1:0] _T_621 = f0val[1] ? f0hist1 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_622 = _T_515 ? _T_620 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] alignhist1 = _T_621 | _T_622; // @[Mux.scala 27:72]
  wire [1:0] _T_633 = {f1hist0[0],f0hist0[0]}; // @[Cat.scala 29:58]
  wire [1:0] _T_634 = f0val[1] ? f0hist0 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_635 = _T_515 ? _T_633 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] alignhist0 = _T_634 | _T_635; // @[Mux.scala 27:72]
  wire [30:0] _T_647 = f0val[1] ? f0pc_plus1 : 31'h0; // @[Mux.scala 27:72]
  wire [30:0] _T_648 = _T_515 ? f1pc : 31'h0; // @[Mux.scala 27:72]
  wire [30:0] secondpc = _T_647 | _T_648; // @[Mux.scala 27:72]
  wire  _T_657 = first4B & alignval[1]; // @[Mux.scala 27:72]
  wire  _T_658 = first2B & alignval[0]; // @[Mux.scala 27:72]
  wire  _T_662 = |alignicaf; // @[ifu_aln_ctl.scala 340:74]
  wire  _T_665 = first4B & _T_662; // @[Mux.scala 27:72]
  wire  _T_666 = first2B & alignicaf[0]; // @[Mux.scala 27:72]
  wire  _T_671 = first4B & _T_513; // @[ifu_aln_ctl.scala 342:54]
  wire  _T_673 = _T_671 & f0val[0]; // @[ifu_aln_ctl.scala 342:66]
  wire  _T_675 = ~alignicaf[0]; // @[ifu_aln_ctl.scala 342:79]
  wire  _T_676 = _T_673 & _T_675; // @[ifu_aln_ctl.scala 342:77]
  wire  _T_678 = ~aligndbecc[0]; // @[ifu_aln_ctl.scala 342:95]
  wire  _T_679 = _T_676 & _T_678; // @[ifu_aln_ctl.scala 342:93]
  wire  icaf_eff = alignicaf[1] | aligndbecc[1]; // @[ifu_aln_ctl.scala 344:31]
  wire  _T_684 = first4B & icaf_eff; // @[ifu_aln_ctl.scala 346:47]
  wire  _T_687 = |aligndbecc; // @[ifu_aln_ctl.scala 348:74]
  wire  _T_690 = first4B & _T_687; // @[Mux.scala 27:72]
  wire  _T_691 = first2B & aligndbecc[0]; // @[Mux.scala 27:72]
  wire [31:0] _T_696 = first4B ? aligndata : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_697 = first2B ? decompressed_io_dout : 32'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_702 = f0pc[8:1] ^ f0pc[16:9]; // @[lib.scala 51:47]
  wire [7:0] firstpc_hash = _T_702 ^ f0pc[24:17]; // @[lib.scala 51:85]
  wire [7:0] _T_706 = secondpc[8:1] ^ secondpc[16:9]; // @[lib.scala 51:47]
  wire [7:0] secondpc_hash = _T_706 ^ secondpc[24:17]; // @[lib.scala 51:85]
  wire [4:0] _T_712 = f0pc[13:9] ^ f0pc[18:14]; // @[lib.scala 42:111]
  wire [4:0] firstbrtag_hash = _T_712 ^ f0pc[23:19]; // @[lib.scala 42:111]
  wire [4:0] _T_717 = secondpc[13:9] ^ secondpc[18:14]; // @[lib.scala 42:111]
  wire [4:0] secondbrtag_hash = _T_717 ^ secondpc[23:19]; // @[lib.scala 42:111]
  wire  _T_719 = first2B & alignbrend[0]; // @[ifu_aln_ctl.scala 365:45]
  wire  _T_721 = first4B & alignbrend[1]; // @[ifu_aln_ctl.scala 365:73]
  wire  _T_722 = _T_719 | _T_721; // @[ifu_aln_ctl.scala 365:62]
  wire  _T_726 = _T_657 & alignbrend[0]; // @[ifu_aln_ctl.scala 365:115]
  wire  _T_729 = first2B & alignret[0]; // @[ifu_aln_ctl.scala 367:49]
  wire  _T_731 = first4B & alignret[1]; // @[ifu_aln_ctl.scala 367:75]
  wire  _T_734 = first2B & alignpc4[0]; // @[ifu_aln_ctl.scala 369:29]
  wire  _T_736 = first4B & alignpc4[1]; // @[ifu_aln_ctl.scala 369:55]
  wire  i0_brp_pc4 = _T_734 | _T_736; // @[ifu_aln_ctl.scala 369:44]
  wire  _T_738 = first2B | alignbrend[0]; // @[ifu_aln_ctl.scala 371:53]
  wire  _T_744 = first2B & alignhist1[0]; // @[ifu_aln_ctl.scala 373:54]
  wire  _T_746 = first4B & alignhist1[1]; // @[ifu_aln_ctl.scala 373:82]
  wire  _T_747 = _T_744 | _T_746; // @[ifu_aln_ctl.scala 373:71]
  wire  _T_749 = first2B & alignhist0[0]; // @[ifu_aln_ctl.scala 374:14]
  wire  _T_751 = first4B & alignhist0[1]; // @[ifu_aln_ctl.scala 374:42]
  wire  _T_752 = _T_749 | _T_751; // @[ifu_aln_ctl.scala 374:31]
  wire  i0_ends_f1 = first4B & _T_515; // @[ifu_aln_ctl.scala 376:28]
  wire  _T_768 = io_dec_aln_aln_ib_i0_brp_valid & i0_brp_pc4; // @[ifu_aln_ctl.scala 385:77]
  wire  _T_769 = _T_768 & first2B; // @[ifu_aln_ctl.scala 385:91]
  wire  _T_770 = ~i0_brp_pc4; // @[ifu_aln_ctl.scala 385:139]
  wire  _T_771 = io_dec_aln_aln_ib_i0_brp_valid & _T_770; // @[ifu_aln_ctl.scala 385:137]
  wire  _T_772 = _T_771 & first4B; // @[ifu_aln_ctl.scala 385:151]
  rvclkhdr rvclkhdr ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_io_l1clk),
    .io_clk(rvclkhdr_io_clk),
    .io_en(rvclkhdr_io_en),
    .io_scan_mode(rvclkhdr_io_scan_mode)
  );
  rvclkhdr rvclkhdr_1 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_1_io_l1clk),
    .io_clk(rvclkhdr_1_io_clk),
    .io_en(rvclkhdr_1_io_en),
    .io_scan_mode(rvclkhdr_1_io_scan_mode)
  );
  rvclkhdr rvclkhdr_2 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_2_io_l1clk),
    .io_clk(rvclkhdr_2_io_clk),
    .io_en(rvclkhdr_2_io_en),
    .io_scan_mode(rvclkhdr_2_io_scan_mode)
  );
  rvclkhdr rvclkhdr_3 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_3_io_l1clk),
    .io_clk(rvclkhdr_3_io_clk),
    .io_en(rvclkhdr_3_io_en),
    .io_scan_mode(rvclkhdr_3_io_scan_mode)
  );
  rvclkhdr rvclkhdr_4 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_4_io_l1clk),
    .io_clk(rvclkhdr_4_io_clk),
    .io_en(rvclkhdr_4_io_en),
    .io_scan_mode(rvclkhdr_4_io_scan_mode)
  );
  rvclkhdr rvclkhdr_5 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_5_io_l1clk),
    .io_clk(rvclkhdr_5_io_clk),
    .io_en(rvclkhdr_5_io_en),
    .io_scan_mode(rvclkhdr_5_io_scan_mode)
  );
  rvclkhdr rvclkhdr_6 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_6_io_l1clk),
    .io_clk(rvclkhdr_6_io_clk),
    .io_en(rvclkhdr_6_io_en),
    .io_scan_mode(rvclkhdr_6_io_scan_mode)
  );
  rvclkhdr rvclkhdr_7 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_7_io_l1clk),
    .io_clk(rvclkhdr_7_io_clk),
    .io_en(rvclkhdr_7_io_en),
    .io_scan_mode(rvclkhdr_7_io_scan_mode)
  );
  rvclkhdr rvclkhdr_8 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_8_io_l1clk),
    .io_clk(rvclkhdr_8_io_clk),
    .io_en(rvclkhdr_8_io_en),
    .io_scan_mode(rvclkhdr_8_io_scan_mode)
  );
  rvclkhdr rvclkhdr_9 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_9_io_l1clk),
    .io_clk(rvclkhdr_9_io_clk),
    .io_en(rvclkhdr_9_io_en),
    .io_scan_mode(rvclkhdr_9_io_scan_mode)
  );
  rvclkhdr rvclkhdr_10 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_10_io_l1clk),
    .io_clk(rvclkhdr_10_io_clk),
    .io_en(rvclkhdr_10_io_en),
    .io_scan_mode(rvclkhdr_10_io_scan_mode)
  );
  rvclkhdr rvclkhdr_11 ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_11_io_l1clk),
    .io_clk(rvclkhdr_11_io_clk),
    .io_en(rvclkhdr_11_io_en),
    .io_scan_mode(rvclkhdr_11_io_scan_mode)
  );
  ifu_compress_ctl decompressed ( // @[ifu_aln_ctl.scala 352:28]
    .io_din(decompressed_io_din),
    .io_dout(decompressed_io_dout)
  );
  assign io_dec_aln_aln_dec_ifu_i0_cinst = aligndata[15:0]; // @[ifu_aln_ctl.scala 331:35]
  assign io_dec_aln_aln_ib_ifu_i0_icaf = _T_665 | _T_666; // @[ifu_aln_ctl.scala 340:33]
  assign io_dec_aln_aln_ib_ifu_i0_icaf_type = _T_679 ? f1ictype : f0ictype; // @[ifu_aln_ctl.scala 342:38]
  assign io_dec_aln_aln_ib_ifu_i0_icaf_f1 = _T_684 & _T_515; // @[ifu_aln_ctl.scala 346:36]
  assign io_dec_aln_aln_ib_ifu_i0_dbecc = _T_690 | _T_691; // @[ifu_aln_ctl.scala 348:34]
  assign io_dec_aln_aln_ib_ifu_i0_bp_index = _T_738 ? firstpc_hash : secondpc_hash; // @[ifu_aln_ctl.scala 387:37]
  assign io_dec_aln_aln_ib_ifu_i0_bp_fghr = i0_ends_f1 ? f1fghr : f0fghr; // @[ifu_aln_ctl.scala 389:36]
  assign io_dec_aln_aln_ib_ifu_i0_bp_btag = _T_738 ? firstbrtag_hash : secondbrtag_hash; // @[ifu_aln_ctl.scala 391:36]
  assign io_dec_aln_aln_ib_ifu_i0_valid = _T_657 | _T_658; // @[ifu_aln_ctl.scala 338:34]
  assign io_dec_aln_aln_ib_ifu_i0_instr = _T_696 | _T_697; // @[ifu_aln_ctl.scala 354:34]
  assign io_dec_aln_aln_ib_ifu_i0_pc = f0pc; // @[ifu_aln_ctl.scala 325:31]
  assign io_dec_aln_aln_ib_ifu_i0_pc4 = aligndata[1:0] == 2'h3; // @[ifu_aln_ctl.scala 329:32]
  assign io_dec_aln_aln_ib_i0_brp_valid = _T_722 | _T_726; // @[ifu_aln_ctl.scala 365:34]
  assign io_dec_aln_aln_ib_i0_brp_bits_toffset = i0_ends_f1 ? f1poffset : f0poffset; // @[ifu_aln_ctl.scala 377:41]
  assign io_dec_aln_aln_ib_i0_brp_bits_hist = {_T_747,_T_752}; // @[ifu_aln_ctl.scala 373:38]
  assign io_dec_aln_aln_ib_i0_brp_bits_br_error = _T_769 | _T_772; // @[ifu_aln_ctl.scala 385:42]
  assign io_dec_aln_aln_ib_i0_brp_bits_br_start_error = _T_657 & alignbrend[0]; // @[ifu_aln_ctl.scala 381:49]
  assign io_dec_aln_aln_ib_i0_brp_bits_bank = _T_738 ? f0pc[0] : secondpc[0]; // @[ifu_aln_ctl.scala 383:49]
  assign io_dec_aln_aln_ib_i0_brp_bits_prett = i0_ends_f1 ? f1prett : f0prett; // @[ifu_aln_ctl.scala 379:39]
  assign io_dec_aln_aln_ib_i0_brp_bits_way = _T_738 ? alignway[0] : alignway[1]; // @[ifu_aln_ctl.scala 371:37]
  assign io_dec_aln_aln_ib_i0_brp_bits_ret = _T_729 | _T_731; // @[ifu_aln_ctl.scala 367:37]
  assign io_dec_aln_ifu_pmu_instr_aligned = io_dec_aln_aln_dec_dec_i0_decode_d & _T_785; // @[ifu_aln_ctl.scala 397:36]
  assign io_ifu_fb_consume1 = _T_312 & _T_1; // @[ifu_aln_ctl.scala 241:22]
  assign io_ifu_fb_consume2 = _T_315 & _T_1; // @[ifu_aln_ctl.scala 242:22]
  assign rvclkhdr_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_io_en = _T_354 | _T_358; // @[lib.scala 371:17]
  assign rvclkhdr_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_1_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_1_io_en = _T_25 | f1_shift_2B; // @[lib.scala 371:17]
  assign rvclkhdr_1_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_2_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_2_io_en = _T_29 | shift_4B; // @[lib.scala 371:17]
  assign rvclkhdr_2_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_3_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_3_io_en = qwen[2]; // @[lib.scala 371:17]
  assign rvclkhdr_3_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_4_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_4_io_en = qwen[1]; // @[lib.scala 371:17]
  assign rvclkhdr_4_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_5_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_5_io_en = qwen[0]; // @[lib.scala 371:17]
  assign rvclkhdr_5_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_6_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_6_io_en = qwen[2]; // @[lib.scala 371:17]
  assign rvclkhdr_6_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_7_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_7_io_en = qwen[1]; // @[lib.scala 371:17]
  assign rvclkhdr_7_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_8_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_8_io_en = qwen[0]; // @[lib.scala 371:17]
  assign rvclkhdr_8_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_9_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_9_io_en = qwen[2]; // @[lib.scala 371:17]
  assign rvclkhdr_9_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_10_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_10_io_en = qwen[1]; // @[lib.scala 371:17]
  assign rvclkhdr_10_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign rvclkhdr_11_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_11_io_en = qwen[0]; // @[lib.scala 371:17]
  assign rvclkhdr_11_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
  assign decompressed_io_din = aligndata[15:0]; // @[ifu_aln_ctl.scala 393:23]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  error_stall = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  wrptr = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  rdptr = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  f2val = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  f1val = _RAND_4[1:0];
  _RAND_5 = {1{`RANDOM}};
  f0val = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  q2off = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  q1off = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  q0off = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  q1 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  q0 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  q2 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  f2pc = _RAND_12[30:0];
  _RAND_13 = {1{`RANDOM}};
  f1pc = _RAND_13[30:0];
  _RAND_14 = {1{`RANDOM}};
  f0pc = _RAND_14[30:0];
  _RAND_15 = {1{`RANDOM}};
  brdata2 = _RAND_15[11:0];
  _RAND_16 = {1{`RANDOM}};
  brdata1 = _RAND_16[11:0];
  _RAND_17 = {1{`RANDOM}};
  brdata0 = _RAND_17[11:0];
  _RAND_18 = {2{`RANDOM}};
  misc2 = _RAND_18[54:0];
  _RAND_19 = {2{`RANDOM}};
  misc1 = _RAND_19[54:0];
  _RAND_20 = {2{`RANDOM}};
  misc0 = _RAND_20[54:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    error_stall = 1'h0;
  end
  if (reset) begin
    wrptr = 2'h0;
  end
  if (reset) begin
    rdptr = 2'h0;
  end
  if (reset) begin
    f2val = 2'h0;
  end
  if (reset) begin
    f1val = 2'h0;
  end
  if (reset) begin
    f0val = 2'h0;
  end
  if (reset) begin
    q2off = 1'h0;
  end
  if (reset) begin
    q1off = 1'h0;
  end
  if (reset) begin
    q0off = 1'h0;
  end
  if (reset) begin
    q1 = 32'h0;
  end
  if (reset) begin
    q0 = 32'h0;
  end
  if (reset) begin
    q2 = 32'h0;
  end
  if (reset) begin
    f2pc = 31'h0;
  end
  if (reset) begin
    f1pc = 31'h0;
  end
  if (reset) begin
    f0pc = 31'h0;
  end
  if (reset) begin
    brdata2 = 12'h0;
  end
  if (reset) begin
    brdata1 = 12'h0;
  end
  if (reset) begin
    brdata0 = 12'h0;
  end
  if (reset) begin
    misc2 = 55'h0;
  end
  if (reset) begin
    misc1 = 55'h0;
  end
  if (reset) begin
    misc0 = 55'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      error_stall <= 1'h0;
    end else begin
      error_stall <= _T & _T_1;
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      wrptr <= 2'h0;
    end else begin
      wrptr <= _T_113 | _T_112;
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      rdptr <= 2'h0;
    end else begin
      rdptr <= _T_90 | _T_85;
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      f2val <= 2'h0;
    end else begin
      f2val <= _T_409 | _T_410;
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      f1val <= 2'h0;
    end else begin
      f1val <= _T_438 | _T_437;
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      f0val <= 2'h0;
    end else begin
      f0val <= _T_474 | _T_472;
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      q2off <= 1'h0;
    end else begin
      q2off <= _T_137 | _T_136;
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      q1off <= 1'h0;
    end else begin
      q1off <= _T_160 | _T_159;
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      q0off <= 1'h0;
    end else begin
      q0off <= _T_183 | _T_182;
    end
  end
  always @(posedge rvclkhdr_10_io_l1clk or posedge reset) begin
    if (reset) begin
      q1 <= 32'h0;
    end else begin
      q1 <= io_ifu_fetch_data_f;
    end
  end
  always @(posedge rvclkhdr_11_io_l1clk or posedge reset) begin
    if (reset) begin
      q0 <= 32'h0;
    end else begin
      q0 <= io_ifu_fetch_data_f;
    end
  end
  always @(posedge rvclkhdr_9_io_l1clk or posedge reset) begin
    if (reset) begin
      q2 <= 32'h0;
    end else begin
      q2 <= io_ifu_fetch_data_f;
    end
  end
  always @(posedge rvclkhdr_io_l1clk or posedge reset) begin
    if (reset) begin
      f2pc <= 31'h0;
    end else begin
      f2pc <= io_ifu_fetch_pc;
    end
  end
  always @(posedge rvclkhdr_1_io_l1clk or posedge reset) begin
    if (reset) begin
      f1pc <= 31'h0;
    end else begin
      f1pc <= _T_378 | _T_377;
    end
  end
  always @(posedge rvclkhdr_2_io_l1clk or posedge reset) begin
    if (reset) begin
      f0pc <= 31'h0;
    end else begin
      f0pc <= _T_395 | _T_393;
    end
  end
  always @(posedge rvclkhdr_3_io_l1clk or posedge reset) begin
    if (reset) begin
      brdata2 <= 12'h0;
    end else begin
      brdata2 <= {_T_246,_T_241};
    end
  end
  always @(posedge rvclkhdr_4_io_l1clk or posedge reset) begin
    if (reset) begin
      brdata1 <= 12'h0;
    end else begin
      brdata1 <= {_T_246,_T_241};
    end
  end
  always @(posedge rvclkhdr_5_io_l1clk or posedge reset) begin
    if (reset) begin
      brdata0 <= 12'h0;
    end else begin
      brdata0 <= {_T_246,_T_241};
    end
  end
  always @(posedge rvclkhdr_6_io_l1clk or posedge reset) begin
    if (reset) begin
      misc2 <= 55'h0;
    end else begin
      misc2 <= {_T_207,_T_205};
    end
  end
  always @(posedge rvclkhdr_7_io_l1clk or posedge reset) begin
    if (reset) begin
      misc1 <= 55'h0;
    end else begin
      misc1 <= {_T_207,_T_205};
    end
  end
  always @(posedge rvclkhdr_8_io_l1clk or posedge reset) begin
    if (reset) begin
      misc0 <= 55'h0;
    end else begin
      misc0 <= {_T_207,_T_205};
    end
  end
endmodule
module ifu_ifc_ctl(
  input         clock,
  input         reset,
  input         io_exu_flush_final,
  input  [30:0] io_exu_flush_path_final,
  input         io_free_clk,
  input         io_active_clk,
  input         io_scan_mode,
  input         io_ic_hit_f,
  input         io_ifu_ic_mb_empty,
  input         io_ifu_fb_consume1,
  input         io_ifu_fb_consume2,
  input         io_ifu_bp_hit_taken_f,
  input  [30:0] io_ifu_bp_btb_target_f,
  input         io_ic_dma_active,
  input         io_ic_write_stall,
  input         io_dec_ifc_dec_tlu_flush_noredir_wb,
  input  [31:0] io_dec_ifc_dec_tlu_mrac_ff,
  output        io_dec_ifc_ifu_pmu_fetch_stall,
  input         io_dma_ifc_dma_iccm_stall_any,
  output [30:0] io_ifc_fetch_addr_f,
  output [30:0] io_ifc_fetch_addr_bf,
  output        io_ifc_fetch_req_f,
  output        io_ifc_fetch_uncacheable_bf,
  output        io_ifc_fetch_req_bf,
  output        io_ifc_fetch_req_bf_raw,
  output        io_ifc_iccm_access_bf,
  output        io_ifc_region_acc_fault_bf,
  output        io_ifc_dma_access_ok
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  wire  rvclkhdr_io_l1clk; // @[lib.scala 368:23]
  wire  rvclkhdr_io_clk; // @[lib.scala 368:23]
  wire  rvclkhdr_io_en; // @[lib.scala 368:23]
  wire  rvclkhdr_io_scan_mode; // @[lib.scala 368:23]
  reg  dma_iccm_stall_any_f; // @[ifu_ifc_ctl.scala 63:58]
  wire  dma_stall = io_ic_dma_active | dma_iccm_stall_any_f; // @[ifu_ifc_ctl.scala 62:36]
  reg  miss_a; // @[ifu_ifc_ctl.scala 65:44]
  wire  _T_2 = ~io_exu_flush_final; // @[ifu_ifc_ctl.scala 67:26]
  wire  _T_3 = ~io_ifc_fetch_req_f; // @[ifu_ifc_ctl.scala 67:49]
  wire  _T_4 = ~io_ic_hit_f; // @[ifu_ifc_ctl.scala 67:71]
  wire  _T_5 = _T_3 | _T_4; // @[ifu_ifc_ctl.scala 67:69]
  wire  sel_last_addr_bf = _T_2 & _T_5; // @[ifu_ifc_ctl.scala 67:46]
  wire  _T_7 = _T_2 & io_ifc_fetch_req_f; // @[ifu_ifc_ctl.scala 68:46]
  wire  _T_8 = _T_7 & io_ifu_bp_hit_taken_f; // @[ifu_ifc_ctl.scala 68:67]
  wire  sel_btb_addr_bf = _T_8 & io_ic_hit_f; // @[ifu_ifc_ctl.scala 68:92]
  wire  _T_11 = ~io_ifu_bp_hit_taken_f; // @[ifu_ifc_ctl.scala 69:69]
  wire  _T_12 = _T_7 & _T_11; // @[ifu_ifc_ctl.scala 69:67]
  wire  sel_next_addr_bf = _T_12 & io_ic_hit_f; // @[ifu_ifc_ctl.scala 69:92]
  wire [30:0] _T_17 = io_exu_flush_final ? io_exu_flush_path_final : 31'h0; // @[Mux.scala 27:72]
  wire [30:0] _T_18 = sel_last_addr_bf ? io_ifc_fetch_addr_f : 31'h0; // @[Mux.scala 27:72]
  wire [30:0] _T_19 = sel_btb_addr_bf ? io_ifu_bp_btb_target_f : 31'h0; // @[Mux.scala 27:72]
  wire [29:0] address_upper = io_ifc_fetch_addr_f[30:1] + 30'h1; // @[ifu_ifc_ctl.scala 78:48]
  wire  _T_29 = address_upper[4] ^ io_ifc_fetch_addr_f[5]; // @[ifu_ifc_ctl.scala 79:63]
  wire  _T_30 = ~_T_29; // @[ifu_ifc_ctl.scala 79:24]
  wire  fetch_addr_next_0 = _T_30 & io_ifc_fetch_addr_f[0]; // @[ifu_ifc_ctl.scala 79:109]
  wire [30:0] fetch_addr_next = {address_upper,fetch_addr_next_0}; // @[Cat.scala 29:58]
  wire [30:0] _T_20 = sel_next_addr_bf ? fetch_addr_next : 31'h0; // @[Mux.scala 27:72]
  wire [30:0] _T_21 = _T_17 | _T_18; // @[Mux.scala 27:72]
  wire [30:0] _T_22 = _T_21 | _T_19; // @[Mux.scala 27:72]
  reg [1:0] state; // @[ifu_ifc_ctl.scala 104:45]
  wire  idle = state == 2'h0; // @[ifu_ifc_ctl.scala 123:17]
  wire  _T_35 = io_ifu_fb_consume2 | io_ifu_fb_consume1; // @[ifu_ifc_ctl.scala 86:91]
  wire  _T_36 = ~_T_35; // @[ifu_ifc_ctl.scala 86:70]
  wire [3:0] _T_121 = io_exu_flush_final ? 4'h1 : 4'h0; // @[Mux.scala 27:72]
  wire  _T_81 = ~io_ifu_fb_consume2; // @[ifu_ifc_ctl.scala 109:38]
  wire  _T_82 = io_ifu_fb_consume1 & _T_81; // @[ifu_ifc_ctl.scala 109:36]
  wire  _T_48 = io_ifc_fetch_req_f & _T_4; // @[ifu_ifc_ctl.scala 91:32]
  wire  miss_f = _T_48 & _T_2; // @[ifu_ifc_ctl.scala 91:47]
  wire  _T_84 = _T_3 | miss_f; // @[ifu_ifc_ctl.scala 109:81]
  wire  _T_85 = _T_82 & _T_84; // @[ifu_ifc_ctl.scala 109:58]
  wire  _T_86 = io_ifu_fb_consume2 & io_ifc_fetch_req_f; // @[ifu_ifc_ctl.scala 110:25]
  wire  fb_right = _T_85 | _T_86; // @[ifu_ifc_ctl.scala 109:92]
  wire  _T_98 = _T_2 & fb_right; // @[ifu_ifc_ctl.scala 117:16]
  reg [3:0] fb_write_f; // @[ifu_ifc_ctl.scala 128:50]
  wire [3:0] _T_101 = {1'h0,fb_write_f[3:1]}; // @[Cat.scala 29:58]
  wire [3:0] _T_122 = _T_98 ? _T_101 : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_126 = _T_121 | _T_122; // @[Mux.scala 27:72]
  wire  fb_right2 = io_ifu_fb_consume2 & _T_84; // @[ifu_ifc_ctl.scala 112:36]
  wire  _T_103 = _T_2 & fb_right2; // @[ifu_ifc_ctl.scala 118:16]
  wire [3:0] _T_106 = {2'h0,fb_write_f[3:2]}; // @[Cat.scala 29:58]
  wire [3:0] _T_123 = _T_103 ? _T_106 : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_127 = _T_126 | _T_123; // @[Mux.scala 27:72]
  wire  _T_91 = io_ifu_fb_consume1 | io_ifu_fb_consume2; // @[ifu_ifc_ctl.scala 113:56]
  wire  _T_92 = ~_T_91; // @[ifu_ifc_ctl.scala 113:35]
  wire  _T_93 = io_ifc_fetch_req_f & _T_92; // @[ifu_ifc_ctl.scala 113:33]
  wire  _T_94 = ~miss_f; // @[ifu_ifc_ctl.scala 113:80]
  wire  fb_left = _T_93 & _T_94; // @[ifu_ifc_ctl.scala 113:78]
  wire  _T_108 = _T_2 & fb_left; // @[ifu_ifc_ctl.scala 119:16]
  wire [3:0] _T_111 = {fb_write_f[2:0],1'h0}; // @[Cat.scala 29:58]
  wire [3:0] _T_124 = _T_108 ? _T_111 : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_128 = _T_127 | _T_124; // @[Mux.scala 27:72]
  wire  _T_113 = ~fb_right; // @[ifu_ifc_ctl.scala 120:18]
  wire  _T_114 = _T_2 & _T_113; // @[ifu_ifc_ctl.scala 120:16]
  wire  _T_115 = ~fb_right2; // @[ifu_ifc_ctl.scala 120:30]
  wire  _T_116 = _T_114 & _T_115; // @[ifu_ifc_ctl.scala 120:28]
  wire  _T_117 = ~fb_left; // @[ifu_ifc_ctl.scala 120:43]
  wire  _T_118 = _T_116 & _T_117; // @[ifu_ifc_ctl.scala 120:41]
  wire [3:0] _T_125 = _T_118 ? fb_write_f : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] fb_write_ns = _T_128 | _T_125; // @[Mux.scala 27:72]
  wire  fb_full_f_ns = fb_write_ns[3]; // @[ifu_ifc_ctl.scala 126:30]
  wire  _T_37 = fb_full_f_ns & _T_36; // @[ifu_ifc_ctl.scala 86:68]
  wire  _T_38 = ~_T_37; // @[ifu_ifc_ctl.scala 86:53]
  wire  _T_39 = io_ifc_fetch_req_bf_raw & _T_38; // @[ifu_ifc_ctl.scala 86:51]
  wire  _T_40 = ~dma_stall; // @[ifu_ifc_ctl.scala 87:5]
  wire  _T_41 = _T_39 & _T_40; // @[ifu_ifc_ctl.scala 86:114]
  wire  _T_42 = ~io_ic_write_stall; // @[ifu_ifc_ctl.scala 87:18]
  wire  _T_43 = _T_41 & _T_42; // @[ifu_ifc_ctl.scala 87:16]
  wire  _T_44 = ~io_dec_ifc_dec_tlu_flush_noredir_wb; // @[ifu_ifc_ctl.scala 87:39]
  wire  _T_51 = io_ifu_ic_mb_empty | io_exu_flush_final; // @[ifu_ifc_ctl.scala 93:39]
  wire  _T_53 = _T_51 & _T_40; // @[ifu_ifc_ctl.scala 93:61]
  wire  _T_55 = _T_53 & _T_94; // @[ifu_ifc_ctl.scala 93:74]
  wire  _T_56 = ~miss_a; // @[ifu_ifc_ctl.scala 93:86]
  wire  mb_empty_mod = _T_55 & _T_56; // @[ifu_ifc_ctl.scala 93:84]
  wire  goto_idle = io_exu_flush_final & io_dec_ifc_dec_tlu_flush_noredir_wb; // @[ifu_ifc_ctl.scala 95:35]
  wire  _T_60 = io_exu_flush_final & _T_44; // @[ifu_ifc_ctl.scala 97:36]
  wire  leave_idle = _T_60 & idle; // @[ifu_ifc_ctl.scala 97:75]
  wire  _T_63 = ~state[1]; // @[ifu_ifc_ctl.scala 99:23]
  wire  _T_65 = _T_63 & state[0]; // @[ifu_ifc_ctl.scala 99:33]
  wire  _T_66 = _T_65 & miss_f; // @[ifu_ifc_ctl.scala 99:44]
  wire  _T_67 = ~goto_idle; // @[ifu_ifc_ctl.scala 99:55]
  wire  _T_68 = _T_66 & _T_67; // @[ifu_ifc_ctl.scala 99:53]
  wire  _T_70 = ~mb_empty_mod; // @[ifu_ifc_ctl.scala 100:17]
  wire  _T_71 = state[1] & _T_70; // @[ifu_ifc_ctl.scala 100:15]
  wire  _T_73 = _T_71 & _T_67; // @[ifu_ifc_ctl.scala 100:31]
  wire  next_state_1 = _T_68 | _T_73; // @[ifu_ifc_ctl.scala 99:67]
  wire  _T_75 = _T_67 & leave_idle; // @[ifu_ifc_ctl.scala 102:34]
  wire  _T_78 = state[0] & _T_67; // @[ifu_ifc_ctl.scala 102:60]
  wire  next_state_0 = _T_75 | _T_78; // @[ifu_ifc_ctl.scala 102:48]
  wire  wfm = state == 2'h3; // @[ifu_ifc_ctl.scala 124:16]
  reg  fb_full_f; // @[ifu_ifc_ctl.scala 127:52]
  wire  _T_136 = _T_35 | io_exu_flush_final; // @[ifu_ifc_ctl.scala 131:61]
  wire  _T_137 = ~_T_136; // @[ifu_ifc_ctl.scala 131:19]
  wire  _T_138 = fb_full_f & _T_137; // @[ifu_ifc_ctl.scala 131:17]
  wire  _T_139 = _T_138 | dma_stall; // @[ifu_ifc_ctl.scala 131:84]
  wire  _T_140 = io_ifc_fetch_req_bf_raw & _T_139; // @[ifu_ifc_ctl.scala 130:68]
  wire [31:0] _T_142 = {io_ifc_fetch_addr_bf,1'h0}; // @[Cat.scala 29:58]
  wire  iccm_acc_in_region_bf = _T_142[31:28] == 4'he; // @[lib.scala 84:47]
  wire  iccm_acc_in_range_bf = _T_142[31:16] == 16'hee00; // @[lib.scala 87:29]
  wire  _T_145 = ~io_ifc_iccm_access_bf; // @[ifu_ifc_ctl.scala 138:30]
  wire  _T_148 = fb_full_f & _T_36; // @[ifu_ifc_ctl.scala 139:16]
  wire  _T_149 = _T_145 | _T_148; // @[ifu_ifc_ctl.scala 138:53]
  wire  _T_150 = ~io_ifc_fetch_req_bf; // @[ifu_ifc_ctl.scala 140:13]
  wire  _T_151 = wfm & _T_150; // @[ifu_ifc_ctl.scala 140:11]
  wire  _T_152 = _T_149 | _T_151; // @[ifu_ifc_ctl.scala 139:62]
  wire  _T_153 = _T_152 | idle; // @[ifu_ifc_ctl.scala 140:35]
  wire  _T_155 = _T_153 & _T_2; // @[ifu_ifc_ctl.scala 140:44]
  wire  _T_157 = ~iccm_acc_in_range_bf; // @[ifu_ifc_ctl.scala 142:33]
  wire [4:0] _T_160 = {io_ifc_fetch_addr_bf[30:27],1'h0}; // @[Cat.scala 29:58]
  wire [31:0] _T_161 = io_dec_ifc_dec_tlu_mrac_ff >> _T_160; // @[ifu_ifc_ctl.scala 143:61]
  reg  _T_164; // @[ifu_ifc_ctl.scala 145:57]
  reg [30:0] _T_166; // @[lib.scala 374:16]
  rvclkhdr rvclkhdr ( // @[lib.scala 368:23]
    .io_l1clk(rvclkhdr_io_l1clk),
    .io_clk(rvclkhdr_io_clk),
    .io_en(rvclkhdr_io_en),
    .io_scan_mode(rvclkhdr_io_scan_mode)
  );
  assign io_dec_ifc_ifu_pmu_fetch_stall = wfm | _T_140; // @[ifu_ifc_ctl.scala 130:34]
  assign io_ifc_fetch_addr_f = _T_166; // @[ifu_ifc_ctl.scala 147:23]
  assign io_ifc_fetch_addr_bf = _T_22 | _T_20; // @[ifu_ifc_ctl.scala 73:24]
  assign io_ifc_fetch_req_f = _T_164; // @[ifu_ifc_ctl.scala 145:22]
  assign io_ifc_fetch_uncacheable_bf = ~_T_161[0]; // @[ifu_ifc_ctl.scala 143:31]
  assign io_ifc_fetch_req_bf = _T_43 & _T_44; // @[ifu_ifc_ctl.scala 86:23]
  assign io_ifc_fetch_req_bf_raw = ~idle; // @[ifu_ifc_ctl.scala 84:27]
  assign io_ifc_iccm_access_bf = _T_142[31:16] == 16'hee00; // @[ifu_ifc_ctl.scala 137:25]
  assign io_ifc_region_acc_fault_bf = _T_157 & iccm_acc_in_region_bf; // @[ifu_ifc_ctl.scala 142:30]
  assign io_ifc_dma_access_ok = _T_155 | dma_iccm_stall_any_f; // @[ifu_ifc_ctl.scala 138:24]
  assign rvclkhdr_io_clk = clock; // @[lib.scala 370:18]
  assign rvclkhdr_io_en = io_exu_flush_final | io_ifc_fetch_req_f; // @[lib.scala 371:17]
  assign rvclkhdr_io_scan_mode = io_scan_mode; // @[lib.scala 372:24]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  dma_iccm_stall_any_f = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  miss_a = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  state = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  fb_write_f = _RAND_3[3:0];
  _RAND_4 = {1{`RANDOM}};
  fb_full_f = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  _T_164 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  _T_166 = _RAND_6[30:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    dma_iccm_stall_any_f = 1'h0;
  end
  if (reset) begin
    miss_a = 1'h0;
  end
  if (reset) begin
    state = 2'h0;
  end
  if (reset) begin
    fb_write_f = 4'h0;
  end
  if (reset) begin
    fb_full_f = 1'h0;
  end
  if (reset) begin
    _T_164 = 1'h0;
  end
  if (reset) begin
    _T_166 = 31'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      dma_iccm_stall_any_f <= 1'h0;
    end else begin
      dma_iccm_stall_any_f <= io_dma_ifc_dma_iccm_stall_any;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      miss_a <= 1'h0;
    end else begin
      miss_a <= _T_48 & _T_2;
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      state <= 2'h0;
    end else begin
      state <= {next_state_1,next_state_0};
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      fb_write_f <= 4'h0;
    end else begin
      fb_write_f <= _T_128 | _T_125;
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      fb_full_f <= 1'h0;
    end else begin
      fb_full_f <= fb_write_ns[3];
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      _T_164 <= 1'h0;
    end else begin
      _T_164 <= io_ifc_fetch_req_bf;
    end
  end
  always @(posedge rvclkhdr_io_l1clk or posedge reset) begin
    if (reset) begin
      _T_166 <= 31'h0;
    end else begin
      _T_166 <= io_ifc_fetch_addr_bf;
    end
  end
endmodule
module ifu(
  input         clock,
  input         reset,
  input         io_exu_flush_final,
  input  [30:0] io_exu_flush_path_final,
  input         io_free_clk,
  input         io_active_clk,
  input         io_ifu_dec_dec_aln_aln_dec_dec_i0_decode_d,
  output [15:0] io_ifu_dec_dec_aln_aln_dec_ifu_i0_cinst,
  output        io_ifu_dec_dec_aln_aln_ib_ifu_i0_icaf,
  output [1:0]  io_ifu_dec_dec_aln_aln_ib_ifu_i0_icaf_type,
  output        io_ifu_dec_dec_aln_aln_ib_ifu_i0_icaf_f1,
  output        io_ifu_dec_dec_aln_aln_ib_ifu_i0_dbecc,
  output [7:0]  io_ifu_dec_dec_aln_aln_ib_ifu_i0_bp_index,
  output [7:0]  io_ifu_dec_dec_aln_aln_ib_ifu_i0_bp_fghr,
  output [4:0]  io_ifu_dec_dec_aln_aln_ib_ifu_i0_bp_btag,
  output        io_ifu_dec_dec_aln_aln_ib_ifu_i0_valid,
  output [31:0] io_ifu_dec_dec_aln_aln_ib_ifu_i0_instr,
  output [30:0] io_ifu_dec_dec_aln_aln_ib_ifu_i0_pc,
  output        io_ifu_dec_dec_aln_aln_ib_ifu_i0_pc4,
  output        io_ifu_dec_dec_aln_aln_ib_i0_brp_valid,
  output [11:0] io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_toffset,
  output [1:0]  io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_hist,
  output        io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_br_error,
  output        io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_br_start_error,
  output        io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_bank,
  output [30:0] io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_prett,
  output        io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_way,
  output        io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_ret,
  output        io_ifu_dec_dec_aln_ifu_pmu_instr_aligned,
  input         io_ifu_dec_dec_mem_ctrl_dec_tlu_flush_err_wb,
  input         io_ifu_dec_dec_mem_ctrl_dec_tlu_i0_commit_cmt,
  input         io_ifu_dec_dec_mem_ctrl_dec_tlu_force_halt,
  input         io_ifu_dec_dec_mem_ctrl_dec_tlu_fence_i_wb,
  input  [70:0] io_ifu_dec_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_wrdata,
  input  [16:0] io_ifu_dec_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_dicawics,
  input         io_ifu_dec_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_rd_valid,
  input         io_ifu_dec_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_wr_valid,
  input         io_ifu_dec_dec_mem_ctrl_dec_tlu_core_ecc_disable,
  output        io_ifu_dec_dec_mem_ctrl_ifu_pmu_ic_miss,
  output        io_ifu_dec_dec_mem_ctrl_ifu_pmu_ic_hit,
  output        io_ifu_dec_dec_mem_ctrl_ifu_pmu_bus_error,
  output        io_ifu_dec_dec_mem_ctrl_ifu_pmu_bus_busy,
  output        io_ifu_dec_dec_mem_ctrl_ifu_pmu_bus_trxn,
  output        io_ifu_dec_dec_mem_ctrl_ifu_ic_error_start,
  output        io_ifu_dec_dec_mem_ctrl_ifu_iccm_rd_ecc_single_err,
  output [70:0] io_ifu_dec_dec_mem_ctrl_ifu_ic_debug_rd_data,
  output        io_ifu_dec_dec_mem_ctrl_ifu_ic_debug_rd_data_valid,
  output        io_ifu_dec_dec_mem_ctrl_ifu_miss_state_idle,
  input         io_ifu_dec_dec_ifc_dec_tlu_flush_noredir_wb,
  input  [31:0] io_ifu_dec_dec_ifc_dec_tlu_mrac_ff,
  output        io_ifu_dec_dec_ifc_ifu_pmu_fetch_stall,
  input         io_ifu_dec_dec_bp_dec_tlu_br0_r_pkt_valid,
  input  [1:0]  io_ifu_dec_dec_bp_dec_tlu_br0_r_pkt_bits_hist,
  input         io_ifu_dec_dec_bp_dec_tlu_br0_r_pkt_bits_br_error,
  input         io_ifu_dec_dec_bp_dec_tlu_br0_r_pkt_bits_br_start_error,
  input         io_ifu_dec_dec_bp_dec_tlu_br0_r_pkt_bits_way,
  input         io_ifu_dec_dec_bp_dec_tlu_br0_r_pkt_bits_middle,
  input         io_ifu_dec_dec_bp_dec_tlu_flush_leak_one_wb,
  input         io_ifu_dec_dec_bp_dec_tlu_bpred_disable,
  input  [7:0]  io_exu_ifu_exu_bp_exu_i0_br_index_r,
  input  [7:0]  io_exu_ifu_exu_bp_exu_i0_br_fghr_r,
  input         io_exu_ifu_exu_bp_exu_i0_br_way_r,
  input         io_exu_ifu_exu_bp_exu_mp_pkt_valid,
  input         io_exu_ifu_exu_bp_exu_mp_pkt_bits_misp,
  input         io_exu_ifu_exu_bp_exu_mp_pkt_bits_ataken,
  input         io_exu_ifu_exu_bp_exu_mp_pkt_bits_boffset,
  input         io_exu_ifu_exu_bp_exu_mp_pkt_bits_pc4,
  input  [1:0]  io_exu_ifu_exu_bp_exu_mp_pkt_bits_hist,
  input  [11:0] io_exu_ifu_exu_bp_exu_mp_pkt_bits_toffset,
  input         io_exu_ifu_exu_bp_exu_mp_pkt_bits_br_error,
  input         io_exu_ifu_exu_bp_exu_mp_pkt_bits_br_start_error,
  input  [30:0] io_exu_ifu_exu_bp_exu_mp_pkt_bits_prett,
  input         io_exu_ifu_exu_bp_exu_mp_pkt_bits_pcall,
  input         io_exu_ifu_exu_bp_exu_mp_pkt_bits_pret,
  input         io_exu_ifu_exu_bp_exu_mp_pkt_bits_pja,
  input         io_exu_ifu_exu_bp_exu_mp_pkt_bits_way,
  input  [7:0]  io_exu_ifu_exu_bp_exu_mp_eghr,
  input  [7:0]  io_exu_ifu_exu_bp_exu_mp_fghr,
  input  [7:0]  io_exu_ifu_exu_bp_exu_mp_index,
  input  [4:0]  io_exu_ifu_exu_bp_exu_mp_btag,
  output [14:0] io_iccm_rw_addr,
  output        io_iccm_buf_correct_ecc,
  output        io_iccm_correction_state,
  output        io_iccm_wren,
  output        io_iccm_rden,
  output [2:0]  io_iccm_wr_size,
  output [77:0] io_iccm_wr_data,
  input  [63:0] io_iccm_rd_data,
  input  [77:0] io_iccm_rd_data_ecc,
  output [30:0] io_ic_rw_addr,
  output [1:0]  io_ic_tag_valid,
  output [1:0]  io_ic_wr_en,
  output        io_ic_rd_en,
  output [70:0] io_ic_wr_data_0,
  output [70:0] io_ic_wr_data_1,
  output [70:0] io_ic_debug_wr_data,
  output [9:0]  io_ic_debug_addr,
  input  [63:0] io_ic_rd_data,
  input  [70:0] io_ic_debug_rd_data,
  input  [25:0] io_ic_tag_debug_rd_data,
  input  [1:0]  io_ic_eccerr,
  input  [1:0]  io_ic_parerr,
  input  [1:0]  io_ic_rd_hit,
  input         io_ic_tag_perr,
  output        io_ic_debug_rd_en,
  output        io_ic_debug_wr_en,
  output        io_ic_debug_tag_array,
  output [1:0]  io_ic_debug_way,
  output [63:0] io_ic_premux_data,
  output        io_ic_sel_premux_data,
  input         io_ifu_aw_ready,
  output        io_ifu_aw_valid,
  output [2:0]  io_ifu_aw_bits_id,
  output [31:0] io_ifu_aw_bits_addr,
  output [3:0]  io_ifu_aw_bits_region,
  output [7:0]  io_ifu_aw_bits_len,
  output [2:0]  io_ifu_aw_bits_size,
  output [1:0]  io_ifu_aw_bits_burst,
  output        io_ifu_aw_bits_lock,
  output [3:0]  io_ifu_aw_bits_cache,
  output [2:0]  io_ifu_aw_bits_prot,
  output [3:0]  io_ifu_aw_bits_qos,
  input         io_ifu_w_ready,
  output        io_ifu_w_valid,
  output [63:0] io_ifu_w_bits_data,
  output [7:0]  io_ifu_w_bits_strb,
  output        io_ifu_w_bits_last,
  output        io_ifu_b_ready,
  input         io_ifu_b_valid,
  input  [1:0]  io_ifu_b_bits_resp,
  input  [2:0]  io_ifu_b_bits_id,
  input         io_ifu_ar_ready,
  output        io_ifu_ar_valid,
  output [2:0]  io_ifu_ar_bits_id,
  output [31:0] io_ifu_ar_bits_addr,
  output [3:0]  io_ifu_ar_bits_region,
  output [7:0]  io_ifu_ar_bits_len,
  output [2:0]  io_ifu_ar_bits_size,
  output [1:0]  io_ifu_ar_bits_burst,
  output        io_ifu_ar_bits_lock,
  output [3:0]  io_ifu_ar_bits_cache,
  output [2:0]  io_ifu_ar_bits_prot,
  output [3:0]  io_ifu_ar_bits_qos,
  output        io_ifu_r_ready,
  input         io_ifu_r_valid,
  input  [2:0]  io_ifu_r_bits_id,
  input  [63:0] io_ifu_r_bits_data,
  input  [1:0]  io_ifu_r_bits_resp,
  input         io_ifu_r_bits_last,
  input         io_ifu_bus_clk_en,
  input         io_ifu_dma_dma_ifc_dma_iccm_stall_any,
  input         io_ifu_dma_dma_mem_ctl_dma_iccm_req,
  input  [31:0] io_ifu_dma_dma_mem_ctl_dma_mem_addr,
  input  [2:0]  io_ifu_dma_dma_mem_ctl_dma_mem_sz,
  input         io_ifu_dma_dma_mem_ctl_dma_mem_write,
  input  [63:0] io_ifu_dma_dma_mem_ctl_dma_mem_wdata,
  input  [2:0]  io_ifu_dma_dma_mem_ctl_dma_mem_tag,
  output        io_iccm_dma_ecc_error,
  output        io_iccm_dma_rvalid,
  output [63:0] io_iccm_dma_rdata,
  output [2:0]  io_iccm_dma_rtag,
  output        io_iccm_ready,
  output        io_iccm_dma_sb_error,
  input         io_dec_tlu_flush_lower_wb,
  input         io_scan_mode
);
  wire  mem_ctl_clock; // @[ifu.scala 34:23]
  wire  mem_ctl_reset; // @[ifu.scala 34:23]
  wire  mem_ctl_io_free_clk; // @[ifu.scala 34:23]
  wire  mem_ctl_io_active_clk; // @[ifu.scala 34:23]
  wire  mem_ctl_io_exu_flush_final; // @[ifu.scala 34:23]
  wire  mem_ctl_io_dec_mem_ctrl_dec_tlu_flush_err_wb; // @[ifu.scala 34:23]
  wire  mem_ctl_io_dec_mem_ctrl_dec_tlu_i0_commit_cmt; // @[ifu.scala 34:23]
  wire  mem_ctl_io_dec_mem_ctrl_dec_tlu_force_halt; // @[ifu.scala 34:23]
  wire  mem_ctl_io_dec_mem_ctrl_dec_tlu_fence_i_wb; // @[ifu.scala 34:23]
  wire [70:0] mem_ctl_io_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_wrdata; // @[ifu.scala 34:23]
  wire [16:0] mem_ctl_io_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_dicawics; // @[ifu.scala 34:23]
  wire  mem_ctl_io_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_rd_valid; // @[ifu.scala 34:23]
  wire  mem_ctl_io_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_wr_valid; // @[ifu.scala 34:23]
  wire  mem_ctl_io_dec_mem_ctrl_dec_tlu_core_ecc_disable; // @[ifu.scala 34:23]
  wire  mem_ctl_io_dec_mem_ctrl_ifu_pmu_ic_miss; // @[ifu.scala 34:23]
  wire  mem_ctl_io_dec_mem_ctrl_ifu_pmu_ic_hit; // @[ifu.scala 34:23]
  wire  mem_ctl_io_dec_mem_ctrl_ifu_pmu_bus_error; // @[ifu.scala 34:23]
  wire  mem_ctl_io_dec_mem_ctrl_ifu_pmu_bus_busy; // @[ifu.scala 34:23]
  wire  mem_ctl_io_dec_mem_ctrl_ifu_pmu_bus_trxn; // @[ifu.scala 34:23]
  wire  mem_ctl_io_dec_mem_ctrl_ifu_ic_error_start; // @[ifu.scala 34:23]
  wire  mem_ctl_io_dec_mem_ctrl_ifu_iccm_rd_ecc_single_err; // @[ifu.scala 34:23]
  wire [70:0] mem_ctl_io_dec_mem_ctrl_ifu_ic_debug_rd_data; // @[ifu.scala 34:23]
  wire  mem_ctl_io_dec_mem_ctrl_ifu_ic_debug_rd_data_valid; // @[ifu.scala 34:23]
  wire  mem_ctl_io_dec_mem_ctrl_ifu_miss_state_idle; // @[ifu.scala 34:23]
  wire [30:0] mem_ctl_io_ifc_fetch_addr_bf; // @[ifu.scala 34:23]
  wire  mem_ctl_io_ifc_fetch_uncacheable_bf; // @[ifu.scala 34:23]
  wire  mem_ctl_io_ifc_fetch_req_bf; // @[ifu.scala 34:23]
  wire  mem_ctl_io_ifc_fetch_req_bf_raw; // @[ifu.scala 34:23]
  wire  mem_ctl_io_ifc_iccm_access_bf; // @[ifu.scala 34:23]
  wire  mem_ctl_io_ifc_region_acc_fault_bf; // @[ifu.scala 34:23]
  wire  mem_ctl_io_ifc_dma_access_ok; // @[ifu.scala 34:23]
  wire  mem_ctl_io_ifu_bp_hit_taken_f; // @[ifu.scala 34:23]
  wire  mem_ctl_io_ifu_bp_inst_mask_f; // @[ifu.scala 34:23]
  wire  mem_ctl_io_ifu_axi_ar_ready; // @[ifu.scala 34:23]
  wire  mem_ctl_io_ifu_axi_ar_valid; // @[ifu.scala 34:23]
  wire [2:0] mem_ctl_io_ifu_axi_ar_bits_id; // @[ifu.scala 34:23]
  wire [31:0] mem_ctl_io_ifu_axi_ar_bits_addr; // @[ifu.scala 34:23]
  wire [3:0] mem_ctl_io_ifu_axi_ar_bits_region; // @[ifu.scala 34:23]
  wire  mem_ctl_io_ifu_axi_r_ready; // @[ifu.scala 34:23]
  wire  mem_ctl_io_ifu_axi_r_valid; // @[ifu.scala 34:23]
  wire [2:0] mem_ctl_io_ifu_axi_r_bits_id; // @[ifu.scala 34:23]
  wire [63:0] mem_ctl_io_ifu_axi_r_bits_data; // @[ifu.scala 34:23]
  wire [1:0] mem_ctl_io_ifu_axi_r_bits_resp; // @[ifu.scala 34:23]
  wire  mem_ctl_io_ifu_bus_clk_en; // @[ifu.scala 34:23]
  wire  mem_ctl_io_dma_mem_ctl_dma_iccm_req; // @[ifu.scala 34:23]
  wire [31:0] mem_ctl_io_dma_mem_ctl_dma_mem_addr; // @[ifu.scala 34:23]
  wire [2:0] mem_ctl_io_dma_mem_ctl_dma_mem_sz; // @[ifu.scala 34:23]
  wire  mem_ctl_io_dma_mem_ctl_dma_mem_write; // @[ifu.scala 34:23]
  wire [63:0] mem_ctl_io_dma_mem_ctl_dma_mem_wdata; // @[ifu.scala 34:23]
  wire [2:0] mem_ctl_io_dma_mem_ctl_dma_mem_tag; // @[ifu.scala 34:23]
  wire [14:0] mem_ctl_io_iccm_rw_addr; // @[ifu.scala 34:23]
  wire  mem_ctl_io_iccm_buf_correct_ecc; // @[ifu.scala 34:23]
  wire  mem_ctl_io_iccm_correction_state; // @[ifu.scala 34:23]
  wire  mem_ctl_io_iccm_wren; // @[ifu.scala 34:23]
  wire  mem_ctl_io_iccm_rden; // @[ifu.scala 34:23]
  wire [2:0] mem_ctl_io_iccm_wr_size; // @[ifu.scala 34:23]
  wire [77:0] mem_ctl_io_iccm_wr_data; // @[ifu.scala 34:23]
  wire [63:0] mem_ctl_io_iccm_rd_data; // @[ifu.scala 34:23]
  wire [77:0] mem_ctl_io_iccm_rd_data_ecc; // @[ifu.scala 34:23]
  wire [30:0] mem_ctl_io_ic_rw_addr; // @[ifu.scala 34:23]
  wire [1:0] mem_ctl_io_ic_tag_valid; // @[ifu.scala 34:23]
  wire [1:0] mem_ctl_io_ic_wr_en; // @[ifu.scala 34:23]
  wire  mem_ctl_io_ic_rd_en; // @[ifu.scala 34:23]
  wire [70:0] mem_ctl_io_ic_wr_data_0; // @[ifu.scala 34:23]
  wire [70:0] mem_ctl_io_ic_wr_data_1; // @[ifu.scala 34:23]
  wire [70:0] mem_ctl_io_ic_debug_wr_data; // @[ifu.scala 34:23]
  wire [9:0] mem_ctl_io_ic_debug_addr; // @[ifu.scala 34:23]
  wire [63:0] mem_ctl_io_ic_rd_data; // @[ifu.scala 34:23]
  wire [70:0] mem_ctl_io_ic_debug_rd_data; // @[ifu.scala 34:23]
  wire [25:0] mem_ctl_io_ic_tag_debug_rd_data; // @[ifu.scala 34:23]
  wire [1:0] mem_ctl_io_ic_eccerr; // @[ifu.scala 34:23]
  wire [1:0] mem_ctl_io_ic_rd_hit; // @[ifu.scala 34:23]
  wire  mem_ctl_io_ic_tag_perr; // @[ifu.scala 34:23]
  wire  mem_ctl_io_ic_debug_rd_en; // @[ifu.scala 34:23]
  wire  mem_ctl_io_ic_debug_wr_en; // @[ifu.scala 34:23]
  wire  mem_ctl_io_ic_debug_tag_array; // @[ifu.scala 34:23]
  wire [1:0] mem_ctl_io_ic_debug_way; // @[ifu.scala 34:23]
  wire [63:0] mem_ctl_io_ic_premux_data; // @[ifu.scala 34:23]
  wire  mem_ctl_io_ic_sel_premux_data; // @[ifu.scala 34:23]
  wire [1:0] mem_ctl_io_ifu_fetch_val; // @[ifu.scala 34:23]
  wire  mem_ctl_io_ifu_ic_mb_empty; // @[ifu.scala 34:23]
  wire  mem_ctl_io_ic_dma_active; // @[ifu.scala 34:23]
  wire  mem_ctl_io_ic_write_stall; // @[ifu.scala 34:23]
  wire  mem_ctl_io_iccm_dma_ecc_error; // @[ifu.scala 34:23]
  wire  mem_ctl_io_iccm_dma_rvalid; // @[ifu.scala 34:23]
  wire [63:0] mem_ctl_io_iccm_dma_rdata; // @[ifu.scala 34:23]
  wire [2:0] mem_ctl_io_iccm_dma_rtag; // @[ifu.scala 34:23]
  wire  mem_ctl_io_iccm_ready; // @[ifu.scala 34:23]
  wire  mem_ctl_io_dec_tlu_flush_lower_wb; // @[ifu.scala 34:23]
  wire  mem_ctl_io_iccm_rd_ecc_double_err; // @[ifu.scala 34:23]
  wire  mem_ctl_io_iccm_dma_sb_error; // @[ifu.scala 34:23]
  wire  mem_ctl_io_ic_hit_f; // @[ifu.scala 34:23]
  wire  mem_ctl_io_ic_access_fault_f; // @[ifu.scala 34:23]
  wire [1:0] mem_ctl_io_ic_access_fault_type_f; // @[ifu.scala 34:23]
  wire  mem_ctl_io_ifu_async_error_start; // @[ifu.scala 34:23]
  wire [1:0] mem_ctl_io_ic_fetch_val_f; // @[ifu.scala 34:23]
  wire [31:0] mem_ctl_io_ic_data_f; // @[ifu.scala 34:23]
  wire  mem_ctl_io_scan_mode; // @[ifu.scala 34:23]
  wire  bp_ctl_clock; // @[ifu.scala 35:22]
  wire  bp_ctl_reset; // @[ifu.scala 35:22]
  wire  bp_ctl_io_active_clk; // @[ifu.scala 35:22]
  wire  bp_ctl_io_ic_hit_f; // @[ifu.scala 35:22]
  wire  bp_ctl_io_exu_flush_final; // @[ifu.scala 35:22]
  wire [30:0] bp_ctl_io_ifc_fetch_addr_f; // @[ifu.scala 35:22]
  wire  bp_ctl_io_ifc_fetch_req_f; // @[ifu.scala 35:22]
  wire  bp_ctl_io_dec_bp_dec_tlu_br0_r_pkt_valid; // @[ifu.scala 35:22]
  wire [1:0] bp_ctl_io_dec_bp_dec_tlu_br0_r_pkt_bits_hist; // @[ifu.scala 35:22]
  wire  bp_ctl_io_dec_bp_dec_tlu_br0_r_pkt_bits_br_error; // @[ifu.scala 35:22]
  wire  bp_ctl_io_dec_bp_dec_tlu_br0_r_pkt_bits_br_start_error; // @[ifu.scala 35:22]
  wire  bp_ctl_io_dec_bp_dec_tlu_br0_r_pkt_bits_way; // @[ifu.scala 35:22]
  wire  bp_ctl_io_dec_bp_dec_tlu_br0_r_pkt_bits_middle; // @[ifu.scala 35:22]
  wire  bp_ctl_io_dec_bp_dec_tlu_flush_leak_one_wb; // @[ifu.scala 35:22]
  wire  bp_ctl_io_dec_bp_dec_tlu_bpred_disable; // @[ifu.scala 35:22]
  wire  bp_ctl_io_dec_tlu_flush_lower_wb; // @[ifu.scala 35:22]
  wire [7:0] bp_ctl_io_exu_bp_exu_i0_br_index_r; // @[ifu.scala 35:22]
  wire [7:0] bp_ctl_io_exu_bp_exu_i0_br_fghr_r; // @[ifu.scala 35:22]
  wire  bp_ctl_io_exu_bp_exu_mp_pkt_bits_misp; // @[ifu.scala 35:22]
  wire  bp_ctl_io_exu_bp_exu_mp_pkt_bits_ataken; // @[ifu.scala 35:22]
  wire  bp_ctl_io_exu_bp_exu_mp_pkt_bits_boffset; // @[ifu.scala 35:22]
  wire  bp_ctl_io_exu_bp_exu_mp_pkt_bits_pc4; // @[ifu.scala 35:22]
  wire [1:0] bp_ctl_io_exu_bp_exu_mp_pkt_bits_hist; // @[ifu.scala 35:22]
  wire [11:0] bp_ctl_io_exu_bp_exu_mp_pkt_bits_toffset; // @[ifu.scala 35:22]
  wire  bp_ctl_io_exu_bp_exu_mp_pkt_bits_pcall; // @[ifu.scala 35:22]
  wire  bp_ctl_io_exu_bp_exu_mp_pkt_bits_pret; // @[ifu.scala 35:22]
  wire  bp_ctl_io_exu_bp_exu_mp_pkt_bits_pja; // @[ifu.scala 35:22]
  wire  bp_ctl_io_exu_bp_exu_mp_pkt_bits_way; // @[ifu.scala 35:22]
  wire [7:0] bp_ctl_io_exu_bp_exu_mp_eghr; // @[ifu.scala 35:22]
  wire [7:0] bp_ctl_io_exu_bp_exu_mp_fghr; // @[ifu.scala 35:22]
  wire [7:0] bp_ctl_io_exu_bp_exu_mp_index; // @[ifu.scala 35:22]
  wire [4:0] bp_ctl_io_exu_bp_exu_mp_btag; // @[ifu.scala 35:22]
  wire  bp_ctl_io_ifu_bp_hit_taken_f; // @[ifu.scala 35:22]
  wire [30:0] bp_ctl_io_ifu_bp_btb_target_f; // @[ifu.scala 35:22]
  wire  bp_ctl_io_ifu_bp_inst_mask_f; // @[ifu.scala 35:22]
  wire [7:0] bp_ctl_io_ifu_bp_fghr_f; // @[ifu.scala 35:22]
  wire [1:0] bp_ctl_io_ifu_bp_way_f; // @[ifu.scala 35:22]
  wire [1:0] bp_ctl_io_ifu_bp_ret_f; // @[ifu.scala 35:22]
  wire [1:0] bp_ctl_io_ifu_bp_hist1_f; // @[ifu.scala 35:22]
  wire [1:0] bp_ctl_io_ifu_bp_hist0_f; // @[ifu.scala 35:22]
  wire [1:0] bp_ctl_io_ifu_bp_pc4_f; // @[ifu.scala 35:22]
  wire [1:0] bp_ctl_io_ifu_bp_valid_f; // @[ifu.scala 35:22]
  wire [11:0] bp_ctl_io_ifu_bp_poffset_f; // @[ifu.scala 35:22]
  wire  bp_ctl_io_scan_mode; // @[ifu.scala 35:22]
  wire  aln_ctl_clock; // @[ifu.scala 36:23]
  wire  aln_ctl_reset; // @[ifu.scala 36:23]
  wire  aln_ctl_io_scan_mode; // @[ifu.scala 36:23]
  wire  aln_ctl_io_active_clk; // @[ifu.scala 36:23]
  wire  aln_ctl_io_ifu_async_error_start; // @[ifu.scala 36:23]
  wire  aln_ctl_io_iccm_rd_ecc_double_err; // @[ifu.scala 36:23]
  wire  aln_ctl_io_ic_access_fault_f; // @[ifu.scala 36:23]
  wire [1:0] aln_ctl_io_ic_access_fault_type_f; // @[ifu.scala 36:23]
  wire [7:0] aln_ctl_io_ifu_bp_fghr_f; // @[ifu.scala 36:23]
  wire [30:0] aln_ctl_io_ifu_bp_btb_target_f; // @[ifu.scala 36:23]
  wire [11:0] aln_ctl_io_ifu_bp_poffset_f; // @[ifu.scala 36:23]
  wire [1:0] aln_ctl_io_ifu_bp_hist0_f; // @[ifu.scala 36:23]
  wire [1:0] aln_ctl_io_ifu_bp_hist1_f; // @[ifu.scala 36:23]
  wire [1:0] aln_ctl_io_ifu_bp_pc4_f; // @[ifu.scala 36:23]
  wire [1:0] aln_ctl_io_ifu_bp_way_f; // @[ifu.scala 36:23]
  wire [1:0] aln_ctl_io_ifu_bp_valid_f; // @[ifu.scala 36:23]
  wire [1:0] aln_ctl_io_ifu_bp_ret_f; // @[ifu.scala 36:23]
  wire  aln_ctl_io_exu_flush_final; // @[ifu.scala 36:23]
  wire  aln_ctl_io_dec_aln_aln_dec_dec_i0_decode_d; // @[ifu.scala 36:23]
  wire [15:0] aln_ctl_io_dec_aln_aln_dec_ifu_i0_cinst; // @[ifu.scala 36:23]
  wire  aln_ctl_io_dec_aln_aln_ib_ifu_i0_icaf; // @[ifu.scala 36:23]
  wire [1:0] aln_ctl_io_dec_aln_aln_ib_ifu_i0_icaf_type; // @[ifu.scala 36:23]
  wire  aln_ctl_io_dec_aln_aln_ib_ifu_i0_icaf_f1; // @[ifu.scala 36:23]
  wire  aln_ctl_io_dec_aln_aln_ib_ifu_i0_dbecc; // @[ifu.scala 36:23]
  wire [7:0] aln_ctl_io_dec_aln_aln_ib_ifu_i0_bp_index; // @[ifu.scala 36:23]
  wire [7:0] aln_ctl_io_dec_aln_aln_ib_ifu_i0_bp_fghr; // @[ifu.scala 36:23]
  wire [4:0] aln_ctl_io_dec_aln_aln_ib_ifu_i0_bp_btag; // @[ifu.scala 36:23]
  wire  aln_ctl_io_dec_aln_aln_ib_ifu_i0_valid; // @[ifu.scala 36:23]
  wire [31:0] aln_ctl_io_dec_aln_aln_ib_ifu_i0_instr; // @[ifu.scala 36:23]
  wire [30:0] aln_ctl_io_dec_aln_aln_ib_ifu_i0_pc; // @[ifu.scala 36:23]
  wire  aln_ctl_io_dec_aln_aln_ib_ifu_i0_pc4; // @[ifu.scala 36:23]
  wire  aln_ctl_io_dec_aln_aln_ib_i0_brp_valid; // @[ifu.scala 36:23]
  wire [11:0] aln_ctl_io_dec_aln_aln_ib_i0_brp_bits_toffset; // @[ifu.scala 36:23]
  wire [1:0] aln_ctl_io_dec_aln_aln_ib_i0_brp_bits_hist; // @[ifu.scala 36:23]
  wire  aln_ctl_io_dec_aln_aln_ib_i0_brp_bits_br_error; // @[ifu.scala 36:23]
  wire  aln_ctl_io_dec_aln_aln_ib_i0_brp_bits_br_start_error; // @[ifu.scala 36:23]
  wire  aln_ctl_io_dec_aln_aln_ib_i0_brp_bits_bank; // @[ifu.scala 36:23]
  wire [30:0] aln_ctl_io_dec_aln_aln_ib_i0_brp_bits_prett; // @[ifu.scala 36:23]
  wire  aln_ctl_io_dec_aln_aln_ib_i0_brp_bits_way; // @[ifu.scala 36:23]
  wire  aln_ctl_io_dec_aln_aln_ib_i0_brp_bits_ret; // @[ifu.scala 36:23]
  wire  aln_ctl_io_dec_aln_ifu_pmu_instr_aligned; // @[ifu.scala 36:23]
  wire [31:0] aln_ctl_io_ifu_fetch_data_f; // @[ifu.scala 36:23]
  wire [1:0] aln_ctl_io_ifu_fetch_val; // @[ifu.scala 36:23]
  wire [30:0] aln_ctl_io_ifu_fetch_pc; // @[ifu.scala 36:23]
  wire  aln_ctl_io_ifu_fb_consume1; // @[ifu.scala 36:23]
  wire  aln_ctl_io_ifu_fb_consume2; // @[ifu.scala 36:23]
  wire  ifc_ctl_clock; // @[ifu.scala 37:23]
  wire  ifc_ctl_reset; // @[ifu.scala 37:23]
  wire  ifc_ctl_io_exu_flush_final; // @[ifu.scala 37:23]
  wire [30:0] ifc_ctl_io_exu_flush_path_final; // @[ifu.scala 37:23]
  wire  ifc_ctl_io_free_clk; // @[ifu.scala 37:23]
  wire  ifc_ctl_io_active_clk; // @[ifu.scala 37:23]
  wire  ifc_ctl_io_scan_mode; // @[ifu.scala 37:23]
  wire  ifc_ctl_io_ic_hit_f; // @[ifu.scala 37:23]
  wire  ifc_ctl_io_ifu_ic_mb_empty; // @[ifu.scala 37:23]
  wire  ifc_ctl_io_ifu_fb_consume1; // @[ifu.scala 37:23]
  wire  ifc_ctl_io_ifu_fb_consume2; // @[ifu.scala 37:23]
  wire  ifc_ctl_io_ifu_bp_hit_taken_f; // @[ifu.scala 37:23]
  wire [30:0] ifc_ctl_io_ifu_bp_btb_target_f; // @[ifu.scala 37:23]
  wire  ifc_ctl_io_ic_dma_active; // @[ifu.scala 37:23]
  wire  ifc_ctl_io_ic_write_stall; // @[ifu.scala 37:23]
  wire  ifc_ctl_io_dec_ifc_dec_tlu_flush_noredir_wb; // @[ifu.scala 37:23]
  wire [31:0] ifc_ctl_io_dec_ifc_dec_tlu_mrac_ff; // @[ifu.scala 37:23]
  wire  ifc_ctl_io_dec_ifc_ifu_pmu_fetch_stall; // @[ifu.scala 37:23]
  wire  ifc_ctl_io_dma_ifc_dma_iccm_stall_any; // @[ifu.scala 37:23]
  wire [30:0] ifc_ctl_io_ifc_fetch_addr_f; // @[ifu.scala 37:23]
  wire [30:0] ifc_ctl_io_ifc_fetch_addr_bf; // @[ifu.scala 37:23]
  wire  ifc_ctl_io_ifc_fetch_req_f; // @[ifu.scala 37:23]
  wire  ifc_ctl_io_ifc_fetch_uncacheable_bf; // @[ifu.scala 37:23]
  wire  ifc_ctl_io_ifc_fetch_req_bf; // @[ifu.scala 37:23]
  wire  ifc_ctl_io_ifc_fetch_req_bf_raw; // @[ifu.scala 37:23]
  wire  ifc_ctl_io_ifc_iccm_access_bf; // @[ifu.scala 37:23]
  wire  ifc_ctl_io_ifc_region_acc_fault_bf; // @[ifu.scala 37:23]
  wire  ifc_ctl_io_ifc_dma_access_ok; // @[ifu.scala 37:23]
  ifu_mem_ctl mem_ctl ( // @[ifu.scala 34:23]
    .clock(mem_ctl_clock),
    .reset(mem_ctl_reset),
    .io_free_clk(mem_ctl_io_free_clk),
    .io_active_clk(mem_ctl_io_active_clk),
    .io_exu_flush_final(mem_ctl_io_exu_flush_final),
    .io_dec_mem_ctrl_dec_tlu_flush_err_wb(mem_ctl_io_dec_mem_ctrl_dec_tlu_flush_err_wb),
    .io_dec_mem_ctrl_dec_tlu_i0_commit_cmt(mem_ctl_io_dec_mem_ctrl_dec_tlu_i0_commit_cmt),
    .io_dec_mem_ctrl_dec_tlu_force_halt(mem_ctl_io_dec_mem_ctrl_dec_tlu_force_halt),
    .io_dec_mem_ctrl_dec_tlu_fence_i_wb(mem_ctl_io_dec_mem_ctrl_dec_tlu_fence_i_wb),
    .io_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_wrdata(mem_ctl_io_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_wrdata),
    .io_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_dicawics(mem_ctl_io_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_dicawics),
    .io_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_rd_valid(mem_ctl_io_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_rd_valid),
    .io_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_wr_valid(mem_ctl_io_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_wr_valid),
    .io_dec_mem_ctrl_dec_tlu_core_ecc_disable(mem_ctl_io_dec_mem_ctrl_dec_tlu_core_ecc_disable),
    .io_dec_mem_ctrl_ifu_pmu_ic_miss(mem_ctl_io_dec_mem_ctrl_ifu_pmu_ic_miss),
    .io_dec_mem_ctrl_ifu_pmu_ic_hit(mem_ctl_io_dec_mem_ctrl_ifu_pmu_ic_hit),
    .io_dec_mem_ctrl_ifu_pmu_bus_error(mem_ctl_io_dec_mem_ctrl_ifu_pmu_bus_error),
    .io_dec_mem_ctrl_ifu_pmu_bus_busy(mem_ctl_io_dec_mem_ctrl_ifu_pmu_bus_busy),
    .io_dec_mem_ctrl_ifu_pmu_bus_trxn(mem_ctl_io_dec_mem_ctrl_ifu_pmu_bus_trxn),
    .io_dec_mem_ctrl_ifu_ic_error_start(mem_ctl_io_dec_mem_ctrl_ifu_ic_error_start),
    .io_dec_mem_ctrl_ifu_iccm_rd_ecc_single_err(mem_ctl_io_dec_mem_ctrl_ifu_iccm_rd_ecc_single_err),
    .io_dec_mem_ctrl_ifu_ic_debug_rd_data(mem_ctl_io_dec_mem_ctrl_ifu_ic_debug_rd_data),
    .io_dec_mem_ctrl_ifu_ic_debug_rd_data_valid(mem_ctl_io_dec_mem_ctrl_ifu_ic_debug_rd_data_valid),
    .io_dec_mem_ctrl_ifu_miss_state_idle(mem_ctl_io_dec_mem_ctrl_ifu_miss_state_idle),
    .io_ifc_fetch_addr_bf(mem_ctl_io_ifc_fetch_addr_bf),
    .io_ifc_fetch_uncacheable_bf(mem_ctl_io_ifc_fetch_uncacheable_bf),
    .io_ifc_fetch_req_bf(mem_ctl_io_ifc_fetch_req_bf),
    .io_ifc_fetch_req_bf_raw(mem_ctl_io_ifc_fetch_req_bf_raw),
    .io_ifc_iccm_access_bf(mem_ctl_io_ifc_iccm_access_bf),
    .io_ifc_region_acc_fault_bf(mem_ctl_io_ifc_region_acc_fault_bf),
    .io_ifc_dma_access_ok(mem_ctl_io_ifc_dma_access_ok),
    .io_ifu_bp_hit_taken_f(mem_ctl_io_ifu_bp_hit_taken_f),
    .io_ifu_bp_inst_mask_f(mem_ctl_io_ifu_bp_inst_mask_f),
    .io_ifu_axi_ar_ready(mem_ctl_io_ifu_axi_ar_ready),
    .io_ifu_axi_ar_valid(mem_ctl_io_ifu_axi_ar_valid),
    .io_ifu_axi_ar_bits_id(mem_ctl_io_ifu_axi_ar_bits_id),
    .io_ifu_axi_ar_bits_addr(mem_ctl_io_ifu_axi_ar_bits_addr),
    .io_ifu_axi_ar_bits_region(mem_ctl_io_ifu_axi_ar_bits_region),
    .io_ifu_axi_r_ready(mem_ctl_io_ifu_axi_r_ready),
    .io_ifu_axi_r_valid(mem_ctl_io_ifu_axi_r_valid),
    .io_ifu_axi_r_bits_id(mem_ctl_io_ifu_axi_r_bits_id),
    .io_ifu_axi_r_bits_data(mem_ctl_io_ifu_axi_r_bits_data),
    .io_ifu_axi_r_bits_resp(mem_ctl_io_ifu_axi_r_bits_resp),
    .io_ifu_bus_clk_en(mem_ctl_io_ifu_bus_clk_en),
    .io_dma_mem_ctl_dma_iccm_req(mem_ctl_io_dma_mem_ctl_dma_iccm_req),
    .io_dma_mem_ctl_dma_mem_addr(mem_ctl_io_dma_mem_ctl_dma_mem_addr),
    .io_dma_mem_ctl_dma_mem_sz(mem_ctl_io_dma_mem_ctl_dma_mem_sz),
    .io_dma_mem_ctl_dma_mem_write(mem_ctl_io_dma_mem_ctl_dma_mem_write),
    .io_dma_mem_ctl_dma_mem_wdata(mem_ctl_io_dma_mem_ctl_dma_mem_wdata),
    .io_dma_mem_ctl_dma_mem_tag(mem_ctl_io_dma_mem_ctl_dma_mem_tag),
    .io_iccm_rw_addr(mem_ctl_io_iccm_rw_addr),
    .io_iccm_buf_correct_ecc(mem_ctl_io_iccm_buf_correct_ecc),
    .io_iccm_correction_state(mem_ctl_io_iccm_correction_state),
    .io_iccm_wren(mem_ctl_io_iccm_wren),
    .io_iccm_rden(mem_ctl_io_iccm_rden),
    .io_iccm_wr_size(mem_ctl_io_iccm_wr_size),
    .io_iccm_wr_data(mem_ctl_io_iccm_wr_data),
    .io_iccm_rd_data(mem_ctl_io_iccm_rd_data),
    .io_iccm_rd_data_ecc(mem_ctl_io_iccm_rd_data_ecc),
    .io_ic_rw_addr(mem_ctl_io_ic_rw_addr),
    .io_ic_tag_valid(mem_ctl_io_ic_tag_valid),
    .io_ic_wr_en(mem_ctl_io_ic_wr_en),
    .io_ic_rd_en(mem_ctl_io_ic_rd_en),
    .io_ic_wr_data_0(mem_ctl_io_ic_wr_data_0),
    .io_ic_wr_data_1(mem_ctl_io_ic_wr_data_1),
    .io_ic_debug_wr_data(mem_ctl_io_ic_debug_wr_data),
    .io_ic_debug_addr(mem_ctl_io_ic_debug_addr),
    .io_ic_rd_data(mem_ctl_io_ic_rd_data),
    .io_ic_debug_rd_data(mem_ctl_io_ic_debug_rd_data),
    .io_ic_tag_debug_rd_data(mem_ctl_io_ic_tag_debug_rd_data),
    .io_ic_eccerr(mem_ctl_io_ic_eccerr),
    .io_ic_rd_hit(mem_ctl_io_ic_rd_hit),
    .io_ic_tag_perr(mem_ctl_io_ic_tag_perr),
    .io_ic_debug_rd_en(mem_ctl_io_ic_debug_rd_en),
    .io_ic_debug_wr_en(mem_ctl_io_ic_debug_wr_en),
    .io_ic_debug_tag_array(mem_ctl_io_ic_debug_tag_array),
    .io_ic_debug_way(mem_ctl_io_ic_debug_way),
    .io_ic_premux_data(mem_ctl_io_ic_premux_data),
    .io_ic_sel_premux_data(mem_ctl_io_ic_sel_premux_data),
    .io_ifu_fetch_val(mem_ctl_io_ifu_fetch_val),
    .io_ifu_ic_mb_empty(mem_ctl_io_ifu_ic_mb_empty),
    .io_ic_dma_active(mem_ctl_io_ic_dma_active),
    .io_ic_write_stall(mem_ctl_io_ic_write_stall),
    .io_iccm_dma_ecc_error(mem_ctl_io_iccm_dma_ecc_error),
    .io_iccm_dma_rvalid(mem_ctl_io_iccm_dma_rvalid),
    .io_iccm_dma_rdata(mem_ctl_io_iccm_dma_rdata),
    .io_iccm_dma_rtag(mem_ctl_io_iccm_dma_rtag),
    .io_iccm_ready(mem_ctl_io_iccm_ready),
    .io_dec_tlu_flush_lower_wb(mem_ctl_io_dec_tlu_flush_lower_wb),
    .io_iccm_rd_ecc_double_err(mem_ctl_io_iccm_rd_ecc_double_err),
    .io_iccm_dma_sb_error(mem_ctl_io_iccm_dma_sb_error),
    .io_ic_hit_f(mem_ctl_io_ic_hit_f),
    .io_ic_access_fault_f(mem_ctl_io_ic_access_fault_f),
    .io_ic_access_fault_type_f(mem_ctl_io_ic_access_fault_type_f),
    .io_ifu_async_error_start(mem_ctl_io_ifu_async_error_start),
    .io_ic_fetch_val_f(mem_ctl_io_ic_fetch_val_f),
    .io_ic_data_f(mem_ctl_io_ic_data_f),
    .io_scan_mode(mem_ctl_io_scan_mode)
  );
  ifu_bp_ctl bp_ctl ( // @[ifu.scala 35:22]
    .clock(bp_ctl_clock),
    .reset(bp_ctl_reset),
    .io_active_clk(bp_ctl_io_active_clk),
    .io_ic_hit_f(bp_ctl_io_ic_hit_f),
    .io_exu_flush_final(bp_ctl_io_exu_flush_final),
    .io_ifc_fetch_addr_f(bp_ctl_io_ifc_fetch_addr_f),
    .io_ifc_fetch_req_f(bp_ctl_io_ifc_fetch_req_f),
    .io_dec_bp_dec_tlu_br0_r_pkt_valid(bp_ctl_io_dec_bp_dec_tlu_br0_r_pkt_valid),
    .io_dec_bp_dec_tlu_br0_r_pkt_bits_hist(bp_ctl_io_dec_bp_dec_tlu_br0_r_pkt_bits_hist),
    .io_dec_bp_dec_tlu_br0_r_pkt_bits_br_error(bp_ctl_io_dec_bp_dec_tlu_br0_r_pkt_bits_br_error),
    .io_dec_bp_dec_tlu_br0_r_pkt_bits_br_start_error(bp_ctl_io_dec_bp_dec_tlu_br0_r_pkt_bits_br_start_error),
    .io_dec_bp_dec_tlu_br0_r_pkt_bits_way(bp_ctl_io_dec_bp_dec_tlu_br0_r_pkt_bits_way),
    .io_dec_bp_dec_tlu_br0_r_pkt_bits_middle(bp_ctl_io_dec_bp_dec_tlu_br0_r_pkt_bits_middle),
    .io_dec_bp_dec_tlu_flush_leak_one_wb(bp_ctl_io_dec_bp_dec_tlu_flush_leak_one_wb),
    .io_dec_bp_dec_tlu_bpred_disable(bp_ctl_io_dec_bp_dec_tlu_bpred_disable),
    .io_dec_tlu_flush_lower_wb(bp_ctl_io_dec_tlu_flush_lower_wb),
    .io_exu_bp_exu_i0_br_index_r(bp_ctl_io_exu_bp_exu_i0_br_index_r),
    .io_exu_bp_exu_i0_br_fghr_r(bp_ctl_io_exu_bp_exu_i0_br_fghr_r),
    .io_exu_bp_exu_mp_pkt_bits_misp(bp_ctl_io_exu_bp_exu_mp_pkt_bits_misp),
    .io_exu_bp_exu_mp_pkt_bits_ataken(bp_ctl_io_exu_bp_exu_mp_pkt_bits_ataken),
    .io_exu_bp_exu_mp_pkt_bits_boffset(bp_ctl_io_exu_bp_exu_mp_pkt_bits_boffset),
    .io_exu_bp_exu_mp_pkt_bits_pc4(bp_ctl_io_exu_bp_exu_mp_pkt_bits_pc4),
    .io_exu_bp_exu_mp_pkt_bits_hist(bp_ctl_io_exu_bp_exu_mp_pkt_bits_hist),
    .io_exu_bp_exu_mp_pkt_bits_toffset(bp_ctl_io_exu_bp_exu_mp_pkt_bits_toffset),
    .io_exu_bp_exu_mp_pkt_bits_pcall(bp_ctl_io_exu_bp_exu_mp_pkt_bits_pcall),
    .io_exu_bp_exu_mp_pkt_bits_pret(bp_ctl_io_exu_bp_exu_mp_pkt_bits_pret),
    .io_exu_bp_exu_mp_pkt_bits_pja(bp_ctl_io_exu_bp_exu_mp_pkt_bits_pja),
    .io_exu_bp_exu_mp_pkt_bits_way(bp_ctl_io_exu_bp_exu_mp_pkt_bits_way),
    .io_exu_bp_exu_mp_eghr(bp_ctl_io_exu_bp_exu_mp_eghr),
    .io_exu_bp_exu_mp_fghr(bp_ctl_io_exu_bp_exu_mp_fghr),
    .io_exu_bp_exu_mp_index(bp_ctl_io_exu_bp_exu_mp_index),
    .io_exu_bp_exu_mp_btag(bp_ctl_io_exu_bp_exu_mp_btag),
    .io_ifu_bp_hit_taken_f(bp_ctl_io_ifu_bp_hit_taken_f),
    .io_ifu_bp_btb_target_f(bp_ctl_io_ifu_bp_btb_target_f),
    .io_ifu_bp_inst_mask_f(bp_ctl_io_ifu_bp_inst_mask_f),
    .io_ifu_bp_fghr_f(bp_ctl_io_ifu_bp_fghr_f),
    .io_ifu_bp_way_f(bp_ctl_io_ifu_bp_way_f),
    .io_ifu_bp_ret_f(bp_ctl_io_ifu_bp_ret_f),
    .io_ifu_bp_hist1_f(bp_ctl_io_ifu_bp_hist1_f),
    .io_ifu_bp_hist0_f(bp_ctl_io_ifu_bp_hist0_f),
    .io_ifu_bp_pc4_f(bp_ctl_io_ifu_bp_pc4_f),
    .io_ifu_bp_valid_f(bp_ctl_io_ifu_bp_valid_f),
    .io_ifu_bp_poffset_f(bp_ctl_io_ifu_bp_poffset_f),
    .io_scan_mode(bp_ctl_io_scan_mode)
  );
  ifu_aln_ctl aln_ctl ( // @[ifu.scala 36:23]
    .clock(aln_ctl_clock),
    .reset(aln_ctl_reset),
    .io_scan_mode(aln_ctl_io_scan_mode),
    .io_active_clk(aln_ctl_io_active_clk),
    .io_ifu_async_error_start(aln_ctl_io_ifu_async_error_start),
    .io_iccm_rd_ecc_double_err(aln_ctl_io_iccm_rd_ecc_double_err),
    .io_ic_access_fault_f(aln_ctl_io_ic_access_fault_f),
    .io_ic_access_fault_type_f(aln_ctl_io_ic_access_fault_type_f),
    .io_ifu_bp_fghr_f(aln_ctl_io_ifu_bp_fghr_f),
    .io_ifu_bp_btb_target_f(aln_ctl_io_ifu_bp_btb_target_f),
    .io_ifu_bp_poffset_f(aln_ctl_io_ifu_bp_poffset_f),
    .io_ifu_bp_hist0_f(aln_ctl_io_ifu_bp_hist0_f),
    .io_ifu_bp_hist1_f(aln_ctl_io_ifu_bp_hist1_f),
    .io_ifu_bp_pc4_f(aln_ctl_io_ifu_bp_pc4_f),
    .io_ifu_bp_way_f(aln_ctl_io_ifu_bp_way_f),
    .io_ifu_bp_valid_f(aln_ctl_io_ifu_bp_valid_f),
    .io_ifu_bp_ret_f(aln_ctl_io_ifu_bp_ret_f),
    .io_exu_flush_final(aln_ctl_io_exu_flush_final),
    .io_dec_aln_aln_dec_dec_i0_decode_d(aln_ctl_io_dec_aln_aln_dec_dec_i0_decode_d),
    .io_dec_aln_aln_dec_ifu_i0_cinst(aln_ctl_io_dec_aln_aln_dec_ifu_i0_cinst),
    .io_dec_aln_aln_ib_ifu_i0_icaf(aln_ctl_io_dec_aln_aln_ib_ifu_i0_icaf),
    .io_dec_aln_aln_ib_ifu_i0_icaf_type(aln_ctl_io_dec_aln_aln_ib_ifu_i0_icaf_type),
    .io_dec_aln_aln_ib_ifu_i0_icaf_f1(aln_ctl_io_dec_aln_aln_ib_ifu_i0_icaf_f1),
    .io_dec_aln_aln_ib_ifu_i0_dbecc(aln_ctl_io_dec_aln_aln_ib_ifu_i0_dbecc),
    .io_dec_aln_aln_ib_ifu_i0_bp_index(aln_ctl_io_dec_aln_aln_ib_ifu_i0_bp_index),
    .io_dec_aln_aln_ib_ifu_i0_bp_fghr(aln_ctl_io_dec_aln_aln_ib_ifu_i0_bp_fghr),
    .io_dec_aln_aln_ib_ifu_i0_bp_btag(aln_ctl_io_dec_aln_aln_ib_ifu_i0_bp_btag),
    .io_dec_aln_aln_ib_ifu_i0_valid(aln_ctl_io_dec_aln_aln_ib_ifu_i0_valid),
    .io_dec_aln_aln_ib_ifu_i0_instr(aln_ctl_io_dec_aln_aln_ib_ifu_i0_instr),
    .io_dec_aln_aln_ib_ifu_i0_pc(aln_ctl_io_dec_aln_aln_ib_ifu_i0_pc),
    .io_dec_aln_aln_ib_ifu_i0_pc4(aln_ctl_io_dec_aln_aln_ib_ifu_i0_pc4),
    .io_dec_aln_aln_ib_i0_brp_valid(aln_ctl_io_dec_aln_aln_ib_i0_brp_valid),
    .io_dec_aln_aln_ib_i0_brp_bits_toffset(aln_ctl_io_dec_aln_aln_ib_i0_brp_bits_toffset),
    .io_dec_aln_aln_ib_i0_brp_bits_hist(aln_ctl_io_dec_aln_aln_ib_i0_brp_bits_hist),
    .io_dec_aln_aln_ib_i0_brp_bits_br_error(aln_ctl_io_dec_aln_aln_ib_i0_brp_bits_br_error),
    .io_dec_aln_aln_ib_i0_brp_bits_br_start_error(aln_ctl_io_dec_aln_aln_ib_i0_brp_bits_br_start_error),
    .io_dec_aln_aln_ib_i0_brp_bits_bank(aln_ctl_io_dec_aln_aln_ib_i0_brp_bits_bank),
    .io_dec_aln_aln_ib_i0_brp_bits_prett(aln_ctl_io_dec_aln_aln_ib_i0_brp_bits_prett),
    .io_dec_aln_aln_ib_i0_brp_bits_way(aln_ctl_io_dec_aln_aln_ib_i0_brp_bits_way),
    .io_dec_aln_aln_ib_i0_brp_bits_ret(aln_ctl_io_dec_aln_aln_ib_i0_brp_bits_ret),
    .io_dec_aln_ifu_pmu_instr_aligned(aln_ctl_io_dec_aln_ifu_pmu_instr_aligned),
    .io_ifu_fetch_data_f(aln_ctl_io_ifu_fetch_data_f),
    .io_ifu_fetch_val(aln_ctl_io_ifu_fetch_val),
    .io_ifu_fetch_pc(aln_ctl_io_ifu_fetch_pc),
    .io_ifu_fb_consume1(aln_ctl_io_ifu_fb_consume1),
    .io_ifu_fb_consume2(aln_ctl_io_ifu_fb_consume2)
  );
  ifu_ifc_ctl ifc_ctl ( // @[ifu.scala 37:23]
    .clock(ifc_ctl_clock),
    .reset(ifc_ctl_reset),
    .io_exu_flush_final(ifc_ctl_io_exu_flush_final),
    .io_exu_flush_path_final(ifc_ctl_io_exu_flush_path_final),
    .io_free_clk(ifc_ctl_io_free_clk),
    .io_active_clk(ifc_ctl_io_active_clk),
    .io_scan_mode(ifc_ctl_io_scan_mode),
    .io_ic_hit_f(ifc_ctl_io_ic_hit_f),
    .io_ifu_ic_mb_empty(ifc_ctl_io_ifu_ic_mb_empty),
    .io_ifu_fb_consume1(ifc_ctl_io_ifu_fb_consume1),
    .io_ifu_fb_consume2(ifc_ctl_io_ifu_fb_consume2),
    .io_ifu_bp_hit_taken_f(ifc_ctl_io_ifu_bp_hit_taken_f),
    .io_ifu_bp_btb_target_f(ifc_ctl_io_ifu_bp_btb_target_f),
    .io_ic_dma_active(ifc_ctl_io_ic_dma_active),
    .io_ic_write_stall(ifc_ctl_io_ic_write_stall),
    .io_dec_ifc_dec_tlu_flush_noredir_wb(ifc_ctl_io_dec_ifc_dec_tlu_flush_noredir_wb),
    .io_dec_ifc_dec_tlu_mrac_ff(ifc_ctl_io_dec_ifc_dec_tlu_mrac_ff),
    .io_dec_ifc_ifu_pmu_fetch_stall(ifc_ctl_io_dec_ifc_ifu_pmu_fetch_stall),
    .io_dma_ifc_dma_iccm_stall_any(ifc_ctl_io_dma_ifc_dma_iccm_stall_any),
    .io_ifc_fetch_addr_f(ifc_ctl_io_ifc_fetch_addr_f),
    .io_ifc_fetch_addr_bf(ifc_ctl_io_ifc_fetch_addr_bf),
    .io_ifc_fetch_req_f(ifc_ctl_io_ifc_fetch_req_f),
    .io_ifc_fetch_uncacheable_bf(ifc_ctl_io_ifc_fetch_uncacheable_bf),
    .io_ifc_fetch_req_bf(ifc_ctl_io_ifc_fetch_req_bf),
    .io_ifc_fetch_req_bf_raw(ifc_ctl_io_ifc_fetch_req_bf_raw),
    .io_ifc_iccm_access_bf(ifc_ctl_io_ifc_iccm_access_bf),
    .io_ifc_region_acc_fault_bf(ifc_ctl_io_ifc_region_acc_fault_bf),
    .io_ifc_dma_access_ok(ifc_ctl_io_ifc_dma_access_ok)
  );
  assign io_ifu_dec_dec_aln_aln_dec_ifu_i0_cinst = aln_ctl_io_dec_aln_aln_dec_ifu_i0_cinst; // @[ifu.scala 73:22]
  assign io_ifu_dec_dec_aln_aln_ib_ifu_i0_icaf = aln_ctl_io_dec_aln_aln_ib_ifu_i0_icaf; // @[ifu.scala 73:22]
  assign io_ifu_dec_dec_aln_aln_ib_ifu_i0_icaf_type = aln_ctl_io_dec_aln_aln_ib_ifu_i0_icaf_type; // @[ifu.scala 73:22]
  assign io_ifu_dec_dec_aln_aln_ib_ifu_i0_icaf_f1 = aln_ctl_io_dec_aln_aln_ib_ifu_i0_icaf_f1; // @[ifu.scala 73:22]
  assign io_ifu_dec_dec_aln_aln_ib_ifu_i0_dbecc = aln_ctl_io_dec_aln_aln_ib_ifu_i0_dbecc; // @[ifu.scala 73:22]
  assign io_ifu_dec_dec_aln_aln_ib_ifu_i0_bp_index = aln_ctl_io_dec_aln_aln_ib_ifu_i0_bp_index; // @[ifu.scala 73:22]
  assign io_ifu_dec_dec_aln_aln_ib_ifu_i0_bp_fghr = aln_ctl_io_dec_aln_aln_ib_ifu_i0_bp_fghr; // @[ifu.scala 73:22]
  assign io_ifu_dec_dec_aln_aln_ib_ifu_i0_bp_btag = aln_ctl_io_dec_aln_aln_ib_ifu_i0_bp_btag; // @[ifu.scala 73:22]
  assign io_ifu_dec_dec_aln_aln_ib_ifu_i0_valid = aln_ctl_io_dec_aln_aln_ib_ifu_i0_valid; // @[ifu.scala 73:22]
  assign io_ifu_dec_dec_aln_aln_ib_ifu_i0_instr = aln_ctl_io_dec_aln_aln_ib_ifu_i0_instr; // @[ifu.scala 73:22]
  assign io_ifu_dec_dec_aln_aln_ib_ifu_i0_pc = aln_ctl_io_dec_aln_aln_ib_ifu_i0_pc; // @[ifu.scala 73:22]
  assign io_ifu_dec_dec_aln_aln_ib_ifu_i0_pc4 = aln_ctl_io_dec_aln_aln_ib_ifu_i0_pc4; // @[ifu.scala 73:22]
  assign io_ifu_dec_dec_aln_aln_ib_i0_brp_valid = aln_ctl_io_dec_aln_aln_ib_i0_brp_valid; // @[ifu.scala 73:22]
  assign io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_toffset = aln_ctl_io_dec_aln_aln_ib_i0_brp_bits_toffset; // @[ifu.scala 73:22]
  assign io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_hist = aln_ctl_io_dec_aln_aln_ib_i0_brp_bits_hist; // @[ifu.scala 73:22]
  assign io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_br_error = aln_ctl_io_dec_aln_aln_ib_i0_brp_bits_br_error; // @[ifu.scala 73:22]
  assign io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_br_start_error = aln_ctl_io_dec_aln_aln_ib_i0_brp_bits_br_start_error; // @[ifu.scala 73:22]
  assign io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_bank = aln_ctl_io_dec_aln_aln_ib_i0_brp_bits_bank; // @[ifu.scala 73:22]
  assign io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_prett = aln_ctl_io_dec_aln_aln_ib_i0_brp_bits_prett; // @[ifu.scala 73:22]
  assign io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_way = aln_ctl_io_dec_aln_aln_ib_i0_brp_bits_way; // @[ifu.scala 73:22]
  assign io_ifu_dec_dec_aln_aln_ib_i0_brp_bits_ret = aln_ctl_io_dec_aln_aln_ib_i0_brp_bits_ret; // @[ifu.scala 73:22]
  assign io_ifu_dec_dec_aln_ifu_pmu_instr_aligned = aln_ctl_io_dec_aln_ifu_pmu_instr_aligned; // @[ifu.scala 73:22]
  assign io_ifu_dec_dec_mem_ctrl_ifu_pmu_ic_miss = mem_ctl_io_dec_mem_ctrl_ifu_pmu_ic_miss; // @[ifu.scala 93:27]
  assign io_ifu_dec_dec_mem_ctrl_ifu_pmu_ic_hit = mem_ctl_io_dec_mem_ctrl_ifu_pmu_ic_hit; // @[ifu.scala 93:27]
  assign io_ifu_dec_dec_mem_ctrl_ifu_pmu_bus_error = mem_ctl_io_dec_mem_ctrl_ifu_pmu_bus_error; // @[ifu.scala 93:27]
  assign io_ifu_dec_dec_mem_ctrl_ifu_pmu_bus_busy = mem_ctl_io_dec_mem_ctrl_ifu_pmu_bus_busy; // @[ifu.scala 93:27]
  assign io_ifu_dec_dec_mem_ctrl_ifu_pmu_bus_trxn = mem_ctl_io_dec_mem_ctrl_ifu_pmu_bus_trxn; // @[ifu.scala 93:27]
  assign io_ifu_dec_dec_mem_ctrl_ifu_ic_error_start = mem_ctl_io_dec_mem_ctrl_ifu_ic_error_start; // @[ifu.scala 93:27]
  assign io_ifu_dec_dec_mem_ctrl_ifu_iccm_rd_ecc_single_err = mem_ctl_io_dec_mem_ctrl_ifu_iccm_rd_ecc_single_err; // @[ifu.scala 93:27]
  assign io_ifu_dec_dec_mem_ctrl_ifu_ic_debug_rd_data = mem_ctl_io_dec_mem_ctrl_ifu_ic_debug_rd_data; // @[ifu.scala 93:27]
  assign io_ifu_dec_dec_mem_ctrl_ifu_ic_debug_rd_data_valid = mem_ctl_io_dec_mem_ctrl_ifu_ic_debug_rd_data_valid; // @[ifu.scala 93:27]
  assign io_ifu_dec_dec_mem_ctrl_ifu_miss_state_idle = mem_ctl_io_dec_mem_ctrl_ifu_miss_state_idle; // @[ifu.scala 93:27]
  assign io_ifu_dec_dec_ifc_ifu_pmu_fetch_stall = ifc_ctl_io_dec_ifc_ifu_pmu_fetch_stall; // @[ifu.scala 46:22]
  assign io_iccm_rw_addr = mem_ctl_io_iccm_rw_addr; // @[ifu.scala 107:19]
  assign io_iccm_buf_correct_ecc = mem_ctl_io_iccm_buf_correct_ecc; // @[ifu.scala 107:19]
  assign io_iccm_correction_state = mem_ctl_io_iccm_correction_state; // @[ifu.scala 107:19]
  assign io_iccm_wren = mem_ctl_io_iccm_wren; // @[ifu.scala 107:19]
  assign io_iccm_rden = mem_ctl_io_iccm_rden; // @[ifu.scala 107:19]
  assign io_iccm_wr_size = mem_ctl_io_iccm_wr_size; // @[ifu.scala 107:19]
  assign io_iccm_wr_data = mem_ctl_io_iccm_wr_data; // @[ifu.scala 107:19]
  assign io_ic_rw_addr = mem_ctl_io_ic_rw_addr; // @[ifu.scala 106:17]
  assign io_ic_tag_valid = mem_ctl_io_ic_tag_valid; // @[ifu.scala 106:17]
  assign io_ic_wr_en = mem_ctl_io_ic_wr_en; // @[ifu.scala 106:17]
  assign io_ic_rd_en = mem_ctl_io_ic_rd_en; // @[ifu.scala 106:17]
  assign io_ic_wr_data_0 = mem_ctl_io_ic_wr_data_0; // @[ifu.scala 106:17]
  assign io_ic_wr_data_1 = mem_ctl_io_ic_wr_data_1; // @[ifu.scala 106:17]
  assign io_ic_debug_wr_data = mem_ctl_io_ic_debug_wr_data; // @[ifu.scala 106:17]
  assign io_ic_debug_addr = mem_ctl_io_ic_debug_addr; // @[ifu.scala 106:17]
  assign io_ic_debug_rd_en = mem_ctl_io_ic_debug_rd_en; // @[ifu.scala 106:17]
  assign io_ic_debug_wr_en = mem_ctl_io_ic_debug_wr_en; // @[ifu.scala 106:17]
  assign io_ic_debug_tag_array = mem_ctl_io_ic_debug_tag_array; // @[ifu.scala 106:17]
  assign io_ic_debug_way = mem_ctl_io_ic_debug_way; // @[ifu.scala 106:17]
  assign io_ic_premux_data = mem_ctl_io_ic_premux_data; // @[ifu.scala 106:17]
  assign io_ic_sel_premux_data = mem_ctl_io_ic_sel_premux_data; // @[ifu.scala 106:17]
  assign io_ifu_aw_valid = 1'h0; // @[ifu.scala 103:22]
  assign io_ifu_aw_bits_id = 3'h0; // @[ifu.scala 103:22]
  assign io_ifu_aw_bits_addr = 32'h0; // @[ifu.scala 103:22]
  assign io_ifu_aw_bits_region = 4'h0; // @[ifu.scala 103:22]
  assign io_ifu_aw_bits_len = 8'h0; // @[ifu.scala 103:22]
  assign io_ifu_aw_bits_size = 3'h0; // @[ifu.scala 103:22]
  assign io_ifu_aw_bits_burst = 2'h0; // @[ifu.scala 103:22]
  assign io_ifu_aw_bits_lock = 1'h0; // @[ifu.scala 103:22]
  assign io_ifu_aw_bits_cache = 4'h0; // @[ifu.scala 103:22]
  assign io_ifu_aw_bits_prot = 3'h0; // @[ifu.scala 103:22]
  assign io_ifu_aw_bits_qos = 4'h0; // @[ifu.scala 103:22]
  assign io_ifu_w_valid = 1'h0; // @[ifu.scala 103:22]
  assign io_ifu_w_bits_data = 64'h0; // @[ifu.scala 103:22]
  assign io_ifu_w_bits_strb = 8'h0; // @[ifu.scala 103:22]
  assign io_ifu_w_bits_last = 1'h0; // @[ifu.scala 103:22]
  assign io_ifu_b_ready = 1'h0; // @[ifu.scala 103:22]
  assign io_ifu_ar_valid = mem_ctl_io_ifu_axi_ar_valid; // @[ifu.scala 103:22]
  assign io_ifu_ar_bits_id = mem_ctl_io_ifu_axi_ar_bits_id; // @[ifu.scala 103:22]
  assign io_ifu_ar_bits_addr = mem_ctl_io_ifu_axi_ar_bits_addr; // @[ifu.scala 103:22]
  assign io_ifu_ar_bits_region = mem_ctl_io_ifu_axi_ar_bits_region; // @[ifu.scala 103:22]
  assign io_ifu_ar_bits_len = 8'h0; // @[ifu.scala 103:22]
  assign io_ifu_ar_bits_size = 3'h3; // @[ifu.scala 103:22]
  assign io_ifu_ar_bits_burst = 2'h1; // @[ifu.scala 103:22]
  assign io_ifu_ar_bits_lock = 1'h0; // @[ifu.scala 103:22]
  assign io_ifu_ar_bits_cache = 4'hf; // @[ifu.scala 103:22]
  assign io_ifu_ar_bits_prot = 3'h0; // @[ifu.scala 103:22]
  assign io_ifu_ar_bits_qos = 4'h0; // @[ifu.scala 103:22]
  assign io_ifu_r_ready = 1'h1; // @[ifu.scala 103:22]
  assign io_iccm_dma_ecc_error = mem_ctl_io_iccm_dma_ecc_error; // @[ifu.scala 113:25]
  assign io_iccm_dma_rvalid = mem_ctl_io_iccm_dma_rvalid; // @[ifu.scala 114:22]
  assign io_iccm_dma_rdata = mem_ctl_io_iccm_dma_rdata; // @[ifu.scala 115:21]
  assign io_iccm_dma_rtag = mem_ctl_io_iccm_dma_rtag; // @[ifu.scala 116:20]
  assign io_iccm_ready = mem_ctl_io_iccm_ready; // @[ifu.scala 117:17]
  assign io_iccm_dma_sb_error = mem_ctl_io_iccm_dma_sb_error; // @[ifu.scala 118:24]
  assign mem_ctl_clock = clock;
  assign mem_ctl_reset = reset;
  assign mem_ctl_io_free_clk = io_free_clk; // @[ifu.scala 90:23]
  assign mem_ctl_io_active_clk = io_active_clk; // @[ifu.scala 91:25]
  assign mem_ctl_io_exu_flush_final = io_exu_flush_final; // @[ifu.scala 92:30]
  assign mem_ctl_io_dec_mem_ctrl_dec_tlu_flush_err_wb = io_ifu_dec_dec_mem_ctrl_dec_tlu_flush_err_wb; // @[ifu.scala 93:27]
  assign mem_ctl_io_dec_mem_ctrl_dec_tlu_i0_commit_cmt = io_ifu_dec_dec_mem_ctrl_dec_tlu_i0_commit_cmt; // @[ifu.scala 93:27]
  assign mem_ctl_io_dec_mem_ctrl_dec_tlu_force_halt = io_ifu_dec_dec_mem_ctrl_dec_tlu_force_halt; // @[ifu.scala 93:27]
  assign mem_ctl_io_dec_mem_ctrl_dec_tlu_fence_i_wb = io_ifu_dec_dec_mem_ctrl_dec_tlu_fence_i_wb; // @[ifu.scala 93:27]
  assign mem_ctl_io_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_wrdata = io_ifu_dec_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_wrdata; // @[ifu.scala 93:27]
  assign mem_ctl_io_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_dicawics = io_ifu_dec_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_dicawics; // @[ifu.scala 93:27]
  assign mem_ctl_io_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_rd_valid = io_ifu_dec_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_rd_valid; // @[ifu.scala 93:27]
  assign mem_ctl_io_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_wr_valid = io_ifu_dec_dec_mem_ctrl_dec_tlu_ic_diag_pkt_icache_wr_valid; // @[ifu.scala 93:27]
  assign mem_ctl_io_dec_mem_ctrl_dec_tlu_core_ecc_disable = io_ifu_dec_dec_mem_ctrl_dec_tlu_core_ecc_disable; // @[ifu.scala 93:27]
  assign mem_ctl_io_ifc_fetch_addr_bf = ifc_ctl_io_ifc_fetch_addr_bf; // @[ifu.scala 94:32]
  assign mem_ctl_io_ifc_fetch_uncacheable_bf = ifc_ctl_io_ifc_fetch_uncacheable_bf; // @[ifu.scala 95:39]
  assign mem_ctl_io_ifc_fetch_req_bf = ifc_ctl_io_ifc_fetch_req_bf; // @[ifu.scala 96:31]
  assign mem_ctl_io_ifc_fetch_req_bf_raw = ifc_ctl_io_ifc_fetch_req_bf_raw; // @[ifu.scala 97:35]
  assign mem_ctl_io_ifc_iccm_access_bf = ifc_ctl_io_ifc_iccm_access_bf; // @[ifu.scala 98:33]
  assign mem_ctl_io_ifc_region_acc_fault_bf = ifc_ctl_io_ifc_region_acc_fault_bf; // @[ifu.scala 99:38]
  assign mem_ctl_io_ifc_dma_access_ok = ifc_ctl_io_ifc_dma_access_ok; // @[ifu.scala 100:32]
  assign mem_ctl_io_ifu_bp_hit_taken_f = bp_ctl_io_ifu_bp_hit_taken_f; // @[ifu.scala 101:33]
  assign mem_ctl_io_ifu_bp_inst_mask_f = bp_ctl_io_ifu_bp_inst_mask_f; // @[ifu.scala 102:33]
  assign mem_ctl_io_ifu_axi_ar_ready = io_ifu_ar_ready; // @[ifu.scala 103:22]
  assign mem_ctl_io_ifu_axi_r_valid = io_ifu_r_valid; // @[ifu.scala 103:22]
  assign mem_ctl_io_ifu_axi_r_bits_id = io_ifu_r_bits_id; // @[ifu.scala 103:22]
  assign mem_ctl_io_ifu_axi_r_bits_data = io_ifu_r_bits_data; // @[ifu.scala 103:22]
  assign mem_ctl_io_ifu_axi_r_bits_resp = io_ifu_r_bits_resp; // @[ifu.scala 103:22]
  assign mem_ctl_io_ifu_bus_clk_en = io_ifu_bus_clk_en; // @[ifu.scala 104:29]
  assign mem_ctl_io_dma_mem_ctl_dma_iccm_req = io_ifu_dma_dma_mem_ctl_dma_iccm_req; // @[ifu.scala 105:26]
  assign mem_ctl_io_dma_mem_ctl_dma_mem_addr = io_ifu_dma_dma_mem_ctl_dma_mem_addr; // @[ifu.scala 105:26]
  assign mem_ctl_io_dma_mem_ctl_dma_mem_sz = io_ifu_dma_dma_mem_ctl_dma_mem_sz; // @[ifu.scala 105:26]
  assign mem_ctl_io_dma_mem_ctl_dma_mem_write = io_ifu_dma_dma_mem_ctl_dma_mem_write; // @[ifu.scala 105:26]
  assign mem_ctl_io_dma_mem_ctl_dma_mem_wdata = io_ifu_dma_dma_mem_ctl_dma_mem_wdata; // @[ifu.scala 105:26]
  assign mem_ctl_io_dma_mem_ctl_dma_mem_tag = io_ifu_dma_dma_mem_ctl_dma_mem_tag; // @[ifu.scala 105:26]
  assign mem_ctl_io_iccm_rd_data = io_iccm_rd_data; // @[ifu.scala 107:19]
  assign mem_ctl_io_iccm_rd_data_ecc = io_iccm_rd_data_ecc; // @[ifu.scala 107:19]
  assign mem_ctl_io_ic_rd_data = io_ic_rd_data; // @[ifu.scala 106:17]
  assign mem_ctl_io_ic_debug_rd_data = io_ic_debug_rd_data; // @[ifu.scala 106:17]
  assign mem_ctl_io_ic_tag_debug_rd_data = io_ic_tag_debug_rd_data; // @[ifu.scala 106:17]
  assign mem_ctl_io_ic_eccerr = io_ic_eccerr; // @[ifu.scala 106:17]
  assign mem_ctl_io_ic_rd_hit = io_ic_rd_hit; // @[ifu.scala 106:17]
  assign mem_ctl_io_ic_tag_perr = io_ic_tag_perr; // @[ifu.scala 106:17]
  assign mem_ctl_io_ifu_fetch_val = mem_ctl_io_ic_fetch_val_f; // @[ifu.scala 108:28]
  assign mem_ctl_io_dec_tlu_flush_lower_wb = io_dec_tlu_flush_lower_wb; // @[ifu.scala 109:37]
  assign mem_ctl_io_scan_mode = io_scan_mode; // @[ifu.scala 110:24]
  assign bp_ctl_clock = clock;
  assign bp_ctl_reset = reset;
  assign bp_ctl_io_active_clk = io_active_clk; // @[ifu.scala 80:24]
  assign bp_ctl_io_ic_hit_f = mem_ctl_io_ic_hit_f; // @[ifu.scala 81:22]
  assign bp_ctl_io_exu_flush_final = io_exu_flush_final; // @[ifu.scala 86:29]
  assign bp_ctl_io_ifc_fetch_addr_f = ifc_ctl_io_ifc_fetch_addr_f; // @[ifu.scala 82:30]
  assign bp_ctl_io_ifc_fetch_req_f = ifc_ctl_io_ifc_fetch_req_f; // @[ifu.scala 83:29]
  assign bp_ctl_io_dec_bp_dec_tlu_br0_r_pkt_valid = io_ifu_dec_dec_bp_dec_tlu_br0_r_pkt_valid; // @[ifu.scala 84:20]
  assign bp_ctl_io_dec_bp_dec_tlu_br0_r_pkt_bits_hist = io_ifu_dec_dec_bp_dec_tlu_br0_r_pkt_bits_hist; // @[ifu.scala 84:20]
  assign bp_ctl_io_dec_bp_dec_tlu_br0_r_pkt_bits_br_error = io_ifu_dec_dec_bp_dec_tlu_br0_r_pkt_bits_br_error; // @[ifu.scala 84:20]
  assign bp_ctl_io_dec_bp_dec_tlu_br0_r_pkt_bits_br_start_error = io_ifu_dec_dec_bp_dec_tlu_br0_r_pkt_bits_br_start_error; // @[ifu.scala 84:20]
  assign bp_ctl_io_dec_bp_dec_tlu_br0_r_pkt_bits_way = io_ifu_dec_dec_bp_dec_tlu_br0_r_pkt_bits_way; // @[ifu.scala 84:20]
  assign bp_ctl_io_dec_bp_dec_tlu_br0_r_pkt_bits_middle = io_ifu_dec_dec_bp_dec_tlu_br0_r_pkt_bits_middle; // @[ifu.scala 84:20]
  assign bp_ctl_io_dec_bp_dec_tlu_flush_leak_one_wb = io_ifu_dec_dec_bp_dec_tlu_flush_leak_one_wb; // @[ifu.scala 84:20]
  assign bp_ctl_io_dec_bp_dec_tlu_bpred_disable = io_ifu_dec_dec_bp_dec_tlu_bpred_disable; // @[ifu.scala 84:20]
  assign bp_ctl_io_dec_tlu_flush_lower_wb = io_dec_tlu_flush_lower_wb; // @[ifu.scala 87:36]
  assign bp_ctl_io_exu_bp_exu_i0_br_index_r = io_exu_ifu_exu_bp_exu_i0_br_index_r; // @[ifu.scala 85:20]
  assign bp_ctl_io_exu_bp_exu_i0_br_fghr_r = io_exu_ifu_exu_bp_exu_i0_br_fghr_r; // @[ifu.scala 85:20]
  assign bp_ctl_io_exu_bp_exu_mp_pkt_bits_misp = io_exu_ifu_exu_bp_exu_mp_pkt_bits_misp; // @[ifu.scala 85:20]
  assign bp_ctl_io_exu_bp_exu_mp_pkt_bits_ataken = io_exu_ifu_exu_bp_exu_mp_pkt_bits_ataken; // @[ifu.scala 85:20]
  assign bp_ctl_io_exu_bp_exu_mp_pkt_bits_boffset = io_exu_ifu_exu_bp_exu_mp_pkt_bits_boffset; // @[ifu.scala 85:20]
  assign bp_ctl_io_exu_bp_exu_mp_pkt_bits_pc4 = io_exu_ifu_exu_bp_exu_mp_pkt_bits_pc4; // @[ifu.scala 85:20]
  assign bp_ctl_io_exu_bp_exu_mp_pkt_bits_hist = io_exu_ifu_exu_bp_exu_mp_pkt_bits_hist; // @[ifu.scala 85:20]
  assign bp_ctl_io_exu_bp_exu_mp_pkt_bits_toffset = io_exu_ifu_exu_bp_exu_mp_pkt_bits_toffset; // @[ifu.scala 85:20]
  assign bp_ctl_io_exu_bp_exu_mp_pkt_bits_pcall = io_exu_ifu_exu_bp_exu_mp_pkt_bits_pcall; // @[ifu.scala 85:20]
  assign bp_ctl_io_exu_bp_exu_mp_pkt_bits_pret = io_exu_ifu_exu_bp_exu_mp_pkt_bits_pret; // @[ifu.scala 85:20]
  assign bp_ctl_io_exu_bp_exu_mp_pkt_bits_pja = io_exu_ifu_exu_bp_exu_mp_pkt_bits_pja; // @[ifu.scala 85:20]
  assign bp_ctl_io_exu_bp_exu_mp_pkt_bits_way = io_exu_ifu_exu_bp_exu_mp_pkt_bits_way; // @[ifu.scala 85:20]
  assign bp_ctl_io_exu_bp_exu_mp_eghr = io_exu_ifu_exu_bp_exu_mp_eghr; // @[ifu.scala 85:20]
  assign bp_ctl_io_exu_bp_exu_mp_fghr = io_exu_ifu_exu_bp_exu_mp_fghr; // @[ifu.scala 85:20]
  assign bp_ctl_io_exu_bp_exu_mp_index = io_exu_ifu_exu_bp_exu_mp_index; // @[ifu.scala 85:20]
  assign bp_ctl_io_exu_bp_exu_mp_btag = io_exu_ifu_exu_bp_exu_mp_btag; // @[ifu.scala 85:20]
  assign bp_ctl_io_scan_mode = io_scan_mode; // @[ifu.scala 79:23]
  assign aln_ctl_clock = clock;
  assign aln_ctl_reset = reset;
  assign aln_ctl_io_scan_mode = io_scan_mode; // @[ifu.scala 57:24]
  assign aln_ctl_io_active_clk = io_active_clk; // @[ifu.scala 58:25]
  assign aln_ctl_io_ifu_async_error_start = mem_ctl_io_ifu_async_error_start; // @[ifu.scala 59:36]
  assign aln_ctl_io_iccm_rd_ecc_double_err = mem_ctl_io_iccm_rd_ecc_double_err; // @[ifu.scala 60:37]
  assign aln_ctl_io_ic_access_fault_f = mem_ctl_io_ic_access_fault_f; // @[ifu.scala 61:32]
  assign aln_ctl_io_ic_access_fault_type_f = mem_ctl_io_ic_access_fault_type_f; // @[ifu.scala 62:37]
  assign aln_ctl_io_ifu_bp_fghr_f = bp_ctl_io_ifu_bp_fghr_f; // @[ifu.scala 63:28]
  assign aln_ctl_io_ifu_bp_btb_target_f = bp_ctl_io_ifu_bp_btb_target_f; // @[ifu.scala 64:34]
  assign aln_ctl_io_ifu_bp_poffset_f = bp_ctl_io_ifu_bp_poffset_f; // @[ifu.scala 65:31]
  assign aln_ctl_io_ifu_bp_hist0_f = bp_ctl_io_ifu_bp_hist0_f; // @[ifu.scala 66:29]
  assign aln_ctl_io_ifu_bp_hist1_f = bp_ctl_io_ifu_bp_hist1_f; // @[ifu.scala 67:29]
  assign aln_ctl_io_ifu_bp_pc4_f = bp_ctl_io_ifu_bp_pc4_f; // @[ifu.scala 68:27]
  assign aln_ctl_io_ifu_bp_way_f = bp_ctl_io_ifu_bp_way_f; // @[ifu.scala 69:27]
  assign aln_ctl_io_ifu_bp_valid_f = bp_ctl_io_ifu_bp_valid_f; // @[ifu.scala 70:29]
  assign aln_ctl_io_ifu_bp_ret_f = bp_ctl_io_ifu_bp_ret_f; // @[ifu.scala 71:27]
  assign aln_ctl_io_exu_flush_final = io_exu_flush_final; // @[ifu.scala 72:30]
  assign aln_ctl_io_dec_aln_aln_dec_dec_i0_decode_d = io_ifu_dec_dec_aln_aln_dec_dec_i0_decode_d; // @[ifu.scala 73:22]
  assign aln_ctl_io_ifu_fetch_data_f = mem_ctl_io_ic_data_f; // @[ifu.scala 74:31]
  assign aln_ctl_io_ifu_fetch_val = mem_ctl_io_ifu_fetch_val; // @[ifu.scala 75:28]
  assign aln_ctl_io_ifu_fetch_pc = ifc_ctl_io_ifc_fetch_addr_f; // @[ifu.scala 76:27]
  assign ifc_ctl_clock = clock;
  assign ifc_ctl_reset = reset;
  assign ifc_ctl_io_exu_flush_final = io_exu_flush_final; // @[ifu.scala 47:30]
  assign ifc_ctl_io_exu_flush_path_final = io_exu_flush_path_final; // @[ifu.scala 54:35]
  assign ifc_ctl_io_free_clk = io_free_clk; // @[ifu.scala 41:23]
  assign ifc_ctl_io_active_clk = io_active_clk; // @[ifu.scala 40:25]
  assign ifc_ctl_io_scan_mode = io_scan_mode; // @[ifu.scala 42:24]
  assign ifc_ctl_io_ic_hit_f = mem_ctl_io_ic_hit_f; // @[ifu.scala 43:23]
  assign ifc_ctl_io_ifu_ic_mb_empty = mem_ctl_io_ifu_ic_mb_empty; // @[ifu.scala 53:30]
  assign ifc_ctl_io_ifu_fb_consume1 = aln_ctl_io_ifu_fb_consume1; // @[ifu.scala 44:30]
  assign ifc_ctl_io_ifu_fb_consume2 = aln_ctl_io_ifu_fb_consume2; // @[ifu.scala 45:30]
  assign ifc_ctl_io_ifu_bp_hit_taken_f = bp_ctl_io_ifu_bp_hit_taken_f; // @[ifu.scala 48:33]
  assign ifc_ctl_io_ifu_bp_btb_target_f = bp_ctl_io_ifu_bp_btb_target_f; // @[ifu.scala 49:34]
  assign ifc_ctl_io_ic_dma_active = mem_ctl_io_ic_dma_active; // @[ifu.scala 50:28]
  assign ifc_ctl_io_ic_write_stall = mem_ctl_io_ic_write_stall; // @[ifu.scala 51:29]
  assign ifc_ctl_io_dec_ifc_dec_tlu_flush_noredir_wb = io_ifu_dec_dec_ifc_dec_tlu_flush_noredir_wb; // @[ifu.scala 46:22]
  assign ifc_ctl_io_dec_ifc_dec_tlu_mrac_ff = io_ifu_dec_dec_ifc_dec_tlu_mrac_ff; // @[ifu.scala 46:22]
  assign ifc_ctl_io_dma_ifc_dma_iccm_stall_any = io_ifu_dma_dma_ifc_dma_iccm_stall_any; // @[ifu.scala 52:22]
endmodule
